module basic_1500_15000_2000_15_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_1290,In_574);
and U1 (N_1,In_1311,In_15);
nor U2 (N_2,In_1190,In_349);
xor U3 (N_3,In_1449,In_930);
xor U4 (N_4,In_1452,In_255);
nor U5 (N_5,In_1416,In_265);
xor U6 (N_6,In_1045,In_1130);
nor U7 (N_7,In_617,In_1430);
nand U8 (N_8,In_205,In_174);
and U9 (N_9,In_308,In_1156);
nand U10 (N_10,In_778,In_852);
or U11 (N_11,In_1063,In_1424);
xnor U12 (N_12,In_1143,In_751);
xnor U13 (N_13,In_515,In_1378);
nand U14 (N_14,In_32,In_467);
and U15 (N_15,In_1056,In_1260);
nand U16 (N_16,In_632,In_61);
and U17 (N_17,In_714,In_779);
or U18 (N_18,In_1080,In_504);
or U19 (N_19,In_1330,In_109);
or U20 (N_20,In_815,In_411);
or U21 (N_21,In_1285,In_7);
nand U22 (N_22,In_301,In_548);
nand U23 (N_23,In_1134,In_837);
nor U24 (N_24,In_802,In_112);
or U25 (N_25,In_219,In_352);
or U26 (N_26,In_280,In_1137);
xnor U27 (N_27,In_323,In_908);
and U28 (N_28,In_1139,In_581);
or U29 (N_29,In_529,In_356);
nor U30 (N_30,In_478,In_1475);
or U31 (N_31,In_1297,In_1404);
and U32 (N_32,In_564,In_1493);
nor U33 (N_33,In_1453,In_596);
or U34 (N_34,In_1046,In_1293);
nand U35 (N_35,In_1103,In_1274);
and U36 (N_36,In_824,In_842);
and U37 (N_37,In_839,In_453);
nand U38 (N_38,In_279,In_995);
xor U39 (N_39,In_1286,In_223);
nor U40 (N_40,In_1494,In_909);
nor U41 (N_41,In_1272,In_1244);
nand U42 (N_42,In_10,In_1210);
nor U43 (N_43,In_106,In_860);
and U44 (N_44,In_388,In_892);
nand U45 (N_45,In_1024,In_1243);
xor U46 (N_46,In_281,In_984);
nand U47 (N_47,In_958,In_706);
nor U48 (N_48,In_1386,In_66);
or U49 (N_49,In_1257,In_787);
or U50 (N_50,In_1444,In_1474);
and U51 (N_51,In_215,In_1002);
nor U52 (N_52,In_9,In_236);
or U53 (N_53,In_641,In_1205);
nand U54 (N_54,In_383,In_364);
nor U55 (N_55,In_1270,In_1218);
nand U56 (N_56,In_677,In_1428);
or U57 (N_57,In_789,In_580);
or U58 (N_58,In_155,In_1202);
nor U59 (N_59,In_756,In_571);
and U60 (N_60,In_702,In_335);
xnor U61 (N_61,In_763,In_1248);
nand U62 (N_62,In_652,In_640);
and U63 (N_63,In_884,In_1402);
nand U64 (N_64,In_907,In_239);
or U65 (N_65,In_931,In_436);
and U66 (N_66,In_158,In_921);
and U67 (N_67,In_748,In_511);
nor U68 (N_68,In_493,In_287);
or U69 (N_69,In_116,In_587);
nand U70 (N_70,In_1390,In_613);
nor U71 (N_71,In_210,In_262);
and U72 (N_72,In_1368,In_363);
nor U73 (N_73,In_101,In_1069);
and U74 (N_74,In_1433,In_1066);
and U75 (N_75,In_822,In_890);
nand U76 (N_76,In_302,In_738);
nor U77 (N_77,In_26,In_711);
and U78 (N_78,In_148,In_694);
and U79 (N_79,In_1194,In_94);
and U80 (N_80,In_774,In_1454);
nand U81 (N_81,In_1085,In_259);
nor U82 (N_82,In_877,In_1089);
and U83 (N_83,In_1229,In_163);
nand U84 (N_84,In_537,In_24);
nand U85 (N_85,In_85,In_807);
and U86 (N_86,In_497,In_875);
or U87 (N_87,In_573,In_570);
nor U88 (N_88,In_403,In_41);
nand U89 (N_89,In_1353,In_235);
nand U90 (N_90,In_1135,In_618);
nor U91 (N_91,In_601,In_326);
or U92 (N_92,In_1015,In_894);
nor U93 (N_93,In_556,In_1017);
or U94 (N_94,In_956,In_568);
nand U95 (N_95,In_1359,In_1414);
nand U96 (N_96,In_18,In_283);
and U97 (N_97,In_1365,In_321);
nand U98 (N_98,In_713,In_462);
nor U99 (N_99,In_635,In_126);
nor U100 (N_100,In_1140,In_91);
nor U101 (N_101,In_737,In_624);
and U102 (N_102,In_656,In_167);
and U103 (N_103,In_594,In_1413);
or U104 (N_104,In_1262,In_1355);
nand U105 (N_105,In_274,In_1049);
and U106 (N_106,In_1060,In_217);
nand U107 (N_107,In_30,In_951);
nand U108 (N_108,In_1282,In_1005);
nor U109 (N_109,In_912,In_1484);
nand U110 (N_110,In_999,In_685);
nand U111 (N_111,In_145,In_535);
or U112 (N_112,In_1079,In_1228);
nand U113 (N_113,In_496,In_809);
or U114 (N_114,In_803,In_676);
or U115 (N_115,In_1022,In_1201);
nor U116 (N_116,In_211,In_128);
nand U117 (N_117,In_1102,In_1332);
xnor U118 (N_118,In_290,In_943);
nand U119 (N_119,In_297,In_608);
or U120 (N_120,In_1233,In_1232);
nor U121 (N_121,In_81,In_1457);
and U122 (N_122,In_20,In_1235);
or U123 (N_123,In_733,In_1356);
nand U124 (N_124,In_143,In_382);
nand U125 (N_125,In_46,In_1168);
and U126 (N_126,In_394,In_992);
and U127 (N_127,In_151,In_147);
or U128 (N_128,In_1059,In_893);
and U129 (N_129,In_1187,In_1048);
and U130 (N_130,In_793,In_589);
and U131 (N_131,In_73,In_65);
nand U132 (N_132,In_567,In_819);
and U133 (N_133,In_1061,In_432);
and U134 (N_134,In_123,In_207);
and U135 (N_135,In_164,In_1068);
nand U136 (N_136,In_75,In_827);
xor U137 (N_137,In_764,In_1468);
and U138 (N_138,In_1411,In_1128);
nand U139 (N_139,In_740,In_649);
and U140 (N_140,In_1223,In_213);
nand U141 (N_141,In_525,In_272);
or U142 (N_142,In_904,In_1379);
or U143 (N_143,In_533,In_1088);
and U144 (N_144,In_555,In_28);
nor U145 (N_145,In_304,In_707);
and U146 (N_146,In_821,In_722);
and U147 (N_147,In_1154,In_410);
nor U148 (N_148,In_43,In_776);
nand U149 (N_149,In_1307,In_362);
or U150 (N_150,In_1276,In_922);
xor U151 (N_151,In_396,In_959);
nor U152 (N_152,In_329,In_476);
or U153 (N_153,In_712,In_704);
nand U154 (N_154,In_437,In_266);
nand U155 (N_155,In_1211,In_1105);
nor U156 (N_156,In_1279,In_332);
nand U157 (N_157,In_448,In_257);
and U158 (N_158,In_103,In_473);
or U159 (N_159,In_1169,In_1072);
and U160 (N_160,In_623,In_784);
xor U161 (N_161,In_683,In_1123);
nor U162 (N_162,In_1148,In_645);
nor U163 (N_163,In_275,In_923);
or U164 (N_164,In_343,In_1343);
and U165 (N_165,In_680,In_34);
xor U166 (N_166,In_1147,In_1398);
and U167 (N_167,In_434,In_267);
or U168 (N_168,In_1497,In_810);
nand U169 (N_169,In_173,In_1462);
nand U170 (N_170,In_626,In_206);
xnor U171 (N_171,In_67,In_871);
nor U172 (N_172,In_709,In_1395);
nand U173 (N_173,In_854,In_340);
xnor U174 (N_174,In_840,In_186);
nor U175 (N_175,In_1142,In_1141);
nor U176 (N_176,In_781,In_1166);
or U177 (N_177,In_138,In_527);
xor U178 (N_178,In_851,In_331);
nor U179 (N_179,In_725,In_643);
or U180 (N_180,In_430,In_818);
xnor U181 (N_181,In_197,In_203);
and U182 (N_182,In_1153,In_1408);
and U183 (N_183,In_228,In_1070);
or U184 (N_184,In_180,In_1363);
xnor U185 (N_185,In_175,In_187);
or U186 (N_186,In_1186,In_455);
and U187 (N_187,In_532,In_1100);
nor U188 (N_188,In_1351,In_928);
nor U189 (N_189,In_687,In_146);
nor U190 (N_190,In_628,In_517);
nand U191 (N_191,In_1062,In_19);
or U192 (N_192,In_1401,In_288);
xor U193 (N_193,In_76,In_1361);
or U194 (N_194,In_1222,In_140);
xor U195 (N_195,In_226,In_440);
nor U196 (N_196,In_1319,In_1393);
xnor U197 (N_197,In_745,In_407);
and U198 (N_198,In_378,In_337);
nand U199 (N_199,In_769,In_1239);
or U200 (N_200,In_51,In_398);
nand U201 (N_201,In_54,In_463);
and U202 (N_202,In_944,In_1426);
or U203 (N_203,In_193,In_154);
and U204 (N_204,In_541,In_873);
nand U205 (N_205,In_625,In_479);
nor U206 (N_206,In_653,In_823);
nor U207 (N_207,In_242,In_1241);
nand U208 (N_208,In_987,In_796);
or U209 (N_209,In_830,In_1008);
nand U210 (N_210,In_744,In_520);
and U211 (N_211,In_289,In_234);
nor U212 (N_212,In_674,In_868);
or U213 (N_213,In_1051,In_710);
nor U214 (N_214,In_1338,In_342);
and U215 (N_215,In_152,In_1138);
and U216 (N_216,In_124,In_1479);
xor U217 (N_217,In_1344,In_572);
and U218 (N_218,In_508,In_499);
nand U219 (N_219,In_661,In_536);
xor U220 (N_220,In_982,In_1380);
nand U221 (N_221,In_545,In_976);
nor U222 (N_222,In_669,In_1224);
nor U223 (N_223,In_450,In_48);
or U224 (N_224,In_277,In_3);
or U225 (N_225,In_948,In_1026);
nor U226 (N_226,In_616,In_954);
and U227 (N_227,In_1461,In_346);
and U228 (N_228,In_178,In_222);
nand U229 (N_229,In_1477,In_129);
xnor U230 (N_230,In_708,In_451);
or U231 (N_231,In_1498,In_1030);
xor U232 (N_232,In_1346,In_35);
xnor U233 (N_233,In_752,In_1055);
nand U234 (N_234,In_1324,In_1388);
nor U235 (N_235,In_528,In_736);
nor U236 (N_236,In_1434,In_421);
nor U237 (N_237,In_916,In_699);
nand U238 (N_238,In_1259,In_629);
or U239 (N_239,In_620,In_972);
nor U240 (N_240,In_507,In_454);
nor U241 (N_241,In_631,In_1432);
xor U242 (N_242,In_978,In_732);
nand U243 (N_243,In_1298,In_208);
and U244 (N_244,In_1458,In_93);
nand U245 (N_245,In_229,In_1001);
or U246 (N_246,In_575,In_719);
xor U247 (N_247,In_874,In_1039);
nand U248 (N_248,In_1418,In_115);
and U249 (N_249,In_171,In_4);
and U250 (N_250,In_1170,In_1409);
nor U251 (N_251,In_934,In_509);
nor U252 (N_252,In_1410,In_1083);
and U253 (N_253,In_953,In_371);
or U254 (N_254,In_731,In_64);
or U255 (N_255,In_1094,In_622);
and U256 (N_256,In_381,In_1372);
and U257 (N_257,In_1250,In_979);
and U258 (N_258,In_829,In_1383);
nand U259 (N_259,In_715,In_1315);
xnor U260 (N_260,In_768,In_1016);
xnor U261 (N_261,In_244,In_241);
and U262 (N_262,In_303,In_986);
or U263 (N_263,In_470,In_159);
nand U264 (N_264,In_1073,In_1289);
and U265 (N_265,In_402,In_602);
nand U266 (N_266,In_552,In_71);
or U267 (N_267,In_718,In_384);
nand U268 (N_268,In_400,In_1172);
and U269 (N_269,In_1028,In_965);
nand U270 (N_270,In_1448,In_232);
or U271 (N_271,In_240,In_1119);
or U272 (N_272,In_1336,In_518);
or U273 (N_273,In_1352,In_578);
nand U274 (N_274,In_1249,In_646);
nand U275 (N_275,In_316,In_1436);
nand U276 (N_276,In_1376,In_1339);
nand U277 (N_277,In_498,In_866);
nand U278 (N_278,In_322,In_2);
and U279 (N_279,In_1165,In_772);
nand U280 (N_280,In_313,In_1482);
nor U281 (N_281,In_1267,In_881);
and U282 (N_282,In_1242,In_1167);
or U283 (N_283,In_1121,In_404);
nor U284 (N_284,In_121,In_1132);
nor U285 (N_285,In_651,In_1082);
or U286 (N_286,In_963,In_831);
xnor U287 (N_287,In_878,In_1440);
nor U288 (N_288,In_896,In_260);
and U289 (N_289,In_834,In_642);
nand U290 (N_290,In_826,In_538);
and U291 (N_291,In_671,In_1120);
nand U292 (N_292,In_937,In_565);
or U293 (N_293,In_856,In_1090);
nor U294 (N_294,In_27,In_513);
nand U295 (N_295,In_1175,In_1313);
nand U296 (N_296,In_424,In_1163);
nor U297 (N_297,In_1360,In_488);
nor U298 (N_298,In_1198,In_734);
nor U299 (N_299,In_443,In_876);
and U300 (N_300,In_862,In_870);
and U301 (N_301,In_87,In_50);
xnor U302 (N_302,In_551,In_1225);
nor U303 (N_303,In_1234,In_735);
or U304 (N_304,In_788,In_561);
nor U305 (N_305,In_315,In_785);
xor U306 (N_306,In_848,In_1450);
and U307 (N_307,In_78,In_659);
or U308 (N_308,In_1397,In_836);
nor U309 (N_309,In_318,In_1369);
or U310 (N_310,In_531,In_347);
and U311 (N_311,In_117,In_1115);
and U312 (N_312,In_294,In_863);
nor U313 (N_313,In_119,In_114);
nor U314 (N_314,In_1320,In_899);
and U315 (N_315,In_1392,In_1111);
or U316 (N_316,In_365,In_1335);
nor U317 (N_317,In_144,In_353);
and U318 (N_318,In_425,In_1269);
nor U319 (N_319,In_29,In_1176);
or U320 (N_320,In_1081,In_1299);
nand U321 (N_321,In_721,In_929);
nand U322 (N_322,In_177,In_1427);
nor U323 (N_323,In_584,In_1020);
nand U324 (N_324,In_780,In_1252);
nor U325 (N_325,In_150,In_729);
and U326 (N_326,In_369,In_585);
nor U327 (N_327,In_1271,In_1181);
or U328 (N_328,In_1192,In_988);
nor U329 (N_329,In_1253,In_549);
and U330 (N_330,In_1464,In_662);
and U331 (N_331,In_1152,In_475);
xor U332 (N_332,In_1441,In_113);
and U333 (N_333,In_761,In_1033);
xor U334 (N_334,In_554,In_1196);
or U335 (N_335,In_942,In_137);
xor U336 (N_336,In_569,In_980);
and U337 (N_337,In_915,In_1263);
and U338 (N_338,In_122,In_981);
or U339 (N_339,In_841,In_1219);
xor U340 (N_340,In_1097,In_975);
or U341 (N_341,In_563,In_1345);
or U342 (N_342,In_136,In_1358);
nor U343 (N_343,In_1291,In_1264);
xor U344 (N_344,In_540,In_654);
nor U345 (N_345,In_1240,In_1326);
xor U346 (N_346,In_926,In_665);
nor U347 (N_347,In_200,In_867);
nor U348 (N_348,In_1419,In_859);
or U349 (N_349,In_273,In_1422);
nor U350 (N_350,In_149,In_547);
or U351 (N_351,In_698,In_750);
or U352 (N_352,In_1389,In_231);
and U353 (N_353,In_1146,In_1483);
nand U354 (N_354,In_1306,In_298);
and U355 (N_355,In_728,In_1273);
nand U356 (N_356,In_345,In_118);
nand U357 (N_357,In_1179,In_1041);
or U358 (N_358,In_647,In_1268);
xnor U359 (N_359,In_947,In_1215);
nand U360 (N_360,In_83,In_1220);
nor U361 (N_361,In_1400,In_1178);
nor U362 (N_362,In_1124,In_1310);
and U363 (N_363,In_832,In_582);
xnor U364 (N_364,In_271,In_247);
nand U365 (N_365,In_162,In_773);
nand U366 (N_366,In_595,In_955);
nand U367 (N_367,In_883,In_1157);
and U368 (N_368,In_757,In_1029);
nor U369 (N_369,In_753,In_1396);
or U370 (N_370,In_1495,In_742);
nand U371 (N_371,In_791,In_330);
nand U372 (N_372,In_477,In_268);
xnor U373 (N_373,In_586,In_293);
and U374 (N_374,In_1478,In_1357);
nand U375 (N_375,In_825,In_361);
nor U376 (N_376,In_1042,In_1321);
xor U377 (N_377,In_389,In_726);
and U378 (N_378,In_605,In_797);
or U379 (N_379,In_1460,In_449);
or U380 (N_380,In_419,In_135);
nand U381 (N_381,In_1074,In_189);
nand U382 (N_382,In_990,In_1496);
and U383 (N_383,In_1314,In_49);
and U384 (N_384,In_1277,In_510);
or U385 (N_385,In_716,In_320);
xnor U386 (N_386,In_47,In_1375);
nand U387 (N_387,In_1000,In_98);
nand U388 (N_388,In_319,In_755);
nand U389 (N_389,In_1305,In_348);
nand U390 (N_390,In_1213,In_392);
nor U391 (N_391,In_58,In_1384);
xor U392 (N_392,In_254,In_458);
or U393 (N_393,In_747,In_1151);
and U394 (N_394,In_486,In_13);
and U395 (N_395,In_1144,In_805);
nor U396 (N_396,In_1447,In_949);
or U397 (N_397,In_427,In_435);
nand U398 (N_398,In_1399,In_1013);
or U399 (N_399,In_633,In_393);
or U400 (N_400,In_77,In_960);
nand U401 (N_401,In_428,In_1471);
nor U402 (N_402,In_355,In_1499);
or U403 (N_403,In_816,In_760);
nor U404 (N_404,In_96,In_366);
and U405 (N_405,In_1387,In_120);
nand U406 (N_406,In_739,In_37);
and U407 (N_407,In_270,In_684);
or U408 (N_408,In_1214,In_553);
xor U409 (N_409,In_246,In_1126);
nor U410 (N_410,In_1117,In_306);
and U411 (N_411,In_1467,In_1431);
nor U412 (N_412,In_1131,In_1221);
nand U413 (N_413,In_1231,In_1304);
and U414 (N_414,In_1093,In_472);
nor U415 (N_415,In_1266,In_1246);
and U416 (N_416,In_172,In_21);
xnor U417 (N_417,In_373,In_1067);
nand U418 (N_418,In_17,In_1300);
nand U419 (N_419,In_190,In_1200);
and U420 (N_420,In_970,In_1364);
nor U421 (N_421,In_406,In_994);
or U422 (N_422,In_317,In_22);
nand U423 (N_423,In_192,In_1287);
xor U424 (N_424,In_813,In_974);
and U425 (N_425,In_1182,In_1108);
and U426 (N_426,In_1018,In_898);
nand U427 (N_427,In_471,In_1295);
nand U428 (N_428,In_847,In_195);
or U429 (N_429,In_1208,In_102);
and U430 (N_430,In_237,In_1366);
nor U431 (N_431,In_940,In_790);
and U432 (N_432,In_689,In_1096);
nand U433 (N_433,In_99,In_166);
or U434 (N_434,In_679,In_559);
nor U435 (N_435,In_1340,In_461);
and U436 (N_436,In_438,In_501);
and U437 (N_437,In_880,In_693);
or U438 (N_438,In_1199,In_1114);
nor U439 (N_439,In_278,In_1036);
or U440 (N_440,In_433,In_184);
nand U441 (N_441,In_957,In_45);
and U442 (N_442,In_1044,In_1207);
xor U443 (N_443,In_74,In_989);
and U444 (N_444,In_638,In_199);
nor U445 (N_445,In_133,In_25);
nor U446 (N_446,In_1382,In_221);
or U447 (N_447,In_1329,In_439);
or U448 (N_448,In_445,In_284);
and U449 (N_449,In_296,In_160);
nor U450 (N_450,In_416,In_1209);
and U451 (N_451,In_194,In_1334);
or U452 (N_452,In_1322,In_1443);
xnor U453 (N_453,In_380,In_606);
or U454 (N_454,In_849,In_1349);
nor U455 (N_455,In_490,In_973);
nand U456 (N_456,In_224,In_249);
nand U457 (N_457,In_1309,In_512);
and U458 (N_458,In_253,In_610);
xor U459 (N_459,In_469,In_985);
nor U460 (N_460,In_614,In_183);
and U461 (N_461,In_991,In_385);
nand U462 (N_462,In_1057,In_1158);
or U463 (N_463,In_1003,In_80);
nor U464 (N_464,In_1227,In_794);
or U465 (N_465,In_933,In_557);
xor U466 (N_466,In_672,In_1116);
nor U467 (N_467,In_59,In_1161);
nand U468 (N_468,In_1405,In_1420);
nor U469 (N_469,In_749,In_1037);
nor U470 (N_470,In_786,In_341);
xor U471 (N_471,In_534,In_946);
nand U472 (N_472,In_983,In_1381);
or U473 (N_473,In_405,In_92);
and U474 (N_474,In_86,In_1183);
or U475 (N_475,In_777,In_359);
xor U476 (N_476,In_452,In_920);
nand U477 (N_477,In_1237,In_544);
nand U478 (N_478,In_727,In_182);
xnor U479 (N_479,In_723,In_492);
nand U480 (N_480,In_579,In_1010);
nand U481 (N_481,In_932,In_324);
nand U482 (N_482,In_607,In_1456);
or U483 (N_483,In_703,In_1367);
nor U484 (N_484,In_1180,In_1446);
nand U485 (N_485,In_351,In_1455);
and U486 (N_486,In_1328,In_724);
nor U487 (N_487,In_741,In_484);
or U488 (N_488,In_1469,In_1058);
or U489 (N_489,In_667,In_1261);
nand U490 (N_490,In_1347,In_168);
nor U491 (N_491,In_397,In_1492);
xnor U492 (N_492,In_619,In_924);
and U493 (N_493,In_339,In_38);
and U494 (N_494,In_127,In_141);
nand U495 (N_495,In_1417,In_717);
nor U496 (N_496,In_169,In_442);
or U497 (N_497,In_52,In_1265);
nand U498 (N_498,In_1312,In_792);
nand U499 (N_499,In_40,In_902);
nor U500 (N_500,In_310,In_901);
and U501 (N_501,In_196,In_1423);
and U502 (N_502,In_1341,In_446);
or U503 (N_503,In_368,In_670);
nor U504 (N_504,In_1323,In_426);
or U505 (N_505,In_686,In_459);
nor U506 (N_506,In_1129,In_1318);
or U507 (N_507,In_97,In_179);
or U508 (N_508,In_105,In_1193);
or U509 (N_509,In_746,In_521);
and U510 (N_510,In_63,In_220);
nand U511 (N_511,In_357,In_691);
and U512 (N_512,In_1155,In_16);
or U513 (N_513,In_1303,In_636);
and U514 (N_514,In_1480,In_634);
nor U515 (N_515,In_576,In_12);
nand U516 (N_516,In_1204,In_1019);
xnor U517 (N_517,In_603,In_648);
nand U518 (N_518,In_82,In_1316);
nor U519 (N_519,In_1333,In_60);
nor U520 (N_520,In_664,In_771);
nand U521 (N_521,In_360,In_1197);
nor U522 (N_522,In_1487,In_358);
nand U523 (N_523,In_925,In_543);
nand U524 (N_524,In_1302,In_887);
nand U525 (N_525,In_165,In_914);
nand U526 (N_526,In_1251,In_524);
or U527 (N_527,In_420,In_95);
nor U528 (N_528,In_869,In_456);
nor U529 (N_529,In_1133,In_1040);
nor U530 (N_530,In_814,In_765);
xnor U531 (N_531,In_198,In_1177);
and U532 (N_532,In_1491,In_1075);
nor U533 (N_533,In_344,In_0);
and U534 (N_534,In_754,In_1439);
nor U535 (N_535,In_1189,In_387);
or U536 (N_536,In_375,In_811);
nand U537 (N_537,In_336,In_374);
or U538 (N_538,In_853,In_377);
or U539 (N_539,In_692,In_441);
xor U540 (N_540,In_1007,In_1226);
nand U541 (N_541,In_828,In_844);
nor U542 (N_542,In_952,In_390);
nor U543 (N_543,In_464,In_1348);
or U544 (N_544,In_526,In_314);
nor U545 (N_545,In_285,In_56);
nand U546 (N_546,In_903,In_225);
and U547 (N_547,In_305,In_615);
nor U548 (N_548,In_62,In_282);
nand U549 (N_549,In_1473,In_1109);
xnor U550 (N_550,In_885,In_1053);
and U551 (N_551,In_855,In_566);
nor U552 (N_552,In_1195,In_245);
nand U553 (N_553,In_1415,In_1113);
nand U554 (N_554,In_977,In_1127);
nor U555 (N_555,In_1486,In_660);
xnor U556 (N_556,In_31,In_964);
nand U557 (N_557,In_1125,In_993);
or U558 (N_558,In_412,In_291);
nor U559 (N_559,In_1403,In_70);
or U560 (N_560,In_1281,In_546);
nor U561 (N_561,In_338,In_1275);
or U562 (N_562,In_1354,In_1006);
nand U563 (N_563,In_422,In_663);
nand U564 (N_564,In_1350,In_637);
nand U565 (N_565,In_759,In_514);
or U566 (N_566,In_139,In_423);
or U567 (N_567,In_72,In_299);
nand U568 (N_568,In_804,In_966);
and U569 (N_569,In_997,In_465);
and U570 (N_570,In_444,In_1301);
nor U571 (N_571,In_838,In_370);
nor U572 (N_572,In_1407,In_1145);
nor U573 (N_573,In_1481,In_417);
and U574 (N_574,In_202,In_1136);
and U575 (N_575,In_882,In_474);
nor U576 (N_576,In_429,In_485);
or U577 (N_577,In_530,In_644);
xor U578 (N_578,In_678,In_230);
or U579 (N_579,In_212,In_906);
nand U580 (N_580,In_1027,In_111);
and U581 (N_581,In_1076,In_650);
nor U582 (N_582,In_812,In_487);
xnor U583 (N_583,In_730,In_658);
xnor U584 (N_584,In_1043,In_57);
or U585 (N_585,In_950,In_481);
or U586 (N_586,In_895,In_1490);
and U587 (N_587,In_775,In_800);
nor U588 (N_588,In_1064,In_269);
nand U589 (N_589,In_612,In_1071);
nand U590 (N_590,In_391,In_1031);
or U591 (N_591,In_483,In_798);
xnor U592 (N_592,In_295,In_592);
xnor U593 (N_593,In_131,In_506);
nand U594 (N_594,In_1374,In_666);
or U595 (N_595,In_379,In_157);
nor U596 (N_596,In_558,In_604);
and U597 (N_597,In_783,In_5);
nor U598 (N_598,In_1283,In_491);
nor U599 (N_599,In_1278,In_132);
or U600 (N_600,In_701,In_1425);
nor U601 (N_601,In_1164,In_44);
or U602 (N_602,In_1445,In_1470);
nand U603 (N_603,In_767,In_597);
and U604 (N_604,In_897,In_1421);
nand U605 (N_605,In_1438,In_1106);
nand U606 (N_606,In_286,In_1203);
nor U607 (N_607,In_100,In_562);
xnor U608 (N_608,In_657,In_1065);
and U609 (N_609,In_399,In_918);
nand U610 (N_610,In_1412,In_1466);
nor U611 (N_611,In_681,In_53);
nor U612 (N_612,In_1451,In_945);
and U613 (N_613,In_516,In_758);
nor U614 (N_614,In_845,In_1485);
nand U615 (N_615,In_1254,In_806);
nor U616 (N_616,In_1038,In_505);
or U617 (N_617,In_1023,In_590);
xor U618 (N_618,In_621,In_996);
or U619 (N_619,In_415,In_1217);
xnor U620 (N_620,In_539,In_1118);
and U621 (N_621,In_191,In_1296);
and U622 (N_622,In_550,In_846);
and U623 (N_623,In_334,In_1212);
nand U624 (N_624,In_1084,In_1337);
nor U625 (N_625,In_204,In_770);
and U626 (N_626,In_256,In_372);
and U627 (N_627,In_913,In_705);
or U628 (N_628,In_872,In_1032);
nand U629 (N_629,In_494,In_1371);
nand U630 (N_630,In_69,In_201);
or U631 (N_631,In_560,In_968);
or U632 (N_632,In_1184,In_327);
nor U633 (N_633,In_248,In_1236);
or U634 (N_634,In_820,In_1391);
or U635 (N_635,In_14,In_107);
and U636 (N_636,In_1160,In_181);
and U637 (N_637,In_176,In_480);
and U638 (N_638,In_1370,In_835);
or U639 (N_639,In_865,In_1034);
and U640 (N_640,In_1047,In_23);
nor U641 (N_641,In_1280,In_905);
or U642 (N_642,In_591,In_1077);
nor U643 (N_643,In_1292,In_598);
nor U644 (N_644,In_682,In_599);
nand U645 (N_645,In_1101,In_697);
and U646 (N_646,In_1054,In_695);
nand U647 (N_647,In_639,In_376);
xnor U648 (N_648,In_690,In_418);
and U649 (N_649,In_495,In_743);
and U650 (N_650,In_1004,In_917);
and U651 (N_651,In_1406,In_90);
nor U652 (N_652,In_1377,In_1238);
nand U653 (N_653,In_888,In_1488);
nand U654 (N_654,In_1206,In_864);
nor U655 (N_655,In_588,In_600);
or U656 (N_656,In_466,In_1191);
nand U657 (N_657,In_89,In_503);
nand U658 (N_658,In_311,In_8);
or U659 (N_659,In_900,In_1112);
or U660 (N_660,In_1091,In_1050);
nor U661 (N_661,In_696,In_1162);
xnor U662 (N_662,In_1325,In_42);
xnor U663 (N_663,In_939,In_457);
nand U664 (N_664,In_542,In_1078);
xor U665 (N_665,In_108,In_1104);
nor U666 (N_666,In_250,In_261);
or U667 (N_667,In_431,In_238);
nand U668 (N_668,In_523,In_68);
nor U669 (N_669,In_276,In_1442);
and U670 (N_670,In_891,In_971);
nand U671 (N_671,In_1173,In_6);
nor U672 (N_672,In_1245,In_627);
nand U673 (N_673,In_482,In_1472);
nor U674 (N_674,In_1342,In_468);
or U675 (N_675,In_833,In_263);
nor U676 (N_676,In_962,In_251);
or U677 (N_677,In_1107,In_401);
and U678 (N_678,In_762,In_1476);
nand U679 (N_679,In_170,In_1284);
nor U680 (N_680,In_1394,In_998);
or U681 (N_681,In_1014,In_1150);
or U682 (N_682,In_500,In_782);
or U683 (N_683,In_1086,In_1465);
or U684 (N_684,In_1437,In_886);
nand U685 (N_685,In_911,In_395);
nor U686 (N_686,In_307,In_1216);
nand U687 (N_687,In_1098,In_583);
nor U688 (N_688,In_1308,In_1362);
and U689 (N_689,In_1122,In_88);
nor U690 (N_690,In_408,In_969);
nand U691 (N_691,In_39,In_312);
nor U692 (N_692,In_214,In_227);
nand U693 (N_693,In_134,In_967);
nor U694 (N_694,In_879,In_209);
nor U695 (N_695,In_153,In_367);
nand U696 (N_696,In_328,In_1052);
nand U697 (N_697,In_1021,In_1463);
and U698 (N_698,In_447,In_325);
xnor U699 (N_699,In_522,In_218);
and U700 (N_700,In_1435,In_808);
or U701 (N_701,In_354,In_33);
and U702 (N_702,In_910,In_188);
or U703 (N_703,In_300,In_1247);
or U704 (N_704,In_216,In_1258);
nor U705 (N_705,In_36,In_795);
and U706 (N_706,In_1331,In_11);
nor U707 (N_707,In_611,In_1317);
nand U708 (N_708,In_1087,In_519);
nor U709 (N_709,In_1095,In_577);
nand U710 (N_710,In_104,In_84);
nand U711 (N_711,In_1429,In_889);
and U712 (N_712,In_292,In_258);
or U713 (N_713,In_688,In_1171);
or U714 (N_714,In_1294,In_55);
nor U715 (N_715,In_673,In_161);
nand U716 (N_716,In_936,In_668);
nand U717 (N_717,In_79,In_413);
nor U718 (N_718,In_386,In_1489);
and U719 (N_719,In_243,In_333);
and U720 (N_720,In_1092,In_1230);
nand U721 (N_721,In_630,In_843);
and U722 (N_722,In_1373,In_799);
or U723 (N_723,In_700,In_1159);
or U724 (N_724,In_1099,In_1385);
and U725 (N_725,In_801,In_264);
nor U726 (N_726,In_414,In_927);
and U727 (N_727,In_938,In_350);
and U728 (N_728,In_850,In_935);
and U729 (N_729,In_861,In_1035);
nand U730 (N_730,In_1011,In_489);
and U731 (N_731,In_142,In_1256);
nand U732 (N_732,In_720,In_675);
and U733 (N_733,In_185,In_1255);
nand U734 (N_734,In_609,In_1185);
nor U735 (N_735,In_130,In_110);
and U736 (N_736,In_1009,In_858);
or U737 (N_737,In_1459,In_1288);
and U738 (N_738,In_125,In_961);
nor U739 (N_739,In_655,In_1110);
xnor U740 (N_740,In_252,In_593);
or U741 (N_741,In_460,In_817);
nand U742 (N_742,In_941,In_1025);
nor U743 (N_743,In_1174,In_766);
or U744 (N_744,In_156,In_1188);
nand U745 (N_745,In_309,In_919);
or U746 (N_746,In_1,In_409);
or U747 (N_747,In_857,In_233);
nor U748 (N_748,In_1012,In_1149);
nor U749 (N_749,In_502,In_1327);
or U750 (N_750,In_849,In_1487);
nor U751 (N_751,In_87,In_1038);
and U752 (N_752,In_177,In_1201);
or U753 (N_753,In_635,In_1109);
and U754 (N_754,In_1224,In_1062);
and U755 (N_755,In_112,In_1314);
nor U756 (N_756,In_376,In_1310);
nor U757 (N_757,In_1494,In_45);
xnor U758 (N_758,In_720,In_48);
or U759 (N_759,In_476,In_955);
or U760 (N_760,In_3,In_585);
nor U761 (N_761,In_486,In_397);
or U762 (N_762,In_243,In_482);
nand U763 (N_763,In_367,In_169);
nor U764 (N_764,In_410,In_528);
and U765 (N_765,In_751,In_1241);
and U766 (N_766,In_212,In_704);
or U767 (N_767,In_337,In_836);
nand U768 (N_768,In_309,In_1485);
xnor U769 (N_769,In_436,In_1208);
nand U770 (N_770,In_271,In_403);
and U771 (N_771,In_894,In_827);
or U772 (N_772,In_925,In_889);
xnor U773 (N_773,In_733,In_1124);
or U774 (N_774,In_531,In_789);
or U775 (N_775,In_1059,In_1065);
and U776 (N_776,In_747,In_1081);
nand U777 (N_777,In_1324,In_862);
nor U778 (N_778,In_1356,In_1277);
nand U779 (N_779,In_806,In_51);
nor U780 (N_780,In_174,In_706);
or U781 (N_781,In_628,In_1029);
xor U782 (N_782,In_59,In_829);
xor U783 (N_783,In_776,In_70);
xnor U784 (N_784,In_550,In_1395);
nor U785 (N_785,In_1239,In_947);
nor U786 (N_786,In_648,In_206);
or U787 (N_787,In_1334,In_1439);
and U788 (N_788,In_795,In_956);
nor U789 (N_789,In_1410,In_1331);
nand U790 (N_790,In_1492,In_1203);
or U791 (N_791,In_420,In_845);
nor U792 (N_792,In_798,In_1061);
xnor U793 (N_793,In_842,In_1125);
and U794 (N_794,In_750,In_591);
nand U795 (N_795,In_581,In_95);
or U796 (N_796,In_1087,In_986);
and U797 (N_797,In_538,In_1189);
nor U798 (N_798,In_630,In_334);
xnor U799 (N_799,In_1164,In_1475);
and U800 (N_800,In_1437,In_874);
nor U801 (N_801,In_1088,In_509);
or U802 (N_802,In_64,In_993);
or U803 (N_803,In_499,In_1307);
nand U804 (N_804,In_36,In_1006);
nor U805 (N_805,In_1177,In_676);
nor U806 (N_806,In_1215,In_1465);
nand U807 (N_807,In_434,In_487);
nor U808 (N_808,In_356,In_189);
nor U809 (N_809,In_630,In_329);
and U810 (N_810,In_1137,In_1104);
nor U811 (N_811,In_131,In_1285);
or U812 (N_812,In_1329,In_301);
and U813 (N_813,In_196,In_1466);
and U814 (N_814,In_1261,In_511);
nand U815 (N_815,In_703,In_45);
or U816 (N_816,In_1221,In_722);
nand U817 (N_817,In_29,In_659);
and U818 (N_818,In_90,In_1254);
nor U819 (N_819,In_383,In_687);
or U820 (N_820,In_915,In_974);
nand U821 (N_821,In_178,In_693);
nor U822 (N_822,In_1024,In_216);
nor U823 (N_823,In_1208,In_29);
xnor U824 (N_824,In_1122,In_215);
xor U825 (N_825,In_904,In_616);
or U826 (N_826,In_1442,In_1106);
nand U827 (N_827,In_1219,In_1081);
or U828 (N_828,In_1197,In_965);
and U829 (N_829,In_93,In_768);
nor U830 (N_830,In_1247,In_673);
nor U831 (N_831,In_266,In_144);
nor U832 (N_832,In_727,In_1156);
and U833 (N_833,In_1156,In_183);
or U834 (N_834,In_342,In_1);
and U835 (N_835,In_1122,In_493);
nand U836 (N_836,In_433,In_1464);
nor U837 (N_837,In_1393,In_1240);
and U838 (N_838,In_487,In_47);
or U839 (N_839,In_1396,In_493);
and U840 (N_840,In_430,In_11);
nor U841 (N_841,In_625,In_1002);
nand U842 (N_842,In_642,In_1467);
nand U843 (N_843,In_660,In_357);
nor U844 (N_844,In_456,In_13);
and U845 (N_845,In_622,In_697);
nand U846 (N_846,In_1463,In_618);
nand U847 (N_847,In_678,In_407);
and U848 (N_848,In_430,In_1089);
and U849 (N_849,In_851,In_140);
nor U850 (N_850,In_478,In_552);
and U851 (N_851,In_1302,In_815);
xor U852 (N_852,In_929,In_521);
xor U853 (N_853,In_226,In_1184);
or U854 (N_854,In_1332,In_880);
and U855 (N_855,In_713,In_646);
nor U856 (N_856,In_1168,In_422);
nand U857 (N_857,In_1211,In_1090);
nor U858 (N_858,In_1157,In_604);
nor U859 (N_859,In_1490,In_359);
nor U860 (N_860,In_578,In_956);
or U861 (N_861,In_879,In_844);
nand U862 (N_862,In_724,In_387);
or U863 (N_863,In_554,In_525);
xnor U864 (N_864,In_1232,In_31);
and U865 (N_865,In_461,In_497);
nor U866 (N_866,In_759,In_1074);
nor U867 (N_867,In_182,In_245);
or U868 (N_868,In_931,In_1184);
nand U869 (N_869,In_873,In_368);
or U870 (N_870,In_95,In_1102);
nand U871 (N_871,In_1455,In_666);
nor U872 (N_872,In_1341,In_544);
xor U873 (N_873,In_548,In_964);
or U874 (N_874,In_995,In_397);
nor U875 (N_875,In_585,In_343);
and U876 (N_876,In_1328,In_46);
xor U877 (N_877,In_1121,In_690);
nand U878 (N_878,In_1033,In_1155);
or U879 (N_879,In_182,In_306);
or U880 (N_880,In_133,In_833);
nand U881 (N_881,In_453,In_1354);
xor U882 (N_882,In_250,In_1129);
nand U883 (N_883,In_701,In_964);
nor U884 (N_884,In_1010,In_20);
or U885 (N_885,In_343,In_1241);
or U886 (N_886,In_61,In_673);
xor U887 (N_887,In_663,In_1137);
or U888 (N_888,In_918,In_29);
nor U889 (N_889,In_1300,In_853);
and U890 (N_890,In_596,In_981);
or U891 (N_891,In_845,In_1029);
nor U892 (N_892,In_48,In_404);
or U893 (N_893,In_1482,In_45);
and U894 (N_894,In_798,In_1416);
nand U895 (N_895,In_1191,In_589);
nand U896 (N_896,In_1260,In_1361);
or U897 (N_897,In_402,In_571);
or U898 (N_898,In_660,In_960);
or U899 (N_899,In_785,In_938);
nor U900 (N_900,In_1151,In_508);
and U901 (N_901,In_745,In_831);
or U902 (N_902,In_316,In_583);
and U903 (N_903,In_283,In_1394);
xnor U904 (N_904,In_917,In_940);
nand U905 (N_905,In_814,In_1224);
or U906 (N_906,In_163,In_686);
or U907 (N_907,In_249,In_1446);
nor U908 (N_908,In_648,In_1001);
nor U909 (N_909,In_834,In_159);
nand U910 (N_910,In_290,In_1255);
nor U911 (N_911,In_778,In_811);
and U912 (N_912,In_734,In_216);
nor U913 (N_913,In_1225,In_1041);
nand U914 (N_914,In_142,In_738);
nand U915 (N_915,In_669,In_940);
and U916 (N_916,In_296,In_1268);
nor U917 (N_917,In_790,In_963);
nand U918 (N_918,In_859,In_55);
or U919 (N_919,In_1367,In_812);
nand U920 (N_920,In_1007,In_702);
and U921 (N_921,In_442,In_328);
nor U922 (N_922,In_1440,In_117);
and U923 (N_923,In_633,In_549);
nor U924 (N_924,In_1215,In_1382);
and U925 (N_925,In_354,In_1183);
nor U926 (N_926,In_780,In_327);
or U927 (N_927,In_1269,In_135);
and U928 (N_928,In_1113,In_1062);
nor U929 (N_929,In_1364,In_1159);
nor U930 (N_930,In_912,In_219);
and U931 (N_931,In_18,In_494);
or U932 (N_932,In_77,In_1135);
and U933 (N_933,In_1015,In_1249);
nand U934 (N_934,In_1187,In_571);
and U935 (N_935,In_126,In_1290);
or U936 (N_936,In_899,In_1479);
or U937 (N_937,In_370,In_933);
and U938 (N_938,In_1214,In_603);
or U939 (N_939,In_1487,In_675);
nand U940 (N_940,In_422,In_210);
xnor U941 (N_941,In_661,In_795);
nand U942 (N_942,In_1053,In_1093);
or U943 (N_943,In_24,In_594);
or U944 (N_944,In_1346,In_1017);
or U945 (N_945,In_1176,In_579);
nor U946 (N_946,In_1391,In_350);
xnor U947 (N_947,In_1147,In_1090);
or U948 (N_948,In_266,In_706);
and U949 (N_949,In_294,In_73);
nand U950 (N_950,In_1246,In_111);
and U951 (N_951,In_1455,In_506);
or U952 (N_952,In_1349,In_308);
nor U953 (N_953,In_675,In_1043);
and U954 (N_954,In_1037,In_164);
nand U955 (N_955,In_738,In_448);
and U956 (N_956,In_932,In_466);
and U957 (N_957,In_433,In_1262);
nand U958 (N_958,In_536,In_1301);
nand U959 (N_959,In_431,In_1415);
nor U960 (N_960,In_1456,In_1275);
nor U961 (N_961,In_1115,In_190);
and U962 (N_962,In_220,In_84);
nor U963 (N_963,In_1007,In_911);
and U964 (N_964,In_1003,In_868);
nand U965 (N_965,In_413,In_1299);
and U966 (N_966,In_252,In_195);
and U967 (N_967,In_1112,In_974);
and U968 (N_968,In_790,In_1084);
or U969 (N_969,In_727,In_846);
nor U970 (N_970,In_888,In_1210);
and U971 (N_971,In_927,In_908);
xnor U972 (N_972,In_284,In_488);
and U973 (N_973,In_338,In_1095);
or U974 (N_974,In_941,In_306);
or U975 (N_975,In_769,In_936);
nand U976 (N_976,In_305,In_581);
nor U977 (N_977,In_831,In_901);
and U978 (N_978,In_352,In_829);
nor U979 (N_979,In_1370,In_341);
nor U980 (N_980,In_1329,In_138);
or U981 (N_981,In_529,In_1090);
nand U982 (N_982,In_1436,In_563);
nor U983 (N_983,In_843,In_970);
or U984 (N_984,In_380,In_856);
xnor U985 (N_985,In_173,In_917);
nor U986 (N_986,In_641,In_440);
xnor U987 (N_987,In_507,In_375);
nand U988 (N_988,In_1158,In_711);
nor U989 (N_989,In_1300,In_205);
or U990 (N_990,In_175,In_240);
nor U991 (N_991,In_856,In_1244);
xnor U992 (N_992,In_205,In_1112);
nand U993 (N_993,In_663,In_667);
nand U994 (N_994,In_11,In_189);
nand U995 (N_995,In_406,In_9);
nand U996 (N_996,In_960,In_380);
nand U997 (N_997,In_1499,In_136);
and U998 (N_998,In_11,In_1182);
and U999 (N_999,In_1282,In_518);
nor U1000 (N_1000,N_144,N_350);
or U1001 (N_1001,N_2,N_419);
and U1002 (N_1002,N_883,N_764);
and U1003 (N_1003,N_200,N_151);
or U1004 (N_1004,N_745,N_576);
and U1005 (N_1005,N_615,N_103);
or U1006 (N_1006,N_335,N_383);
or U1007 (N_1007,N_125,N_153);
nor U1008 (N_1008,N_311,N_773);
or U1009 (N_1009,N_270,N_435);
nor U1010 (N_1010,N_947,N_436);
nor U1011 (N_1011,N_616,N_645);
xnor U1012 (N_1012,N_849,N_664);
nor U1013 (N_1013,N_681,N_845);
and U1014 (N_1014,N_635,N_267);
nand U1015 (N_1015,N_77,N_646);
and U1016 (N_1016,N_826,N_708);
xnor U1017 (N_1017,N_361,N_688);
or U1018 (N_1018,N_366,N_900);
xor U1019 (N_1019,N_266,N_997);
nand U1020 (N_1020,N_956,N_416);
xor U1021 (N_1021,N_902,N_400);
nand U1022 (N_1022,N_299,N_985);
xnor U1023 (N_1023,N_491,N_272);
or U1024 (N_1024,N_740,N_560);
and U1025 (N_1025,N_188,N_458);
or U1026 (N_1026,N_921,N_980);
nor U1027 (N_1027,N_60,N_940);
and U1028 (N_1028,N_717,N_57);
xor U1029 (N_1029,N_225,N_808);
nand U1030 (N_1030,N_755,N_661);
or U1031 (N_1031,N_329,N_164);
nand U1032 (N_1032,N_523,N_608);
nand U1033 (N_1033,N_514,N_539);
or U1034 (N_1034,N_493,N_170);
nand U1035 (N_1035,N_48,N_589);
and U1036 (N_1036,N_71,N_369);
nor U1037 (N_1037,N_246,N_104);
nand U1038 (N_1038,N_18,N_332);
and U1039 (N_1039,N_224,N_27);
or U1040 (N_1040,N_247,N_127);
xnor U1041 (N_1041,N_248,N_898);
nor U1042 (N_1042,N_882,N_472);
nand U1043 (N_1043,N_524,N_265);
and U1044 (N_1044,N_169,N_111);
nand U1045 (N_1045,N_67,N_769);
nor U1046 (N_1046,N_916,N_237);
or U1047 (N_1047,N_308,N_199);
and U1048 (N_1048,N_438,N_802);
and U1049 (N_1049,N_494,N_544);
nand U1050 (N_1050,N_675,N_205);
and U1051 (N_1051,N_919,N_279);
nand U1052 (N_1052,N_610,N_991);
or U1053 (N_1053,N_149,N_886);
or U1054 (N_1054,N_952,N_218);
nand U1055 (N_1055,N_621,N_622);
nor U1056 (N_1056,N_0,N_154);
nand U1057 (N_1057,N_552,N_896);
nor U1058 (N_1058,N_639,N_146);
or U1059 (N_1059,N_23,N_823);
and U1060 (N_1060,N_770,N_547);
or U1061 (N_1061,N_291,N_709);
and U1062 (N_1062,N_47,N_126);
nand U1063 (N_1063,N_602,N_938);
nor U1064 (N_1064,N_935,N_25);
or U1065 (N_1065,N_724,N_322);
nand U1066 (N_1066,N_190,N_293);
nor U1067 (N_1067,N_964,N_692);
or U1068 (N_1068,N_393,N_100);
nor U1069 (N_1069,N_577,N_506);
nor U1070 (N_1070,N_413,N_428);
nand U1071 (N_1071,N_390,N_12);
or U1072 (N_1072,N_797,N_668);
or U1073 (N_1073,N_926,N_452);
nor U1074 (N_1074,N_92,N_160);
or U1075 (N_1075,N_580,N_286);
or U1076 (N_1076,N_582,N_88);
nand U1077 (N_1077,N_949,N_695);
or U1078 (N_1078,N_349,N_798);
nor U1079 (N_1079,N_939,N_777);
nand U1080 (N_1080,N_139,N_716);
nor U1081 (N_1081,N_933,N_564);
and U1082 (N_1082,N_888,N_482);
nand U1083 (N_1083,N_175,N_113);
nor U1084 (N_1084,N_663,N_288);
nand U1085 (N_1085,N_780,N_852);
nand U1086 (N_1086,N_213,N_52);
nor U1087 (N_1087,N_98,N_843);
or U1088 (N_1088,N_387,N_904);
nand U1089 (N_1089,N_410,N_33);
or U1090 (N_1090,N_243,N_121);
nor U1091 (N_1091,N_346,N_987);
and U1092 (N_1092,N_459,N_466);
nor U1093 (N_1093,N_557,N_891);
nor U1094 (N_1094,N_925,N_330);
or U1095 (N_1095,N_747,N_893);
and U1096 (N_1096,N_261,N_269);
and U1097 (N_1097,N_219,N_347);
nand U1098 (N_1098,N_217,N_39);
and U1099 (N_1099,N_207,N_359);
nor U1100 (N_1100,N_22,N_763);
nand U1101 (N_1101,N_385,N_696);
nor U1102 (N_1102,N_173,N_42);
nand U1103 (N_1103,N_930,N_29);
or U1104 (N_1104,N_344,N_44);
or U1105 (N_1105,N_63,N_495);
nor U1106 (N_1106,N_572,N_80);
and U1107 (N_1107,N_944,N_827);
and U1108 (N_1108,N_28,N_325);
and U1109 (N_1109,N_599,N_147);
or U1110 (N_1110,N_855,N_978);
nor U1111 (N_1111,N_233,N_297);
nand U1112 (N_1112,N_611,N_937);
nor U1113 (N_1113,N_508,N_640);
nand U1114 (N_1114,N_525,N_690);
or U1115 (N_1115,N_365,N_856);
or U1116 (N_1116,N_409,N_873);
and U1117 (N_1117,N_473,N_184);
or U1118 (N_1118,N_249,N_848);
or U1119 (N_1119,N_503,N_627);
xor U1120 (N_1120,N_737,N_965);
or U1121 (N_1121,N_376,N_15);
nor U1122 (N_1122,N_487,N_162);
or U1123 (N_1123,N_596,N_180);
nand U1124 (N_1124,N_791,N_296);
or U1125 (N_1125,N_734,N_700);
or U1126 (N_1126,N_110,N_631);
or U1127 (N_1127,N_415,N_538);
nor U1128 (N_1128,N_370,N_658);
nand U1129 (N_1129,N_21,N_394);
xor U1130 (N_1130,N_927,N_634);
nor U1131 (N_1131,N_836,N_283);
and U1132 (N_1132,N_194,N_697);
nor U1133 (N_1133,N_74,N_398);
nand U1134 (N_1134,N_941,N_439);
or U1135 (N_1135,N_784,N_26);
nor U1136 (N_1136,N_278,N_263);
nand U1137 (N_1137,N_301,N_327);
nor U1138 (N_1138,N_356,N_253);
nand U1139 (N_1139,N_474,N_399);
nor U1140 (N_1140,N_943,N_559);
nand U1141 (N_1141,N_381,N_603);
nand U1142 (N_1142,N_594,N_567);
or U1143 (N_1143,N_316,N_442);
xnor U1144 (N_1144,N_542,N_885);
nor U1145 (N_1145,N_620,N_352);
xor U1146 (N_1146,N_223,N_793);
nand U1147 (N_1147,N_584,N_711);
nor U1148 (N_1148,N_533,N_446);
or U1149 (N_1149,N_806,N_264);
xnor U1150 (N_1150,N_55,N_448);
or U1151 (N_1151,N_723,N_707);
or U1152 (N_1152,N_537,N_295);
nand U1153 (N_1153,N_928,N_226);
nor U1154 (N_1154,N_159,N_816);
nand U1155 (N_1155,N_231,N_426);
nand U1156 (N_1156,N_768,N_13);
nor U1157 (N_1157,N_858,N_644);
xnor U1158 (N_1158,N_331,N_4);
or U1159 (N_1159,N_983,N_592);
nand U1160 (N_1160,N_321,N_846);
nand U1161 (N_1161,N_251,N_315);
and U1162 (N_1162,N_586,N_570);
nor U1163 (N_1163,N_285,N_871);
or U1164 (N_1164,N_429,N_682);
nand U1165 (N_1165,N_629,N_698);
nor U1166 (N_1166,N_833,N_216);
nand U1167 (N_1167,N_483,N_14);
or U1168 (N_1168,N_142,N_591);
nor U1169 (N_1169,N_766,N_617);
nand U1170 (N_1170,N_877,N_931);
nand U1171 (N_1171,N_179,N_371);
nor U1172 (N_1172,N_450,N_756);
or U1173 (N_1173,N_500,N_804);
nor U1174 (N_1174,N_715,N_579);
and U1175 (N_1175,N_585,N_929);
or U1176 (N_1176,N_529,N_782);
and U1177 (N_1177,N_678,N_84);
and U1178 (N_1178,N_862,N_718);
or U1179 (N_1179,N_509,N_484);
nor U1180 (N_1180,N_202,N_890);
and U1181 (N_1181,N_517,N_624);
and U1182 (N_1182,N_951,N_519);
and U1183 (N_1183,N_545,N_722);
and U1184 (N_1184,N_684,N_172);
or U1185 (N_1185,N_659,N_320);
and U1186 (N_1186,N_914,N_401);
nor U1187 (N_1187,N_772,N_676);
or U1188 (N_1188,N_865,N_56);
nor U1189 (N_1189,N_779,N_606);
xnor U1190 (N_1190,N_1,N_367);
nor U1191 (N_1191,N_837,N_386);
or U1192 (N_1192,N_748,N_957);
or U1193 (N_1193,N_260,N_66);
nand U1194 (N_1194,N_274,N_986);
nor U1195 (N_1195,N_730,N_553);
nand U1196 (N_1196,N_960,N_62);
xnor U1197 (N_1197,N_106,N_362);
or U1198 (N_1198,N_569,N_895);
nand U1199 (N_1199,N_568,N_280);
xnor U1200 (N_1200,N_481,N_775);
or U1201 (N_1201,N_203,N_314);
nor U1202 (N_1202,N_795,N_447);
or U1203 (N_1203,N_727,N_600);
nand U1204 (N_1204,N_7,N_339);
and U1205 (N_1205,N_750,N_345);
nor U1206 (N_1206,N_854,N_465);
or U1207 (N_1207,N_936,N_543);
nand U1208 (N_1208,N_424,N_887);
xnor U1209 (N_1209,N_832,N_8);
nand U1210 (N_1210,N_408,N_762);
nand U1211 (N_1211,N_397,N_469);
and U1212 (N_1212,N_417,N_189);
and U1213 (N_1213,N_742,N_463);
or U1214 (N_1214,N_423,N_945);
xor U1215 (N_1215,N_999,N_876);
or U1216 (N_1216,N_701,N_598);
nand U1217 (N_1217,N_702,N_488);
nor U1218 (N_1218,N_825,N_215);
and U1219 (N_1219,N_421,N_889);
nand U1220 (N_1220,N_872,N_312);
or U1221 (N_1221,N_300,N_504);
nand U1222 (N_1222,N_130,N_443);
nor U1223 (N_1223,N_357,N_648);
and U1224 (N_1224,N_3,N_794);
and U1225 (N_1225,N_323,N_735);
nor U1226 (N_1226,N_49,N_68);
xnor U1227 (N_1227,N_562,N_554);
and U1228 (N_1228,N_120,N_510);
nor U1229 (N_1229,N_108,N_556);
and U1230 (N_1230,N_196,N_94);
and U1231 (N_1231,N_35,N_241);
or U1232 (N_1232,N_19,N_526);
nor U1233 (N_1233,N_105,N_181);
nor U1234 (N_1234,N_183,N_185);
nand U1235 (N_1235,N_112,N_412);
nor U1236 (N_1236,N_751,N_384);
and U1237 (N_1237,N_875,N_354);
or U1238 (N_1238,N_96,N_788);
nand U1239 (N_1239,N_140,N_642);
nor U1240 (N_1240,N_210,N_815);
nand U1241 (N_1241,N_101,N_461);
and U1242 (N_1242,N_674,N_990);
and U1243 (N_1243,N_122,N_456);
nor U1244 (N_1244,N_683,N_275);
and U1245 (N_1245,N_981,N_842);
xor U1246 (N_1246,N_761,N_10);
and U1247 (N_1247,N_479,N_505);
nor U1248 (N_1248,N_649,N_50);
and U1249 (N_1249,N_238,N_908);
nor U1250 (N_1250,N_619,N_168);
xor U1251 (N_1251,N_289,N_379);
nor U1252 (N_1252,N_731,N_395);
and U1253 (N_1253,N_433,N_427);
or U1254 (N_1254,N_662,N_116);
or U1255 (N_1255,N_31,N_341);
or U1256 (N_1256,N_628,N_430);
or U1257 (N_1257,N_9,N_637);
nand U1258 (N_1258,N_85,N_382);
and U1259 (N_1259,N_489,N_565);
nor U1260 (N_1260,N_966,N_258);
nand U1261 (N_1261,N_901,N_502);
and U1262 (N_1262,N_971,N_499);
nand U1263 (N_1263,N_209,N_135);
nor U1264 (N_1264,N_656,N_753);
and U1265 (N_1265,N_899,N_24);
or U1266 (N_1266,N_37,N_820);
and U1267 (N_1267,N_738,N_497);
and U1268 (N_1268,N_437,N_630);
or U1269 (N_1269,N_853,N_32);
nor U1270 (N_1270,N_968,N_680);
and U1271 (N_1271,N_982,N_364);
and U1272 (N_1272,N_287,N_208);
xnor U1273 (N_1273,N_198,N_6);
nand U1274 (N_1274,N_652,N_530);
nor U1275 (N_1275,N_571,N_819);
or U1276 (N_1276,N_691,N_911);
and U1277 (N_1277,N_641,N_158);
and U1278 (N_1278,N_176,N_273);
or U1279 (N_1279,N_245,N_374);
or U1280 (N_1280,N_211,N_30);
nand U1281 (N_1281,N_633,N_989);
nand U1282 (N_1282,N_913,N_403);
nand U1283 (N_1283,N_392,N_182);
nand U1284 (N_1284,N_262,N_654);
nand U1285 (N_1285,N_59,N_752);
xor U1286 (N_1286,N_623,N_699);
xnor U1287 (N_1287,N_667,N_89);
nand U1288 (N_1288,N_857,N_522);
nand U1289 (N_1289,N_282,N_64);
nand U1290 (N_1290,N_632,N_636);
or U1291 (N_1291,N_792,N_133);
or U1292 (N_1292,N_771,N_741);
nand U1293 (N_1293,N_292,N_490);
nor U1294 (N_1294,N_705,N_992);
nor U1295 (N_1295,N_760,N_977);
and U1296 (N_1296,N_587,N_774);
nor U1297 (N_1297,N_425,N_869);
or U1298 (N_1298,N_498,N_134);
and U1299 (N_1299,N_230,N_192);
nor U1300 (N_1300,N_254,N_831);
nor U1301 (N_1301,N_870,N_710);
nand U1302 (N_1302,N_732,N_174);
nand U1303 (N_1303,N_726,N_787);
nand U1304 (N_1304,N_259,N_157);
or U1305 (N_1305,N_746,N_454);
nand U1306 (N_1306,N_475,N_478);
or U1307 (N_1307,N_575,N_881);
xnor U1308 (N_1308,N_643,N_924);
nand U1309 (N_1309,N_758,N_536);
xor U1310 (N_1310,N_95,N_467);
nor U1311 (N_1311,N_725,N_665);
and U1312 (N_1312,N_204,N_138);
nand U1313 (N_1313,N_907,N_706);
and U1314 (N_1314,N_444,N_534);
nand U1315 (N_1315,N_810,N_595);
nor U1316 (N_1316,N_17,N_767);
nor U1317 (N_1317,N_970,N_141);
nand U1318 (N_1318,N_340,N_834);
or U1319 (N_1319,N_821,N_470);
nor U1320 (N_1320,N_516,N_822);
nor U1321 (N_1321,N_389,N_445);
or U1322 (N_1322,N_551,N_460);
nand U1323 (N_1323,N_161,N_82);
or U1324 (N_1324,N_918,N_720);
nor U1325 (N_1325,N_388,N_178);
nand U1326 (N_1326,N_829,N_593);
nand U1327 (N_1327,N_306,N_609);
nor U1328 (N_1328,N_626,N_65);
or U1329 (N_1329,N_714,N_897);
nor U1330 (N_1330,N_377,N_136);
nand U1331 (N_1331,N_109,N_670);
and U1332 (N_1332,N_486,N_840);
nor U1333 (N_1333,N_781,N_229);
or U1334 (N_1334,N_812,N_800);
xor U1335 (N_1335,N_239,N_830);
or U1336 (N_1336,N_948,N_449);
and U1337 (N_1337,N_880,N_235);
nand U1338 (N_1338,N_492,N_36);
and U1339 (N_1339,N_647,N_342);
nand U1340 (N_1340,N_480,N_431);
and U1341 (N_1341,N_757,N_613);
or U1342 (N_1342,N_256,N_729);
or U1343 (N_1343,N_550,N_932);
nor U1344 (N_1344,N_90,N_693);
and U1345 (N_1345,N_276,N_268);
nand U1346 (N_1346,N_97,N_236);
and U1347 (N_1347,N_197,N_114);
and U1348 (N_1348,N_411,N_220);
or U1349 (N_1349,N_541,N_549);
and U1350 (N_1350,N_372,N_5);
or U1351 (N_1351,N_420,N_257);
and U1352 (N_1352,N_561,N_581);
or U1353 (N_1353,N_343,N_511);
nor U1354 (N_1354,N_650,N_863);
or U1355 (N_1355,N_453,N_719);
nand U1356 (N_1356,N_671,N_573);
or U1357 (N_1357,N_778,N_324);
and U1358 (N_1358,N_625,N_689);
or U1359 (N_1359,N_471,N_242);
xnor U1360 (N_1360,N_58,N_51);
or U1361 (N_1361,N_563,N_809);
nor U1362 (N_1362,N_79,N_102);
nor U1363 (N_1363,N_993,N_785);
or U1364 (N_1364,N_574,N_326);
and U1365 (N_1365,N_588,N_405);
and U1366 (N_1366,N_685,N_638);
nand U1367 (N_1367,N_920,N_790);
xnor U1368 (N_1368,N_171,N_614);
nor U1369 (N_1369,N_462,N_422);
or U1370 (N_1370,N_337,N_165);
nand U1371 (N_1371,N_546,N_686);
nand U1372 (N_1372,N_123,N_866);
and U1373 (N_1373,N_950,N_860);
nor U1374 (N_1374,N_660,N_783);
nor U1375 (N_1375,N_368,N_255);
nor U1376 (N_1376,N_507,N_281);
or U1377 (N_1377,N_532,N_76);
and U1378 (N_1378,N_477,N_418);
nand U1379 (N_1379,N_905,N_378);
nor U1380 (N_1380,N_129,N_191);
and U1381 (N_1381,N_975,N_380);
or U1382 (N_1382,N_132,N_73);
nand U1383 (N_1383,N_406,N_455);
or U1384 (N_1384,N_277,N_290);
nand U1385 (N_1385,N_441,N_404);
and U1386 (N_1386,N_396,N_16);
or U1387 (N_1387,N_527,N_850);
and U1388 (N_1388,N_704,N_669);
nor U1389 (N_1389,N_319,N_228);
or U1390 (N_1390,N_958,N_535);
xor U1391 (N_1391,N_923,N_468);
or U1392 (N_1392,N_451,N_961);
nor U1393 (N_1393,N_861,N_375);
and U1394 (N_1394,N_45,N_578);
nor U1395 (N_1395,N_518,N_607);
nor U1396 (N_1396,N_967,N_694);
nand U1397 (N_1397,N_119,N_867);
or U1398 (N_1398,N_252,N_83);
nand U1399 (N_1399,N_736,N_879);
and U1400 (N_1400,N_744,N_884);
nand U1401 (N_1401,N_868,N_234);
and U1402 (N_1402,N_942,N_328);
and U1403 (N_1403,N_152,N_712);
and U1404 (N_1404,N_107,N_995);
or U1405 (N_1405,N_847,N_811);
and U1406 (N_1406,N_310,N_214);
nor U1407 (N_1407,N_984,N_733);
and U1408 (N_1408,N_612,N_894);
and U1409 (N_1409,N_655,N_835);
nor U1410 (N_1410,N_313,N_759);
or U1411 (N_1411,N_43,N_959);
or U1412 (N_1412,N_34,N_167);
nand U1413 (N_1413,N_605,N_555);
xnor U1414 (N_1414,N_687,N_903);
or U1415 (N_1415,N_776,N_355);
and U1416 (N_1416,N_221,N_851);
nor U1417 (N_1417,N_115,N_976);
nand U1418 (N_1418,N_227,N_20);
nor U1419 (N_1419,N_72,N_360);
and U1420 (N_1420,N_131,N_250);
nor U1421 (N_1421,N_601,N_206);
or U1422 (N_1422,N_953,N_358);
or U1423 (N_1423,N_40,N_212);
and U1424 (N_1424,N_294,N_128);
or U1425 (N_1425,N_521,N_240);
and U1426 (N_1426,N_803,N_307);
xnor U1427 (N_1427,N_163,N_839);
nor U1428 (N_1428,N_402,N_651);
nor U1429 (N_1429,N_590,N_118);
and U1430 (N_1430,N_910,N_222);
nand U1431 (N_1431,N_351,N_679);
nand U1432 (N_1432,N_11,N_998);
xnor U1433 (N_1433,N_177,N_117);
nand U1434 (N_1434,N_457,N_972);
nor U1435 (N_1435,N_677,N_187);
nor U1436 (N_1436,N_807,N_548);
nand U1437 (N_1437,N_922,N_721);
xor U1438 (N_1438,N_786,N_70);
and U1439 (N_1439,N_193,N_909);
nand U1440 (N_1440,N_874,N_244);
and U1441 (N_1441,N_155,N_520);
or U1442 (N_1442,N_618,N_912);
xor U1443 (N_1443,N_137,N_955);
nor U1444 (N_1444,N_512,N_302);
nor U1445 (N_1445,N_391,N_333);
nand U1446 (N_1446,N_353,N_996);
or U1447 (N_1447,N_962,N_906);
nand U1448 (N_1448,N_61,N_994);
and U1449 (N_1449,N_817,N_841);
and U1450 (N_1450,N_813,N_99);
and U1451 (N_1451,N_653,N_878);
nand U1452 (N_1452,N_304,N_41);
or U1453 (N_1453,N_407,N_38);
xor U1454 (N_1454,N_46,N_974);
and U1455 (N_1455,N_69,N_828);
nor U1456 (N_1456,N_796,N_566);
nor U1457 (N_1457,N_988,N_583);
and U1458 (N_1458,N_143,N_373);
xnor U1459 (N_1459,N_528,N_814);
nand U1460 (N_1460,N_973,N_78);
and U1461 (N_1461,N_789,N_476);
nand U1462 (N_1462,N_91,N_336);
nand U1463 (N_1463,N_513,N_334);
or U1464 (N_1464,N_186,N_824);
and U1465 (N_1465,N_284,N_309);
nor U1466 (N_1466,N_338,N_838);
nor U1467 (N_1467,N_271,N_892);
nor U1468 (N_1468,N_979,N_749);
and U1469 (N_1469,N_298,N_801);
nand U1470 (N_1470,N_844,N_963);
and U1471 (N_1471,N_501,N_597);
nand U1472 (N_1472,N_124,N_156);
xnor U1473 (N_1473,N_434,N_54);
or U1474 (N_1474,N_917,N_317);
nand U1475 (N_1475,N_305,N_496);
and U1476 (N_1476,N_805,N_145);
nor U1477 (N_1477,N_432,N_864);
nor U1478 (N_1478,N_53,N_166);
nor U1479 (N_1479,N_303,N_87);
nor U1480 (N_1480,N_954,N_739);
xor U1481 (N_1481,N_348,N_934);
and U1482 (N_1482,N_440,N_485);
xnor U1483 (N_1483,N_195,N_743);
nand U1484 (N_1484,N_363,N_232);
nor U1485 (N_1485,N_540,N_765);
nor U1486 (N_1486,N_754,N_318);
nor U1487 (N_1487,N_81,N_86);
and U1488 (N_1488,N_703,N_558);
nor U1489 (N_1489,N_666,N_464);
nand U1490 (N_1490,N_946,N_515);
and U1491 (N_1491,N_859,N_969);
or U1492 (N_1492,N_657,N_414);
xnor U1493 (N_1493,N_531,N_604);
nand U1494 (N_1494,N_673,N_150);
xor U1495 (N_1495,N_75,N_148);
or U1496 (N_1496,N_93,N_799);
and U1497 (N_1497,N_728,N_201);
nand U1498 (N_1498,N_713,N_915);
nand U1499 (N_1499,N_672,N_818);
nand U1500 (N_1500,N_846,N_978);
nand U1501 (N_1501,N_492,N_977);
and U1502 (N_1502,N_372,N_682);
xnor U1503 (N_1503,N_336,N_656);
or U1504 (N_1504,N_813,N_647);
nand U1505 (N_1505,N_259,N_575);
nor U1506 (N_1506,N_329,N_459);
nor U1507 (N_1507,N_33,N_283);
nor U1508 (N_1508,N_15,N_487);
or U1509 (N_1509,N_589,N_455);
and U1510 (N_1510,N_52,N_419);
or U1511 (N_1511,N_53,N_507);
xnor U1512 (N_1512,N_961,N_487);
and U1513 (N_1513,N_676,N_17);
and U1514 (N_1514,N_717,N_653);
or U1515 (N_1515,N_172,N_933);
nand U1516 (N_1516,N_567,N_90);
and U1517 (N_1517,N_458,N_770);
nor U1518 (N_1518,N_831,N_708);
and U1519 (N_1519,N_391,N_371);
and U1520 (N_1520,N_56,N_201);
nor U1521 (N_1521,N_915,N_145);
nand U1522 (N_1522,N_762,N_588);
and U1523 (N_1523,N_137,N_414);
and U1524 (N_1524,N_236,N_73);
and U1525 (N_1525,N_855,N_834);
or U1526 (N_1526,N_369,N_434);
nand U1527 (N_1527,N_68,N_445);
or U1528 (N_1528,N_342,N_270);
and U1529 (N_1529,N_939,N_334);
or U1530 (N_1530,N_834,N_604);
nor U1531 (N_1531,N_210,N_206);
and U1532 (N_1532,N_336,N_270);
or U1533 (N_1533,N_62,N_715);
nor U1534 (N_1534,N_385,N_255);
nand U1535 (N_1535,N_474,N_918);
nor U1536 (N_1536,N_788,N_73);
nor U1537 (N_1537,N_421,N_290);
nor U1538 (N_1538,N_368,N_685);
nor U1539 (N_1539,N_663,N_865);
or U1540 (N_1540,N_489,N_394);
nor U1541 (N_1541,N_730,N_628);
nand U1542 (N_1542,N_436,N_860);
xnor U1543 (N_1543,N_636,N_354);
nand U1544 (N_1544,N_57,N_966);
nor U1545 (N_1545,N_929,N_327);
xnor U1546 (N_1546,N_832,N_596);
and U1547 (N_1547,N_185,N_490);
nand U1548 (N_1548,N_847,N_464);
and U1549 (N_1549,N_642,N_598);
nor U1550 (N_1550,N_75,N_322);
nand U1551 (N_1551,N_759,N_859);
nor U1552 (N_1552,N_571,N_850);
nand U1553 (N_1553,N_485,N_293);
nand U1554 (N_1554,N_692,N_157);
xnor U1555 (N_1555,N_92,N_63);
and U1556 (N_1556,N_180,N_830);
nand U1557 (N_1557,N_438,N_230);
and U1558 (N_1558,N_547,N_739);
or U1559 (N_1559,N_435,N_859);
or U1560 (N_1560,N_56,N_580);
nor U1561 (N_1561,N_555,N_720);
nor U1562 (N_1562,N_121,N_999);
nor U1563 (N_1563,N_417,N_963);
and U1564 (N_1564,N_214,N_313);
and U1565 (N_1565,N_15,N_665);
nand U1566 (N_1566,N_544,N_790);
or U1567 (N_1567,N_565,N_666);
xnor U1568 (N_1568,N_145,N_742);
and U1569 (N_1569,N_369,N_42);
xor U1570 (N_1570,N_613,N_780);
or U1571 (N_1571,N_243,N_582);
and U1572 (N_1572,N_154,N_271);
nand U1573 (N_1573,N_662,N_418);
or U1574 (N_1574,N_142,N_739);
or U1575 (N_1575,N_364,N_838);
nand U1576 (N_1576,N_302,N_215);
and U1577 (N_1577,N_941,N_972);
nand U1578 (N_1578,N_106,N_395);
nand U1579 (N_1579,N_222,N_602);
and U1580 (N_1580,N_458,N_648);
nor U1581 (N_1581,N_239,N_226);
and U1582 (N_1582,N_265,N_49);
nand U1583 (N_1583,N_351,N_556);
nand U1584 (N_1584,N_711,N_836);
nor U1585 (N_1585,N_275,N_444);
and U1586 (N_1586,N_105,N_923);
xor U1587 (N_1587,N_86,N_766);
nor U1588 (N_1588,N_296,N_448);
nor U1589 (N_1589,N_656,N_202);
xor U1590 (N_1590,N_163,N_462);
or U1591 (N_1591,N_363,N_872);
or U1592 (N_1592,N_566,N_489);
nor U1593 (N_1593,N_731,N_773);
or U1594 (N_1594,N_900,N_901);
and U1595 (N_1595,N_227,N_799);
nand U1596 (N_1596,N_504,N_223);
and U1597 (N_1597,N_521,N_148);
nor U1598 (N_1598,N_184,N_470);
and U1599 (N_1599,N_793,N_7);
nand U1600 (N_1600,N_975,N_659);
and U1601 (N_1601,N_586,N_134);
or U1602 (N_1602,N_67,N_81);
nand U1603 (N_1603,N_712,N_956);
nor U1604 (N_1604,N_321,N_9);
nand U1605 (N_1605,N_351,N_669);
and U1606 (N_1606,N_934,N_962);
xnor U1607 (N_1607,N_623,N_299);
and U1608 (N_1608,N_267,N_694);
nor U1609 (N_1609,N_263,N_481);
nand U1610 (N_1610,N_937,N_265);
nand U1611 (N_1611,N_328,N_59);
nor U1612 (N_1612,N_236,N_171);
nor U1613 (N_1613,N_542,N_895);
nor U1614 (N_1614,N_259,N_499);
xor U1615 (N_1615,N_848,N_449);
or U1616 (N_1616,N_259,N_38);
nand U1617 (N_1617,N_780,N_860);
or U1618 (N_1618,N_151,N_150);
xor U1619 (N_1619,N_924,N_554);
and U1620 (N_1620,N_967,N_333);
nand U1621 (N_1621,N_283,N_259);
and U1622 (N_1622,N_710,N_157);
xor U1623 (N_1623,N_406,N_886);
nor U1624 (N_1624,N_762,N_998);
or U1625 (N_1625,N_425,N_896);
nand U1626 (N_1626,N_159,N_510);
and U1627 (N_1627,N_743,N_394);
and U1628 (N_1628,N_905,N_84);
xor U1629 (N_1629,N_47,N_40);
nand U1630 (N_1630,N_557,N_654);
nor U1631 (N_1631,N_207,N_550);
and U1632 (N_1632,N_334,N_3);
nor U1633 (N_1633,N_528,N_33);
nor U1634 (N_1634,N_857,N_187);
and U1635 (N_1635,N_976,N_303);
or U1636 (N_1636,N_326,N_957);
and U1637 (N_1637,N_770,N_86);
nor U1638 (N_1638,N_907,N_820);
or U1639 (N_1639,N_939,N_672);
or U1640 (N_1640,N_39,N_545);
nand U1641 (N_1641,N_223,N_785);
xor U1642 (N_1642,N_595,N_946);
nand U1643 (N_1643,N_812,N_260);
and U1644 (N_1644,N_788,N_610);
and U1645 (N_1645,N_201,N_738);
nand U1646 (N_1646,N_658,N_737);
and U1647 (N_1647,N_880,N_73);
xnor U1648 (N_1648,N_814,N_729);
nand U1649 (N_1649,N_583,N_130);
nor U1650 (N_1650,N_171,N_380);
and U1651 (N_1651,N_797,N_732);
nor U1652 (N_1652,N_707,N_210);
nand U1653 (N_1653,N_454,N_511);
nor U1654 (N_1654,N_558,N_800);
nand U1655 (N_1655,N_3,N_883);
nand U1656 (N_1656,N_815,N_732);
and U1657 (N_1657,N_224,N_49);
xnor U1658 (N_1658,N_511,N_99);
and U1659 (N_1659,N_964,N_992);
nor U1660 (N_1660,N_73,N_847);
nand U1661 (N_1661,N_651,N_252);
or U1662 (N_1662,N_955,N_529);
or U1663 (N_1663,N_969,N_3);
nor U1664 (N_1664,N_61,N_78);
or U1665 (N_1665,N_353,N_558);
xor U1666 (N_1666,N_778,N_895);
xor U1667 (N_1667,N_734,N_395);
nor U1668 (N_1668,N_109,N_0);
or U1669 (N_1669,N_777,N_908);
and U1670 (N_1670,N_110,N_607);
nor U1671 (N_1671,N_193,N_4);
nor U1672 (N_1672,N_188,N_470);
and U1673 (N_1673,N_375,N_754);
nand U1674 (N_1674,N_204,N_200);
nor U1675 (N_1675,N_633,N_365);
xnor U1676 (N_1676,N_960,N_473);
nand U1677 (N_1677,N_368,N_950);
or U1678 (N_1678,N_367,N_492);
nor U1679 (N_1679,N_435,N_474);
or U1680 (N_1680,N_509,N_536);
nand U1681 (N_1681,N_443,N_773);
or U1682 (N_1682,N_38,N_715);
nor U1683 (N_1683,N_105,N_387);
or U1684 (N_1684,N_558,N_253);
and U1685 (N_1685,N_816,N_207);
nand U1686 (N_1686,N_812,N_445);
or U1687 (N_1687,N_356,N_665);
or U1688 (N_1688,N_513,N_580);
and U1689 (N_1689,N_526,N_897);
nand U1690 (N_1690,N_286,N_116);
or U1691 (N_1691,N_915,N_656);
or U1692 (N_1692,N_671,N_699);
nor U1693 (N_1693,N_679,N_893);
and U1694 (N_1694,N_250,N_900);
nor U1695 (N_1695,N_606,N_741);
and U1696 (N_1696,N_335,N_236);
and U1697 (N_1697,N_750,N_913);
and U1698 (N_1698,N_667,N_59);
nand U1699 (N_1699,N_891,N_252);
nor U1700 (N_1700,N_778,N_1);
xor U1701 (N_1701,N_386,N_746);
nand U1702 (N_1702,N_24,N_768);
or U1703 (N_1703,N_522,N_753);
or U1704 (N_1704,N_217,N_49);
nor U1705 (N_1705,N_815,N_152);
nor U1706 (N_1706,N_515,N_233);
and U1707 (N_1707,N_31,N_600);
or U1708 (N_1708,N_313,N_256);
and U1709 (N_1709,N_956,N_14);
or U1710 (N_1710,N_576,N_66);
or U1711 (N_1711,N_189,N_59);
or U1712 (N_1712,N_915,N_737);
or U1713 (N_1713,N_324,N_772);
nor U1714 (N_1714,N_806,N_112);
or U1715 (N_1715,N_489,N_923);
or U1716 (N_1716,N_961,N_529);
or U1717 (N_1717,N_270,N_810);
nand U1718 (N_1718,N_276,N_396);
and U1719 (N_1719,N_25,N_22);
or U1720 (N_1720,N_646,N_662);
and U1721 (N_1721,N_329,N_70);
nor U1722 (N_1722,N_493,N_271);
and U1723 (N_1723,N_738,N_118);
and U1724 (N_1724,N_798,N_358);
xor U1725 (N_1725,N_343,N_356);
nand U1726 (N_1726,N_290,N_539);
and U1727 (N_1727,N_209,N_466);
and U1728 (N_1728,N_816,N_477);
nand U1729 (N_1729,N_174,N_87);
or U1730 (N_1730,N_427,N_566);
or U1731 (N_1731,N_765,N_90);
or U1732 (N_1732,N_834,N_935);
and U1733 (N_1733,N_180,N_508);
nor U1734 (N_1734,N_571,N_977);
xnor U1735 (N_1735,N_442,N_255);
and U1736 (N_1736,N_581,N_329);
or U1737 (N_1737,N_945,N_86);
nand U1738 (N_1738,N_693,N_716);
and U1739 (N_1739,N_280,N_503);
nor U1740 (N_1740,N_23,N_217);
or U1741 (N_1741,N_865,N_19);
nand U1742 (N_1742,N_327,N_322);
and U1743 (N_1743,N_486,N_411);
nand U1744 (N_1744,N_398,N_811);
nor U1745 (N_1745,N_614,N_359);
and U1746 (N_1746,N_50,N_979);
nor U1747 (N_1747,N_805,N_285);
nor U1748 (N_1748,N_340,N_596);
nor U1749 (N_1749,N_330,N_393);
nor U1750 (N_1750,N_757,N_765);
and U1751 (N_1751,N_608,N_41);
nand U1752 (N_1752,N_900,N_834);
nand U1753 (N_1753,N_62,N_267);
nor U1754 (N_1754,N_179,N_969);
and U1755 (N_1755,N_868,N_370);
or U1756 (N_1756,N_477,N_601);
or U1757 (N_1757,N_169,N_624);
xor U1758 (N_1758,N_82,N_943);
nand U1759 (N_1759,N_495,N_325);
and U1760 (N_1760,N_191,N_566);
nand U1761 (N_1761,N_805,N_617);
xnor U1762 (N_1762,N_260,N_921);
nor U1763 (N_1763,N_71,N_182);
or U1764 (N_1764,N_170,N_380);
and U1765 (N_1765,N_721,N_397);
xor U1766 (N_1766,N_775,N_178);
or U1767 (N_1767,N_93,N_792);
nand U1768 (N_1768,N_99,N_531);
nand U1769 (N_1769,N_829,N_206);
nand U1770 (N_1770,N_377,N_18);
and U1771 (N_1771,N_917,N_377);
nor U1772 (N_1772,N_829,N_141);
nor U1773 (N_1773,N_926,N_69);
nand U1774 (N_1774,N_422,N_57);
and U1775 (N_1775,N_148,N_823);
and U1776 (N_1776,N_160,N_53);
or U1777 (N_1777,N_142,N_797);
nand U1778 (N_1778,N_197,N_856);
and U1779 (N_1779,N_936,N_588);
nor U1780 (N_1780,N_242,N_831);
or U1781 (N_1781,N_343,N_829);
or U1782 (N_1782,N_192,N_752);
and U1783 (N_1783,N_730,N_824);
nand U1784 (N_1784,N_276,N_314);
or U1785 (N_1785,N_748,N_113);
or U1786 (N_1786,N_277,N_417);
or U1787 (N_1787,N_311,N_21);
or U1788 (N_1788,N_743,N_912);
nor U1789 (N_1789,N_421,N_794);
nand U1790 (N_1790,N_630,N_839);
xnor U1791 (N_1791,N_470,N_730);
or U1792 (N_1792,N_295,N_439);
nand U1793 (N_1793,N_283,N_227);
nand U1794 (N_1794,N_40,N_214);
or U1795 (N_1795,N_709,N_703);
nand U1796 (N_1796,N_381,N_899);
or U1797 (N_1797,N_333,N_594);
nor U1798 (N_1798,N_392,N_468);
nand U1799 (N_1799,N_55,N_407);
and U1800 (N_1800,N_826,N_919);
or U1801 (N_1801,N_762,N_117);
and U1802 (N_1802,N_330,N_470);
and U1803 (N_1803,N_841,N_221);
or U1804 (N_1804,N_87,N_634);
nand U1805 (N_1805,N_161,N_213);
nor U1806 (N_1806,N_691,N_199);
nor U1807 (N_1807,N_466,N_658);
nand U1808 (N_1808,N_27,N_499);
nand U1809 (N_1809,N_780,N_760);
nand U1810 (N_1810,N_568,N_950);
nand U1811 (N_1811,N_539,N_251);
or U1812 (N_1812,N_222,N_331);
and U1813 (N_1813,N_707,N_749);
nor U1814 (N_1814,N_444,N_435);
or U1815 (N_1815,N_392,N_367);
or U1816 (N_1816,N_755,N_915);
or U1817 (N_1817,N_855,N_536);
xnor U1818 (N_1818,N_756,N_183);
or U1819 (N_1819,N_1,N_691);
and U1820 (N_1820,N_951,N_409);
nor U1821 (N_1821,N_414,N_654);
and U1822 (N_1822,N_641,N_427);
xor U1823 (N_1823,N_179,N_213);
and U1824 (N_1824,N_487,N_301);
or U1825 (N_1825,N_251,N_213);
and U1826 (N_1826,N_836,N_346);
xnor U1827 (N_1827,N_605,N_47);
or U1828 (N_1828,N_918,N_543);
nand U1829 (N_1829,N_673,N_525);
nor U1830 (N_1830,N_274,N_229);
and U1831 (N_1831,N_545,N_931);
or U1832 (N_1832,N_79,N_944);
or U1833 (N_1833,N_935,N_382);
nand U1834 (N_1834,N_252,N_813);
or U1835 (N_1835,N_979,N_624);
xor U1836 (N_1836,N_858,N_948);
nor U1837 (N_1837,N_424,N_894);
and U1838 (N_1838,N_327,N_468);
nor U1839 (N_1839,N_690,N_101);
and U1840 (N_1840,N_805,N_335);
nand U1841 (N_1841,N_611,N_845);
or U1842 (N_1842,N_418,N_740);
nor U1843 (N_1843,N_560,N_869);
or U1844 (N_1844,N_942,N_256);
or U1845 (N_1845,N_460,N_230);
nor U1846 (N_1846,N_198,N_117);
or U1847 (N_1847,N_720,N_824);
nor U1848 (N_1848,N_160,N_818);
and U1849 (N_1849,N_41,N_698);
nand U1850 (N_1850,N_992,N_431);
nor U1851 (N_1851,N_631,N_387);
nand U1852 (N_1852,N_208,N_360);
or U1853 (N_1853,N_117,N_448);
nor U1854 (N_1854,N_42,N_552);
nand U1855 (N_1855,N_406,N_197);
and U1856 (N_1856,N_168,N_146);
nand U1857 (N_1857,N_390,N_14);
or U1858 (N_1858,N_496,N_152);
nor U1859 (N_1859,N_598,N_872);
and U1860 (N_1860,N_941,N_263);
nand U1861 (N_1861,N_461,N_653);
nand U1862 (N_1862,N_76,N_415);
nor U1863 (N_1863,N_712,N_483);
or U1864 (N_1864,N_660,N_397);
or U1865 (N_1865,N_587,N_228);
and U1866 (N_1866,N_749,N_150);
nor U1867 (N_1867,N_695,N_9);
nand U1868 (N_1868,N_186,N_129);
nor U1869 (N_1869,N_842,N_352);
and U1870 (N_1870,N_529,N_481);
or U1871 (N_1871,N_358,N_486);
nor U1872 (N_1872,N_546,N_60);
nor U1873 (N_1873,N_255,N_771);
nor U1874 (N_1874,N_958,N_977);
nand U1875 (N_1875,N_669,N_681);
nand U1876 (N_1876,N_776,N_710);
and U1877 (N_1877,N_515,N_381);
nand U1878 (N_1878,N_366,N_213);
or U1879 (N_1879,N_962,N_660);
and U1880 (N_1880,N_690,N_297);
or U1881 (N_1881,N_490,N_682);
nand U1882 (N_1882,N_445,N_56);
or U1883 (N_1883,N_701,N_885);
or U1884 (N_1884,N_612,N_817);
and U1885 (N_1885,N_960,N_125);
nand U1886 (N_1886,N_601,N_761);
or U1887 (N_1887,N_610,N_888);
nor U1888 (N_1888,N_783,N_802);
and U1889 (N_1889,N_377,N_795);
and U1890 (N_1890,N_93,N_506);
and U1891 (N_1891,N_96,N_442);
nor U1892 (N_1892,N_667,N_906);
and U1893 (N_1893,N_449,N_343);
or U1894 (N_1894,N_52,N_348);
nor U1895 (N_1895,N_234,N_583);
or U1896 (N_1896,N_554,N_311);
nand U1897 (N_1897,N_489,N_225);
nor U1898 (N_1898,N_226,N_801);
or U1899 (N_1899,N_309,N_447);
xnor U1900 (N_1900,N_406,N_160);
nor U1901 (N_1901,N_779,N_654);
nor U1902 (N_1902,N_325,N_721);
nand U1903 (N_1903,N_994,N_148);
and U1904 (N_1904,N_450,N_555);
nand U1905 (N_1905,N_396,N_223);
nand U1906 (N_1906,N_751,N_397);
nand U1907 (N_1907,N_384,N_980);
or U1908 (N_1908,N_777,N_566);
nor U1909 (N_1909,N_546,N_711);
nand U1910 (N_1910,N_833,N_380);
nor U1911 (N_1911,N_189,N_407);
nor U1912 (N_1912,N_722,N_636);
and U1913 (N_1913,N_882,N_935);
or U1914 (N_1914,N_270,N_729);
and U1915 (N_1915,N_409,N_513);
xor U1916 (N_1916,N_584,N_913);
xor U1917 (N_1917,N_36,N_773);
nor U1918 (N_1918,N_804,N_736);
nand U1919 (N_1919,N_69,N_607);
xor U1920 (N_1920,N_814,N_925);
or U1921 (N_1921,N_21,N_222);
nand U1922 (N_1922,N_343,N_716);
or U1923 (N_1923,N_199,N_643);
nand U1924 (N_1924,N_61,N_734);
nor U1925 (N_1925,N_62,N_397);
xnor U1926 (N_1926,N_133,N_491);
xor U1927 (N_1927,N_801,N_892);
or U1928 (N_1928,N_223,N_322);
nor U1929 (N_1929,N_672,N_41);
and U1930 (N_1930,N_59,N_650);
or U1931 (N_1931,N_409,N_152);
and U1932 (N_1932,N_505,N_560);
or U1933 (N_1933,N_486,N_266);
nor U1934 (N_1934,N_493,N_312);
or U1935 (N_1935,N_914,N_883);
or U1936 (N_1936,N_872,N_377);
nor U1937 (N_1937,N_691,N_517);
or U1938 (N_1938,N_496,N_30);
and U1939 (N_1939,N_852,N_124);
and U1940 (N_1940,N_677,N_542);
and U1941 (N_1941,N_101,N_88);
nand U1942 (N_1942,N_128,N_580);
nor U1943 (N_1943,N_898,N_603);
xnor U1944 (N_1944,N_709,N_946);
xor U1945 (N_1945,N_783,N_449);
or U1946 (N_1946,N_266,N_263);
nor U1947 (N_1947,N_566,N_850);
nor U1948 (N_1948,N_48,N_476);
xor U1949 (N_1949,N_373,N_221);
or U1950 (N_1950,N_120,N_142);
nand U1951 (N_1951,N_325,N_418);
nor U1952 (N_1952,N_352,N_723);
or U1953 (N_1953,N_580,N_159);
and U1954 (N_1954,N_931,N_23);
and U1955 (N_1955,N_757,N_728);
or U1956 (N_1956,N_701,N_162);
or U1957 (N_1957,N_81,N_624);
nand U1958 (N_1958,N_248,N_752);
nor U1959 (N_1959,N_279,N_670);
nand U1960 (N_1960,N_537,N_532);
nor U1961 (N_1961,N_277,N_981);
nand U1962 (N_1962,N_591,N_585);
and U1963 (N_1963,N_570,N_34);
nor U1964 (N_1964,N_351,N_125);
nor U1965 (N_1965,N_618,N_634);
nor U1966 (N_1966,N_741,N_393);
or U1967 (N_1967,N_995,N_220);
nand U1968 (N_1968,N_38,N_884);
and U1969 (N_1969,N_31,N_847);
and U1970 (N_1970,N_349,N_891);
or U1971 (N_1971,N_151,N_800);
nand U1972 (N_1972,N_187,N_717);
and U1973 (N_1973,N_347,N_598);
nand U1974 (N_1974,N_782,N_637);
or U1975 (N_1975,N_185,N_854);
nand U1976 (N_1976,N_64,N_10);
nor U1977 (N_1977,N_604,N_454);
nor U1978 (N_1978,N_366,N_950);
and U1979 (N_1979,N_340,N_575);
nand U1980 (N_1980,N_484,N_540);
xnor U1981 (N_1981,N_217,N_645);
xnor U1982 (N_1982,N_502,N_6);
nor U1983 (N_1983,N_76,N_698);
xnor U1984 (N_1984,N_148,N_147);
and U1985 (N_1985,N_58,N_229);
and U1986 (N_1986,N_221,N_624);
and U1987 (N_1987,N_176,N_186);
or U1988 (N_1988,N_262,N_282);
or U1989 (N_1989,N_502,N_715);
nand U1990 (N_1990,N_983,N_423);
xnor U1991 (N_1991,N_540,N_588);
nor U1992 (N_1992,N_998,N_285);
and U1993 (N_1993,N_274,N_397);
nor U1994 (N_1994,N_86,N_603);
nand U1995 (N_1995,N_258,N_790);
or U1996 (N_1996,N_583,N_697);
nand U1997 (N_1997,N_151,N_676);
nor U1998 (N_1998,N_225,N_507);
and U1999 (N_1999,N_498,N_665);
or U2000 (N_2000,N_1833,N_1948);
nor U2001 (N_2001,N_1643,N_1990);
or U2002 (N_2002,N_1563,N_1575);
and U2003 (N_2003,N_1526,N_1440);
xnor U2004 (N_2004,N_1172,N_1959);
nor U2005 (N_2005,N_1475,N_1284);
nor U2006 (N_2006,N_1272,N_1546);
xor U2007 (N_2007,N_1862,N_1216);
and U2008 (N_2008,N_1908,N_1049);
nor U2009 (N_2009,N_1950,N_1285);
or U2010 (N_2010,N_1421,N_1616);
xnor U2011 (N_2011,N_1792,N_1749);
or U2012 (N_2012,N_1168,N_1112);
nand U2013 (N_2013,N_1394,N_1263);
and U2014 (N_2014,N_1785,N_1422);
nor U2015 (N_2015,N_1859,N_1732);
and U2016 (N_2016,N_1283,N_1254);
nor U2017 (N_2017,N_1371,N_1884);
xnor U2018 (N_2018,N_1712,N_1387);
and U2019 (N_2019,N_1495,N_1138);
nor U2020 (N_2020,N_1695,N_1032);
nor U2021 (N_2021,N_1095,N_1404);
and U2022 (N_2022,N_1600,N_1516);
nand U2023 (N_2023,N_1758,N_1364);
and U2024 (N_2024,N_1152,N_1562);
or U2025 (N_2025,N_1971,N_1150);
nand U2026 (N_2026,N_1092,N_1524);
or U2027 (N_2027,N_1123,N_1228);
or U2028 (N_2028,N_1299,N_1343);
or U2029 (N_2029,N_1824,N_1587);
nand U2030 (N_2030,N_1718,N_1273);
nor U2031 (N_2031,N_1504,N_1076);
or U2032 (N_2032,N_1756,N_1435);
and U2033 (N_2033,N_1484,N_1264);
nand U2034 (N_2034,N_1480,N_1182);
or U2035 (N_2035,N_1117,N_1292);
or U2036 (N_2036,N_1115,N_1847);
or U2037 (N_2037,N_1790,N_1459);
or U2038 (N_2038,N_1019,N_1669);
nand U2039 (N_2039,N_1752,N_1428);
or U2040 (N_2040,N_1318,N_1518);
nand U2041 (N_2041,N_1417,N_1881);
and U2042 (N_2042,N_1736,N_1259);
or U2043 (N_2043,N_1572,N_1576);
and U2044 (N_2044,N_1864,N_1287);
nor U2045 (N_2045,N_1485,N_1746);
nor U2046 (N_2046,N_1072,N_1844);
nand U2047 (N_2047,N_1629,N_1193);
or U2048 (N_2048,N_1674,N_1458);
and U2049 (N_2049,N_1224,N_1532);
xnor U2050 (N_2050,N_1602,N_1125);
and U2051 (N_2051,N_1256,N_1826);
or U2052 (N_2052,N_1769,N_1313);
xor U2053 (N_2053,N_1953,N_1728);
or U2054 (N_2054,N_1657,N_1385);
or U2055 (N_2055,N_1090,N_1091);
or U2056 (N_2056,N_1678,N_1099);
or U2057 (N_2057,N_1347,N_1561);
or U2058 (N_2058,N_1337,N_1835);
xor U2059 (N_2059,N_1604,N_1325);
nor U2060 (N_2060,N_1455,N_1799);
xor U2061 (N_2061,N_1593,N_1231);
nor U2062 (N_2062,N_1633,N_1613);
nor U2063 (N_2063,N_1734,N_1836);
and U2064 (N_2064,N_1995,N_1900);
or U2065 (N_2065,N_1582,N_1101);
nand U2066 (N_2066,N_1146,N_1567);
nand U2067 (N_2067,N_1609,N_1490);
and U2068 (N_2068,N_1447,N_1324);
or U2069 (N_2069,N_1743,N_1830);
nand U2070 (N_2070,N_1926,N_1724);
or U2071 (N_2071,N_1437,N_1492);
or U2072 (N_2072,N_1828,N_1584);
or U2073 (N_2073,N_1260,N_1751);
and U2074 (N_2074,N_1628,N_1442);
or U2075 (N_2075,N_1787,N_1288);
or U2076 (N_2076,N_1329,N_1837);
nand U2077 (N_2077,N_1086,N_1088);
nand U2078 (N_2078,N_1491,N_1244);
and U2079 (N_2079,N_1658,N_1432);
or U2080 (N_2080,N_1187,N_1396);
nand U2081 (N_2081,N_1986,N_1973);
xor U2082 (N_2082,N_1006,N_1649);
and U2083 (N_2083,N_1477,N_1391);
or U2084 (N_2084,N_1365,N_1931);
and U2085 (N_2085,N_1652,N_1411);
nand U2086 (N_2086,N_1850,N_1321);
nor U2087 (N_2087,N_1191,N_1543);
nor U2088 (N_2088,N_1098,N_1741);
nor U2089 (N_2089,N_1975,N_1726);
or U2090 (N_2090,N_1399,N_1816);
xnor U2091 (N_2091,N_1974,N_1109);
nand U2092 (N_2092,N_1819,N_1426);
and U2093 (N_2093,N_1834,N_1009);
and U2094 (N_2094,N_1498,N_1813);
and U2095 (N_2095,N_1661,N_1320);
and U2096 (N_2096,N_1965,N_1692);
xnor U2097 (N_2097,N_1290,N_1755);
nand U2098 (N_2098,N_1598,N_1463);
nand U2099 (N_2099,N_1552,N_1048);
and U2100 (N_2100,N_1814,N_1199);
or U2101 (N_2101,N_1248,N_1467);
or U2102 (N_2102,N_1856,N_1858);
nand U2103 (N_2103,N_1877,N_1470);
nor U2104 (N_2104,N_1512,N_1868);
and U2105 (N_2105,N_1945,N_1219);
nand U2106 (N_2106,N_1849,N_1777);
nand U2107 (N_2107,N_1345,N_1988);
nand U2108 (N_2108,N_1348,N_1664);
and U2109 (N_2109,N_1124,N_1876);
nor U2110 (N_2110,N_1209,N_1653);
xnor U2111 (N_2111,N_1855,N_1829);
nand U2112 (N_2112,N_1686,N_1185);
and U2113 (N_2113,N_1153,N_1240);
nand U2114 (N_2114,N_1111,N_1780);
nor U2115 (N_2115,N_1748,N_1427);
nor U2116 (N_2116,N_1719,N_1118);
and U2117 (N_2117,N_1433,N_1760);
nor U2118 (N_2118,N_1171,N_1960);
nand U2119 (N_2119,N_1169,N_1625);
nor U2120 (N_2120,N_1984,N_1978);
nor U2121 (N_2121,N_1818,N_1204);
and U2122 (N_2122,N_1599,N_1201);
and U2123 (N_2123,N_1456,N_1805);
and U2124 (N_2124,N_1899,N_1367);
and U2125 (N_2125,N_1632,N_1671);
and U2126 (N_2126,N_1815,N_1865);
nor U2127 (N_2127,N_1061,N_1142);
nand U2128 (N_2128,N_1523,N_1885);
and U2129 (N_2129,N_1810,N_1392);
and U2130 (N_2130,N_1670,N_1703);
nor U2131 (N_2131,N_1772,N_1537);
nand U2132 (N_2132,N_1175,N_1449);
nor U2133 (N_2133,N_1872,N_1226);
and U2134 (N_2134,N_1497,N_1461);
xnor U2135 (N_2135,N_1473,N_1326);
or U2136 (N_2136,N_1615,N_1162);
xnor U2137 (N_2137,N_1566,N_1745);
xnor U2138 (N_2138,N_1667,N_1972);
xor U2139 (N_2139,N_1544,N_1301);
and U2140 (N_2140,N_1921,N_1358);
nor U2141 (N_2141,N_1909,N_1237);
xor U2142 (N_2142,N_1050,N_1603);
xnor U2143 (N_2143,N_1932,N_1639);
nand U2144 (N_2144,N_1549,N_1383);
and U2145 (N_2145,N_1608,N_1571);
xor U2146 (N_2146,N_1779,N_1373);
nor U2147 (N_2147,N_1957,N_1462);
nand U2148 (N_2148,N_1937,N_1481);
nand U2149 (N_2149,N_1964,N_1400);
nand U2150 (N_2150,N_1378,N_1514);
nor U2151 (N_2151,N_1419,N_1155);
nand U2152 (N_2152,N_1701,N_1023);
nor U2153 (N_2153,N_1406,N_1483);
or U2154 (N_2154,N_1954,N_1793);
nor U2155 (N_2155,N_1531,N_1731);
and U2156 (N_2156,N_1360,N_1113);
nor U2157 (N_2157,N_1100,N_1520);
nor U2158 (N_2158,N_1807,N_1194);
or U2159 (N_2159,N_1918,N_1294);
nor U2160 (N_2160,N_1474,N_1160);
or U2161 (N_2161,N_1716,N_1782);
and U2162 (N_2162,N_1870,N_1302);
nor U2163 (N_2163,N_1528,N_1203);
nor U2164 (N_2164,N_1243,N_1108);
or U2165 (N_2165,N_1103,N_1460);
nand U2166 (N_2166,N_1725,N_1840);
nor U2167 (N_2167,N_1466,N_1135);
or U2168 (N_2168,N_1660,N_1941);
nand U2169 (N_2169,N_1179,N_1992);
or U2170 (N_2170,N_1943,N_1143);
and U2171 (N_2171,N_1246,N_1403);
and U2172 (N_2172,N_1409,N_1554);
and U2173 (N_2173,N_1936,N_1129);
or U2174 (N_2174,N_1457,N_1611);
xnor U2175 (N_2175,N_1017,N_1890);
nand U2176 (N_2176,N_1407,N_1940);
nor U2177 (N_2177,N_1277,N_1683);
nand U2178 (N_2178,N_1097,N_1647);
or U2179 (N_2179,N_1910,N_1158);
nor U2180 (N_2180,N_1083,N_1357);
xor U2181 (N_2181,N_1105,N_1798);
or U2182 (N_2182,N_1797,N_1375);
or U2183 (N_2183,N_1355,N_1700);
and U2184 (N_2184,N_1454,N_1882);
nor U2185 (N_2185,N_1672,N_1778);
nand U2186 (N_2186,N_1036,N_1699);
nor U2187 (N_2187,N_1052,N_1525);
or U2188 (N_2188,N_1156,N_1080);
nand U2189 (N_2189,N_1096,N_1744);
or U2190 (N_2190,N_1223,N_1874);
xor U2191 (N_2191,N_1126,N_1222);
and U2192 (N_2192,N_1202,N_1676);
nand U2193 (N_2193,N_1916,N_1236);
nor U2194 (N_2194,N_1641,N_1585);
nand U2195 (N_2195,N_1693,N_1315);
xnor U2196 (N_2196,N_1705,N_1892);
or U2197 (N_2197,N_1586,N_1107);
and U2198 (N_2198,N_1879,N_1128);
nor U2199 (N_2199,N_1564,N_1691);
or U2200 (N_2200,N_1255,N_1843);
and U2201 (N_2201,N_1891,N_1211);
and U2202 (N_2202,N_1607,N_1328);
nor U2203 (N_2203,N_1188,N_1165);
nand U2204 (N_2204,N_1293,N_1003);
and U2205 (N_2205,N_1073,N_1178);
or U2206 (N_2206,N_1210,N_1962);
and U2207 (N_2207,N_1522,N_1077);
nor U2208 (N_2208,N_1521,N_1413);
nand U2209 (N_2209,N_1689,N_1687);
or U2210 (N_2210,N_1920,N_1763);
nand U2211 (N_2211,N_1527,N_1684);
nand U2212 (N_2212,N_1180,N_1359);
nor U2213 (N_2213,N_1637,N_1913);
nor U2214 (N_2214,N_1742,N_1055);
nor U2215 (N_2215,N_1043,N_1016);
nor U2216 (N_2216,N_1606,N_1853);
nand U2217 (N_2217,N_1468,N_1140);
nand U2218 (N_2218,N_1651,N_1279);
nor U2219 (N_2219,N_1266,N_1548);
xnor U2220 (N_2220,N_1331,N_1645);
and U2221 (N_2221,N_1738,N_1808);
and U2222 (N_2222,N_1297,N_1114);
or U2223 (N_2223,N_1912,N_1247);
nor U2224 (N_2224,N_1542,N_1154);
and U2225 (N_2225,N_1577,N_1754);
nand U2226 (N_2226,N_1996,N_1698);
nand U2227 (N_2227,N_1389,N_1919);
and U2228 (N_2228,N_1070,N_1045);
and U2229 (N_2229,N_1866,N_1192);
nor U2230 (N_2230,N_1911,N_1638);
or U2231 (N_2231,N_1424,N_1679);
nand U2232 (N_2232,N_1614,N_1361);
nor U2233 (N_2233,N_1106,N_1878);
or U2234 (N_2234,N_1452,N_1104);
or U2235 (N_2235,N_1028,N_1008);
nor U2236 (N_2236,N_1570,N_1282);
nand U2237 (N_2237,N_1014,N_1081);
nand U2238 (N_2238,N_1905,N_1875);
xnor U2239 (N_2239,N_1267,N_1377);
nand U2240 (N_2240,N_1323,N_1047);
or U2241 (N_2241,N_1958,N_1886);
nor U2242 (N_2242,N_1565,N_1517);
and U2243 (N_2243,N_1997,N_1478);
and U2244 (N_2244,N_1136,N_1225);
nand U2245 (N_2245,N_1949,N_1341);
and U2246 (N_2246,N_1704,N_1644);
and U2247 (N_2247,N_1583,N_1213);
nor U2248 (N_2248,N_1665,N_1416);
and U2249 (N_2249,N_1821,N_1601);
xor U2250 (N_2250,N_1472,N_1852);
nand U2251 (N_2251,N_1306,N_1464);
or U2252 (N_2252,N_1708,N_1507);
or U2253 (N_2253,N_1229,N_1386);
nand U2254 (N_2254,N_1854,N_1783);
and U2255 (N_2255,N_1027,N_1983);
nand U2256 (N_2256,N_1740,N_1038);
or U2257 (N_2257,N_1308,N_1515);
xnor U2258 (N_2258,N_1354,N_1873);
nor U2259 (N_2259,N_1093,N_1506);
or U2260 (N_2260,N_1084,N_1541);
or U2261 (N_2261,N_1794,N_1057);
or U2262 (N_2262,N_1502,N_1771);
nor U2263 (N_2263,N_1619,N_1977);
nor U2264 (N_2264,N_1144,N_1902);
nand U2265 (N_2265,N_1271,N_1163);
nor U2266 (N_2266,N_1773,N_1967);
or U2267 (N_2267,N_1924,N_1767);
nor U2268 (N_2268,N_1309,N_1976);
nand U2269 (N_2269,N_1888,N_1883);
nand U2270 (N_2270,N_1690,N_1446);
or U2271 (N_2271,N_1078,N_1650);
and U2272 (N_2272,N_1401,N_1476);
nor U2273 (N_2273,N_1319,N_1946);
nor U2274 (N_2274,N_1827,N_1774);
and U2275 (N_2275,N_1519,N_1018);
nor U2276 (N_2276,N_1594,N_1089);
nor U2277 (N_2277,N_1901,N_1344);
or U2278 (N_2278,N_1781,N_1654);
and U2279 (N_2279,N_1534,N_1333);
and U2280 (N_2280,N_1711,N_1044);
nor U2281 (N_2281,N_1167,N_1961);
or U2282 (N_2282,N_1300,N_1925);
and U2283 (N_2283,N_1035,N_1021);
nand U2284 (N_2284,N_1212,N_1764);
nand U2285 (N_2285,N_1147,N_1860);
nor U2286 (N_2286,N_1494,N_1304);
nand U2287 (N_2287,N_1381,N_1249);
nand U2288 (N_2288,N_1697,N_1176);
and U2289 (N_2289,N_1710,N_1930);
or U2290 (N_2290,N_1227,N_1568);
xnor U2291 (N_2291,N_1635,N_1803);
or U2292 (N_2292,N_1831,N_1039);
xnor U2293 (N_2293,N_1806,N_1370);
and U2294 (N_2294,N_1947,N_1423);
xor U2295 (N_2295,N_1183,N_1617);
or U2296 (N_2296,N_1120,N_1897);
nor U2297 (N_2297,N_1336,N_1938);
xor U2298 (N_2298,N_1620,N_1677);
nor U2299 (N_2299,N_1591,N_1757);
nor U2300 (N_2300,N_1317,N_1922);
nand U2301 (N_2301,N_1513,N_1753);
or U2302 (N_2302,N_1075,N_1245);
nand U2303 (N_2303,N_1031,N_1966);
or U2304 (N_2304,N_1714,N_1007);
nor U2305 (N_2305,N_1206,N_1904);
nand U2306 (N_2306,N_1332,N_1215);
xnor U2307 (N_2307,N_1342,N_1270);
or U2308 (N_2308,N_1362,N_1241);
and U2309 (N_2309,N_1207,N_1857);
nor U2310 (N_2310,N_1715,N_1917);
xor U2311 (N_2311,N_1012,N_1968);
nand U2312 (N_2312,N_1707,N_1436);
nand U2313 (N_2313,N_1379,N_1776);
or U2314 (N_2314,N_1041,N_1220);
or U2315 (N_2315,N_1274,N_1559);
nand U2316 (N_2316,N_1157,N_1214);
nor U2317 (N_2317,N_1952,N_1574);
nand U2318 (N_2318,N_1186,N_1907);
nand U2319 (N_2319,N_1750,N_1388);
and U2320 (N_2320,N_1982,N_1702);
and U2321 (N_2321,N_1251,N_1955);
xor U2322 (N_2322,N_1051,N_1685);
or U2323 (N_2323,N_1346,N_1311);
and U2324 (N_2324,N_1863,N_1681);
or U2325 (N_2325,N_1933,N_1762);
nand U2326 (N_2326,N_1479,N_1682);
xnor U2327 (N_2327,N_1327,N_1026);
nand U2328 (N_2328,N_1030,N_1141);
or U2329 (N_2329,N_1139,N_1405);
or U2330 (N_2330,N_1706,N_1987);
nand U2331 (N_2331,N_1130,N_1727);
and U2332 (N_2332,N_1296,N_1801);
and U2333 (N_2333,N_1253,N_1448);
nor U2334 (N_2334,N_1942,N_1232);
nor U2335 (N_2335,N_1087,N_1981);
nand U2336 (N_2336,N_1197,N_1894);
xnor U2337 (N_2337,N_1286,N_1013);
and U2338 (N_2338,N_1024,N_1796);
nor U2339 (N_2339,N_1802,N_1074);
nor U2340 (N_2340,N_1970,N_1597);
or U2341 (N_2341,N_1250,N_1149);
xnor U2342 (N_2342,N_1791,N_1914);
xor U2343 (N_2343,N_1334,N_1867);
nand U2344 (N_2344,N_1208,N_1861);
or U2345 (N_2345,N_1845,N_1842);
nand U2346 (N_2346,N_1261,N_1486);
or U2347 (N_2347,N_1001,N_1636);
and U2348 (N_2348,N_1005,N_1372);
or U2349 (N_2349,N_1289,N_1058);
or U2350 (N_2350,N_1848,N_1322);
xnor U2351 (N_2351,N_1989,N_1065);
nand U2352 (N_2352,N_1985,N_1280);
or U2353 (N_2353,N_1316,N_1596);
nand U2354 (N_2354,N_1713,N_1430);
nor U2355 (N_2355,N_1717,N_1042);
or U2356 (N_2356,N_1553,N_1369);
nand U2357 (N_2357,N_1631,N_1376);
or U2358 (N_2358,N_1173,N_1438);
nor U2359 (N_2359,N_1735,N_1656);
and U2360 (N_2360,N_1127,N_1268);
and U2361 (N_2361,N_1662,N_1994);
nand U2362 (N_2362,N_1605,N_1465);
nand U2363 (N_2363,N_1257,N_1122);
nand U2364 (N_2364,N_1906,N_1339);
or U2365 (N_2365,N_1999,N_1159);
xor U2366 (N_2366,N_1443,N_1721);
xor U2367 (N_2367,N_1094,N_1121);
and U2368 (N_2368,N_1295,N_1846);
or U2369 (N_2369,N_1589,N_1530);
nor U2370 (N_2370,N_1063,N_1189);
or U2371 (N_2371,N_1812,N_1281);
and U2372 (N_2372,N_1896,N_1184);
and U2373 (N_2373,N_1062,N_1418);
and U2374 (N_2374,N_1694,N_1927);
or U2375 (N_2375,N_1618,N_1759);
or U2376 (N_2376,N_1451,N_1547);
nor U2377 (N_2377,N_1439,N_1696);
or U2378 (N_2378,N_1545,N_1068);
nor U2379 (N_2379,N_1174,N_1923);
nand U2380 (N_2380,N_1034,N_1434);
or U2381 (N_2381,N_1397,N_1119);
nor U2382 (N_2382,N_1276,N_1823);
nor U2383 (N_2383,N_1022,N_1310);
nor U2384 (N_2384,N_1059,N_1148);
nor U2385 (N_2385,N_1487,N_1217);
nor U2386 (N_2386,N_1993,N_1181);
xnor U2387 (N_2387,N_1053,N_1800);
xor U2388 (N_2388,N_1675,N_1822);
xor U2389 (N_2389,N_1258,N_1221);
or U2390 (N_2390,N_1511,N_1166);
nor U2391 (N_2391,N_1010,N_1588);
nand U2392 (N_2392,N_1770,N_1500);
and U2393 (N_2393,N_1402,N_1415);
nand U2394 (N_2394,N_1196,N_1839);
and U2395 (N_2395,N_1356,N_1889);
and U2396 (N_2396,N_1929,N_1811);
and U2397 (N_2397,N_1275,N_1131);
and U2398 (N_2398,N_1569,N_1556);
nor U2399 (N_2399,N_1505,N_1020);
nand U2400 (N_2400,N_1789,N_1000);
nor U2401 (N_2401,N_1841,N_1085);
nor U2402 (N_2402,N_1340,N_1151);
or U2403 (N_2403,N_1659,N_1979);
nor U2404 (N_2404,N_1538,N_1765);
and U2405 (N_2405,N_1015,N_1352);
nand U2406 (N_2406,N_1382,N_1626);
and U2407 (N_2407,N_1627,N_1335);
or U2408 (N_2408,N_1412,N_1508);
nand U2409 (N_2409,N_1624,N_1642);
or U2410 (N_2410,N_1238,N_1673);
xor U2411 (N_2411,N_1558,N_1775);
or U2412 (N_2412,N_1262,N_1723);
nor U2413 (N_2413,N_1116,N_1205);
nor U2414 (N_2414,N_1488,N_1011);
nand U2415 (N_2415,N_1134,N_1366);
nand U2416 (N_2416,N_1145,N_1398);
or U2417 (N_2417,N_1234,N_1655);
nand U2418 (N_2418,N_1529,N_1198);
nor U2419 (N_2419,N_1539,N_1298);
nor U2420 (N_2420,N_1969,N_1832);
or U2421 (N_2421,N_1869,N_1838);
and U2422 (N_2422,N_1503,N_1557);
or U2423 (N_2423,N_1935,N_1349);
nor U2424 (N_2424,N_1580,N_1200);
xnor U2425 (N_2425,N_1560,N_1368);
or U2426 (N_2426,N_1510,N_1766);
or U2427 (N_2427,N_1177,N_1795);
nor U2428 (N_2428,N_1786,N_1420);
or U2429 (N_2429,N_1393,N_1688);
nand U2430 (N_2430,N_1573,N_1610);
nor U2431 (N_2431,N_1509,N_1110);
or U2432 (N_2432,N_1056,N_1944);
or U2433 (N_2433,N_1002,N_1265);
or U2434 (N_2434,N_1501,N_1825);
or U2435 (N_2435,N_1278,N_1425);
nor U2436 (N_2436,N_1729,N_1761);
or U2437 (N_2437,N_1893,N_1046);
nor U2438 (N_2438,N_1195,N_1312);
or U2439 (N_2439,N_1330,N_1351);
xnor U2440 (N_2440,N_1132,N_1747);
nand U2441 (N_2441,N_1064,N_1029);
xnor U2442 (N_2442,N_1668,N_1471);
xnor U2443 (N_2443,N_1499,N_1071);
nor U2444 (N_2444,N_1784,N_1380);
and U2445 (N_2445,N_1956,N_1303);
nor U2446 (N_2446,N_1663,N_1535);
or U2447 (N_2447,N_1579,N_1350);
nand U2448 (N_2448,N_1739,N_1737);
or U2449 (N_2449,N_1429,N_1252);
xnor U2450 (N_2450,N_1581,N_1450);
or U2451 (N_2451,N_1037,N_1934);
nand U2452 (N_2452,N_1733,N_1060);
and U2453 (N_2453,N_1998,N_1666);
and U2454 (N_2454,N_1242,N_1493);
nand U2455 (N_2455,N_1218,N_1305);
nor U2456 (N_2456,N_1079,N_1054);
nor U2457 (N_2457,N_1623,N_1871);
nor U2458 (N_2458,N_1768,N_1851);
nand U2459 (N_2459,N_1040,N_1536);
nor U2460 (N_2460,N_1338,N_1991);
and U2461 (N_2461,N_1307,N_1069);
or U2462 (N_2462,N_1887,N_1489);
and U2463 (N_2463,N_1395,N_1314);
xor U2464 (N_2464,N_1550,N_1555);
nor U2465 (N_2465,N_1578,N_1033);
xor U2466 (N_2466,N_1809,N_1137);
xor U2467 (N_2467,N_1634,N_1190);
and U2468 (N_2468,N_1648,N_1431);
nor U2469 (N_2469,N_1592,N_1533);
and U2470 (N_2470,N_1353,N_1363);
nor U2471 (N_2471,N_1408,N_1164);
nor U2472 (N_2472,N_1170,N_1709);
xor U2473 (N_2473,N_1239,N_1939);
xnor U2474 (N_2474,N_1482,N_1898);
xnor U2475 (N_2475,N_1233,N_1680);
nand U2476 (N_2476,N_1067,N_1230);
nand U2477 (N_2477,N_1082,N_1595);
nand U2478 (N_2478,N_1469,N_1880);
nor U2479 (N_2479,N_1730,N_1903);
and U2480 (N_2480,N_1820,N_1928);
or U2481 (N_2481,N_1025,N_1788);
nor U2482 (N_2482,N_1590,N_1004);
nor U2483 (N_2483,N_1630,N_1804);
nand U2484 (N_2484,N_1817,N_1640);
nor U2485 (N_2485,N_1269,N_1414);
nand U2486 (N_2486,N_1720,N_1980);
nand U2487 (N_2487,N_1410,N_1540);
nand U2488 (N_2488,N_1622,N_1612);
nor U2489 (N_2489,N_1963,N_1621);
nand U2490 (N_2490,N_1390,N_1102);
nor U2491 (N_2491,N_1161,N_1551);
or U2492 (N_2492,N_1895,N_1441);
nor U2493 (N_2493,N_1444,N_1235);
or U2494 (N_2494,N_1646,N_1951);
nand U2495 (N_2495,N_1133,N_1915);
or U2496 (N_2496,N_1445,N_1066);
or U2497 (N_2497,N_1384,N_1453);
nor U2498 (N_2498,N_1291,N_1496);
xor U2499 (N_2499,N_1722,N_1374);
nand U2500 (N_2500,N_1902,N_1602);
and U2501 (N_2501,N_1382,N_1852);
or U2502 (N_2502,N_1679,N_1537);
or U2503 (N_2503,N_1876,N_1345);
nor U2504 (N_2504,N_1300,N_1531);
and U2505 (N_2505,N_1804,N_1077);
or U2506 (N_2506,N_1908,N_1489);
nor U2507 (N_2507,N_1839,N_1799);
nand U2508 (N_2508,N_1711,N_1331);
and U2509 (N_2509,N_1741,N_1825);
nand U2510 (N_2510,N_1400,N_1910);
xor U2511 (N_2511,N_1873,N_1194);
nor U2512 (N_2512,N_1763,N_1314);
nor U2513 (N_2513,N_1845,N_1743);
nor U2514 (N_2514,N_1260,N_1684);
or U2515 (N_2515,N_1369,N_1321);
nand U2516 (N_2516,N_1434,N_1025);
nor U2517 (N_2517,N_1507,N_1954);
nor U2518 (N_2518,N_1797,N_1145);
nand U2519 (N_2519,N_1928,N_1089);
and U2520 (N_2520,N_1669,N_1947);
and U2521 (N_2521,N_1467,N_1217);
nor U2522 (N_2522,N_1769,N_1833);
and U2523 (N_2523,N_1932,N_1059);
and U2524 (N_2524,N_1656,N_1937);
nand U2525 (N_2525,N_1597,N_1020);
or U2526 (N_2526,N_1479,N_1041);
and U2527 (N_2527,N_1457,N_1810);
nor U2528 (N_2528,N_1473,N_1968);
nand U2529 (N_2529,N_1414,N_1223);
nand U2530 (N_2530,N_1504,N_1910);
or U2531 (N_2531,N_1546,N_1017);
or U2532 (N_2532,N_1963,N_1713);
nand U2533 (N_2533,N_1502,N_1344);
or U2534 (N_2534,N_1647,N_1665);
nor U2535 (N_2535,N_1889,N_1765);
nand U2536 (N_2536,N_1470,N_1191);
nor U2537 (N_2537,N_1119,N_1746);
and U2538 (N_2538,N_1808,N_1948);
nor U2539 (N_2539,N_1225,N_1032);
nand U2540 (N_2540,N_1625,N_1791);
nand U2541 (N_2541,N_1507,N_1996);
nor U2542 (N_2542,N_1167,N_1193);
and U2543 (N_2543,N_1501,N_1148);
xnor U2544 (N_2544,N_1010,N_1025);
and U2545 (N_2545,N_1971,N_1115);
nand U2546 (N_2546,N_1422,N_1086);
nor U2547 (N_2547,N_1211,N_1312);
nor U2548 (N_2548,N_1494,N_1138);
or U2549 (N_2549,N_1497,N_1079);
nor U2550 (N_2550,N_1010,N_1639);
and U2551 (N_2551,N_1181,N_1537);
nand U2552 (N_2552,N_1815,N_1262);
or U2553 (N_2553,N_1670,N_1642);
nand U2554 (N_2554,N_1066,N_1745);
nand U2555 (N_2555,N_1269,N_1904);
or U2556 (N_2556,N_1938,N_1047);
xnor U2557 (N_2557,N_1469,N_1499);
nand U2558 (N_2558,N_1201,N_1500);
nand U2559 (N_2559,N_1091,N_1049);
or U2560 (N_2560,N_1603,N_1218);
nor U2561 (N_2561,N_1616,N_1027);
nor U2562 (N_2562,N_1050,N_1015);
nor U2563 (N_2563,N_1112,N_1777);
or U2564 (N_2564,N_1545,N_1129);
nand U2565 (N_2565,N_1651,N_1444);
nor U2566 (N_2566,N_1554,N_1021);
or U2567 (N_2567,N_1712,N_1634);
nor U2568 (N_2568,N_1837,N_1195);
nor U2569 (N_2569,N_1932,N_1655);
or U2570 (N_2570,N_1681,N_1888);
and U2571 (N_2571,N_1571,N_1003);
and U2572 (N_2572,N_1495,N_1924);
nand U2573 (N_2573,N_1267,N_1633);
or U2574 (N_2574,N_1654,N_1297);
or U2575 (N_2575,N_1202,N_1427);
nor U2576 (N_2576,N_1058,N_1627);
nand U2577 (N_2577,N_1261,N_1702);
and U2578 (N_2578,N_1821,N_1842);
nand U2579 (N_2579,N_1948,N_1096);
and U2580 (N_2580,N_1298,N_1698);
and U2581 (N_2581,N_1730,N_1928);
and U2582 (N_2582,N_1330,N_1129);
nor U2583 (N_2583,N_1067,N_1135);
and U2584 (N_2584,N_1796,N_1686);
or U2585 (N_2585,N_1389,N_1969);
or U2586 (N_2586,N_1092,N_1416);
and U2587 (N_2587,N_1717,N_1704);
nor U2588 (N_2588,N_1617,N_1996);
nor U2589 (N_2589,N_1655,N_1306);
or U2590 (N_2590,N_1727,N_1650);
nor U2591 (N_2591,N_1739,N_1461);
or U2592 (N_2592,N_1792,N_1884);
nand U2593 (N_2593,N_1551,N_1786);
and U2594 (N_2594,N_1720,N_1223);
nand U2595 (N_2595,N_1045,N_1196);
xor U2596 (N_2596,N_1329,N_1404);
and U2597 (N_2597,N_1523,N_1897);
nand U2598 (N_2598,N_1704,N_1981);
xnor U2599 (N_2599,N_1701,N_1922);
and U2600 (N_2600,N_1668,N_1394);
nor U2601 (N_2601,N_1189,N_1400);
or U2602 (N_2602,N_1710,N_1580);
nor U2603 (N_2603,N_1477,N_1990);
and U2604 (N_2604,N_1495,N_1491);
and U2605 (N_2605,N_1292,N_1313);
nand U2606 (N_2606,N_1766,N_1216);
nor U2607 (N_2607,N_1283,N_1587);
nor U2608 (N_2608,N_1543,N_1163);
nor U2609 (N_2609,N_1008,N_1479);
nor U2610 (N_2610,N_1834,N_1065);
and U2611 (N_2611,N_1325,N_1428);
and U2612 (N_2612,N_1926,N_1949);
nor U2613 (N_2613,N_1083,N_1628);
and U2614 (N_2614,N_1705,N_1311);
xnor U2615 (N_2615,N_1888,N_1424);
and U2616 (N_2616,N_1408,N_1825);
nor U2617 (N_2617,N_1388,N_1714);
or U2618 (N_2618,N_1922,N_1290);
nand U2619 (N_2619,N_1148,N_1097);
and U2620 (N_2620,N_1161,N_1361);
and U2621 (N_2621,N_1813,N_1565);
nor U2622 (N_2622,N_1369,N_1926);
nand U2623 (N_2623,N_1399,N_1321);
and U2624 (N_2624,N_1538,N_1130);
nand U2625 (N_2625,N_1237,N_1123);
xnor U2626 (N_2626,N_1349,N_1254);
nor U2627 (N_2627,N_1959,N_1124);
nor U2628 (N_2628,N_1426,N_1067);
or U2629 (N_2629,N_1417,N_1046);
or U2630 (N_2630,N_1851,N_1907);
or U2631 (N_2631,N_1177,N_1294);
xnor U2632 (N_2632,N_1347,N_1817);
xor U2633 (N_2633,N_1650,N_1465);
or U2634 (N_2634,N_1591,N_1053);
nor U2635 (N_2635,N_1035,N_1729);
and U2636 (N_2636,N_1197,N_1520);
and U2637 (N_2637,N_1095,N_1311);
and U2638 (N_2638,N_1087,N_1285);
nand U2639 (N_2639,N_1186,N_1663);
or U2640 (N_2640,N_1054,N_1855);
and U2641 (N_2641,N_1208,N_1489);
or U2642 (N_2642,N_1346,N_1978);
nor U2643 (N_2643,N_1155,N_1099);
nor U2644 (N_2644,N_1745,N_1225);
nand U2645 (N_2645,N_1959,N_1726);
or U2646 (N_2646,N_1186,N_1281);
and U2647 (N_2647,N_1971,N_1021);
and U2648 (N_2648,N_1595,N_1774);
nor U2649 (N_2649,N_1837,N_1110);
nor U2650 (N_2650,N_1922,N_1062);
xnor U2651 (N_2651,N_1751,N_1762);
and U2652 (N_2652,N_1266,N_1625);
nor U2653 (N_2653,N_1269,N_1678);
nor U2654 (N_2654,N_1710,N_1977);
xnor U2655 (N_2655,N_1268,N_1375);
or U2656 (N_2656,N_1835,N_1840);
and U2657 (N_2657,N_1530,N_1609);
or U2658 (N_2658,N_1800,N_1982);
or U2659 (N_2659,N_1173,N_1996);
nand U2660 (N_2660,N_1263,N_1786);
or U2661 (N_2661,N_1091,N_1289);
nand U2662 (N_2662,N_1297,N_1187);
or U2663 (N_2663,N_1059,N_1954);
nand U2664 (N_2664,N_1056,N_1702);
nand U2665 (N_2665,N_1636,N_1147);
and U2666 (N_2666,N_1231,N_1056);
nor U2667 (N_2667,N_1284,N_1634);
xnor U2668 (N_2668,N_1388,N_1543);
nor U2669 (N_2669,N_1982,N_1124);
or U2670 (N_2670,N_1866,N_1194);
and U2671 (N_2671,N_1200,N_1579);
xnor U2672 (N_2672,N_1952,N_1336);
or U2673 (N_2673,N_1357,N_1926);
and U2674 (N_2674,N_1117,N_1681);
xor U2675 (N_2675,N_1918,N_1270);
nor U2676 (N_2676,N_1646,N_1293);
or U2677 (N_2677,N_1976,N_1954);
or U2678 (N_2678,N_1215,N_1565);
or U2679 (N_2679,N_1243,N_1441);
and U2680 (N_2680,N_1903,N_1532);
nor U2681 (N_2681,N_1055,N_1657);
nand U2682 (N_2682,N_1388,N_1351);
nand U2683 (N_2683,N_1970,N_1366);
or U2684 (N_2684,N_1425,N_1633);
or U2685 (N_2685,N_1692,N_1801);
and U2686 (N_2686,N_1517,N_1558);
nand U2687 (N_2687,N_1028,N_1804);
nor U2688 (N_2688,N_1955,N_1927);
or U2689 (N_2689,N_1219,N_1064);
nand U2690 (N_2690,N_1469,N_1825);
nand U2691 (N_2691,N_1293,N_1860);
or U2692 (N_2692,N_1579,N_1960);
or U2693 (N_2693,N_1775,N_1432);
nand U2694 (N_2694,N_1751,N_1694);
or U2695 (N_2695,N_1392,N_1692);
or U2696 (N_2696,N_1630,N_1097);
and U2697 (N_2697,N_1935,N_1766);
and U2698 (N_2698,N_1518,N_1049);
nand U2699 (N_2699,N_1202,N_1131);
and U2700 (N_2700,N_1797,N_1853);
or U2701 (N_2701,N_1678,N_1025);
or U2702 (N_2702,N_1297,N_1143);
and U2703 (N_2703,N_1381,N_1063);
and U2704 (N_2704,N_1467,N_1718);
or U2705 (N_2705,N_1255,N_1958);
nor U2706 (N_2706,N_1876,N_1700);
xor U2707 (N_2707,N_1964,N_1231);
nand U2708 (N_2708,N_1001,N_1152);
nand U2709 (N_2709,N_1108,N_1168);
nand U2710 (N_2710,N_1212,N_1590);
xor U2711 (N_2711,N_1819,N_1795);
and U2712 (N_2712,N_1014,N_1133);
and U2713 (N_2713,N_1094,N_1104);
and U2714 (N_2714,N_1661,N_1999);
nand U2715 (N_2715,N_1099,N_1734);
nand U2716 (N_2716,N_1732,N_1153);
nor U2717 (N_2717,N_1133,N_1413);
or U2718 (N_2718,N_1648,N_1194);
nor U2719 (N_2719,N_1024,N_1149);
or U2720 (N_2720,N_1313,N_1245);
nor U2721 (N_2721,N_1689,N_1782);
nand U2722 (N_2722,N_1142,N_1216);
nand U2723 (N_2723,N_1015,N_1729);
nor U2724 (N_2724,N_1847,N_1741);
nand U2725 (N_2725,N_1841,N_1237);
nand U2726 (N_2726,N_1167,N_1428);
or U2727 (N_2727,N_1143,N_1082);
or U2728 (N_2728,N_1246,N_1250);
nor U2729 (N_2729,N_1469,N_1404);
nand U2730 (N_2730,N_1260,N_1042);
nor U2731 (N_2731,N_1427,N_1670);
or U2732 (N_2732,N_1165,N_1776);
and U2733 (N_2733,N_1758,N_1398);
nand U2734 (N_2734,N_1468,N_1752);
nor U2735 (N_2735,N_1335,N_1083);
xnor U2736 (N_2736,N_1751,N_1265);
or U2737 (N_2737,N_1469,N_1896);
or U2738 (N_2738,N_1021,N_1318);
or U2739 (N_2739,N_1731,N_1384);
nand U2740 (N_2740,N_1818,N_1077);
or U2741 (N_2741,N_1630,N_1115);
or U2742 (N_2742,N_1143,N_1892);
xnor U2743 (N_2743,N_1715,N_1108);
and U2744 (N_2744,N_1357,N_1047);
and U2745 (N_2745,N_1103,N_1786);
nor U2746 (N_2746,N_1821,N_1477);
nor U2747 (N_2747,N_1007,N_1267);
nor U2748 (N_2748,N_1472,N_1684);
and U2749 (N_2749,N_1479,N_1775);
nor U2750 (N_2750,N_1593,N_1018);
or U2751 (N_2751,N_1100,N_1687);
nor U2752 (N_2752,N_1274,N_1832);
and U2753 (N_2753,N_1049,N_1559);
xor U2754 (N_2754,N_1840,N_1405);
nand U2755 (N_2755,N_1518,N_1019);
or U2756 (N_2756,N_1012,N_1720);
nor U2757 (N_2757,N_1802,N_1665);
xor U2758 (N_2758,N_1811,N_1541);
nand U2759 (N_2759,N_1548,N_1930);
or U2760 (N_2760,N_1506,N_1053);
or U2761 (N_2761,N_1988,N_1226);
nor U2762 (N_2762,N_1739,N_1658);
nor U2763 (N_2763,N_1613,N_1101);
and U2764 (N_2764,N_1685,N_1795);
nand U2765 (N_2765,N_1130,N_1146);
and U2766 (N_2766,N_1710,N_1940);
nor U2767 (N_2767,N_1184,N_1843);
or U2768 (N_2768,N_1839,N_1336);
nor U2769 (N_2769,N_1457,N_1995);
nand U2770 (N_2770,N_1979,N_1062);
nand U2771 (N_2771,N_1483,N_1329);
nand U2772 (N_2772,N_1403,N_1108);
nor U2773 (N_2773,N_1419,N_1824);
nor U2774 (N_2774,N_1610,N_1864);
nand U2775 (N_2775,N_1691,N_1579);
nor U2776 (N_2776,N_1231,N_1605);
nand U2777 (N_2777,N_1284,N_1389);
or U2778 (N_2778,N_1101,N_1482);
nor U2779 (N_2779,N_1797,N_1945);
nand U2780 (N_2780,N_1541,N_1638);
nand U2781 (N_2781,N_1186,N_1991);
and U2782 (N_2782,N_1199,N_1335);
and U2783 (N_2783,N_1930,N_1878);
and U2784 (N_2784,N_1642,N_1826);
or U2785 (N_2785,N_1768,N_1723);
xor U2786 (N_2786,N_1703,N_1626);
nor U2787 (N_2787,N_1483,N_1390);
nand U2788 (N_2788,N_1448,N_1203);
and U2789 (N_2789,N_1906,N_1466);
or U2790 (N_2790,N_1955,N_1531);
nor U2791 (N_2791,N_1787,N_1221);
and U2792 (N_2792,N_1533,N_1504);
nor U2793 (N_2793,N_1192,N_1489);
or U2794 (N_2794,N_1413,N_1938);
or U2795 (N_2795,N_1475,N_1380);
nand U2796 (N_2796,N_1030,N_1351);
nand U2797 (N_2797,N_1414,N_1157);
or U2798 (N_2798,N_1442,N_1860);
xnor U2799 (N_2799,N_1431,N_1278);
nor U2800 (N_2800,N_1755,N_1947);
or U2801 (N_2801,N_1375,N_1339);
or U2802 (N_2802,N_1293,N_1960);
and U2803 (N_2803,N_1721,N_1771);
or U2804 (N_2804,N_1270,N_1030);
or U2805 (N_2805,N_1794,N_1010);
xor U2806 (N_2806,N_1603,N_1804);
and U2807 (N_2807,N_1860,N_1081);
nand U2808 (N_2808,N_1706,N_1738);
and U2809 (N_2809,N_1500,N_1288);
or U2810 (N_2810,N_1942,N_1641);
and U2811 (N_2811,N_1647,N_1117);
nor U2812 (N_2812,N_1589,N_1283);
nor U2813 (N_2813,N_1010,N_1479);
nor U2814 (N_2814,N_1669,N_1741);
or U2815 (N_2815,N_1245,N_1052);
and U2816 (N_2816,N_1254,N_1821);
nor U2817 (N_2817,N_1429,N_1929);
or U2818 (N_2818,N_1349,N_1842);
nor U2819 (N_2819,N_1573,N_1763);
and U2820 (N_2820,N_1965,N_1991);
and U2821 (N_2821,N_1728,N_1265);
and U2822 (N_2822,N_1143,N_1202);
nor U2823 (N_2823,N_1024,N_1435);
and U2824 (N_2824,N_1108,N_1571);
nor U2825 (N_2825,N_1170,N_1669);
nor U2826 (N_2826,N_1433,N_1642);
nor U2827 (N_2827,N_1411,N_1306);
nand U2828 (N_2828,N_1773,N_1757);
or U2829 (N_2829,N_1384,N_1643);
nand U2830 (N_2830,N_1462,N_1514);
nand U2831 (N_2831,N_1783,N_1218);
xnor U2832 (N_2832,N_1248,N_1704);
xnor U2833 (N_2833,N_1993,N_1898);
and U2834 (N_2834,N_1480,N_1526);
and U2835 (N_2835,N_1999,N_1662);
or U2836 (N_2836,N_1720,N_1991);
xnor U2837 (N_2837,N_1589,N_1091);
nand U2838 (N_2838,N_1210,N_1479);
or U2839 (N_2839,N_1700,N_1118);
and U2840 (N_2840,N_1978,N_1047);
or U2841 (N_2841,N_1782,N_1207);
or U2842 (N_2842,N_1016,N_1507);
nor U2843 (N_2843,N_1711,N_1620);
nor U2844 (N_2844,N_1832,N_1735);
nand U2845 (N_2845,N_1205,N_1069);
and U2846 (N_2846,N_1692,N_1581);
nand U2847 (N_2847,N_1605,N_1155);
and U2848 (N_2848,N_1495,N_1724);
nand U2849 (N_2849,N_1603,N_1013);
or U2850 (N_2850,N_1397,N_1806);
nand U2851 (N_2851,N_1421,N_1935);
nand U2852 (N_2852,N_1633,N_1760);
and U2853 (N_2853,N_1710,N_1289);
or U2854 (N_2854,N_1116,N_1534);
nor U2855 (N_2855,N_1287,N_1226);
and U2856 (N_2856,N_1504,N_1742);
and U2857 (N_2857,N_1823,N_1046);
nand U2858 (N_2858,N_1889,N_1748);
nand U2859 (N_2859,N_1512,N_1174);
nand U2860 (N_2860,N_1406,N_1808);
or U2861 (N_2861,N_1531,N_1155);
nand U2862 (N_2862,N_1074,N_1911);
nor U2863 (N_2863,N_1430,N_1924);
or U2864 (N_2864,N_1411,N_1168);
xor U2865 (N_2865,N_1740,N_1608);
nand U2866 (N_2866,N_1083,N_1511);
and U2867 (N_2867,N_1986,N_1393);
and U2868 (N_2868,N_1027,N_1364);
nand U2869 (N_2869,N_1050,N_1536);
nand U2870 (N_2870,N_1875,N_1233);
or U2871 (N_2871,N_1643,N_1680);
and U2872 (N_2872,N_1701,N_1857);
nand U2873 (N_2873,N_1631,N_1227);
nor U2874 (N_2874,N_1426,N_1973);
nor U2875 (N_2875,N_1927,N_1894);
nor U2876 (N_2876,N_1419,N_1254);
or U2877 (N_2877,N_1745,N_1432);
or U2878 (N_2878,N_1573,N_1722);
nor U2879 (N_2879,N_1013,N_1949);
and U2880 (N_2880,N_1780,N_1259);
nor U2881 (N_2881,N_1105,N_1414);
or U2882 (N_2882,N_1998,N_1099);
nand U2883 (N_2883,N_1671,N_1818);
nor U2884 (N_2884,N_1797,N_1975);
nor U2885 (N_2885,N_1698,N_1425);
and U2886 (N_2886,N_1078,N_1229);
nand U2887 (N_2887,N_1947,N_1168);
or U2888 (N_2888,N_1233,N_1617);
nand U2889 (N_2889,N_1620,N_1092);
xor U2890 (N_2890,N_1190,N_1104);
and U2891 (N_2891,N_1479,N_1090);
nor U2892 (N_2892,N_1965,N_1966);
or U2893 (N_2893,N_1617,N_1352);
xnor U2894 (N_2894,N_1237,N_1593);
nor U2895 (N_2895,N_1494,N_1890);
nand U2896 (N_2896,N_1918,N_1822);
nand U2897 (N_2897,N_1362,N_1409);
nor U2898 (N_2898,N_1928,N_1639);
or U2899 (N_2899,N_1452,N_1394);
and U2900 (N_2900,N_1768,N_1380);
nor U2901 (N_2901,N_1766,N_1093);
nor U2902 (N_2902,N_1634,N_1219);
or U2903 (N_2903,N_1228,N_1357);
xor U2904 (N_2904,N_1698,N_1510);
nand U2905 (N_2905,N_1496,N_1230);
and U2906 (N_2906,N_1524,N_1073);
or U2907 (N_2907,N_1413,N_1325);
xor U2908 (N_2908,N_1299,N_1662);
nand U2909 (N_2909,N_1660,N_1128);
nor U2910 (N_2910,N_1660,N_1500);
nand U2911 (N_2911,N_1373,N_1472);
nand U2912 (N_2912,N_1122,N_1479);
nor U2913 (N_2913,N_1254,N_1290);
nor U2914 (N_2914,N_1616,N_1842);
nand U2915 (N_2915,N_1722,N_1189);
nand U2916 (N_2916,N_1393,N_1206);
nor U2917 (N_2917,N_1043,N_1440);
nor U2918 (N_2918,N_1222,N_1397);
nand U2919 (N_2919,N_1680,N_1644);
nand U2920 (N_2920,N_1974,N_1061);
nand U2921 (N_2921,N_1658,N_1577);
or U2922 (N_2922,N_1079,N_1637);
or U2923 (N_2923,N_1201,N_1642);
nand U2924 (N_2924,N_1454,N_1500);
nor U2925 (N_2925,N_1094,N_1764);
xnor U2926 (N_2926,N_1216,N_1911);
nor U2927 (N_2927,N_1832,N_1173);
and U2928 (N_2928,N_1948,N_1003);
nand U2929 (N_2929,N_1668,N_1030);
or U2930 (N_2930,N_1367,N_1447);
or U2931 (N_2931,N_1713,N_1591);
or U2932 (N_2932,N_1035,N_1272);
or U2933 (N_2933,N_1238,N_1898);
nand U2934 (N_2934,N_1831,N_1313);
nor U2935 (N_2935,N_1599,N_1351);
and U2936 (N_2936,N_1958,N_1140);
nor U2937 (N_2937,N_1925,N_1836);
xor U2938 (N_2938,N_1284,N_1450);
xnor U2939 (N_2939,N_1621,N_1231);
nand U2940 (N_2940,N_1446,N_1966);
or U2941 (N_2941,N_1920,N_1801);
or U2942 (N_2942,N_1005,N_1520);
nand U2943 (N_2943,N_1742,N_1481);
or U2944 (N_2944,N_1908,N_1104);
or U2945 (N_2945,N_1511,N_1913);
and U2946 (N_2946,N_1454,N_1078);
nand U2947 (N_2947,N_1377,N_1496);
nand U2948 (N_2948,N_1142,N_1215);
and U2949 (N_2949,N_1857,N_1889);
nor U2950 (N_2950,N_1947,N_1313);
nor U2951 (N_2951,N_1555,N_1531);
and U2952 (N_2952,N_1581,N_1679);
and U2953 (N_2953,N_1721,N_1749);
nor U2954 (N_2954,N_1812,N_1016);
or U2955 (N_2955,N_1469,N_1440);
and U2956 (N_2956,N_1253,N_1949);
nor U2957 (N_2957,N_1944,N_1046);
xor U2958 (N_2958,N_1200,N_1269);
or U2959 (N_2959,N_1689,N_1655);
nand U2960 (N_2960,N_1329,N_1185);
nand U2961 (N_2961,N_1915,N_1836);
or U2962 (N_2962,N_1321,N_1656);
xnor U2963 (N_2963,N_1242,N_1799);
nand U2964 (N_2964,N_1357,N_1709);
or U2965 (N_2965,N_1774,N_1281);
xnor U2966 (N_2966,N_1470,N_1986);
nand U2967 (N_2967,N_1647,N_1996);
or U2968 (N_2968,N_1952,N_1880);
or U2969 (N_2969,N_1191,N_1902);
or U2970 (N_2970,N_1617,N_1614);
nand U2971 (N_2971,N_1006,N_1013);
xnor U2972 (N_2972,N_1038,N_1182);
nor U2973 (N_2973,N_1457,N_1381);
nand U2974 (N_2974,N_1387,N_1101);
nand U2975 (N_2975,N_1070,N_1609);
nor U2976 (N_2976,N_1541,N_1830);
and U2977 (N_2977,N_1817,N_1219);
and U2978 (N_2978,N_1770,N_1964);
or U2979 (N_2979,N_1726,N_1499);
xnor U2980 (N_2980,N_1337,N_1069);
nand U2981 (N_2981,N_1288,N_1631);
nor U2982 (N_2982,N_1020,N_1172);
xnor U2983 (N_2983,N_1041,N_1366);
nor U2984 (N_2984,N_1541,N_1235);
or U2985 (N_2985,N_1464,N_1004);
nor U2986 (N_2986,N_1335,N_1490);
or U2987 (N_2987,N_1744,N_1325);
and U2988 (N_2988,N_1083,N_1718);
nand U2989 (N_2989,N_1978,N_1307);
nand U2990 (N_2990,N_1005,N_1000);
or U2991 (N_2991,N_1149,N_1113);
nand U2992 (N_2992,N_1322,N_1412);
xnor U2993 (N_2993,N_1805,N_1895);
or U2994 (N_2994,N_1397,N_1079);
or U2995 (N_2995,N_1387,N_1958);
xor U2996 (N_2996,N_1945,N_1284);
or U2997 (N_2997,N_1460,N_1941);
nand U2998 (N_2998,N_1105,N_1555);
nand U2999 (N_2999,N_1615,N_1283);
nor U3000 (N_3000,N_2022,N_2240);
nand U3001 (N_3001,N_2998,N_2598);
and U3002 (N_3002,N_2366,N_2800);
or U3003 (N_3003,N_2061,N_2378);
nor U3004 (N_3004,N_2138,N_2114);
or U3005 (N_3005,N_2658,N_2889);
nand U3006 (N_3006,N_2261,N_2445);
nand U3007 (N_3007,N_2473,N_2190);
or U3008 (N_3008,N_2915,N_2469);
or U3009 (N_3009,N_2568,N_2880);
nor U3010 (N_3010,N_2287,N_2657);
or U3011 (N_3011,N_2257,N_2596);
or U3012 (N_3012,N_2735,N_2095);
and U3013 (N_3013,N_2862,N_2235);
and U3014 (N_3014,N_2036,N_2802);
xnor U3015 (N_3015,N_2982,N_2638);
or U3016 (N_3016,N_2843,N_2818);
and U3017 (N_3017,N_2985,N_2957);
or U3018 (N_3018,N_2230,N_2444);
nand U3019 (N_3019,N_2952,N_2438);
and U3020 (N_3020,N_2056,N_2478);
xor U3021 (N_3021,N_2318,N_2447);
nand U3022 (N_3022,N_2728,N_2667);
or U3023 (N_3023,N_2365,N_2292);
nor U3024 (N_3024,N_2648,N_2085);
and U3025 (N_3025,N_2496,N_2009);
nor U3026 (N_3026,N_2961,N_2726);
nand U3027 (N_3027,N_2031,N_2514);
or U3028 (N_3028,N_2389,N_2908);
and U3029 (N_3029,N_2427,N_2500);
nand U3030 (N_3030,N_2168,N_2015);
nor U3031 (N_3031,N_2200,N_2238);
nand U3032 (N_3032,N_2197,N_2781);
or U3033 (N_3033,N_2105,N_2038);
nor U3034 (N_3034,N_2760,N_2334);
and U3035 (N_3035,N_2441,N_2739);
nand U3036 (N_3036,N_2079,N_2160);
and U3037 (N_3037,N_2356,N_2388);
nand U3038 (N_3038,N_2472,N_2703);
and U3039 (N_3039,N_2350,N_2124);
or U3040 (N_3040,N_2731,N_2923);
and U3041 (N_3041,N_2978,N_2316);
nor U3042 (N_3042,N_2440,N_2903);
or U3043 (N_3043,N_2089,N_2225);
nand U3044 (N_3044,N_2698,N_2680);
xor U3045 (N_3045,N_2593,N_2629);
or U3046 (N_3046,N_2819,N_2494);
and U3047 (N_3047,N_2814,N_2758);
nor U3048 (N_3048,N_2492,N_2100);
or U3049 (N_3049,N_2987,N_2590);
or U3050 (N_3050,N_2752,N_2834);
and U3051 (N_3051,N_2591,N_2154);
nor U3052 (N_3052,N_2142,N_2204);
nor U3053 (N_3053,N_2376,N_2176);
nand U3054 (N_3054,N_2361,N_2264);
and U3055 (N_3055,N_2610,N_2763);
nor U3056 (N_3056,N_2305,N_2931);
nor U3057 (N_3057,N_2359,N_2448);
or U3058 (N_3058,N_2443,N_2548);
nand U3059 (N_3059,N_2996,N_2258);
nand U3060 (N_3060,N_2169,N_2929);
nor U3061 (N_3061,N_2970,N_2701);
nand U3062 (N_3062,N_2161,N_2796);
and U3063 (N_3063,N_2520,N_2381);
nor U3064 (N_3064,N_2326,N_2363);
or U3065 (N_3065,N_2072,N_2665);
and U3066 (N_3066,N_2250,N_2824);
and U3067 (N_3067,N_2704,N_2139);
or U3068 (N_3068,N_2127,N_2642);
and U3069 (N_3069,N_2832,N_2362);
or U3070 (N_3070,N_2630,N_2575);
nor U3071 (N_3071,N_2508,N_2733);
and U3072 (N_3072,N_2829,N_2799);
and U3073 (N_3073,N_2001,N_2586);
nor U3074 (N_3074,N_2858,N_2717);
xnor U3075 (N_3075,N_2049,N_2259);
xor U3076 (N_3076,N_2963,N_2157);
and U3077 (N_3077,N_2347,N_2003);
xor U3078 (N_3078,N_2660,N_2120);
and U3079 (N_3079,N_2331,N_2067);
or U3080 (N_3080,N_2725,N_2954);
nor U3081 (N_3081,N_2689,N_2664);
nand U3082 (N_3082,N_2865,N_2827);
nor U3083 (N_3083,N_2984,N_2416);
nand U3084 (N_3084,N_2737,N_2408);
and U3085 (N_3085,N_2718,N_2368);
nand U3086 (N_3086,N_2644,N_2504);
nor U3087 (N_3087,N_2609,N_2918);
and U3088 (N_3088,N_2897,N_2219);
or U3089 (N_3089,N_2811,N_2246);
or U3090 (N_3090,N_2309,N_2652);
nor U3091 (N_3091,N_2470,N_2828);
nand U3092 (N_3092,N_2775,N_2750);
nand U3093 (N_3093,N_2171,N_2322);
nor U3094 (N_3094,N_2046,N_2086);
and U3095 (N_3095,N_2479,N_2551);
xnor U3096 (N_3096,N_2497,N_2097);
and U3097 (N_3097,N_2608,N_2450);
nor U3098 (N_3098,N_2765,N_2772);
nor U3099 (N_3099,N_2545,N_2274);
and U3100 (N_3100,N_2659,N_2851);
or U3101 (N_3101,N_2794,N_2021);
nor U3102 (N_3102,N_2439,N_2393);
nor U3103 (N_3103,N_2044,N_2084);
nand U3104 (N_3104,N_2353,N_2011);
xnor U3105 (N_3105,N_2375,N_2815);
nor U3106 (N_3106,N_2613,N_2354);
or U3107 (N_3107,N_2513,N_2301);
nand U3108 (N_3108,N_2921,N_2195);
nand U3109 (N_3109,N_2189,N_2339);
nor U3110 (N_3110,N_2569,N_2213);
and U3111 (N_3111,N_2065,N_2501);
and U3112 (N_3112,N_2747,N_2276);
and U3113 (N_3113,N_2993,N_2421);
or U3114 (N_3114,N_2340,N_2398);
nand U3115 (N_3115,N_2692,N_2966);
or U3116 (N_3116,N_2282,N_2349);
nor U3117 (N_3117,N_2749,N_2974);
nor U3118 (N_3118,N_2005,N_2143);
or U3119 (N_3119,N_2620,N_2959);
and U3120 (N_3120,N_2275,N_2938);
nor U3121 (N_3121,N_2288,N_2615);
xnor U3122 (N_3122,N_2911,N_2175);
and U3123 (N_3123,N_2646,N_2283);
nand U3124 (N_3124,N_2730,N_2502);
and U3125 (N_3125,N_2564,N_2116);
nor U3126 (N_3126,N_2101,N_2268);
nor U3127 (N_3127,N_2655,N_2767);
xor U3128 (N_3128,N_2806,N_2380);
nand U3129 (N_3129,N_2119,N_2023);
or U3130 (N_3130,N_2302,N_2635);
nor U3131 (N_3131,N_2994,N_2297);
and U3132 (N_3132,N_2228,N_2191);
nand U3133 (N_3133,N_2488,N_2988);
and U3134 (N_3134,N_2778,N_2820);
or U3135 (N_3135,N_2543,N_2188);
and U3136 (N_3136,N_2631,N_2449);
nor U3137 (N_3137,N_2248,N_2262);
nand U3138 (N_3138,N_2144,N_2239);
nand U3139 (N_3139,N_2847,N_2841);
nand U3140 (N_3140,N_2060,N_2577);
xor U3141 (N_3141,N_2226,N_2266);
nor U3142 (N_3142,N_2149,N_2404);
and U3143 (N_3143,N_2383,N_2163);
and U3144 (N_3144,N_2104,N_2294);
nand U3145 (N_3145,N_2173,N_2342);
or U3146 (N_3146,N_2184,N_2669);
or U3147 (N_3147,N_2306,N_2333);
nand U3148 (N_3148,N_2418,N_2357);
and U3149 (N_3149,N_2122,N_2420);
and U3150 (N_3150,N_2822,N_2976);
or U3151 (N_3151,N_2691,N_2556);
nor U3152 (N_3152,N_2958,N_2770);
and U3153 (N_3153,N_2177,N_2284);
nand U3154 (N_3154,N_2695,N_2083);
and U3155 (N_3155,N_2094,N_2587);
and U3156 (N_3156,N_2872,N_2483);
or U3157 (N_3157,N_2076,N_2267);
nand U3158 (N_3158,N_2845,N_2400);
and U3159 (N_3159,N_2583,N_2134);
nor U3160 (N_3160,N_2563,N_2905);
nor U3161 (N_3161,N_2341,N_2312);
nand U3162 (N_3162,N_2199,N_2111);
nor U3163 (N_3163,N_2410,N_2415);
nor U3164 (N_3164,N_2927,N_2227);
nor U3165 (N_3165,N_2837,N_2485);
nor U3166 (N_3166,N_2759,N_2973);
and U3167 (N_3167,N_2016,N_2979);
or U3168 (N_3168,N_2618,N_2888);
nand U3169 (N_3169,N_2201,N_2458);
nor U3170 (N_3170,N_2599,N_2899);
and U3171 (N_3171,N_2842,N_2627);
or U3172 (N_3172,N_2768,N_2956);
nor U3173 (N_3173,N_2152,N_2771);
and U3174 (N_3174,N_2930,N_2481);
nand U3175 (N_3175,N_2140,N_2935);
and U3176 (N_3176,N_2741,N_2917);
or U3177 (N_3177,N_2052,N_2928);
and U3178 (N_3178,N_2512,N_2178);
nand U3179 (N_3179,N_2051,N_2037);
nor U3180 (N_3180,N_2185,N_2162);
nand U3181 (N_3181,N_2992,N_2466);
or U3182 (N_3182,N_2130,N_2249);
and U3183 (N_3183,N_2937,N_2603);
nand U3184 (N_3184,N_2541,N_2311);
and U3185 (N_3185,N_2358,N_2537);
or U3186 (N_3186,N_2078,N_2417);
or U3187 (N_3187,N_2108,N_2990);
and U3188 (N_3188,N_2732,N_2172);
or U3189 (N_3189,N_2224,N_2476);
or U3190 (N_3190,N_2401,N_2547);
and U3191 (N_3191,N_2251,N_2237);
nand U3192 (N_3192,N_2636,N_2271);
xnor U3193 (N_3193,N_2619,N_2430);
and U3194 (N_3194,N_2645,N_2308);
and U3195 (N_3195,N_2696,N_2431);
nor U3196 (N_3196,N_2456,N_2403);
and U3197 (N_3197,N_2343,N_2286);
nand U3198 (N_3198,N_2017,N_2209);
nor U3199 (N_3199,N_2682,N_2714);
and U3200 (N_3200,N_2164,N_2407);
or U3201 (N_3201,N_2857,N_2746);
nor U3202 (N_3202,N_2040,N_2112);
or U3203 (N_3203,N_2572,N_2711);
nand U3204 (N_3204,N_2616,N_2907);
nand U3205 (N_3205,N_2662,N_2678);
nor U3206 (N_3206,N_2886,N_2700);
xor U3207 (N_3207,N_2774,N_2207);
and U3208 (N_3208,N_2482,N_2352);
nand U3209 (N_3209,N_2018,N_2327);
and U3210 (N_3210,N_2203,N_2675);
or U3211 (N_3211,N_2495,N_2882);
nand U3212 (N_3212,N_2121,N_2032);
and U3213 (N_3213,N_2584,N_2621);
or U3214 (N_3214,N_2805,N_2756);
nor U3215 (N_3215,N_2877,N_2158);
or U3216 (N_3216,N_2091,N_2372);
nand U3217 (N_3217,N_2394,N_2428);
and U3218 (N_3218,N_2791,N_2137);
or U3219 (N_3219,N_2883,N_2451);
or U3220 (N_3220,N_2891,N_2136);
nor U3221 (N_3221,N_2000,N_2853);
or U3222 (N_3222,N_2864,N_2058);
nor U3223 (N_3223,N_2565,N_2355);
nor U3224 (N_3224,N_2873,N_2523);
or U3225 (N_3225,N_2098,N_2133);
or U3226 (N_3226,N_2521,N_2594);
and U3227 (N_3227,N_2838,N_2159);
and U3228 (N_3228,N_2848,N_2382);
or U3229 (N_3229,N_2123,N_2869);
nand U3230 (N_3230,N_2740,N_2041);
nor U3231 (N_3231,N_2310,N_2919);
nand U3232 (N_3232,N_2345,N_2429);
nand U3233 (N_3233,N_2890,N_2221);
xor U3234 (N_3234,N_2167,N_2825);
and U3235 (N_3235,N_2859,N_2020);
nor U3236 (N_3236,N_2922,N_2007);
nor U3237 (N_3237,N_2462,N_2314);
nand U3238 (N_3238,N_2307,N_2464);
nor U3239 (N_3239,N_2411,N_2379);
nand U3240 (N_3240,N_2526,N_2792);
xnor U3241 (N_3241,N_2045,N_2953);
xnor U3242 (N_3242,N_2220,N_2006);
xnor U3243 (N_3243,N_2839,N_2503);
or U3244 (N_3244,N_2141,N_2600);
nand U3245 (N_3245,N_2894,N_2955);
or U3246 (N_3246,N_2384,N_2087);
and U3247 (N_3247,N_2742,N_2773);
nor U3248 (N_3248,N_2835,N_2868);
nor U3249 (N_3249,N_2107,N_2975);
nor U3250 (N_3250,N_2117,N_2332);
nor U3251 (N_3251,N_2474,N_2968);
nor U3252 (N_3252,N_2335,N_2622);
nand U3253 (N_3253,N_2181,N_2743);
xor U3254 (N_3254,N_2509,N_2280);
nor U3255 (N_3255,N_2135,N_2515);
and U3256 (N_3256,N_2278,N_2281);
nand U3257 (N_3257,N_2304,N_2673);
nand U3258 (N_3258,N_2480,N_2454);
nor U3259 (N_3259,N_2807,N_2723);
and U3260 (N_3260,N_2785,N_2212);
nand U3261 (N_3261,N_2786,N_2313);
and U3262 (N_3262,N_2683,N_2578);
and U3263 (N_3263,N_2180,N_2777);
nor U3264 (N_3264,N_2560,N_2183);
and U3265 (N_3265,N_2528,N_2153);
xnor U3266 (N_3266,N_2933,N_2193);
xor U3267 (N_3267,N_2272,N_2831);
nor U3268 (N_3268,N_2323,N_2298);
xor U3269 (N_3269,N_2677,N_2782);
or U3270 (N_3270,N_2518,N_2099);
and U3271 (N_3271,N_2024,N_2113);
or U3272 (N_3272,N_2950,N_2236);
xor U3273 (N_3273,N_2672,N_2406);
and U3274 (N_3274,N_2385,N_2944);
nand U3275 (N_3275,N_2885,N_2849);
nor U3276 (N_3276,N_2914,N_2187);
and U3277 (N_3277,N_2423,N_2075);
xnor U3278 (N_3278,N_2793,N_2446);
nor U3279 (N_3279,N_2370,N_2716);
nor U3280 (N_3280,N_2054,N_2971);
and U3281 (N_3281,N_2866,N_2002);
nand U3282 (N_3282,N_2255,N_2924);
nand U3283 (N_3283,N_2486,N_2433);
or U3284 (N_3284,N_2592,N_2198);
and U3285 (N_3285,N_2895,N_2290);
nor U3286 (N_3286,N_2442,N_2604);
and U3287 (N_3287,N_2625,N_2260);
nand U3288 (N_3288,N_2748,N_2337);
nand U3289 (N_3289,N_2132,N_2395);
nor U3290 (N_3290,N_2096,N_2724);
nor U3291 (N_3291,N_2090,N_2540);
and U3292 (N_3292,N_2906,N_2901);
nor U3293 (N_3293,N_2374,N_2269);
or U3294 (N_3294,N_2150,N_2055);
and U3295 (N_3295,N_2289,N_2852);
nor U3296 (N_3296,N_2721,N_2795);
and U3297 (N_3297,N_2809,N_2720);
and U3298 (N_3298,N_2939,N_2524);
nor U3299 (N_3299,N_2863,N_2606);
or U3300 (N_3300,N_2202,N_2436);
nor U3301 (N_3301,N_2319,N_2684);
or U3302 (N_3302,N_2064,N_2926);
nand U3303 (N_3303,N_2229,N_2707);
and U3304 (N_3304,N_2761,N_2387);
nor U3305 (N_3305,N_2110,N_2241);
and U3306 (N_3306,N_2457,N_2535);
xor U3307 (N_3307,N_2424,N_2463);
or U3308 (N_3308,N_2364,N_2798);
and U3309 (N_3309,N_2062,N_2783);
and U3310 (N_3310,N_2900,N_2641);
nor U3311 (N_3311,N_2639,N_2223);
nand U3312 (N_3312,N_2030,N_2790);
nor U3313 (N_3313,N_2234,N_2147);
nor U3314 (N_3314,N_2296,N_2115);
xor U3315 (N_3315,N_2686,N_2208);
or U3316 (N_3316,N_2059,N_2371);
nand U3317 (N_3317,N_2557,N_2554);
or U3318 (N_3318,N_2581,N_2538);
nor U3319 (N_3319,N_2103,N_2881);
or U3320 (N_3320,N_2624,N_2705);
and U3321 (N_3321,N_2053,N_2047);
nor U3322 (N_3322,N_2048,N_2391);
or U3323 (N_3323,N_2126,N_2634);
and U3324 (N_3324,N_2027,N_2817);
nor U3325 (N_3325,N_2567,N_2043);
and U3326 (N_3326,N_2833,N_2887);
or U3327 (N_3327,N_2329,N_2517);
or U3328 (N_3328,N_2855,N_2344);
nand U3329 (N_3329,N_2546,N_2348);
or U3330 (N_3330,N_2702,N_2788);
nor U3331 (N_3331,N_2602,N_2012);
nand U3332 (N_3332,N_2605,N_2836);
nand U3333 (N_3333,N_2066,N_2654);
and U3334 (N_3334,N_2293,N_2109);
nor U3335 (N_3335,N_2623,N_2025);
and U3336 (N_3336,N_2505,N_2812);
nor U3337 (N_3337,N_2409,N_2650);
and U3338 (N_3338,N_2668,N_2934);
nand U3339 (N_3339,N_2081,N_2803);
nand U3340 (N_3340,N_2490,N_2779);
or U3341 (N_3341,N_2688,N_2576);
and U3342 (N_3342,N_2516,N_2070);
xnor U3343 (N_3343,N_2338,N_2008);
nand U3344 (N_3344,N_2697,N_2151);
nand U3345 (N_3345,N_2367,N_2166);
nand U3346 (N_3346,N_2561,N_2532);
xnor U3347 (N_3347,N_2870,N_2425);
or U3348 (N_3348,N_2910,N_2247);
xnor U3349 (N_3349,N_2713,N_2965);
and U3350 (N_3350,N_2039,N_2875);
and U3351 (N_3351,N_2597,N_2754);
nand U3352 (N_3352,N_2983,N_2148);
nand U3353 (N_3353,N_2542,N_2493);
nand U3354 (N_3354,N_2414,N_2690);
nor U3355 (N_3355,N_2093,N_2816);
nor U3356 (N_3356,N_2484,N_2265);
xnor U3357 (N_3357,N_2980,N_2253);
nor U3358 (N_3358,N_2320,N_2670);
nor U3359 (N_3359,N_2653,N_2218);
nor U3360 (N_3360,N_2736,N_2527);
nand U3361 (N_3361,N_2981,N_2874);
nor U3362 (N_3362,N_2751,N_2467);
and U3363 (N_3363,N_2242,N_2489);
xor U3364 (N_3364,N_2912,N_2589);
and U3365 (N_3365,N_2533,N_2215);
nand U3366 (N_3366,N_2898,N_2582);
nand U3367 (N_3367,N_2263,N_2324);
nor U3368 (N_3368,N_2035,N_2434);
and U3369 (N_3369,N_2744,N_2346);
nor U3370 (N_3370,N_2534,N_2951);
xor U3371 (N_3371,N_2997,N_2155);
nand U3372 (N_3372,N_2491,N_2932);
or U3373 (N_3373,N_2536,N_2455);
nand U3374 (N_3374,N_2315,N_2475);
nor U3375 (N_3375,N_2063,N_2402);
nor U3376 (N_3376,N_2813,N_2468);
nor U3377 (N_3377,N_2823,N_2131);
or U3378 (N_3378,N_2727,N_2205);
nand U3379 (N_3379,N_2571,N_2465);
and U3380 (N_3380,N_2562,N_2471);
nand U3381 (N_3381,N_2633,N_2073);
nor U3382 (N_3382,N_2102,N_2077);
nor U3383 (N_3383,N_2632,N_2369);
nand U3384 (N_3384,N_2902,N_2511);
or U3385 (N_3385,N_2867,N_2506);
or U3386 (N_3386,N_2570,N_2373);
nand U3387 (N_3387,N_2579,N_2734);
nor U3388 (N_3388,N_2245,N_2614);
xnor U3389 (N_3389,N_2846,N_2129);
and U3390 (N_3390,N_2214,N_2753);
xor U3391 (N_3391,N_2766,N_2967);
nor U3392 (N_3392,N_2580,N_2745);
or U3393 (N_3393,N_2757,N_2738);
and U3394 (N_3394,N_2679,N_2461);
and U3395 (N_3395,N_2422,N_2936);
xor U3396 (N_3396,N_2676,N_2940);
nand U3397 (N_3397,N_2328,N_2611);
nor U3398 (N_3398,N_2871,N_2913);
nor U3399 (N_3399,N_2004,N_2671);
or U3400 (N_3400,N_2270,N_2057);
and U3401 (N_3401,N_2661,N_2397);
nand U3402 (N_3402,N_2128,N_2507);
nand U3403 (N_3403,N_2946,N_2019);
nor U3404 (N_3404,N_2244,N_2206);
nor U3405 (N_3405,N_2273,N_2941);
or U3406 (N_3406,N_2170,N_2068);
or U3407 (N_3407,N_2013,N_2896);
nor U3408 (N_3408,N_2459,N_2573);
and U3409 (N_3409,N_2186,N_2092);
xnor U3410 (N_3410,N_2074,N_2558);
xor U3411 (N_3411,N_2709,N_2909);
or U3412 (N_3412,N_2377,N_2844);
and U3413 (N_3413,N_2291,N_2519);
and U3414 (N_3414,N_2192,N_2687);
and U3415 (N_3415,N_2972,N_2830);
nand U3416 (N_3416,N_2964,N_2336);
and U3417 (N_3417,N_2962,N_2681);
and U3418 (N_3418,N_2719,N_2574);
and U3419 (N_3419,N_2317,N_2106);
nor U3420 (N_3420,N_2810,N_2588);
nor U3421 (N_3421,N_2525,N_2499);
or U3422 (N_3422,N_2071,N_2712);
and U3423 (N_3423,N_2626,N_2165);
nor U3424 (N_3424,N_2196,N_2028);
and U3425 (N_3425,N_2330,N_2999);
xnor U3426 (N_3426,N_2784,N_2549);
nand U3427 (N_3427,N_2850,N_2252);
nand U3428 (N_3428,N_2014,N_2413);
or U3429 (N_3429,N_2892,N_2453);
and U3430 (N_3430,N_2390,N_2295);
nand U3431 (N_3431,N_2948,N_2656);
and U3432 (N_3432,N_2797,N_2585);
nand U3433 (N_3433,N_2729,N_2437);
nand U3434 (N_3434,N_2925,N_2601);
xor U3435 (N_3435,N_2351,N_2995);
nor U3436 (N_3436,N_2647,N_2945);
nand U3437 (N_3437,N_2042,N_2145);
nand U3438 (N_3438,N_2531,N_2801);
nor U3439 (N_3439,N_2211,N_2780);
nand U3440 (N_3440,N_2498,N_2663);
nor U3441 (N_3441,N_2082,N_2510);
nor U3442 (N_3442,N_2256,N_2989);
nor U3443 (N_3443,N_2426,N_2555);
or U3444 (N_3444,N_2452,N_2435);
nor U3445 (N_3445,N_2460,N_2789);
xnor U3446 (N_3446,N_2685,N_2231);
or U3447 (N_3447,N_2916,N_2217);
nor U3448 (N_3448,N_2530,N_2386);
nand U3449 (N_3449,N_2708,N_2860);
nand U3450 (N_3450,N_2787,N_2861);
or U3451 (N_3451,N_2666,N_2764);
nor U3452 (N_3452,N_2949,N_2854);
or U3453 (N_3453,N_2088,N_2826);
or U3454 (N_3454,N_2325,N_2986);
xor U3455 (N_3455,N_2182,N_2285);
and U3456 (N_3456,N_2303,N_2392);
or U3457 (N_3457,N_2710,N_2960);
or U3458 (N_3458,N_2477,N_2222);
or U3459 (N_3459,N_2808,N_2878);
and U3460 (N_3460,N_2080,N_2405);
nand U3461 (N_3461,N_2879,N_2769);
nor U3462 (N_3462,N_2884,N_2550);
or U3463 (N_3463,N_2706,N_2755);
or U3464 (N_3464,N_2321,N_2034);
nor U3465 (N_3465,N_2607,N_2942);
nor U3466 (N_3466,N_2553,N_2432);
or U3467 (N_3467,N_2920,N_2254);
nand U3468 (N_3468,N_2522,N_2300);
nor U3469 (N_3469,N_2694,N_2194);
nor U3470 (N_3470,N_2243,N_2396);
and U3471 (N_3471,N_2893,N_2156);
xnor U3472 (N_3472,N_2821,N_2699);
nand U3473 (N_3473,N_2210,N_2010);
nand U3474 (N_3474,N_2232,N_2529);
and U3475 (N_3475,N_2146,N_2412);
nor U3476 (N_3476,N_2559,N_2637);
nand U3477 (N_3477,N_2943,N_2643);
and U3478 (N_3478,N_2840,N_2674);
and U3479 (N_3479,N_2299,N_2279);
nor U3480 (N_3480,N_2566,N_2539);
and U3481 (N_3481,N_2544,N_2233);
or U3482 (N_3482,N_2617,N_2649);
and U3483 (N_3483,N_2174,N_2029);
and U3484 (N_3484,N_2033,N_2947);
and U3485 (N_3485,N_2762,N_2651);
xnor U3486 (N_3486,N_2977,N_2715);
nor U3487 (N_3487,N_2118,N_2904);
or U3488 (N_3488,N_2360,N_2876);
or U3489 (N_3489,N_2069,N_2487);
and U3490 (N_3490,N_2419,N_2179);
nand U3491 (N_3491,N_2277,N_2856);
and U3492 (N_3492,N_2050,N_2612);
and U3493 (N_3493,N_2595,N_2026);
xnor U3494 (N_3494,N_2722,N_2969);
nor U3495 (N_3495,N_2125,N_2628);
nand U3496 (N_3496,N_2552,N_2693);
and U3497 (N_3497,N_2804,N_2640);
nand U3498 (N_3498,N_2776,N_2216);
nor U3499 (N_3499,N_2991,N_2399);
or U3500 (N_3500,N_2753,N_2903);
nor U3501 (N_3501,N_2685,N_2472);
or U3502 (N_3502,N_2655,N_2913);
nand U3503 (N_3503,N_2887,N_2841);
nor U3504 (N_3504,N_2888,N_2811);
nor U3505 (N_3505,N_2925,N_2281);
xor U3506 (N_3506,N_2421,N_2377);
and U3507 (N_3507,N_2418,N_2554);
or U3508 (N_3508,N_2598,N_2450);
or U3509 (N_3509,N_2998,N_2892);
or U3510 (N_3510,N_2431,N_2566);
or U3511 (N_3511,N_2706,N_2796);
and U3512 (N_3512,N_2110,N_2202);
and U3513 (N_3513,N_2725,N_2814);
nor U3514 (N_3514,N_2304,N_2808);
nand U3515 (N_3515,N_2540,N_2534);
xnor U3516 (N_3516,N_2342,N_2821);
or U3517 (N_3517,N_2560,N_2124);
or U3518 (N_3518,N_2855,N_2890);
nor U3519 (N_3519,N_2304,N_2423);
nor U3520 (N_3520,N_2139,N_2293);
or U3521 (N_3521,N_2150,N_2074);
nand U3522 (N_3522,N_2886,N_2122);
or U3523 (N_3523,N_2868,N_2877);
or U3524 (N_3524,N_2938,N_2583);
nor U3525 (N_3525,N_2451,N_2849);
nand U3526 (N_3526,N_2023,N_2324);
nor U3527 (N_3527,N_2559,N_2536);
nand U3528 (N_3528,N_2314,N_2637);
or U3529 (N_3529,N_2143,N_2503);
nor U3530 (N_3530,N_2495,N_2922);
or U3531 (N_3531,N_2305,N_2191);
nand U3532 (N_3532,N_2531,N_2656);
and U3533 (N_3533,N_2880,N_2879);
nor U3534 (N_3534,N_2458,N_2749);
or U3535 (N_3535,N_2494,N_2846);
and U3536 (N_3536,N_2768,N_2054);
or U3537 (N_3537,N_2934,N_2113);
nor U3538 (N_3538,N_2413,N_2736);
nand U3539 (N_3539,N_2758,N_2318);
nand U3540 (N_3540,N_2194,N_2920);
and U3541 (N_3541,N_2310,N_2586);
nand U3542 (N_3542,N_2089,N_2298);
nor U3543 (N_3543,N_2398,N_2763);
and U3544 (N_3544,N_2979,N_2875);
nand U3545 (N_3545,N_2004,N_2527);
or U3546 (N_3546,N_2245,N_2158);
or U3547 (N_3547,N_2044,N_2123);
nand U3548 (N_3548,N_2490,N_2247);
nand U3549 (N_3549,N_2109,N_2095);
or U3550 (N_3550,N_2865,N_2690);
nand U3551 (N_3551,N_2124,N_2450);
or U3552 (N_3552,N_2261,N_2474);
nand U3553 (N_3553,N_2918,N_2626);
and U3554 (N_3554,N_2075,N_2487);
nand U3555 (N_3555,N_2223,N_2389);
nand U3556 (N_3556,N_2981,N_2797);
nand U3557 (N_3557,N_2885,N_2829);
nor U3558 (N_3558,N_2377,N_2758);
and U3559 (N_3559,N_2928,N_2340);
nor U3560 (N_3560,N_2580,N_2266);
nand U3561 (N_3561,N_2926,N_2360);
and U3562 (N_3562,N_2093,N_2488);
nor U3563 (N_3563,N_2830,N_2381);
nor U3564 (N_3564,N_2596,N_2728);
nand U3565 (N_3565,N_2967,N_2566);
and U3566 (N_3566,N_2732,N_2502);
nor U3567 (N_3567,N_2880,N_2652);
and U3568 (N_3568,N_2341,N_2524);
or U3569 (N_3569,N_2870,N_2400);
nor U3570 (N_3570,N_2335,N_2680);
nor U3571 (N_3571,N_2043,N_2785);
xnor U3572 (N_3572,N_2107,N_2816);
nor U3573 (N_3573,N_2900,N_2466);
or U3574 (N_3574,N_2788,N_2154);
xnor U3575 (N_3575,N_2242,N_2171);
and U3576 (N_3576,N_2112,N_2099);
and U3577 (N_3577,N_2515,N_2107);
nor U3578 (N_3578,N_2844,N_2938);
xnor U3579 (N_3579,N_2073,N_2707);
nand U3580 (N_3580,N_2688,N_2855);
or U3581 (N_3581,N_2790,N_2624);
nand U3582 (N_3582,N_2517,N_2797);
nor U3583 (N_3583,N_2701,N_2543);
xnor U3584 (N_3584,N_2916,N_2168);
or U3585 (N_3585,N_2991,N_2555);
or U3586 (N_3586,N_2051,N_2280);
or U3587 (N_3587,N_2016,N_2044);
nor U3588 (N_3588,N_2351,N_2693);
and U3589 (N_3589,N_2333,N_2548);
and U3590 (N_3590,N_2428,N_2373);
nor U3591 (N_3591,N_2056,N_2324);
nand U3592 (N_3592,N_2010,N_2381);
or U3593 (N_3593,N_2471,N_2552);
nor U3594 (N_3594,N_2122,N_2742);
or U3595 (N_3595,N_2408,N_2237);
and U3596 (N_3596,N_2482,N_2049);
nand U3597 (N_3597,N_2424,N_2184);
nor U3598 (N_3598,N_2282,N_2309);
nor U3599 (N_3599,N_2211,N_2744);
nor U3600 (N_3600,N_2848,N_2154);
nand U3601 (N_3601,N_2705,N_2044);
nor U3602 (N_3602,N_2856,N_2330);
nor U3603 (N_3603,N_2301,N_2847);
nand U3604 (N_3604,N_2894,N_2876);
or U3605 (N_3605,N_2209,N_2743);
and U3606 (N_3606,N_2356,N_2445);
and U3607 (N_3607,N_2608,N_2684);
nand U3608 (N_3608,N_2219,N_2242);
nor U3609 (N_3609,N_2083,N_2779);
nand U3610 (N_3610,N_2074,N_2184);
nand U3611 (N_3611,N_2489,N_2996);
xnor U3612 (N_3612,N_2478,N_2250);
xor U3613 (N_3613,N_2150,N_2488);
nand U3614 (N_3614,N_2218,N_2687);
or U3615 (N_3615,N_2098,N_2677);
nor U3616 (N_3616,N_2847,N_2051);
or U3617 (N_3617,N_2060,N_2910);
or U3618 (N_3618,N_2280,N_2681);
xor U3619 (N_3619,N_2111,N_2913);
and U3620 (N_3620,N_2261,N_2829);
or U3621 (N_3621,N_2815,N_2574);
and U3622 (N_3622,N_2333,N_2012);
and U3623 (N_3623,N_2213,N_2129);
xnor U3624 (N_3624,N_2423,N_2251);
nor U3625 (N_3625,N_2537,N_2962);
nand U3626 (N_3626,N_2090,N_2382);
and U3627 (N_3627,N_2460,N_2857);
nor U3628 (N_3628,N_2670,N_2732);
and U3629 (N_3629,N_2133,N_2396);
or U3630 (N_3630,N_2508,N_2239);
xnor U3631 (N_3631,N_2791,N_2776);
nand U3632 (N_3632,N_2557,N_2365);
nor U3633 (N_3633,N_2815,N_2343);
nor U3634 (N_3634,N_2066,N_2521);
xnor U3635 (N_3635,N_2310,N_2315);
nand U3636 (N_3636,N_2073,N_2691);
or U3637 (N_3637,N_2269,N_2023);
nor U3638 (N_3638,N_2559,N_2474);
or U3639 (N_3639,N_2232,N_2772);
xor U3640 (N_3640,N_2117,N_2972);
nand U3641 (N_3641,N_2912,N_2054);
and U3642 (N_3642,N_2283,N_2351);
or U3643 (N_3643,N_2402,N_2650);
nand U3644 (N_3644,N_2522,N_2572);
nand U3645 (N_3645,N_2751,N_2098);
nor U3646 (N_3646,N_2661,N_2777);
xor U3647 (N_3647,N_2237,N_2808);
and U3648 (N_3648,N_2014,N_2743);
nor U3649 (N_3649,N_2313,N_2082);
nor U3650 (N_3650,N_2193,N_2230);
nand U3651 (N_3651,N_2023,N_2283);
and U3652 (N_3652,N_2527,N_2896);
and U3653 (N_3653,N_2405,N_2412);
or U3654 (N_3654,N_2360,N_2628);
or U3655 (N_3655,N_2683,N_2321);
or U3656 (N_3656,N_2965,N_2223);
nand U3657 (N_3657,N_2622,N_2177);
nor U3658 (N_3658,N_2318,N_2949);
or U3659 (N_3659,N_2123,N_2776);
nand U3660 (N_3660,N_2801,N_2399);
or U3661 (N_3661,N_2848,N_2681);
nor U3662 (N_3662,N_2048,N_2359);
or U3663 (N_3663,N_2326,N_2086);
and U3664 (N_3664,N_2067,N_2236);
and U3665 (N_3665,N_2478,N_2100);
or U3666 (N_3666,N_2801,N_2540);
nand U3667 (N_3667,N_2877,N_2049);
and U3668 (N_3668,N_2796,N_2986);
nand U3669 (N_3669,N_2697,N_2054);
or U3670 (N_3670,N_2345,N_2452);
or U3671 (N_3671,N_2934,N_2268);
nand U3672 (N_3672,N_2605,N_2825);
and U3673 (N_3673,N_2823,N_2815);
nand U3674 (N_3674,N_2000,N_2087);
and U3675 (N_3675,N_2704,N_2234);
xnor U3676 (N_3676,N_2562,N_2570);
and U3677 (N_3677,N_2165,N_2658);
nor U3678 (N_3678,N_2799,N_2636);
nor U3679 (N_3679,N_2309,N_2754);
nand U3680 (N_3680,N_2609,N_2674);
and U3681 (N_3681,N_2364,N_2488);
or U3682 (N_3682,N_2088,N_2261);
and U3683 (N_3683,N_2503,N_2119);
nand U3684 (N_3684,N_2397,N_2450);
or U3685 (N_3685,N_2230,N_2955);
and U3686 (N_3686,N_2374,N_2424);
and U3687 (N_3687,N_2318,N_2225);
nand U3688 (N_3688,N_2433,N_2298);
or U3689 (N_3689,N_2168,N_2836);
or U3690 (N_3690,N_2388,N_2733);
xor U3691 (N_3691,N_2740,N_2602);
xnor U3692 (N_3692,N_2639,N_2009);
xnor U3693 (N_3693,N_2428,N_2408);
xor U3694 (N_3694,N_2223,N_2586);
or U3695 (N_3695,N_2699,N_2883);
or U3696 (N_3696,N_2397,N_2144);
and U3697 (N_3697,N_2938,N_2431);
and U3698 (N_3698,N_2797,N_2779);
nor U3699 (N_3699,N_2588,N_2181);
and U3700 (N_3700,N_2023,N_2338);
xor U3701 (N_3701,N_2838,N_2901);
nand U3702 (N_3702,N_2844,N_2417);
nor U3703 (N_3703,N_2475,N_2564);
and U3704 (N_3704,N_2230,N_2214);
or U3705 (N_3705,N_2940,N_2061);
and U3706 (N_3706,N_2372,N_2649);
or U3707 (N_3707,N_2981,N_2452);
or U3708 (N_3708,N_2346,N_2482);
or U3709 (N_3709,N_2029,N_2072);
nand U3710 (N_3710,N_2292,N_2504);
and U3711 (N_3711,N_2425,N_2937);
nand U3712 (N_3712,N_2982,N_2351);
nand U3713 (N_3713,N_2249,N_2598);
and U3714 (N_3714,N_2658,N_2661);
xor U3715 (N_3715,N_2828,N_2643);
nand U3716 (N_3716,N_2115,N_2262);
nor U3717 (N_3717,N_2087,N_2690);
xnor U3718 (N_3718,N_2277,N_2479);
nand U3719 (N_3719,N_2831,N_2922);
nand U3720 (N_3720,N_2167,N_2750);
nor U3721 (N_3721,N_2818,N_2796);
and U3722 (N_3722,N_2290,N_2907);
nand U3723 (N_3723,N_2160,N_2337);
or U3724 (N_3724,N_2105,N_2448);
xor U3725 (N_3725,N_2056,N_2885);
and U3726 (N_3726,N_2843,N_2994);
nand U3727 (N_3727,N_2724,N_2984);
nor U3728 (N_3728,N_2236,N_2506);
and U3729 (N_3729,N_2439,N_2406);
nor U3730 (N_3730,N_2707,N_2996);
nor U3731 (N_3731,N_2483,N_2704);
or U3732 (N_3732,N_2837,N_2855);
and U3733 (N_3733,N_2696,N_2082);
xnor U3734 (N_3734,N_2376,N_2478);
nor U3735 (N_3735,N_2096,N_2551);
nand U3736 (N_3736,N_2611,N_2537);
and U3737 (N_3737,N_2723,N_2442);
nor U3738 (N_3738,N_2916,N_2411);
xnor U3739 (N_3739,N_2923,N_2445);
nor U3740 (N_3740,N_2705,N_2538);
nor U3741 (N_3741,N_2729,N_2409);
or U3742 (N_3742,N_2683,N_2537);
nand U3743 (N_3743,N_2651,N_2600);
and U3744 (N_3744,N_2880,N_2475);
and U3745 (N_3745,N_2361,N_2788);
and U3746 (N_3746,N_2019,N_2822);
nand U3747 (N_3747,N_2735,N_2041);
nand U3748 (N_3748,N_2372,N_2743);
and U3749 (N_3749,N_2152,N_2871);
nand U3750 (N_3750,N_2448,N_2741);
or U3751 (N_3751,N_2335,N_2655);
or U3752 (N_3752,N_2910,N_2828);
nand U3753 (N_3753,N_2112,N_2328);
nand U3754 (N_3754,N_2250,N_2949);
and U3755 (N_3755,N_2450,N_2862);
and U3756 (N_3756,N_2417,N_2959);
nor U3757 (N_3757,N_2698,N_2852);
or U3758 (N_3758,N_2822,N_2425);
nand U3759 (N_3759,N_2644,N_2860);
nand U3760 (N_3760,N_2148,N_2894);
nor U3761 (N_3761,N_2185,N_2020);
nor U3762 (N_3762,N_2710,N_2566);
or U3763 (N_3763,N_2518,N_2484);
or U3764 (N_3764,N_2225,N_2907);
nand U3765 (N_3765,N_2453,N_2458);
and U3766 (N_3766,N_2756,N_2892);
nor U3767 (N_3767,N_2027,N_2371);
and U3768 (N_3768,N_2845,N_2638);
nor U3769 (N_3769,N_2098,N_2207);
xor U3770 (N_3770,N_2134,N_2400);
nand U3771 (N_3771,N_2930,N_2051);
nor U3772 (N_3772,N_2284,N_2403);
nor U3773 (N_3773,N_2398,N_2599);
nor U3774 (N_3774,N_2184,N_2443);
and U3775 (N_3775,N_2216,N_2038);
nor U3776 (N_3776,N_2533,N_2976);
and U3777 (N_3777,N_2982,N_2251);
nor U3778 (N_3778,N_2981,N_2673);
nor U3779 (N_3779,N_2432,N_2793);
and U3780 (N_3780,N_2832,N_2436);
and U3781 (N_3781,N_2863,N_2936);
nand U3782 (N_3782,N_2637,N_2931);
or U3783 (N_3783,N_2941,N_2623);
nor U3784 (N_3784,N_2464,N_2171);
or U3785 (N_3785,N_2700,N_2444);
nor U3786 (N_3786,N_2433,N_2314);
nand U3787 (N_3787,N_2261,N_2929);
or U3788 (N_3788,N_2249,N_2463);
xor U3789 (N_3789,N_2390,N_2099);
nand U3790 (N_3790,N_2123,N_2775);
or U3791 (N_3791,N_2619,N_2239);
nand U3792 (N_3792,N_2319,N_2611);
nor U3793 (N_3793,N_2039,N_2520);
nand U3794 (N_3794,N_2249,N_2423);
nor U3795 (N_3795,N_2751,N_2324);
nor U3796 (N_3796,N_2284,N_2629);
or U3797 (N_3797,N_2134,N_2171);
nand U3798 (N_3798,N_2095,N_2345);
or U3799 (N_3799,N_2773,N_2782);
nand U3800 (N_3800,N_2379,N_2417);
or U3801 (N_3801,N_2518,N_2441);
nand U3802 (N_3802,N_2508,N_2271);
xnor U3803 (N_3803,N_2357,N_2526);
xnor U3804 (N_3804,N_2281,N_2188);
and U3805 (N_3805,N_2745,N_2122);
xor U3806 (N_3806,N_2403,N_2120);
nand U3807 (N_3807,N_2132,N_2135);
and U3808 (N_3808,N_2328,N_2473);
nor U3809 (N_3809,N_2029,N_2584);
or U3810 (N_3810,N_2975,N_2240);
or U3811 (N_3811,N_2939,N_2865);
nor U3812 (N_3812,N_2186,N_2629);
and U3813 (N_3813,N_2071,N_2823);
nor U3814 (N_3814,N_2534,N_2077);
nor U3815 (N_3815,N_2196,N_2772);
nor U3816 (N_3816,N_2331,N_2017);
nand U3817 (N_3817,N_2023,N_2032);
nand U3818 (N_3818,N_2440,N_2309);
nor U3819 (N_3819,N_2179,N_2151);
nand U3820 (N_3820,N_2176,N_2274);
nor U3821 (N_3821,N_2888,N_2608);
or U3822 (N_3822,N_2340,N_2265);
nand U3823 (N_3823,N_2244,N_2537);
or U3824 (N_3824,N_2678,N_2766);
or U3825 (N_3825,N_2809,N_2687);
nand U3826 (N_3826,N_2489,N_2372);
xnor U3827 (N_3827,N_2666,N_2374);
nor U3828 (N_3828,N_2405,N_2733);
and U3829 (N_3829,N_2624,N_2847);
or U3830 (N_3830,N_2100,N_2727);
nor U3831 (N_3831,N_2422,N_2821);
and U3832 (N_3832,N_2620,N_2893);
and U3833 (N_3833,N_2985,N_2448);
nor U3834 (N_3834,N_2430,N_2003);
xnor U3835 (N_3835,N_2992,N_2598);
and U3836 (N_3836,N_2971,N_2484);
or U3837 (N_3837,N_2271,N_2386);
nor U3838 (N_3838,N_2123,N_2899);
nand U3839 (N_3839,N_2993,N_2700);
nor U3840 (N_3840,N_2774,N_2763);
and U3841 (N_3841,N_2738,N_2611);
and U3842 (N_3842,N_2347,N_2791);
nand U3843 (N_3843,N_2091,N_2110);
and U3844 (N_3844,N_2333,N_2111);
or U3845 (N_3845,N_2636,N_2683);
nor U3846 (N_3846,N_2900,N_2577);
nor U3847 (N_3847,N_2408,N_2126);
xnor U3848 (N_3848,N_2499,N_2532);
nor U3849 (N_3849,N_2123,N_2737);
nand U3850 (N_3850,N_2802,N_2832);
nor U3851 (N_3851,N_2293,N_2275);
or U3852 (N_3852,N_2808,N_2356);
and U3853 (N_3853,N_2624,N_2356);
and U3854 (N_3854,N_2301,N_2717);
and U3855 (N_3855,N_2000,N_2956);
and U3856 (N_3856,N_2818,N_2299);
or U3857 (N_3857,N_2202,N_2773);
nor U3858 (N_3858,N_2550,N_2797);
and U3859 (N_3859,N_2948,N_2341);
and U3860 (N_3860,N_2047,N_2481);
or U3861 (N_3861,N_2579,N_2410);
or U3862 (N_3862,N_2581,N_2663);
and U3863 (N_3863,N_2167,N_2695);
and U3864 (N_3864,N_2885,N_2248);
nand U3865 (N_3865,N_2210,N_2826);
nand U3866 (N_3866,N_2280,N_2340);
nor U3867 (N_3867,N_2721,N_2064);
nand U3868 (N_3868,N_2940,N_2430);
nand U3869 (N_3869,N_2330,N_2452);
nor U3870 (N_3870,N_2498,N_2436);
nor U3871 (N_3871,N_2537,N_2116);
nor U3872 (N_3872,N_2908,N_2205);
nand U3873 (N_3873,N_2082,N_2756);
nand U3874 (N_3874,N_2004,N_2449);
nand U3875 (N_3875,N_2544,N_2288);
nand U3876 (N_3876,N_2794,N_2384);
and U3877 (N_3877,N_2987,N_2816);
nor U3878 (N_3878,N_2865,N_2601);
and U3879 (N_3879,N_2031,N_2876);
nor U3880 (N_3880,N_2729,N_2854);
nor U3881 (N_3881,N_2579,N_2226);
nand U3882 (N_3882,N_2140,N_2792);
nor U3883 (N_3883,N_2711,N_2369);
xor U3884 (N_3884,N_2476,N_2147);
or U3885 (N_3885,N_2052,N_2710);
nand U3886 (N_3886,N_2693,N_2993);
nor U3887 (N_3887,N_2143,N_2617);
and U3888 (N_3888,N_2934,N_2292);
and U3889 (N_3889,N_2902,N_2237);
or U3890 (N_3890,N_2135,N_2186);
xor U3891 (N_3891,N_2401,N_2866);
nand U3892 (N_3892,N_2858,N_2555);
and U3893 (N_3893,N_2540,N_2492);
or U3894 (N_3894,N_2809,N_2618);
and U3895 (N_3895,N_2876,N_2674);
and U3896 (N_3896,N_2864,N_2710);
nand U3897 (N_3897,N_2221,N_2371);
nor U3898 (N_3898,N_2981,N_2426);
and U3899 (N_3899,N_2629,N_2934);
and U3900 (N_3900,N_2466,N_2458);
or U3901 (N_3901,N_2723,N_2536);
xor U3902 (N_3902,N_2557,N_2045);
nor U3903 (N_3903,N_2812,N_2842);
and U3904 (N_3904,N_2028,N_2052);
xor U3905 (N_3905,N_2120,N_2432);
nand U3906 (N_3906,N_2140,N_2606);
or U3907 (N_3907,N_2479,N_2463);
nand U3908 (N_3908,N_2106,N_2728);
nor U3909 (N_3909,N_2061,N_2458);
and U3910 (N_3910,N_2233,N_2053);
nor U3911 (N_3911,N_2145,N_2624);
and U3912 (N_3912,N_2110,N_2907);
nand U3913 (N_3913,N_2254,N_2624);
and U3914 (N_3914,N_2605,N_2250);
nor U3915 (N_3915,N_2626,N_2171);
xor U3916 (N_3916,N_2353,N_2783);
and U3917 (N_3917,N_2249,N_2607);
or U3918 (N_3918,N_2272,N_2145);
nor U3919 (N_3919,N_2318,N_2386);
nand U3920 (N_3920,N_2594,N_2344);
xnor U3921 (N_3921,N_2085,N_2330);
or U3922 (N_3922,N_2695,N_2579);
and U3923 (N_3923,N_2397,N_2974);
xnor U3924 (N_3924,N_2122,N_2502);
nand U3925 (N_3925,N_2737,N_2245);
nand U3926 (N_3926,N_2876,N_2646);
nor U3927 (N_3927,N_2766,N_2295);
and U3928 (N_3928,N_2742,N_2674);
nor U3929 (N_3929,N_2266,N_2605);
nor U3930 (N_3930,N_2914,N_2459);
or U3931 (N_3931,N_2886,N_2212);
nor U3932 (N_3932,N_2014,N_2020);
and U3933 (N_3933,N_2764,N_2828);
or U3934 (N_3934,N_2719,N_2499);
nor U3935 (N_3935,N_2980,N_2544);
and U3936 (N_3936,N_2836,N_2449);
nand U3937 (N_3937,N_2259,N_2809);
xor U3938 (N_3938,N_2057,N_2549);
or U3939 (N_3939,N_2548,N_2247);
xnor U3940 (N_3940,N_2243,N_2882);
nor U3941 (N_3941,N_2867,N_2210);
or U3942 (N_3942,N_2421,N_2382);
nor U3943 (N_3943,N_2901,N_2365);
nand U3944 (N_3944,N_2145,N_2298);
nand U3945 (N_3945,N_2440,N_2511);
or U3946 (N_3946,N_2971,N_2906);
nor U3947 (N_3947,N_2467,N_2611);
nor U3948 (N_3948,N_2166,N_2517);
nand U3949 (N_3949,N_2859,N_2346);
or U3950 (N_3950,N_2691,N_2331);
nor U3951 (N_3951,N_2129,N_2341);
or U3952 (N_3952,N_2403,N_2372);
nor U3953 (N_3953,N_2483,N_2396);
and U3954 (N_3954,N_2309,N_2642);
nor U3955 (N_3955,N_2575,N_2794);
or U3956 (N_3956,N_2764,N_2840);
nor U3957 (N_3957,N_2920,N_2963);
or U3958 (N_3958,N_2363,N_2506);
or U3959 (N_3959,N_2252,N_2750);
and U3960 (N_3960,N_2162,N_2262);
xor U3961 (N_3961,N_2699,N_2588);
nand U3962 (N_3962,N_2140,N_2295);
or U3963 (N_3963,N_2698,N_2470);
nand U3964 (N_3964,N_2070,N_2885);
or U3965 (N_3965,N_2624,N_2735);
nor U3966 (N_3966,N_2324,N_2927);
nor U3967 (N_3967,N_2911,N_2373);
nand U3968 (N_3968,N_2362,N_2436);
and U3969 (N_3969,N_2476,N_2409);
xnor U3970 (N_3970,N_2801,N_2146);
or U3971 (N_3971,N_2441,N_2461);
or U3972 (N_3972,N_2421,N_2554);
and U3973 (N_3973,N_2906,N_2414);
nand U3974 (N_3974,N_2419,N_2629);
or U3975 (N_3975,N_2788,N_2216);
nand U3976 (N_3976,N_2354,N_2286);
and U3977 (N_3977,N_2157,N_2341);
xor U3978 (N_3978,N_2115,N_2422);
xnor U3979 (N_3979,N_2291,N_2448);
and U3980 (N_3980,N_2299,N_2347);
or U3981 (N_3981,N_2947,N_2294);
and U3982 (N_3982,N_2793,N_2560);
and U3983 (N_3983,N_2325,N_2350);
nor U3984 (N_3984,N_2443,N_2038);
and U3985 (N_3985,N_2655,N_2785);
nor U3986 (N_3986,N_2333,N_2592);
nor U3987 (N_3987,N_2106,N_2307);
nand U3988 (N_3988,N_2209,N_2156);
or U3989 (N_3989,N_2742,N_2085);
xor U3990 (N_3990,N_2927,N_2901);
or U3991 (N_3991,N_2822,N_2323);
nand U3992 (N_3992,N_2655,N_2129);
or U3993 (N_3993,N_2497,N_2870);
and U3994 (N_3994,N_2498,N_2537);
or U3995 (N_3995,N_2286,N_2184);
or U3996 (N_3996,N_2456,N_2490);
and U3997 (N_3997,N_2026,N_2436);
and U3998 (N_3998,N_2485,N_2947);
or U3999 (N_3999,N_2128,N_2538);
or U4000 (N_4000,N_3477,N_3825);
xnor U4001 (N_4001,N_3503,N_3898);
nor U4002 (N_4002,N_3808,N_3348);
nor U4003 (N_4003,N_3134,N_3890);
or U4004 (N_4004,N_3499,N_3698);
or U4005 (N_4005,N_3545,N_3066);
xor U4006 (N_4006,N_3551,N_3256);
and U4007 (N_4007,N_3979,N_3332);
nand U4008 (N_4008,N_3307,N_3687);
or U4009 (N_4009,N_3353,N_3373);
and U4010 (N_4010,N_3925,N_3516);
or U4011 (N_4011,N_3905,N_3127);
xor U4012 (N_4012,N_3575,N_3234);
and U4013 (N_4013,N_3467,N_3835);
and U4014 (N_4014,N_3676,N_3514);
and U4015 (N_4015,N_3889,N_3419);
or U4016 (N_4016,N_3966,N_3100);
nor U4017 (N_4017,N_3781,N_3543);
nor U4018 (N_4018,N_3088,N_3400);
or U4019 (N_4019,N_3039,N_3357);
and U4020 (N_4020,N_3518,N_3047);
or U4021 (N_4021,N_3011,N_3365);
nand U4022 (N_4022,N_3466,N_3061);
nor U4023 (N_4023,N_3085,N_3236);
and U4024 (N_4024,N_3582,N_3857);
nand U4025 (N_4025,N_3157,N_3622);
nand U4026 (N_4026,N_3691,N_3570);
xnor U4027 (N_4027,N_3382,N_3787);
nand U4028 (N_4028,N_3405,N_3488);
and U4029 (N_4029,N_3663,N_3867);
nor U4030 (N_4030,N_3693,N_3305);
nand U4031 (N_4031,N_3831,N_3786);
and U4032 (N_4032,N_3126,N_3653);
xor U4033 (N_4033,N_3189,N_3214);
and U4034 (N_4034,N_3866,N_3123);
or U4035 (N_4035,N_3121,N_3681);
nand U4036 (N_4036,N_3945,N_3447);
and U4037 (N_4037,N_3186,N_3745);
nor U4038 (N_4038,N_3022,N_3480);
nand U4039 (N_4039,N_3069,N_3221);
and U4040 (N_4040,N_3721,N_3457);
nor U4041 (N_4041,N_3815,N_3832);
nor U4042 (N_4042,N_3573,N_3602);
nor U4043 (N_4043,N_3208,N_3362);
xnor U4044 (N_4044,N_3046,N_3374);
and U4045 (N_4045,N_3963,N_3548);
nor U4046 (N_4046,N_3107,N_3692);
or U4047 (N_4047,N_3559,N_3398);
nand U4048 (N_4048,N_3724,N_3198);
and U4049 (N_4049,N_3395,N_3145);
xor U4050 (N_4050,N_3428,N_3555);
nand U4051 (N_4051,N_3961,N_3689);
nand U4052 (N_4052,N_3836,N_3279);
nor U4053 (N_4053,N_3713,N_3420);
nor U4054 (N_4054,N_3772,N_3408);
or U4055 (N_4055,N_3792,N_3810);
or U4056 (N_4056,N_3727,N_3601);
or U4057 (N_4057,N_3885,N_3344);
nor U4058 (N_4058,N_3747,N_3049);
nor U4059 (N_4059,N_3132,N_3768);
nor U4060 (N_4060,N_3935,N_3036);
or U4061 (N_4061,N_3274,N_3504);
and U4062 (N_4062,N_3986,N_3980);
and U4063 (N_4063,N_3245,N_3042);
xnor U4064 (N_4064,N_3782,N_3795);
and U4065 (N_4065,N_3656,N_3811);
nor U4066 (N_4066,N_3062,N_3052);
nand U4067 (N_4067,N_3872,N_3006);
or U4068 (N_4068,N_3718,N_3759);
nand U4069 (N_4069,N_3094,N_3226);
and U4070 (N_4070,N_3711,N_3156);
nand U4071 (N_4071,N_3129,N_3669);
nand U4072 (N_4072,N_3369,N_3677);
and U4073 (N_4073,N_3306,N_3024);
nand U4074 (N_4074,N_3003,N_3794);
nand U4075 (N_4075,N_3170,N_3084);
nor U4076 (N_4076,N_3078,N_3426);
xor U4077 (N_4077,N_3192,N_3865);
and U4078 (N_4078,N_3101,N_3947);
nand U4079 (N_4079,N_3137,N_3363);
and U4080 (N_4080,N_3233,N_3299);
nor U4081 (N_4081,N_3922,N_3526);
xnor U4082 (N_4082,N_3859,N_3005);
and U4083 (N_4083,N_3125,N_3641);
or U4084 (N_4084,N_3584,N_3934);
and U4085 (N_4085,N_3148,N_3250);
and U4086 (N_4086,N_3197,N_3339);
nand U4087 (N_4087,N_3478,N_3139);
xnor U4088 (N_4088,N_3613,N_3605);
and U4089 (N_4089,N_3273,N_3318);
or U4090 (N_4090,N_3871,N_3141);
or U4091 (N_4091,N_3425,N_3291);
nand U4092 (N_4092,N_3846,N_3805);
nand U4093 (N_4093,N_3690,N_3349);
nand U4094 (N_4094,N_3124,N_3591);
nand U4095 (N_4095,N_3886,N_3163);
and U4096 (N_4096,N_3410,N_3512);
nand U4097 (N_4097,N_3701,N_3229);
and U4098 (N_4098,N_3965,N_3056);
and U4099 (N_4099,N_3596,N_3450);
nor U4100 (N_4100,N_3709,N_3762);
xor U4101 (N_4101,N_3235,N_3699);
nand U4102 (N_4102,N_3660,N_3975);
nor U4103 (N_4103,N_3538,N_3902);
or U4104 (N_4104,N_3059,N_3485);
nor U4105 (N_4105,N_3744,N_3376);
nand U4106 (N_4106,N_3443,N_3916);
or U4107 (N_4107,N_3923,N_3719);
and U4108 (N_4108,N_3414,N_3817);
nand U4109 (N_4109,N_3300,N_3267);
and U4110 (N_4110,N_3589,N_3638);
or U4111 (N_4111,N_3496,N_3015);
or U4112 (N_4112,N_3280,N_3623);
nand U4113 (N_4113,N_3804,N_3160);
nor U4114 (N_4114,N_3377,N_3619);
or U4115 (N_4115,N_3714,N_3430);
nand U4116 (N_4116,N_3568,N_3284);
or U4117 (N_4117,N_3972,N_3493);
nand U4118 (N_4118,N_3595,N_3682);
nor U4119 (N_4119,N_3448,N_3833);
and U4120 (N_4120,N_3283,N_3295);
nor U4121 (N_4121,N_3278,N_3440);
or U4122 (N_4122,N_3055,N_3816);
xor U4123 (N_4123,N_3571,N_3281);
or U4124 (N_4124,N_3521,N_3712);
xor U4125 (N_4125,N_3065,N_3976);
and U4126 (N_4126,N_3556,N_3812);
nor U4127 (N_4127,N_3684,N_3996);
or U4128 (N_4128,N_3436,N_3341);
xnor U4129 (N_4129,N_3176,N_3708);
and U4130 (N_4130,N_3847,N_3057);
nand U4131 (N_4131,N_3607,N_3862);
nand U4132 (N_4132,N_3385,N_3809);
xor U4133 (N_4133,N_3704,N_3199);
xor U4134 (N_4134,N_3020,N_3603);
xor U4135 (N_4135,N_3325,N_3914);
and U4136 (N_4136,N_3298,N_3726);
xnor U4137 (N_4137,N_3232,N_3658);
and U4138 (N_4138,N_3824,N_3883);
nand U4139 (N_4139,N_3820,N_3322);
nand U4140 (N_4140,N_3111,N_3814);
xnor U4141 (N_4141,N_3608,N_3860);
xor U4142 (N_4142,N_3995,N_3268);
nor U4143 (N_4143,N_3407,N_3540);
nor U4144 (N_4144,N_3371,N_3722);
and U4145 (N_4145,N_3557,N_3984);
xnor U4146 (N_4146,N_3928,N_3948);
nand U4147 (N_4147,N_3943,N_3444);
or U4148 (N_4148,N_3051,N_3949);
nor U4149 (N_4149,N_3741,N_3252);
and U4150 (N_4150,N_3523,N_3579);
xnor U4151 (N_4151,N_3293,N_3218);
and U4152 (N_4152,N_3610,N_3451);
and U4153 (N_4153,N_3565,N_3618);
and U4154 (N_4154,N_3505,N_3520);
xnor U4155 (N_4155,N_3191,N_3275);
nand U4156 (N_4156,N_3265,N_3894);
xor U4157 (N_4157,N_3841,N_3182);
nand U4158 (N_4158,N_3981,N_3577);
nand U4159 (N_4159,N_3880,N_3277);
and U4160 (N_4160,N_3650,N_3799);
nor U4161 (N_4161,N_3219,N_3239);
nor U4162 (N_4162,N_3875,N_3616);
or U4163 (N_4163,N_3432,N_3155);
nand U4164 (N_4164,N_3924,N_3585);
and U4165 (N_4165,N_3490,N_3651);
nand U4166 (N_4166,N_3509,N_3884);
nand U4167 (N_4167,N_3133,N_3533);
nor U4168 (N_4168,N_3458,N_3159);
nand U4169 (N_4169,N_3368,N_3175);
nor U4170 (N_4170,N_3498,N_3674);
or U4171 (N_4171,N_3931,N_3661);
or U4172 (N_4172,N_3876,N_3639);
or U4173 (N_4173,N_3383,N_3738);
nand U4174 (N_4174,N_3647,N_3827);
and U4175 (N_4175,N_3461,N_3891);
nor U4176 (N_4176,N_3586,N_3850);
nand U4177 (N_4177,N_3528,N_3287);
and U4178 (N_4178,N_3413,N_3750);
or U4179 (N_4179,N_3029,N_3169);
or U4180 (N_4180,N_3072,N_3513);
and U4181 (N_4181,N_3248,N_3249);
nor U4182 (N_4182,N_3359,N_3522);
and U4183 (N_4183,N_3671,N_3725);
nor U4184 (N_4184,N_3933,N_3845);
nand U4185 (N_4185,N_3347,N_3379);
nand U4186 (N_4186,N_3920,N_3899);
and U4187 (N_4187,N_3043,N_3355);
nor U4188 (N_4188,N_3999,N_3896);
nand U4189 (N_4189,N_3659,N_3957);
nand U4190 (N_4190,N_3097,N_3225);
nand U4191 (N_4191,N_3956,N_3893);
nor U4192 (N_4192,N_3761,N_3646);
nor U4193 (N_4193,N_3828,N_3764);
nand U4194 (N_4194,N_3212,N_3580);
or U4195 (N_4195,N_3858,N_3630);
and U4196 (N_4196,N_3755,N_3384);
and U4197 (N_4197,N_3624,N_3746);
and U4198 (N_4198,N_3168,N_3113);
and U4199 (N_4199,N_3913,N_3813);
and U4200 (N_4200,N_3678,N_3951);
or U4201 (N_4201,N_3779,N_3146);
nor U4202 (N_4202,N_3184,N_3282);
or U4203 (N_4203,N_3465,N_3853);
or U4204 (N_4204,N_3769,N_3209);
nor U4205 (N_4205,N_3370,N_3271);
and U4206 (N_4206,N_3936,N_3797);
and U4207 (N_4207,N_3452,N_3844);
or U4208 (N_4208,N_3083,N_3262);
and U4209 (N_4209,N_3435,N_3544);
and U4210 (N_4210,N_3380,N_3753);
and U4211 (N_4211,N_3574,N_3806);
or U4212 (N_4212,N_3007,N_3227);
xor U4213 (N_4213,N_3328,N_3662);
nor U4214 (N_4214,N_3144,N_3321);
nand U4215 (N_4215,N_3688,N_3908);
nor U4216 (N_4216,N_3946,N_3877);
or U4217 (N_4217,N_3930,N_3354);
nand U4218 (N_4218,N_3429,N_3732);
nand U4219 (N_4219,N_3897,N_3257);
and U4220 (N_4220,N_3723,N_3290);
or U4221 (N_4221,N_3801,N_3600);
nor U4222 (N_4222,N_3937,N_3092);
nand U4223 (N_4223,N_3323,N_3968);
or U4224 (N_4224,N_3918,N_3849);
or U4225 (N_4225,N_3469,N_3592);
nand U4226 (N_4226,N_3629,N_3120);
nor U4227 (N_4227,N_3785,N_3459);
nand U4228 (N_4228,N_3422,N_3479);
xor U4229 (N_4229,N_3783,N_3237);
xor U4230 (N_4230,N_3453,N_3040);
or U4231 (N_4231,N_3238,N_3912);
or U4232 (N_4232,N_3864,N_3734);
nor U4233 (N_4233,N_3386,N_3438);
xor U4234 (N_4234,N_3462,N_3188);
nor U4235 (N_4235,N_3330,N_3054);
and U4236 (N_4236,N_3955,N_3567);
or U4237 (N_4237,N_3736,N_3320);
or U4238 (N_4238,N_3507,N_3626);
nand U4239 (N_4239,N_3473,N_3973);
nand U4240 (N_4240,N_3977,N_3843);
nand U4241 (N_4241,N_3686,N_3631);
and U4242 (N_4242,N_3529,N_3077);
or U4243 (N_4243,N_3308,N_3775);
and U4244 (N_4244,N_3441,N_3439);
nand U4245 (N_4245,N_3103,N_3494);
xor U4246 (N_4246,N_3154,N_3789);
or U4247 (N_4247,N_3643,N_3185);
nand U4248 (N_4248,N_3166,N_3487);
nor U4249 (N_4249,N_3076,N_3645);
nor U4250 (N_4250,N_3878,N_3378);
nand U4251 (N_4251,N_3991,N_3819);
nand U4252 (N_4252,N_3165,N_3666);
and U4253 (N_4253,N_3840,N_3285);
nor U4254 (N_4254,N_3838,N_3672);
or U4255 (N_4255,N_3336,N_3404);
or U4256 (N_4256,N_3401,N_3969);
or U4257 (N_4257,N_3988,N_3879);
or U4258 (N_4258,N_3151,N_3118);
nand U4259 (N_4259,N_3338,N_3563);
nor U4260 (N_4260,N_3941,N_3068);
nand U4261 (N_4261,N_3959,N_3392);
nor U4262 (N_4262,N_3763,N_3437);
or U4263 (N_4263,N_3652,N_3826);
and U4264 (N_4264,N_3263,N_3823);
and U4265 (N_4265,N_3220,N_3486);
and U4266 (N_4266,N_3205,N_3201);
xnor U4267 (N_4267,N_3707,N_3576);
nor U4268 (N_4268,N_3492,N_3352);
nand U4269 (N_4269,N_3294,N_3906);
or U4270 (N_4270,N_3030,N_3446);
or U4271 (N_4271,N_3770,N_3096);
nor U4272 (N_4272,N_3694,N_3754);
nor U4273 (N_4273,N_3390,N_3019);
or U4274 (N_4274,N_3014,N_3167);
nor U4275 (N_4275,N_3997,N_3416);
nand U4276 (N_4276,N_3900,N_3442);
or U4277 (N_4277,N_3793,N_3715);
xor U4278 (N_4278,N_3970,N_3919);
nor U4279 (N_4279,N_3194,N_3621);
nor U4280 (N_4280,N_3177,N_3842);
and U4281 (N_4281,N_3091,N_3756);
nand U4282 (N_4282,N_3983,N_3153);
and U4283 (N_4283,N_3105,N_3181);
nand U4284 (N_4284,N_3319,N_3978);
nand U4285 (N_4285,N_3481,N_3861);
or U4286 (N_4286,N_3010,N_3818);
nand U4287 (N_4287,N_3086,N_3482);
nand U4288 (N_4288,N_3475,N_3501);
and U4289 (N_4289,N_3588,N_3207);
or U4290 (N_4290,N_3260,N_3335);
nand U4291 (N_4291,N_3391,N_3637);
and U4292 (N_4292,N_3800,N_3106);
xnor U4293 (N_4293,N_3270,N_3032);
or U4294 (N_4294,N_3748,N_3033);
and U4295 (N_4295,N_3953,N_3216);
nand U4296 (N_4296,N_3561,N_3038);
nor U4297 (N_4297,N_3028,N_3854);
nand U4298 (N_4298,N_3244,N_3735);
and U4299 (N_4299,N_3259,N_3484);
or U4300 (N_4300,N_3640,N_3733);
or U4301 (N_4301,N_3173,N_3697);
nor U4302 (N_4302,N_3751,N_3449);
and U4303 (N_4303,N_3366,N_3670);
nor U4304 (N_4304,N_3989,N_3381);
xor U4305 (N_4305,N_3519,N_3655);
and U4306 (N_4306,N_3471,N_3312);
xor U4307 (N_4307,N_3445,N_3074);
or U4308 (N_4308,N_3767,N_3717);
nor U4309 (N_4309,N_3803,N_3415);
xnor U4310 (N_4310,N_3668,N_3675);
and U4311 (N_4311,N_3881,N_3140);
and U4312 (N_4312,N_3050,N_3037);
nand U4313 (N_4313,N_3739,N_3327);
nand U4314 (N_4314,N_3217,N_3851);
nor U4315 (N_4315,N_3149,N_3648);
nand U4316 (N_4316,N_3784,N_3636);
xor U4317 (N_4317,N_3228,N_3009);
and U4318 (N_4318,N_3903,N_3927);
or U4319 (N_4319,N_3994,N_3546);
nor U4320 (N_4320,N_3583,N_3604);
or U4321 (N_4321,N_3939,N_3508);
xor U4322 (N_4322,N_3635,N_3642);
nand U4323 (N_4323,N_3350,N_3578);
or U4324 (N_4324,N_3387,N_3231);
nand U4325 (N_4325,N_3564,N_3644);
xnor U4326 (N_4326,N_3064,N_3255);
nor U4327 (N_4327,N_3830,N_3301);
nand U4328 (N_4328,N_3628,N_3004);
nand U4329 (N_4329,N_3292,N_3915);
nor U4330 (N_4330,N_3119,N_3837);
or U4331 (N_4331,N_3324,N_3780);
nand U4332 (N_4332,N_3539,N_3992);
xor U4333 (N_4333,N_3702,N_3164);
nand U4334 (N_4334,N_3073,N_3873);
or U4335 (N_4335,N_3460,N_3476);
or U4336 (N_4336,N_3614,N_3740);
nor U4337 (N_4337,N_3152,N_3612);
or U4338 (N_4338,N_3852,N_3720);
nand U4339 (N_4339,N_3109,N_3547);
xnor U4340 (N_4340,N_3456,N_3537);
nor U4341 (N_4341,N_3314,N_3215);
nand U4342 (N_4342,N_3468,N_3510);
nand U4343 (N_4343,N_3625,N_3397);
nor U4344 (N_4344,N_3193,N_3269);
nand U4345 (N_4345,N_3863,N_3790);
nand U4346 (N_4346,N_3634,N_3394);
nand U4347 (N_4347,N_3026,N_3230);
nor U4348 (N_4348,N_3749,N_3087);
or U4349 (N_4349,N_3206,N_3243);
nand U4350 (N_4350,N_3333,N_3700);
nand U4351 (N_4351,N_3210,N_3599);
nand U4352 (N_4352,N_3904,N_3572);
nand U4353 (N_4353,N_3778,N_3388);
or U4354 (N_4354,N_3093,N_3195);
and U4355 (N_4355,N_3654,N_3337);
and U4356 (N_4356,N_3023,N_3921);
xor U4357 (N_4357,N_3822,N_3590);
or U4358 (N_4358,N_3553,N_3649);
or U4359 (N_4359,N_3421,N_3587);
or U4360 (N_4360,N_3550,N_3502);
nor U4361 (N_4361,N_3423,N_3855);
or U4362 (N_4362,N_3211,N_3190);
or U4363 (N_4363,N_3174,N_3895);
nor U4364 (N_4364,N_3705,N_3266);
and U4365 (N_4365,N_3346,N_3315);
or U4366 (N_4366,N_3581,N_3673);
nor U4367 (N_4367,N_3296,N_3679);
or U4368 (N_4368,N_3760,N_3560);
nand U4369 (N_4369,N_3807,N_3090);
or U4370 (N_4370,N_3424,N_3311);
nor U4371 (N_4371,N_3489,N_3773);
or U4372 (N_4372,N_3982,N_3632);
or U4373 (N_4373,N_3002,N_3147);
nand U4374 (N_4374,N_3060,N_3431);
and U4375 (N_4375,N_3964,N_3901);
or U4376 (N_4376,N_3246,N_3798);
nor U4377 (N_4377,N_3788,N_3117);
nor U4378 (N_4378,N_3351,N_3954);
xnor U4379 (N_4379,N_3500,N_3716);
nor U4380 (N_4380,N_3549,N_3909);
xnor U4381 (N_4381,N_3834,N_3515);
nor U4382 (N_4382,N_3597,N_3455);
xnor U4383 (N_4383,N_3776,N_3554);
nor U4384 (N_4384,N_3372,N_3114);
nand U4385 (N_4385,N_3535,N_3247);
nand U4386 (N_4386,N_3288,N_3310);
and U4387 (N_4387,N_3075,N_3839);
nor U4388 (N_4388,N_3329,N_3021);
nor U4389 (N_4389,N_3829,N_3987);
and U4390 (N_4390,N_3360,N_3342);
or U4391 (N_4391,N_3869,N_3758);
nand U4392 (N_4392,N_3095,N_3730);
and U4393 (N_4393,N_3258,N_3929);
or U4394 (N_4394,N_3304,N_3356);
and U4395 (N_4395,N_3598,N_3178);
nand U4396 (N_4396,N_3874,N_3402);
nor U4397 (N_4397,N_3364,N_3187);
or U4398 (N_4398,N_3017,N_3998);
or U4399 (N_4399,N_3771,N_3375);
nor U4400 (N_4400,N_3868,N_3034);
and U4401 (N_4401,N_3737,N_3491);
or U4402 (N_4402,N_3196,N_3665);
or U4403 (N_4403,N_3534,N_3361);
and U4404 (N_4404,N_3393,N_3286);
or U4405 (N_4405,N_3222,N_3944);
nand U4406 (N_4406,N_3474,N_3962);
nand U4407 (N_4407,N_3958,N_3203);
nand U4408 (N_4408,N_3765,N_3495);
nand U4409 (N_4409,N_3082,N_3035);
xor U4410 (N_4410,N_3566,N_3728);
and U4411 (N_4411,N_3766,N_3223);
nor U4412 (N_4412,N_3008,N_3031);
nand U4413 (N_4413,N_3541,N_3367);
nand U4414 (N_4414,N_3742,N_3142);
or U4415 (N_4415,N_3264,N_3112);
or U4416 (N_4416,N_3752,N_3552);
or U4417 (N_4417,N_3411,N_3303);
and U4418 (N_4418,N_3940,N_3044);
nand U4419 (N_4419,N_3706,N_3358);
or U4420 (N_4420,N_3606,N_3213);
nand U4421 (N_4421,N_3696,N_3942);
nand U4422 (N_4422,N_3136,N_3135);
xor U4423 (N_4423,N_3483,N_3048);
nand U4424 (N_4424,N_3172,N_3657);
and U4425 (N_4425,N_3932,N_3202);
nand U4426 (N_4426,N_3888,N_3907);
and U4427 (N_4427,N_3870,N_3013);
or U4428 (N_4428,N_3045,N_3911);
nand U4429 (N_4429,N_3558,N_3887);
xor U4430 (N_4430,N_3403,N_3434);
or U4431 (N_4431,N_3001,N_3856);
nor U4432 (N_4432,N_3594,N_3396);
and U4433 (N_4433,N_3345,N_3729);
nand U4434 (N_4434,N_3180,N_3297);
nand U4435 (N_4435,N_3240,N_3241);
nor U4436 (N_4436,N_3012,N_3016);
nand U4437 (N_4437,N_3000,N_3882);
nor U4438 (N_4438,N_3081,N_3971);
xnor U4439 (N_4439,N_3974,N_3796);
and U4440 (N_4440,N_3938,N_3162);
and U4441 (N_4441,N_3161,N_3470);
nor U4442 (N_4442,N_3777,N_3289);
and U4443 (N_4443,N_3317,N_3389);
xor U4444 (N_4444,N_3326,N_3276);
nor U4445 (N_4445,N_3695,N_3967);
nor U4446 (N_4446,N_3417,N_3108);
nand U4447 (N_4447,N_3399,N_3183);
nand U4448 (N_4448,N_3418,N_3609);
nor U4449 (N_4449,N_3562,N_3633);
and U4450 (N_4450,N_3116,N_3089);
nand U4451 (N_4451,N_3150,N_3667);
or U4452 (N_4452,N_3179,N_3427);
and U4453 (N_4453,N_3224,N_3316);
and U4454 (N_4454,N_3952,N_3536);
xor U4455 (N_4455,N_3615,N_3334);
nand U4456 (N_4456,N_3079,N_3527);
or U4457 (N_4457,N_3593,N_3703);
xnor U4458 (N_4458,N_3497,N_3985);
nor U4459 (N_4459,N_3517,N_3104);
and U4460 (N_4460,N_3532,N_3506);
and U4461 (N_4461,N_3821,N_3454);
nand U4462 (N_4462,N_3018,N_3524);
and U4463 (N_4463,N_3710,N_3058);
nor U4464 (N_4464,N_3071,N_3343);
nand U4465 (N_4465,N_3313,N_3960);
xor U4466 (N_4466,N_3892,N_3433);
nand U4467 (N_4467,N_3917,N_3251);
nor U4468 (N_4468,N_3110,N_3993);
or U4469 (N_4469,N_3412,N_3261);
or U4470 (N_4470,N_3743,N_3530);
nand U4471 (N_4471,N_3254,N_3627);
xor U4472 (N_4472,N_3158,N_3302);
xnor U4473 (N_4473,N_3067,N_3683);
nand U4474 (N_4474,N_3620,N_3531);
nand U4475 (N_4475,N_3063,N_3926);
nand U4476 (N_4476,N_3406,N_3115);
xor U4477 (N_4477,N_3053,N_3472);
and U4478 (N_4478,N_3542,N_3143);
nor U4479 (N_4479,N_3025,N_3731);
nand U4480 (N_4480,N_3409,N_3130);
and U4481 (N_4481,N_3027,N_3664);
nand U4482 (N_4482,N_3525,N_3138);
or U4483 (N_4483,N_3171,N_3774);
nor U4484 (N_4484,N_3950,N_3309);
and U4485 (N_4485,N_3102,N_3910);
nand U4486 (N_4486,N_3331,N_3802);
xor U4487 (N_4487,N_3041,N_3272);
nand U4488 (N_4488,N_3340,N_3122);
or U4489 (N_4489,N_3680,N_3204);
or U4490 (N_4490,N_3253,N_3611);
nor U4491 (N_4491,N_3242,N_3080);
nand U4492 (N_4492,N_3848,N_3791);
or U4493 (N_4493,N_3569,N_3990);
and U4494 (N_4494,N_3098,N_3128);
nand U4495 (N_4495,N_3617,N_3464);
xor U4496 (N_4496,N_3099,N_3511);
xor U4497 (N_4497,N_3757,N_3463);
and U4498 (N_4498,N_3685,N_3131);
nor U4499 (N_4499,N_3200,N_3070);
or U4500 (N_4500,N_3176,N_3425);
nand U4501 (N_4501,N_3909,N_3593);
and U4502 (N_4502,N_3676,N_3253);
or U4503 (N_4503,N_3963,N_3809);
or U4504 (N_4504,N_3140,N_3647);
or U4505 (N_4505,N_3565,N_3707);
nand U4506 (N_4506,N_3258,N_3809);
or U4507 (N_4507,N_3258,N_3004);
nor U4508 (N_4508,N_3577,N_3301);
nand U4509 (N_4509,N_3641,N_3311);
or U4510 (N_4510,N_3981,N_3313);
and U4511 (N_4511,N_3756,N_3962);
or U4512 (N_4512,N_3049,N_3672);
and U4513 (N_4513,N_3015,N_3754);
nand U4514 (N_4514,N_3009,N_3819);
xor U4515 (N_4515,N_3210,N_3186);
and U4516 (N_4516,N_3198,N_3684);
and U4517 (N_4517,N_3478,N_3030);
nor U4518 (N_4518,N_3280,N_3478);
and U4519 (N_4519,N_3699,N_3630);
or U4520 (N_4520,N_3807,N_3553);
nor U4521 (N_4521,N_3160,N_3411);
or U4522 (N_4522,N_3906,N_3152);
and U4523 (N_4523,N_3184,N_3463);
nor U4524 (N_4524,N_3247,N_3003);
and U4525 (N_4525,N_3021,N_3941);
and U4526 (N_4526,N_3996,N_3729);
nand U4527 (N_4527,N_3106,N_3693);
and U4528 (N_4528,N_3456,N_3839);
nor U4529 (N_4529,N_3843,N_3490);
or U4530 (N_4530,N_3851,N_3934);
or U4531 (N_4531,N_3717,N_3904);
or U4532 (N_4532,N_3021,N_3636);
nor U4533 (N_4533,N_3328,N_3765);
or U4534 (N_4534,N_3352,N_3449);
nand U4535 (N_4535,N_3006,N_3644);
nor U4536 (N_4536,N_3565,N_3598);
nor U4537 (N_4537,N_3182,N_3875);
xnor U4538 (N_4538,N_3252,N_3315);
xnor U4539 (N_4539,N_3430,N_3588);
nor U4540 (N_4540,N_3291,N_3545);
or U4541 (N_4541,N_3893,N_3911);
nand U4542 (N_4542,N_3030,N_3486);
or U4543 (N_4543,N_3032,N_3798);
nor U4544 (N_4544,N_3622,N_3603);
or U4545 (N_4545,N_3955,N_3173);
nor U4546 (N_4546,N_3052,N_3899);
nor U4547 (N_4547,N_3295,N_3973);
or U4548 (N_4548,N_3745,N_3188);
nor U4549 (N_4549,N_3535,N_3950);
and U4550 (N_4550,N_3968,N_3717);
and U4551 (N_4551,N_3441,N_3290);
and U4552 (N_4552,N_3798,N_3632);
or U4553 (N_4553,N_3670,N_3961);
nand U4554 (N_4554,N_3603,N_3988);
and U4555 (N_4555,N_3203,N_3795);
nor U4556 (N_4556,N_3734,N_3310);
and U4557 (N_4557,N_3007,N_3034);
nand U4558 (N_4558,N_3492,N_3504);
nand U4559 (N_4559,N_3466,N_3623);
and U4560 (N_4560,N_3206,N_3904);
nand U4561 (N_4561,N_3888,N_3103);
nand U4562 (N_4562,N_3393,N_3631);
nor U4563 (N_4563,N_3659,N_3402);
or U4564 (N_4564,N_3047,N_3705);
or U4565 (N_4565,N_3408,N_3249);
nand U4566 (N_4566,N_3131,N_3066);
nor U4567 (N_4567,N_3049,N_3973);
nand U4568 (N_4568,N_3913,N_3265);
or U4569 (N_4569,N_3788,N_3582);
nor U4570 (N_4570,N_3907,N_3327);
nor U4571 (N_4571,N_3792,N_3676);
nand U4572 (N_4572,N_3690,N_3698);
nor U4573 (N_4573,N_3577,N_3965);
nor U4574 (N_4574,N_3668,N_3920);
or U4575 (N_4575,N_3294,N_3313);
and U4576 (N_4576,N_3237,N_3966);
nor U4577 (N_4577,N_3758,N_3637);
and U4578 (N_4578,N_3759,N_3632);
nor U4579 (N_4579,N_3218,N_3601);
nor U4580 (N_4580,N_3983,N_3002);
nand U4581 (N_4581,N_3100,N_3787);
nand U4582 (N_4582,N_3108,N_3647);
nor U4583 (N_4583,N_3864,N_3684);
and U4584 (N_4584,N_3158,N_3449);
nor U4585 (N_4585,N_3177,N_3508);
nand U4586 (N_4586,N_3312,N_3154);
nor U4587 (N_4587,N_3829,N_3656);
or U4588 (N_4588,N_3674,N_3977);
nand U4589 (N_4589,N_3769,N_3973);
and U4590 (N_4590,N_3426,N_3332);
nor U4591 (N_4591,N_3667,N_3176);
nor U4592 (N_4592,N_3774,N_3919);
or U4593 (N_4593,N_3163,N_3838);
xnor U4594 (N_4594,N_3953,N_3309);
and U4595 (N_4595,N_3887,N_3424);
nand U4596 (N_4596,N_3562,N_3342);
or U4597 (N_4597,N_3349,N_3212);
nor U4598 (N_4598,N_3539,N_3167);
nor U4599 (N_4599,N_3405,N_3632);
or U4600 (N_4600,N_3149,N_3447);
or U4601 (N_4601,N_3059,N_3487);
and U4602 (N_4602,N_3542,N_3674);
nor U4603 (N_4603,N_3247,N_3491);
nor U4604 (N_4604,N_3435,N_3844);
nor U4605 (N_4605,N_3142,N_3546);
nand U4606 (N_4606,N_3946,N_3561);
or U4607 (N_4607,N_3652,N_3434);
nor U4608 (N_4608,N_3295,N_3040);
or U4609 (N_4609,N_3716,N_3570);
and U4610 (N_4610,N_3760,N_3884);
or U4611 (N_4611,N_3173,N_3023);
nor U4612 (N_4612,N_3076,N_3459);
nand U4613 (N_4613,N_3152,N_3317);
or U4614 (N_4614,N_3332,N_3720);
nor U4615 (N_4615,N_3146,N_3557);
or U4616 (N_4616,N_3145,N_3196);
nand U4617 (N_4617,N_3015,N_3618);
nand U4618 (N_4618,N_3133,N_3152);
and U4619 (N_4619,N_3318,N_3130);
or U4620 (N_4620,N_3516,N_3620);
nand U4621 (N_4621,N_3715,N_3766);
and U4622 (N_4622,N_3162,N_3044);
xor U4623 (N_4623,N_3494,N_3986);
nor U4624 (N_4624,N_3915,N_3451);
nor U4625 (N_4625,N_3014,N_3921);
nor U4626 (N_4626,N_3744,N_3055);
and U4627 (N_4627,N_3634,N_3028);
nor U4628 (N_4628,N_3711,N_3716);
or U4629 (N_4629,N_3307,N_3674);
nand U4630 (N_4630,N_3248,N_3703);
and U4631 (N_4631,N_3473,N_3741);
nand U4632 (N_4632,N_3132,N_3916);
nor U4633 (N_4633,N_3642,N_3613);
nand U4634 (N_4634,N_3446,N_3122);
xnor U4635 (N_4635,N_3165,N_3586);
xnor U4636 (N_4636,N_3404,N_3836);
nand U4637 (N_4637,N_3980,N_3180);
nand U4638 (N_4638,N_3873,N_3434);
nor U4639 (N_4639,N_3754,N_3385);
and U4640 (N_4640,N_3703,N_3083);
or U4641 (N_4641,N_3260,N_3792);
nand U4642 (N_4642,N_3903,N_3719);
nand U4643 (N_4643,N_3215,N_3637);
or U4644 (N_4644,N_3838,N_3239);
xor U4645 (N_4645,N_3073,N_3421);
nor U4646 (N_4646,N_3327,N_3428);
nand U4647 (N_4647,N_3410,N_3967);
nor U4648 (N_4648,N_3739,N_3193);
nand U4649 (N_4649,N_3467,N_3382);
and U4650 (N_4650,N_3741,N_3895);
or U4651 (N_4651,N_3155,N_3436);
nor U4652 (N_4652,N_3485,N_3879);
and U4653 (N_4653,N_3576,N_3953);
xor U4654 (N_4654,N_3279,N_3930);
or U4655 (N_4655,N_3963,N_3768);
or U4656 (N_4656,N_3799,N_3328);
or U4657 (N_4657,N_3047,N_3977);
nor U4658 (N_4658,N_3122,N_3736);
xor U4659 (N_4659,N_3239,N_3590);
or U4660 (N_4660,N_3894,N_3247);
nand U4661 (N_4661,N_3046,N_3867);
or U4662 (N_4662,N_3620,N_3440);
or U4663 (N_4663,N_3216,N_3214);
or U4664 (N_4664,N_3490,N_3521);
nor U4665 (N_4665,N_3993,N_3476);
and U4666 (N_4666,N_3457,N_3361);
and U4667 (N_4667,N_3799,N_3598);
nor U4668 (N_4668,N_3532,N_3112);
nor U4669 (N_4669,N_3438,N_3062);
nand U4670 (N_4670,N_3765,N_3789);
xor U4671 (N_4671,N_3225,N_3228);
and U4672 (N_4672,N_3266,N_3895);
nor U4673 (N_4673,N_3339,N_3657);
nor U4674 (N_4674,N_3043,N_3817);
xor U4675 (N_4675,N_3365,N_3852);
nor U4676 (N_4676,N_3529,N_3614);
and U4677 (N_4677,N_3404,N_3251);
nor U4678 (N_4678,N_3321,N_3482);
or U4679 (N_4679,N_3324,N_3365);
or U4680 (N_4680,N_3173,N_3149);
xor U4681 (N_4681,N_3557,N_3062);
nor U4682 (N_4682,N_3846,N_3000);
nand U4683 (N_4683,N_3925,N_3296);
or U4684 (N_4684,N_3909,N_3418);
or U4685 (N_4685,N_3154,N_3751);
nand U4686 (N_4686,N_3520,N_3255);
xor U4687 (N_4687,N_3877,N_3262);
and U4688 (N_4688,N_3361,N_3043);
nor U4689 (N_4689,N_3865,N_3798);
nor U4690 (N_4690,N_3072,N_3434);
nor U4691 (N_4691,N_3640,N_3327);
or U4692 (N_4692,N_3852,N_3152);
xor U4693 (N_4693,N_3511,N_3787);
and U4694 (N_4694,N_3932,N_3607);
or U4695 (N_4695,N_3848,N_3724);
nand U4696 (N_4696,N_3542,N_3124);
and U4697 (N_4697,N_3561,N_3216);
nor U4698 (N_4698,N_3590,N_3543);
and U4699 (N_4699,N_3673,N_3598);
and U4700 (N_4700,N_3027,N_3015);
and U4701 (N_4701,N_3327,N_3415);
and U4702 (N_4702,N_3844,N_3172);
xnor U4703 (N_4703,N_3651,N_3900);
xor U4704 (N_4704,N_3272,N_3988);
and U4705 (N_4705,N_3534,N_3664);
nand U4706 (N_4706,N_3419,N_3965);
nand U4707 (N_4707,N_3271,N_3995);
nor U4708 (N_4708,N_3682,N_3001);
nor U4709 (N_4709,N_3848,N_3967);
nand U4710 (N_4710,N_3552,N_3021);
and U4711 (N_4711,N_3681,N_3097);
nand U4712 (N_4712,N_3002,N_3715);
and U4713 (N_4713,N_3899,N_3128);
or U4714 (N_4714,N_3801,N_3441);
nor U4715 (N_4715,N_3050,N_3479);
and U4716 (N_4716,N_3702,N_3097);
and U4717 (N_4717,N_3387,N_3433);
xor U4718 (N_4718,N_3666,N_3901);
xnor U4719 (N_4719,N_3070,N_3089);
nand U4720 (N_4720,N_3812,N_3184);
and U4721 (N_4721,N_3858,N_3519);
and U4722 (N_4722,N_3203,N_3110);
xor U4723 (N_4723,N_3153,N_3289);
or U4724 (N_4724,N_3710,N_3465);
and U4725 (N_4725,N_3596,N_3889);
nand U4726 (N_4726,N_3575,N_3724);
or U4727 (N_4727,N_3840,N_3850);
and U4728 (N_4728,N_3014,N_3876);
xnor U4729 (N_4729,N_3746,N_3218);
or U4730 (N_4730,N_3706,N_3958);
nand U4731 (N_4731,N_3787,N_3659);
nand U4732 (N_4732,N_3051,N_3092);
or U4733 (N_4733,N_3428,N_3910);
nand U4734 (N_4734,N_3228,N_3059);
nand U4735 (N_4735,N_3831,N_3809);
or U4736 (N_4736,N_3631,N_3465);
nor U4737 (N_4737,N_3350,N_3071);
and U4738 (N_4738,N_3386,N_3756);
and U4739 (N_4739,N_3510,N_3968);
nand U4740 (N_4740,N_3188,N_3373);
and U4741 (N_4741,N_3489,N_3642);
nand U4742 (N_4742,N_3385,N_3435);
nor U4743 (N_4743,N_3495,N_3804);
nor U4744 (N_4744,N_3661,N_3901);
nor U4745 (N_4745,N_3224,N_3652);
and U4746 (N_4746,N_3569,N_3841);
and U4747 (N_4747,N_3073,N_3356);
nor U4748 (N_4748,N_3906,N_3277);
and U4749 (N_4749,N_3790,N_3931);
and U4750 (N_4750,N_3053,N_3635);
or U4751 (N_4751,N_3562,N_3621);
nor U4752 (N_4752,N_3032,N_3088);
and U4753 (N_4753,N_3528,N_3407);
and U4754 (N_4754,N_3595,N_3753);
or U4755 (N_4755,N_3448,N_3351);
nand U4756 (N_4756,N_3729,N_3771);
nand U4757 (N_4757,N_3106,N_3572);
nand U4758 (N_4758,N_3423,N_3780);
nor U4759 (N_4759,N_3652,N_3246);
or U4760 (N_4760,N_3183,N_3703);
nor U4761 (N_4761,N_3723,N_3997);
xor U4762 (N_4762,N_3992,N_3735);
xor U4763 (N_4763,N_3863,N_3032);
or U4764 (N_4764,N_3777,N_3234);
and U4765 (N_4765,N_3073,N_3847);
and U4766 (N_4766,N_3494,N_3924);
or U4767 (N_4767,N_3273,N_3058);
and U4768 (N_4768,N_3343,N_3333);
or U4769 (N_4769,N_3688,N_3715);
and U4770 (N_4770,N_3475,N_3595);
xnor U4771 (N_4771,N_3031,N_3909);
xnor U4772 (N_4772,N_3954,N_3216);
xor U4773 (N_4773,N_3366,N_3078);
and U4774 (N_4774,N_3080,N_3251);
or U4775 (N_4775,N_3180,N_3086);
nand U4776 (N_4776,N_3436,N_3346);
and U4777 (N_4777,N_3620,N_3686);
xnor U4778 (N_4778,N_3523,N_3850);
nand U4779 (N_4779,N_3888,N_3468);
xnor U4780 (N_4780,N_3093,N_3662);
nor U4781 (N_4781,N_3054,N_3942);
and U4782 (N_4782,N_3376,N_3419);
nand U4783 (N_4783,N_3654,N_3605);
or U4784 (N_4784,N_3565,N_3354);
or U4785 (N_4785,N_3270,N_3200);
nand U4786 (N_4786,N_3436,N_3638);
nor U4787 (N_4787,N_3757,N_3358);
or U4788 (N_4788,N_3511,N_3882);
nand U4789 (N_4789,N_3807,N_3044);
or U4790 (N_4790,N_3376,N_3638);
nand U4791 (N_4791,N_3873,N_3451);
and U4792 (N_4792,N_3489,N_3820);
xnor U4793 (N_4793,N_3864,N_3633);
xor U4794 (N_4794,N_3062,N_3427);
nand U4795 (N_4795,N_3612,N_3028);
xor U4796 (N_4796,N_3280,N_3861);
and U4797 (N_4797,N_3157,N_3652);
nor U4798 (N_4798,N_3095,N_3651);
and U4799 (N_4799,N_3264,N_3060);
nor U4800 (N_4800,N_3114,N_3988);
nor U4801 (N_4801,N_3242,N_3886);
nand U4802 (N_4802,N_3328,N_3512);
xnor U4803 (N_4803,N_3478,N_3480);
nand U4804 (N_4804,N_3936,N_3790);
or U4805 (N_4805,N_3894,N_3366);
nand U4806 (N_4806,N_3929,N_3343);
nor U4807 (N_4807,N_3876,N_3492);
nor U4808 (N_4808,N_3667,N_3844);
and U4809 (N_4809,N_3847,N_3711);
nand U4810 (N_4810,N_3957,N_3340);
or U4811 (N_4811,N_3555,N_3022);
nand U4812 (N_4812,N_3686,N_3719);
or U4813 (N_4813,N_3023,N_3148);
nor U4814 (N_4814,N_3179,N_3597);
nand U4815 (N_4815,N_3441,N_3563);
and U4816 (N_4816,N_3799,N_3624);
nor U4817 (N_4817,N_3064,N_3813);
nor U4818 (N_4818,N_3078,N_3138);
nand U4819 (N_4819,N_3496,N_3106);
nand U4820 (N_4820,N_3405,N_3238);
or U4821 (N_4821,N_3825,N_3927);
nand U4822 (N_4822,N_3384,N_3754);
nand U4823 (N_4823,N_3000,N_3103);
nand U4824 (N_4824,N_3714,N_3489);
or U4825 (N_4825,N_3786,N_3609);
nand U4826 (N_4826,N_3866,N_3048);
nand U4827 (N_4827,N_3071,N_3863);
nor U4828 (N_4828,N_3564,N_3570);
nand U4829 (N_4829,N_3695,N_3101);
nor U4830 (N_4830,N_3787,N_3678);
nor U4831 (N_4831,N_3668,N_3782);
nand U4832 (N_4832,N_3773,N_3983);
or U4833 (N_4833,N_3705,N_3638);
or U4834 (N_4834,N_3838,N_3503);
nor U4835 (N_4835,N_3960,N_3831);
or U4836 (N_4836,N_3880,N_3008);
or U4837 (N_4837,N_3510,N_3134);
and U4838 (N_4838,N_3528,N_3084);
nor U4839 (N_4839,N_3673,N_3662);
nand U4840 (N_4840,N_3174,N_3943);
and U4841 (N_4841,N_3620,N_3359);
or U4842 (N_4842,N_3807,N_3970);
and U4843 (N_4843,N_3890,N_3686);
and U4844 (N_4844,N_3401,N_3932);
or U4845 (N_4845,N_3331,N_3075);
xor U4846 (N_4846,N_3033,N_3806);
nand U4847 (N_4847,N_3559,N_3485);
nand U4848 (N_4848,N_3979,N_3386);
xor U4849 (N_4849,N_3849,N_3766);
or U4850 (N_4850,N_3956,N_3227);
nand U4851 (N_4851,N_3472,N_3396);
and U4852 (N_4852,N_3992,N_3725);
xnor U4853 (N_4853,N_3143,N_3452);
or U4854 (N_4854,N_3366,N_3442);
nor U4855 (N_4855,N_3512,N_3036);
nand U4856 (N_4856,N_3874,N_3743);
nor U4857 (N_4857,N_3869,N_3594);
nand U4858 (N_4858,N_3396,N_3536);
and U4859 (N_4859,N_3202,N_3233);
nand U4860 (N_4860,N_3680,N_3294);
nor U4861 (N_4861,N_3386,N_3791);
nor U4862 (N_4862,N_3336,N_3825);
or U4863 (N_4863,N_3870,N_3716);
nand U4864 (N_4864,N_3714,N_3781);
or U4865 (N_4865,N_3508,N_3936);
nand U4866 (N_4866,N_3109,N_3839);
nand U4867 (N_4867,N_3489,N_3249);
xnor U4868 (N_4868,N_3397,N_3448);
and U4869 (N_4869,N_3971,N_3985);
and U4870 (N_4870,N_3062,N_3775);
or U4871 (N_4871,N_3323,N_3844);
or U4872 (N_4872,N_3804,N_3716);
nand U4873 (N_4873,N_3290,N_3286);
and U4874 (N_4874,N_3156,N_3622);
nand U4875 (N_4875,N_3989,N_3555);
nor U4876 (N_4876,N_3066,N_3606);
nor U4877 (N_4877,N_3197,N_3416);
nor U4878 (N_4878,N_3212,N_3093);
nor U4879 (N_4879,N_3583,N_3407);
nor U4880 (N_4880,N_3737,N_3837);
nand U4881 (N_4881,N_3500,N_3074);
nand U4882 (N_4882,N_3554,N_3115);
or U4883 (N_4883,N_3881,N_3117);
and U4884 (N_4884,N_3298,N_3300);
nor U4885 (N_4885,N_3118,N_3862);
nor U4886 (N_4886,N_3690,N_3789);
nand U4887 (N_4887,N_3613,N_3100);
or U4888 (N_4888,N_3424,N_3310);
or U4889 (N_4889,N_3664,N_3596);
and U4890 (N_4890,N_3590,N_3495);
nor U4891 (N_4891,N_3010,N_3874);
or U4892 (N_4892,N_3538,N_3627);
and U4893 (N_4893,N_3785,N_3206);
or U4894 (N_4894,N_3585,N_3706);
nor U4895 (N_4895,N_3335,N_3816);
nand U4896 (N_4896,N_3099,N_3631);
and U4897 (N_4897,N_3146,N_3128);
and U4898 (N_4898,N_3591,N_3916);
or U4899 (N_4899,N_3038,N_3912);
nand U4900 (N_4900,N_3857,N_3162);
nor U4901 (N_4901,N_3964,N_3022);
and U4902 (N_4902,N_3284,N_3403);
and U4903 (N_4903,N_3947,N_3709);
or U4904 (N_4904,N_3274,N_3312);
or U4905 (N_4905,N_3385,N_3567);
and U4906 (N_4906,N_3260,N_3119);
and U4907 (N_4907,N_3354,N_3094);
nand U4908 (N_4908,N_3770,N_3093);
or U4909 (N_4909,N_3157,N_3470);
nand U4910 (N_4910,N_3650,N_3132);
nand U4911 (N_4911,N_3355,N_3554);
and U4912 (N_4912,N_3144,N_3207);
nor U4913 (N_4913,N_3885,N_3982);
xnor U4914 (N_4914,N_3048,N_3736);
nand U4915 (N_4915,N_3784,N_3986);
and U4916 (N_4916,N_3369,N_3352);
nand U4917 (N_4917,N_3650,N_3764);
and U4918 (N_4918,N_3331,N_3757);
xnor U4919 (N_4919,N_3719,N_3519);
and U4920 (N_4920,N_3099,N_3473);
nand U4921 (N_4921,N_3127,N_3672);
and U4922 (N_4922,N_3443,N_3653);
nand U4923 (N_4923,N_3002,N_3010);
xor U4924 (N_4924,N_3976,N_3245);
xor U4925 (N_4925,N_3701,N_3006);
and U4926 (N_4926,N_3968,N_3278);
nor U4927 (N_4927,N_3312,N_3991);
and U4928 (N_4928,N_3200,N_3358);
xnor U4929 (N_4929,N_3068,N_3088);
nand U4930 (N_4930,N_3596,N_3576);
nand U4931 (N_4931,N_3713,N_3233);
nor U4932 (N_4932,N_3710,N_3487);
or U4933 (N_4933,N_3137,N_3767);
or U4934 (N_4934,N_3913,N_3361);
or U4935 (N_4935,N_3689,N_3985);
nand U4936 (N_4936,N_3776,N_3579);
nor U4937 (N_4937,N_3704,N_3643);
or U4938 (N_4938,N_3157,N_3992);
nand U4939 (N_4939,N_3682,N_3660);
nor U4940 (N_4940,N_3828,N_3939);
xor U4941 (N_4941,N_3381,N_3795);
nand U4942 (N_4942,N_3027,N_3627);
or U4943 (N_4943,N_3211,N_3497);
or U4944 (N_4944,N_3588,N_3677);
xor U4945 (N_4945,N_3760,N_3499);
nand U4946 (N_4946,N_3553,N_3733);
nand U4947 (N_4947,N_3684,N_3582);
nand U4948 (N_4948,N_3877,N_3700);
and U4949 (N_4949,N_3145,N_3738);
nand U4950 (N_4950,N_3638,N_3477);
nor U4951 (N_4951,N_3867,N_3945);
nor U4952 (N_4952,N_3159,N_3323);
and U4953 (N_4953,N_3439,N_3261);
nand U4954 (N_4954,N_3756,N_3659);
nor U4955 (N_4955,N_3705,N_3037);
nor U4956 (N_4956,N_3456,N_3477);
nand U4957 (N_4957,N_3494,N_3577);
nor U4958 (N_4958,N_3718,N_3070);
nand U4959 (N_4959,N_3105,N_3393);
nor U4960 (N_4960,N_3339,N_3707);
nand U4961 (N_4961,N_3700,N_3412);
nor U4962 (N_4962,N_3345,N_3840);
and U4963 (N_4963,N_3317,N_3556);
or U4964 (N_4964,N_3518,N_3934);
nor U4965 (N_4965,N_3763,N_3244);
xnor U4966 (N_4966,N_3261,N_3494);
or U4967 (N_4967,N_3464,N_3936);
nand U4968 (N_4968,N_3368,N_3740);
or U4969 (N_4969,N_3076,N_3783);
nor U4970 (N_4970,N_3304,N_3452);
xnor U4971 (N_4971,N_3142,N_3402);
xor U4972 (N_4972,N_3697,N_3107);
nand U4973 (N_4973,N_3110,N_3398);
xnor U4974 (N_4974,N_3039,N_3922);
or U4975 (N_4975,N_3729,N_3809);
nand U4976 (N_4976,N_3147,N_3027);
xnor U4977 (N_4977,N_3705,N_3339);
nor U4978 (N_4978,N_3071,N_3028);
or U4979 (N_4979,N_3294,N_3971);
xor U4980 (N_4980,N_3588,N_3291);
nor U4981 (N_4981,N_3128,N_3366);
nor U4982 (N_4982,N_3670,N_3033);
and U4983 (N_4983,N_3470,N_3350);
xor U4984 (N_4984,N_3045,N_3116);
and U4985 (N_4985,N_3732,N_3832);
nand U4986 (N_4986,N_3991,N_3976);
nor U4987 (N_4987,N_3482,N_3947);
nand U4988 (N_4988,N_3401,N_3541);
nand U4989 (N_4989,N_3386,N_3642);
nand U4990 (N_4990,N_3568,N_3262);
or U4991 (N_4991,N_3489,N_3672);
and U4992 (N_4992,N_3399,N_3983);
or U4993 (N_4993,N_3492,N_3949);
and U4994 (N_4994,N_3977,N_3896);
and U4995 (N_4995,N_3838,N_3846);
nor U4996 (N_4996,N_3498,N_3973);
nand U4997 (N_4997,N_3221,N_3093);
or U4998 (N_4998,N_3978,N_3062);
nor U4999 (N_4999,N_3139,N_3718);
or U5000 (N_5000,N_4674,N_4397);
or U5001 (N_5001,N_4317,N_4227);
and U5002 (N_5002,N_4382,N_4771);
nand U5003 (N_5003,N_4727,N_4838);
or U5004 (N_5004,N_4273,N_4339);
nand U5005 (N_5005,N_4873,N_4686);
nand U5006 (N_5006,N_4801,N_4582);
nor U5007 (N_5007,N_4409,N_4604);
nand U5008 (N_5008,N_4244,N_4598);
nor U5009 (N_5009,N_4495,N_4275);
nor U5010 (N_5010,N_4204,N_4767);
xor U5011 (N_5011,N_4590,N_4892);
nor U5012 (N_5012,N_4084,N_4831);
nor U5013 (N_5013,N_4781,N_4913);
xor U5014 (N_5014,N_4836,N_4312);
and U5015 (N_5015,N_4743,N_4333);
xor U5016 (N_5016,N_4652,N_4923);
or U5017 (N_5017,N_4436,N_4370);
nor U5018 (N_5018,N_4944,N_4504);
and U5019 (N_5019,N_4295,N_4281);
nand U5020 (N_5020,N_4931,N_4797);
xor U5021 (N_5021,N_4092,N_4109);
and U5022 (N_5022,N_4262,N_4565);
nand U5023 (N_5023,N_4145,N_4950);
or U5024 (N_5024,N_4734,N_4747);
xnor U5025 (N_5025,N_4525,N_4406);
and U5026 (N_5026,N_4815,N_4830);
nor U5027 (N_5027,N_4825,N_4167);
and U5028 (N_5028,N_4940,N_4818);
or U5029 (N_5029,N_4803,N_4443);
and U5030 (N_5030,N_4776,N_4459);
or U5031 (N_5031,N_4354,N_4570);
or U5032 (N_5032,N_4435,N_4659);
or U5033 (N_5033,N_4680,N_4041);
nand U5034 (N_5034,N_4143,N_4912);
nand U5035 (N_5035,N_4543,N_4507);
or U5036 (N_5036,N_4728,N_4720);
nand U5037 (N_5037,N_4121,N_4695);
nand U5038 (N_5038,N_4186,N_4454);
or U5039 (N_5039,N_4025,N_4744);
or U5040 (N_5040,N_4179,N_4226);
nor U5041 (N_5041,N_4019,N_4497);
xnor U5042 (N_5042,N_4501,N_4661);
or U5043 (N_5043,N_4424,N_4534);
and U5044 (N_5044,N_4717,N_4641);
nor U5045 (N_5045,N_4033,N_4420);
xor U5046 (N_5046,N_4779,N_4160);
xnor U5047 (N_5047,N_4144,N_4919);
and U5048 (N_5048,N_4219,N_4045);
xnor U5049 (N_5049,N_4673,N_4391);
nand U5050 (N_5050,N_4172,N_4897);
nor U5051 (N_5051,N_4692,N_4231);
nor U5052 (N_5052,N_4955,N_4533);
xnor U5053 (N_5053,N_4136,N_4889);
and U5054 (N_5054,N_4321,N_4489);
and U5055 (N_5055,N_4289,N_4702);
or U5056 (N_5056,N_4948,N_4899);
nand U5057 (N_5057,N_4957,N_4483);
nand U5058 (N_5058,N_4412,N_4643);
nand U5059 (N_5059,N_4970,N_4085);
and U5060 (N_5060,N_4866,N_4098);
and U5061 (N_5061,N_4705,N_4097);
and U5062 (N_5062,N_4065,N_4294);
nor U5063 (N_5063,N_4183,N_4434);
nand U5064 (N_5064,N_4515,N_4153);
nand U5065 (N_5065,N_4539,N_4920);
or U5066 (N_5066,N_4987,N_4693);
nand U5067 (N_5067,N_4263,N_4319);
xor U5068 (N_5068,N_4168,N_4799);
nand U5069 (N_5069,N_4625,N_4173);
nand U5070 (N_5070,N_4928,N_4672);
xnor U5071 (N_5071,N_4649,N_4017);
nor U5072 (N_5072,N_4117,N_4917);
xor U5073 (N_5073,N_4959,N_4701);
or U5074 (N_5074,N_4184,N_4079);
and U5075 (N_5075,N_4812,N_4318);
nor U5076 (N_5076,N_4552,N_4845);
and U5077 (N_5077,N_4934,N_4675);
nor U5078 (N_5078,N_4764,N_4556);
nand U5079 (N_5079,N_4574,N_4983);
nand U5080 (N_5080,N_4973,N_4522);
or U5081 (N_5081,N_4827,N_4795);
nand U5082 (N_5082,N_4239,N_4510);
and U5083 (N_5083,N_4069,N_4133);
and U5084 (N_5084,N_4207,N_4667);
or U5085 (N_5085,N_4629,N_4320);
nor U5086 (N_5086,N_4607,N_4031);
nand U5087 (N_5087,N_4954,N_4621);
xor U5088 (N_5088,N_4765,N_4698);
nor U5089 (N_5089,N_4502,N_4660);
xnor U5090 (N_5090,N_4199,N_4224);
nand U5091 (N_5091,N_4044,N_4740);
xor U5092 (N_5092,N_4202,N_4964);
nor U5093 (N_5093,N_4030,N_4300);
or U5094 (N_5094,N_4494,N_4834);
nand U5095 (N_5095,N_4829,N_4863);
and U5096 (N_5096,N_4596,N_4938);
nand U5097 (N_5097,N_4915,N_4428);
nor U5098 (N_5098,N_4786,N_4580);
and U5099 (N_5099,N_4373,N_4372);
nor U5100 (N_5100,N_4439,N_4241);
nor U5101 (N_5101,N_4430,N_4392);
nand U5102 (N_5102,N_4427,N_4056);
nor U5103 (N_5103,N_4936,N_4345);
nand U5104 (N_5104,N_4111,N_4557);
xor U5105 (N_5105,N_4689,N_4042);
and U5106 (N_5106,N_4324,N_4684);
or U5107 (N_5107,N_4415,N_4127);
nand U5108 (N_5108,N_4004,N_4894);
nand U5109 (N_5109,N_4448,N_4752);
or U5110 (N_5110,N_4176,N_4194);
nor U5111 (N_5111,N_4662,N_4218);
nand U5112 (N_5112,N_4737,N_4826);
and U5113 (N_5113,N_4368,N_4909);
or U5114 (N_5114,N_4986,N_4389);
nand U5115 (N_5115,N_4791,N_4178);
and U5116 (N_5116,N_4385,N_4648);
nor U5117 (N_5117,N_4956,N_4891);
or U5118 (N_5118,N_4146,N_4837);
xor U5119 (N_5119,N_4361,N_4225);
xnor U5120 (N_5120,N_4542,N_4843);
nand U5121 (N_5121,N_4518,N_4256);
nor U5122 (N_5122,N_4364,N_4792);
or U5123 (N_5123,N_4282,N_4335);
nand U5124 (N_5124,N_4161,N_4022);
nand U5125 (N_5125,N_4418,N_4212);
nor U5126 (N_5126,N_4935,N_4141);
nand U5127 (N_5127,N_4992,N_4119);
or U5128 (N_5128,N_4278,N_4969);
nand U5129 (N_5129,N_4887,N_4575);
and U5130 (N_5130,N_4960,N_4038);
xnor U5131 (N_5131,N_4293,N_4709);
and U5132 (N_5132,N_4578,N_4358);
nand U5133 (N_5133,N_4441,N_4214);
nand U5134 (N_5134,N_4187,N_4614);
or U5135 (N_5135,N_4835,N_4820);
nor U5136 (N_5136,N_4733,N_4620);
or U5137 (N_5137,N_4139,N_4669);
nor U5138 (N_5138,N_4794,N_4157);
and U5139 (N_5139,N_4024,N_4601);
nand U5140 (N_5140,N_4402,N_4375);
nand U5141 (N_5141,N_4298,N_4793);
or U5142 (N_5142,N_4156,N_4859);
nand U5143 (N_5143,N_4591,N_4057);
or U5144 (N_5144,N_4087,N_4841);
or U5145 (N_5145,N_4589,N_4035);
or U5146 (N_5146,N_4393,N_4636);
nand U5147 (N_5147,N_4433,N_4061);
or U5148 (N_5148,N_4266,N_4325);
and U5149 (N_5149,N_4624,N_4788);
or U5150 (N_5150,N_4094,N_4639);
xor U5151 (N_5151,N_4399,N_4381);
nand U5152 (N_5152,N_4164,N_4129);
or U5153 (N_5153,N_4509,N_4585);
xnor U5154 (N_5154,N_4777,N_4376);
xnor U5155 (N_5155,N_4817,N_4857);
and U5156 (N_5156,N_4754,N_4713);
or U5157 (N_5157,N_4645,N_4076);
xnor U5158 (N_5158,N_4100,N_4880);
or U5159 (N_5159,N_4222,N_4088);
nand U5160 (N_5160,N_4491,N_4458);
or U5161 (N_5161,N_4126,N_4002);
xor U5162 (N_5162,N_4657,N_4751);
or U5163 (N_5163,N_4677,N_4271);
nor U5164 (N_5164,N_4310,N_4058);
or U5165 (N_5165,N_4559,N_4461);
nor U5166 (N_5166,N_4664,N_4150);
nor U5167 (N_5167,N_4537,N_4895);
and U5168 (N_5168,N_4425,N_4949);
xnor U5169 (N_5169,N_4650,N_4472);
nand U5170 (N_5170,N_4498,N_4592);
or U5171 (N_5171,N_4029,N_4758);
nor U5172 (N_5172,N_4584,N_4930);
xor U5173 (N_5173,N_4484,N_4807);
and U5174 (N_5174,N_4422,N_4229);
nand U5175 (N_5175,N_4520,N_4982);
and U5176 (N_5176,N_4452,N_4663);
and U5177 (N_5177,N_4579,N_4927);
or U5178 (N_5178,N_4074,N_4910);
xor U5179 (N_5179,N_4103,N_4798);
and U5180 (N_5180,N_4429,N_4622);
nor U5181 (N_5181,N_4216,N_4706);
and U5182 (N_5182,N_4488,N_4140);
and U5183 (N_5183,N_4438,N_4616);
nand U5184 (N_5184,N_4658,N_4419);
or U5185 (N_5185,N_4608,N_4309);
nand U5186 (N_5186,N_4196,N_4540);
xor U5187 (N_5187,N_4619,N_4359);
nor U5188 (N_5188,N_4450,N_4943);
or U5189 (N_5189,N_4993,N_4242);
nand U5190 (N_5190,N_4963,N_4095);
or U5191 (N_5191,N_4761,N_4277);
nand U5192 (N_5192,N_4444,N_4588);
or U5193 (N_5193,N_4729,N_4211);
nor U5194 (N_5194,N_4985,N_4260);
or U5195 (N_5195,N_4334,N_4130);
nor U5196 (N_5196,N_4205,N_4174);
nor U5197 (N_5197,N_4286,N_4383);
and U5198 (N_5198,N_4347,N_4678);
nor U5199 (N_5199,N_4162,N_4975);
xor U5200 (N_5200,N_4432,N_4503);
nand U5201 (N_5201,N_4978,N_4006);
or U5202 (N_5202,N_4043,N_4355);
or U5203 (N_5203,N_4081,N_4093);
xnor U5204 (N_5204,N_4916,N_4269);
or U5205 (N_5205,N_4267,N_4055);
nor U5206 (N_5206,N_4896,N_4426);
or U5207 (N_5207,N_4201,N_4314);
xor U5208 (N_5208,N_4464,N_4554);
xnor U5209 (N_5209,N_4685,N_4340);
nand U5210 (N_5210,N_4462,N_4280);
nand U5211 (N_5211,N_4423,N_4351);
nor U5212 (N_5212,N_4431,N_4809);
nor U5213 (N_5213,N_4165,N_4228);
and U5214 (N_5214,N_4555,N_4971);
nand U5215 (N_5215,N_4617,N_4569);
and U5216 (N_5216,N_4465,N_4305);
or U5217 (N_5217,N_4387,N_4154);
and U5218 (N_5218,N_4250,N_4341);
or U5219 (N_5219,N_4769,N_4731);
or U5220 (N_5220,N_4152,N_4220);
or U5221 (N_5221,N_4724,N_4470);
and U5222 (N_5222,N_4466,N_4530);
nor U5223 (N_5223,N_4384,N_4989);
and U5224 (N_5224,N_4463,N_4716);
and U5225 (N_5225,N_4099,N_4711);
xnor U5226 (N_5226,N_4247,N_4775);
or U5227 (N_5227,N_4182,N_4712);
nor U5228 (N_5228,N_4929,N_4846);
and U5229 (N_5229,N_4925,N_4191);
nor U5230 (N_5230,N_4704,N_4203);
and U5231 (N_5231,N_4521,N_4493);
or U5232 (N_5232,N_4922,N_4632);
xnor U5233 (N_5233,N_4886,N_4638);
nor U5234 (N_5234,N_4666,N_4064);
or U5235 (N_5235,N_4356,N_4599);
nand U5236 (N_5236,N_4404,N_4301);
or U5237 (N_5237,N_4148,N_4135);
nand U5238 (N_5238,N_4288,N_4519);
or U5239 (N_5239,N_4805,N_4911);
and U5240 (N_5240,N_4481,N_4067);
nand U5241 (N_5241,N_4311,N_4732);
nor U5242 (N_5242,N_4471,N_4457);
nor U5243 (N_5243,N_4445,N_4511);
xor U5244 (N_5244,N_4597,N_4933);
nor U5245 (N_5245,N_4332,N_4968);
or U5246 (N_5246,N_4040,N_4115);
and U5247 (N_5247,N_4068,N_4122);
nor U5248 (N_5248,N_4655,N_4166);
or U5249 (N_5249,N_4603,N_4535);
xor U5250 (N_5250,N_4486,N_4197);
and U5251 (N_5251,N_4369,N_4362);
nor U5252 (N_5252,N_4773,N_4583);
or U5253 (N_5253,N_4958,N_4531);
nand U5254 (N_5254,N_4814,N_4742);
nor U5255 (N_5255,N_4871,N_4527);
or U5256 (N_5256,N_4550,N_4114);
nand U5257 (N_5257,N_4644,N_4746);
and U5258 (N_5258,N_4901,N_4396);
nor U5259 (N_5259,N_4721,N_4903);
and U5260 (N_5260,N_4110,N_4366);
nor U5261 (N_5261,N_4772,N_4234);
and U5262 (N_5262,N_4487,N_4646);
or U5263 (N_5263,N_4352,N_4342);
nor U5264 (N_5264,N_4046,N_4524);
nand U5265 (N_5265,N_4236,N_4855);
nand U5266 (N_5266,N_4051,N_4240);
nor U5267 (N_5267,N_4177,N_4086);
or U5268 (N_5268,N_4408,N_4175);
or U5269 (N_5269,N_4651,N_4905);
xor U5270 (N_5270,N_4755,N_4566);
nand U5271 (N_5271,N_4365,N_4181);
and U5272 (N_5272,N_4823,N_4215);
nor U5273 (N_5273,N_4995,N_4888);
nor U5274 (N_5274,N_4749,N_4979);
or U5275 (N_5275,N_4882,N_4163);
nand U5276 (N_5276,N_4039,N_4326);
or U5277 (N_5277,N_4138,N_4821);
nor U5278 (N_5278,N_4453,N_4102);
nand U5279 (N_5279,N_4008,N_4800);
and U5280 (N_5280,N_4101,N_4832);
nand U5281 (N_5281,N_4485,N_4852);
and U5282 (N_5282,N_4571,N_4237);
nor U5283 (N_5283,N_4548,N_4842);
nor U5284 (N_5284,N_4654,N_4467);
nor U5285 (N_5285,N_4839,N_4516);
and U5286 (N_5286,N_4595,N_4208);
nor U5287 (N_5287,N_4386,N_4316);
nor U5288 (N_5288,N_4499,N_4473);
nor U5289 (N_5289,N_4049,N_4123);
nor U5290 (N_5290,N_4806,N_4718);
and U5291 (N_5291,N_4627,N_4193);
nor U5292 (N_5292,N_4082,N_4676);
and U5293 (N_5293,N_4926,N_4546);
nor U5294 (N_5294,N_4151,N_4900);
nand U5295 (N_5295,N_4508,N_4131);
or U5296 (N_5296,N_4988,N_4885);
nor U5297 (N_5297,N_4070,N_4346);
nor U5298 (N_5298,N_4563,N_4254);
nor U5299 (N_5299,N_4991,N_4587);
xnor U5300 (N_5300,N_4967,N_4190);
and U5301 (N_5301,N_4159,N_4750);
or U5302 (N_5302,N_4034,N_4544);
nand U5303 (N_5303,N_4116,N_4052);
and U5304 (N_5304,N_4395,N_4517);
nand U5305 (N_5305,N_4020,N_4016);
nor U5306 (N_5306,N_4884,N_4822);
nor U5307 (N_5307,N_4343,N_4577);
xnor U5308 (N_5308,N_4653,N_4252);
and U5309 (N_5309,N_4877,N_4059);
xnor U5310 (N_5310,N_4628,N_4865);
nand U5311 (N_5311,N_4864,N_4403);
or U5312 (N_5312,N_4071,N_4405);
and U5313 (N_5313,N_4715,N_4108);
nand U5314 (N_5314,N_4671,N_4562);
nand U5315 (N_5315,N_4753,N_4748);
nor U5316 (N_5316,N_4736,N_4500);
and U5317 (N_5317,N_4075,N_4966);
or U5318 (N_5318,N_4407,N_4953);
nand U5319 (N_5319,N_4918,N_4951);
and U5320 (N_5320,N_4394,N_4694);
nor U5321 (N_5321,N_4290,N_4687);
nand U5322 (N_5322,N_4819,N_4490);
or U5323 (N_5323,N_4688,N_4072);
nor U5324 (N_5324,N_4626,N_4907);
or U5325 (N_5325,N_4937,N_4532);
nand U5326 (N_5326,N_4411,N_4854);
or U5327 (N_5327,N_4810,N_4947);
and U5328 (N_5328,N_4482,N_4875);
and U5329 (N_5329,N_4681,N_4447);
and U5330 (N_5330,N_4506,N_4840);
nor U5331 (N_5331,N_4784,N_4440);
nor U5332 (N_5332,N_4914,N_4185);
and U5333 (N_5333,N_4344,N_4613);
and U5334 (N_5334,N_4939,N_4703);
xor U5335 (N_5335,N_4990,N_4719);
nand U5336 (N_5336,N_4248,N_4107);
nor U5337 (N_5337,N_4379,N_4328);
nor U5338 (N_5338,N_4763,N_4670);
nand U5339 (N_5339,N_4745,N_4551);
and U5340 (N_5340,N_4856,N_4633);
and U5341 (N_5341,N_4813,N_4780);
or U5342 (N_5342,N_4270,N_4999);
nor U5343 (N_5343,N_4155,N_4353);
nand U5344 (N_5344,N_4195,N_4634);
or U5345 (N_5345,N_4259,N_4106);
nor U5346 (N_5346,N_4083,N_4390);
nand U5347 (N_5347,N_4924,N_4421);
nor U5348 (N_5348,N_4526,N_4981);
xnor U5349 (N_5349,N_4512,N_4547);
or U5350 (N_5350,N_4089,N_4018);
nand U5351 (N_5351,N_4848,N_4665);
and U5352 (N_5352,N_4505,N_4572);
and U5353 (N_5353,N_4861,N_4460);
and U5354 (N_5354,N_4066,N_4946);
nand U5355 (N_5355,N_4125,N_4050);
or U5356 (N_5356,N_4456,N_4233);
nand U5357 (N_5357,N_4860,N_4630);
xnor U5358 (N_5358,N_4330,N_4388);
or U5359 (N_5359,N_4299,N_4850);
nand U5360 (N_5360,N_4513,N_4398);
nor U5361 (N_5361,N_4210,N_4442);
or U5362 (N_5362,N_4477,N_4009);
and U5363 (N_5363,N_4774,N_4170);
nand U5364 (N_5364,N_4881,N_4446);
and U5365 (N_5365,N_4054,N_4974);
or U5366 (N_5366,N_4400,N_4378);
nand U5367 (N_5367,N_4682,N_4028);
or U5368 (N_5368,N_4158,N_4610);
or U5369 (N_5369,N_4357,N_4545);
nand U5370 (N_5370,N_4576,N_4245);
or U5371 (N_5371,N_4553,N_4272);
nor U5372 (N_5372,N_4893,N_4707);
nand U5373 (N_5373,N_4833,N_4573);
xnor U5374 (N_5374,N_4246,N_4679);
and U5375 (N_5375,N_4479,N_4962);
nand U5376 (N_5376,N_4735,N_4104);
or U5377 (N_5377,N_4708,N_4036);
or U5378 (N_5378,N_4206,N_4062);
xor U5379 (N_5379,N_4249,N_4605);
nor U5380 (N_5380,N_4437,N_4722);
nor U5381 (N_5381,N_4015,N_4455);
xnor U5382 (N_5382,N_4528,N_4238);
and U5383 (N_5383,N_4331,N_4862);
nor U5384 (N_5384,N_4091,N_4696);
and U5385 (N_5385,N_4476,N_4642);
or U5386 (N_5386,N_4714,N_4315);
and U5387 (N_5387,N_4984,N_4451);
nand U5388 (N_5388,N_4232,N_4327);
and U5389 (N_5389,N_4869,N_4010);
xnor U5390 (N_5390,N_4243,N_4802);
and U5391 (N_5391,N_4380,N_4996);
and U5392 (N_5392,N_4416,N_4700);
and U5393 (N_5393,N_4053,N_4902);
and U5394 (N_5394,N_4149,N_4623);
or U5395 (N_5395,N_4611,N_4741);
or U5396 (N_5396,N_4338,N_4297);
or U5397 (N_5397,N_4759,N_4618);
or U5398 (N_5398,N_4377,N_4292);
xor U5399 (N_5399,N_4561,N_4096);
or U5400 (N_5400,N_4189,N_4307);
and U5401 (N_5401,N_4268,N_4198);
and U5402 (N_5402,N_4105,N_4048);
and U5403 (N_5403,N_4770,N_4235);
nor U5404 (N_5404,N_4783,N_4258);
xnor U5405 (N_5405,N_4014,N_4756);
xnor U5406 (N_5406,N_4980,N_4112);
and U5407 (N_5407,N_4007,N_4602);
nand U5408 (N_5408,N_4874,N_4027);
and U5409 (N_5409,N_4337,N_4323);
or U5410 (N_5410,N_4538,N_4171);
nor U5411 (N_5411,N_4348,N_4253);
xor U5412 (N_5412,N_4192,N_4941);
nand U5413 (N_5413,N_4001,N_4615);
and U5414 (N_5414,N_4997,N_4047);
nor U5415 (N_5415,N_4230,N_4858);
and U5416 (N_5416,N_4853,N_4594);
xor U5417 (N_5417,N_4942,N_4213);
nand U5418 (N_5418,N_4011,N_4593);
nor U5419 (N_5419,N_4492,N_4363);
nand U5420 (N_5420,N_4549,N_4514);
and U5421 (N_5421,N_4080,N_4142);
nor U5422 (N_5422,N_4291,N_4828);
or U5423 (N_5423,N_4000,N_4762);
nor U5424 (N_5424,N_4609,N_4303);
or U5425 (N_5425,N_4257,N_4564);
nor U5426 (N_5426,N_4137,N_4322);
and U5427 (N_5427,N_4876,N_4870);
or U5428 (N_5428,N_4690,N_4872);
nand U5429 (N_5429,N_4804,N_4200);
and U5430 (N_5430,N_4283,N_4284);
or U5431 (N_5431,N_4349,N_4906);
nor U5432 (N_5432,N_4306,N_4413);
nor U5433 (N_5433,N_4581,N_4723);
xor U5434 (N_5434,N_4710,N_4904);
or U5435 (N_5435,N_4849,N_4032);
or U5436 (N_5436,N_4945,N_4132);
nand U5437 (N_5437,N_4128,N_4401);
nor U5438 (N_5438,N_4739,N_4026);
and U5439 (N_5439,N_4134,N_4113);
or U5440 (N_5440,N_4118,N_4668);
nor U5441 (N_5441,N_4478,N_4414);
and U5442 (N_5442,N_4635,N_4077);
xor U5443 (N_5443,N_4188,N_4560);
nor U5444 (N_5444,N_4255,N_4867);
xnor U5445 (N_5445,N_4060,N_4037);
nor U5446 (N_5446,N_4612,N_4790);
and U5447 (N_5447,N_4785,N_4725);
nor U5448 (N_5448,N_4816,N_4012);
and U5449 (N_5449,N_4367,N_4568);
or U5450 (N_5450,N_4013,N_4757);
nor U5451 (N_5451,N_4371,N_4285);
nand U5452 (N_5452,N_4374,N_4217);
and U5453 (N_5453,N_4782,N_4647);
xnor U5454 (N_5454,N_4023,N_4878);
or U5455 (N_5455,N_4417,N_4656);
nand U5456 (N_5456,N_4586,N_4265);
nor U5457 (N_5457,N_4223,N_4844);
or U5458 (N_5458,N_4276,N_4449);
nand U5459 (N_5459,N_4637,N_4683);
and U5460 (N_5460,N_4063,N_4261);
nand U5461 (N_5461,N_4078,N_4169);
and U5462 (N_5462,N_4691,N_4811);
xor U5463 (N_5463,N_4496,N_4961);
xnor U5464 (N_5464,N_4965,N_4868);
and U5465 (N_5465,N_4977,N_4541);
nor U5466 (N_5466,N_4697,N_4766);
xor U5467 (N_5467,N_4536,N_4274);
or U5468 (N_5468,N_4475,N_4336);
nor U5469 (N_5469,N_4808,N_4279);
nand U5470 (N_5470,N_4124,N_4005);
and U5471 (N_5471,N_4302,N_4738);
and U5472 (N_5472,N_4787,N_4640);
xor U5473 (N_5473,N_4824,N_4890);
nand U5474 (N_5474,N_4567,N_4469);
or U5475 (N_5475,N_4468,N_4529);
and U5476 (N_5476,N_4264,N_4908);
or U5477 (N_5477,N_4120,N_4480);
nor U5478 (N_5478,N_4350,N_4523);
nand U5479 (N_5479,N_4606,N_4221);
nand U5480 (N_5480,N_4313,N_4768);
nor U5481 (N_5481,N_4021,N_4994);
xor U5482 (N_5482,N_4251,N_4730);
nand U5483 (N_5483,N_4921,N_4296);
and U5484 (N_5484,N_4329,N_4147);
nor U5485 (N_5485,N_4631,N_4972);
or U5486 (N_5486,N_4287,N_4090);
nand U5487 (N_5487,N_4883,N_4898);
nand U5488 (N_5488,N_4796,N_4699);
nand U5489 (N_5489,N_4998,N_4976);
and U5490 (N_5490,N_4726,N_4847);
nand U5491 (N_5491,N_4410,N_4474);
or U5492 (N_5492,N_4209,N_4932);
nand U5493 (N_5493,N_4879,N_4789);
or U5494 (N_5494,N_4760,N_4600);
and U5495 (N_5495,N_4360,N_4304);
and U5496 (N_5496,N_4778,N_4003);
or U5497 (N_5497,N_4073,N_4308);
nor U5498 (N_5498,N_4558,N_4851);
nand U5499 (N_5499,N_4180,N_4952);
and U5500 (N_5500,N_4135,N_4639);
nand U5501 (N_5501,N_4953,N_4195);
nor U5502 (N_5502,N_4033,N_4120);
nor U5503 (N_5503,N_4945,N_4193);
nand U5504 (N_5504,N_4795,N_4488);
and U5505 (N_5505,N_4682,N_4837);
nor U5506 (N_5506,N_4862,N_4355);
xor U5507 (N_5507,N_4048,N_4827);
nand U5508 (N_5508,N_4439,N_4714);
and U5509 (N_5509,N_4046,N_4105);
or U5510 (N_5510,N_4327,N_4007);
nand U5511 (N_5511,N_4096,N_4685);
or U5512 (N_5512,N_4726,N_4478);
and U5513 (N_5513,N_4982,N_4918);
or U5514 (N_5514,N_4149,N_4110);
xor U5515 (N_5515,N_4013,N_4096);
nor U5516 (N_5516,N_4722,N_4658);
nor U5517 (N_5517,N_4831,N_4254);
and U5518 (N_5518,N_4691,N_4237);
nand U5519 (N_5519,N_4189,N_4798);
xnor U5520 (N_5520,N_4988,N_4870);
nand U5521 (N_5521,N_4778,N_4898);
or U5522 (N_5522,N_4622,N_4165);
nor U5523 (N_5523,N_4245,N_4238);
xor U5524 (N_5524,N_4856,N_4138);
xnor U5525 (N_5525,N_4405,N_4978);
nand U5526 (N_5526,N_4677,N_4207);
or U5527 (N_5527,N_4067,N_4144);
nand U5528 (N_5528,N_4174,N_4248);
nor U5529 (N_5529,N_4076,N_4380);
and U5530 (N_5530,N_4509,N_4855);
or U5531 (N_5531,N_4255,N_4631);
and U5532 (N_5532,N_4292,N_4058);
and U5533 (N_5533,N_4945,N_4482);
nand U5534 (N_5534,N_4696,N_4936);
nor U5535 (N_5535,N_4015,N_4195);
or U5536 (N_5536,N_4781,N_4982);
nand U5537 (N_5537,N_4350,N_4682);
and U5538 (N_5538,N_4680,N_4301);
nand U5539 (N_5539,N_4796,N_4025);
and U5540 (N_5540,N_4816,N_4159);
or U5541 (N_5541,N_4442,N_4634);
nor U5542 (N_5542,N_4858,N_4220);
or U5543 (N_5543,N_4056,N_4863);
and U5544 (N_5544,N_4498,N_4082);
nand U5545 (N_5545,N_4510,N_4467);
nor U5546 (N_5546,N_4930,N_4088);
or U5547 (N_5547,N_4973,N_4376);
nand U5548 (N_5548,N_4036,N_4744);
nor U5549 (N_5549,N_4741,N_4801);
nor U5550 (N_5550,N_4083,N_4867);
nand U5551 (N_5551,N_4925,N_4883);
and U5552 (N_5552,N_4192,N_4665);
nand U5553 (N_5553,N_4122,N_4694);
or U5554 (N_5554,N_4093,N_4348);
or U5555 (N_5555,N_4493,N_4149);
or U5556 (N_5556,N_4805,N_4328);
and U5557 (N_5557,N_4837,N_4024);
or U5558 (N_5558,N_4135,N_4701);
nand U5559 (N_5559,N_4647,N_4572);
or U5560 (N_5560,N_4058,N_4035);
nand U5561 (N_5561,N_4799,N_4640);
nor U5562 (N_5562,N_4733,N_4308);
nor U5563 (N_5563,N_4828,N_4073);
or U5564 (N_5564,N_4656,N_4594);
nand U5565 (N_5565,N_4678,N_4284);
nand U5566 (N_5566,N_4252,N_4330);
nand U5567 (N_5567,N_4211,N_4308);
and U5568 (N_5568,N_4772,N_4082);
nand U5569 (N_5569,N_4020,N_4445);
nand U5570 (N_5570,N_4996,N_4382);
and U5571 (N_5571,N_4824,N_4071);
and U5572 (N_5572,N_4623,N_4341);
and U5573 (N_5573,N_4131,N_4622);
nor U5574 (N_5574,N_4023,N_4283);
xnor U5575 (N_5575,N_4840,N_4492);
and U5576 (N_5576,N_4445,N_4621);
nand U5577 (N_5577,N_4247,N_4086);
xor U5578 (N_5578,N_4114,N_4320);
xor U5579 (N_5579,N_4219,N_4592);
nor U5580 (N_5580,N_4583,N_4687);
nor U5581 (N_5581,N_4729,N_4045);
nor U5582 (N_5582,N_4168,N_4134);
nor U5583 (N_5583,N_4533,N_4558);
or U5584 (N_5584,N_4439,N_4863);
and U5585 (N_5585,N_4580,N_4546);
or U5586 (N_5586,N_4239,N_4664);
nor U5587 (N_5587,N_4264,N_4452);
nand U5588 (N_5588,N_4655,N_4505);
nand U5589 (N_5589,N_4633,N_4363);
and U5590 (N_5590,N_4278,N_4237);
or U5591 (N_5591,N_4933,N_4342);
xnor U5592 (N_5592,N_4799,N_4873);
or U5593 (N_5593,N_4282,N_4292);
nor U5594 (N_5594,N_4723,N_4625);
nand U5595 (N_5595,N_4944,N_4176);
nand U5596 (N_5596,N_4615,N_4100);
nand U5597 (N_5597,N_4008,N_4058);
and U5598 (N_5598,N_4753,N_4678);
or U5599 (N_5599,N_4496,N_4678);
or U5600 (N_5600,N_4270,N_4475);
nand U5601 (N_5601,N_4063,N_4239);
nor U5602 (N_5602,N_4951,N_4489);
nor U5603 (N_5603,N_4306,N_4327);
or U5604 (N_5604,N_4302,N_4823);
nor U5605 (N_5605,N_4375,N_4841);
or U5606 (N_5606,N_4436,N_4076);
or U5607 (N_5607,N_4747,N_4468);
nand U5608 (N_5608,N_4069,N_4086);
or U5609 (N_5609,N_4384,N_4034);
nor U5610 (N_5610,N_4142,N_4228);
nand U5611 (N_5611,N_4197,N_4618);
and U5612 (N_5612,N_4007,N_4181);
or U5613 (N_5613,N_4227,N_4130);
nand U5614 (N_5614,N_4255,N_4871);
or U5615 (N_5615,N_4310,N_4143);
or U5616 (N_5616,N_4873,N_4403);
nand U5617 (N_5617,N_4080,N_4832);
or U5618 (N_5618,N_4770,N_4557);
or U5619 (N_5619,N_4501,N_4258);
or U5620 (N_5620,N_4708,N_4820);
xor U5621 (N_5621,N_4463,N_4340);
nand U5622 (N_5622,N_4075,N_4106);
nand U5623 (N_5623,N_4446,N_4663);
and U5624 (N_5624,N_4959,N_4180);
and U5625 (N_5625,N_4249,N_4282);
nand U5626 (N_5626,N_4160,N_4198);
nand U5627 (N_5627,N_4806,N_4693);
nor U5628 (N_5628,N_4454,N_4792);
and U5629 (N_5629,N_4265,N_4522);
nor U5630 (N_5630,N_4845,N_4623);
nand U5631 (N_5631,N_4647,N_4759);
nand U5632 (N_5632,N_4489,N_4065);
or U5633 (N_5633,N_4584,N_4508);
nand U5634 (N_5634,N_4482,N_4189);
and U5635 (N_5635,N_4822,N_4289);
nor U5636 (N_5636,N_4471,N_4018);
and U5637 (N_5637,N_4355,N_4170);
nor U5638 (N_5638,N_4445,N_4282);
or U5639 (N_5639,N_4872,N_4693);
nand U5640 (N_5640,N_4301,N_4944);
nand U5641 (N_5641,N_4067,N_4567);
and U5642 (N_5642,N_4785,N_4185);
and U5643 (N_5643,N_4780,N_4231);
and U5644 (N_5644,N_4043,N_4258);
nor U5645 (N_5645,N_4184,N_4344);
nor U5646 (N_5646,N_4284,N_4797);
or U5647 (N_5647,N_4957,N_4586);
and U5648 (N_5648,N_4145,N_4401);
or U5649 (N_5649,N_4514,N_4327);
and U5650 (N_5650,N_4468,N_4202);
nand U5651 (N_5651,N_4674,N_4610);
and U5652 (N_5652,N_4393,N_4705);
nand U5653 (N_5653,N_4220,N_4579);
or U5654 (N_5654,N_4838,N_4994);
or U5655 (N_5655,N_4554,N_4168);
and U5656 (N_5656,N_4998,N_4540);
nand U5657 (N_5657,N_4422,N_4144);
nand U5658 (N_5658,N_4805,N_4244);
nand U5659 (N_5659,N_4557,N_4029);
xnor U5660 (N_5660,N_4038,N_4465);
xor U5661 (N_5661,N_4330,N_4391);
or U5662 (N_5662,N_4863,N_4303);
and U5663 (N_5663,N_4251,N_4785);
nor U5664 (N_5664,N_4991,N_4486);
or U5665 (N_5665,N_4839,N_4370);
nand U5666 (N_5666,N_4791,N_4748);
and U5667 (N_5667,N_4575,N_4585);
and U5668 (N_5668,N_4713,N_4976);
or U5669 (N_5669,N_4399,N_4036);
xnor U5670 (N_5670,N_4792,N_4439);
nand U5671 (N_5671,N_4884,N_4593);
or U5672 (N_5672,N_4205,N_4414);
xnor U5673 (N_5673,N_4311,N_4868);
and U5674 (N_5674,N_4866,N_4892);
nand U5675 (N_5675,N_4375,N_4753);
or U5676 (N_5676,N_4628,N_4487);
nand U5677 (N_5677,N_4368,N_4421);
nor U5678 (N_5678,N_4658,N_4831);
and U5679 (N_5679,N_4195,N_4772);
or U5680 (N_5680,N_4834,N_4608);
nand U5681 (N_5681,N_4502,N_4118);
and U5682 (N_5682,N_4934,N_4988);
or U5683 (N_5683,N_4212,N_4723);
and U5684 (N_5684,N_4646,N_4951);
and U5685 (N_5685,N_4644,N_4496);
nor U5686 (N_5686,N_4130,N_4404);
nand U5687 (N_5687,N_4081,N_4131);
and U5688 (N_5688,N_4335,N_4919);
nand U5689 (N_5689,N_4397,N_4175);
and U5690 (N_5690,N_4846,N_4346);
nand U5691 (N_5691,N_4964,N_4819);
nand U5692 (N_5692,N_4628,N_4046);
nand U5693 (N_5693,N_4438,N_4620);
and U5694 (N_5694,N_4834,N_4261);
or U5695 (N_5695,N_4649,N_4248);
nor U5696 (N_5696,N_4632,N_4234);
or U5697 (N_5697,N_4286,N_4061);
or U5698 (N_5698,N_4158,N_4836);
and U5699 (N_5699,N_4626,N_4800);
or U5700 (N_5700,N_4500,N_4715);
nand U5701 (N_5701,N_4309,N_4636);
or U5702 (N_5702,N_4173,N_4416);
or U5703 (N_5703,N_4421,N_4073);
and U5704 (N_5704,N_4910,N_4983);
xnor U5705 (N_5705,N_4136,N_4251);
nand U5706 (N_5706,N_4276,N_4495);
or U5707 (N_5707,N_4089,N_4016);
or U5708 (N_5708,N_4954,N_4720);
nand U5709 (N_5709,N_4073,N_4948);
and U5710 (N_5710,N_4697,N_4091);
or U5711 (N_5711,N_4444,N_4594);
nor U5712 (N_5712,N_4574,N_4099);
xor U5713 (N_5713,N_4221,N_4675);
xor U5714 (N_5714,N_4737,N_4386);
nand U5715 (N_5715,N_4852,N_4787);
or U5716 (N_5716,N_4425,N_4940);
and U5717 (N_5717,N_4119,N_4762);
or U5718 (N_5718,N_4871,N_4463);
and U5719 (N_5719,N_4332,N_4660);
xnor U5720 (N_5720,N_4410,N_4073);
xnor U5721 (N_5721,N_4354,N_4187);
nand U5722 (N_5722,N_4623,N_4376);
nor U5723 (N_5723,N_4547,N_4424);
nor U5724 (N_5724,N_4093,N_4560);
nand U5725 (N_5725,N_4181,N_4260);
nor U5726 (N_5726,N_4041,N_4132);
nand U5727 (N_5727,N_4946,N_4415);
or U5728 (N_5728,N_4572,N_4691);
or U5729 (N_5729,N_4989,N_4884);
and U5730 (N_5730,N_4576,N_4677);
and U5731 (N_5731,N_4819,N_4546);
nand U5732 (N_5732,N_4514,N_4624);
and U5733 (N_5733,N_4562,N_4893);
and U5734 (N_5734,N_4933,N_4375);
xnor U5735 (N_5735,N_4659,N_4393);
and U5736 (N_5736,N_4116,N_4794);
nand U5737 (N_5737,N_4232,N_4009);
nor U5738 (N_5738,N_4113,N_4893);
or U5739 (N_5739,N_4154,N_4184);
or U5740 (N_5740,N_4196,N_4976);
or U5741 (N_5741,N_4713,N_4235);
and U5742 (N_5742,N_4932,N_4114);
and U5743 (N_5743,N_4938,N_4731);
nor U5744 (N_5744,N_4639,N_4173);
nand U5745 (N_5745,N_4520,N_4804);
nor U5746 (N_5746,N_4629,N_4375);
nor U5747 (N_5747,N_4608,N_4116);
xnor U5748 (N_5748,N_4898,N_4580);
and U5749 (N_5749,N_4322,N_4600);
nand U5750 (N_5750,N_4508,N_4596);
and U5751 (N_5751,N_4611,N_4972);
nand U5752 (N_5752,N_4974,N_4169);
nand U5753 (N_5753,N_4919,N_4707);
nor U5754 (N_5754,N_4160,N_4652);
or U5755 (N_5755,N_4689,N_4473);
nand U5756 (N_5756,N_4170,N_4414);
xor U5757 (N_5757,N_4399,N_4237);
nand U5758 (N_5758,N_4811,N_4746);
xnor U5759 (N_5759,N_4533,N_4484);
nor U5760 (N_5760,N_4499,N_4847);
or U5761 (N_5761,N_4900,N_4408);
and U5762 (N_5762,N_4193,N_4682);
nand U5763 (N_5763,N_4656,N_4351);
nor U5764 (N_5764,N_4711,N_4718);
xor U5765 (N_5765,N_4473,N_4750);
xor U5766 (N_5766,N_4913,N_4777);
and U5767 (N_5767,N_4313,N_4145);
and U5768 (N_5768,N_4016,N_4212);
or U5769 (N_5769,N_4272,N_4482);
nor U5770 (N_5770,N_4675,N_4716);
or U5771 (N_5771,N_4676,N_4559);
nand U5772 (N_5772,N_4904,N_4919);
nand U5773 (N_5773,N_4955,N_4192);
or U5774 (N_5774,N_4996,N_4704);
nand U5775 (N_5775,N_4077,N_4547);
and U5776 (N_5776,N_4561,N_4008);
nand U5777 (N_5777,N_4815,N_4077);
xor U5778 (N_5778,N_4956,N_4360);
and U5779 (N_5779,N_4653,N_4441);
nand U5780 (N_5780,N_4703,N_4043);
or U5781 (N_5781,N_4304,N_4185);
or U5782 (N_5782,N_4556,N_4660);
nand U5783 (N_5783,N_4112,N_4266);
nand U5784 (N_5784,N_4550,N_4597);
nor U5785 (N_5785,N_4710,N_4777);
nand U5786 (N_5786,N_4443,N_4753);
nor U5787 (N_5787,N_4413,N_4056);
xnor U5788 (N_5788,N_4121,N_4397);
nand U5789 (N_5789,N_4189,N_4089);
or U5790 (N_5790,N_4540,N_4954);
or U5791 (N_5791,N_4572,N_4863);
and U5792 (N_5792,N_4246,N_4187);
nand U5793 (N_5793,N_4464,N_4144);
xnor U5794 (N_5794,N_4455,N_4153);
and U5795 (N_5795,N_4430,N_4981);
nor U5796 (N_5796,N_4097,N_4833);
nand U5797 (N_5797,N_4649,N_4868);
nor U5798 (N_5798,N_4954,N_4021);
or U5799 (N_5799,N_4553,N_4588);
nor U5800 (N_5800,N_4924,N_4319);
nand U5801 (N_5801,N_4371,N_4752);
or U5802 (N_5802,N_4963,N_4808);
and U5803 (N_5803,N_4598,N_4709);
nor U5804 (N_5804,N_4716,N_4241);
and U5805 (N_5805,N_4586,N_4578);
nor U5806 (N_5806,N_4884,N_4328);
nor U5807 (N_5807,N_4925,N_4913);
xnor U5808 (N_5808,N_4349,N_4773);
xor U5809 (N_5809,N_4562,N_4822);
or U5810 (N_5810,N_4129,N_4481);
and U5811 (N_5811,N_4818,N_4880);
xnor U5812 (N_5812,N_4973,N_4716);
nor U5813 (N_5813,N_4325,N_4753);
nand U5814 (N_5814,N_4915,N_4744);
and U5815 (N_5815,N_4065,N_4897);
and U5816 (N_5816,N_4298,N_4838);
nor U5817 (N_5817,N_4987,N_4496);
nand U5818 (N_5818,N_4654,N_4195);
or U5819 (N_5819,N_4706,N_4522);
or U5820 (N_5820,N_4692,N_4180);
or U5821 (N_5821,N_4188,N_4296);
nor U5822 (N_5822,N_4651,N_4254);
and U5823 (N_5823,N_4195,N_4935);
nand U5824 (N_5824,N_4502,N_4125);
and U5825 (N_5825,N_4005,N_4617);
nand U5826 (N_5826,N_4712,N_4694);
and U5827 (N_5827,N_4004,N_4114);
nand U5828 (N_5828,N_4836,N_4336);
or U5829 (N_5829,N_4337,N_4373);
and U5830 (N_5830,N_4985,N_4299);
and U5831 (N_5831,N_4858,N_4825);
or U5832 (N_5832,N_4563,N_4435);
and U5833 (N_5833,N_4100,N_4498);
nor U5834 (N_5834,N_4636,N_4834);
nor U5835 (N_5835,N_4895,N_4942);
or U5836 (N_5836,N_4637,N_4461);
or U5837 (N_5837,N_4550,N_4191);
nor U5838 (N_5838,N_4530,N_4903);
or U5839 (N_5839,N_4843,N_4488);
nor U5840 (N_5840,N_4669,N_4413);
and U5841 (N_5841,N_4370,N_4754);
or U5842 (N_5842,N_4764,N_4813);
nor U5843 (N_5843,N_4921,N_4514);
or U5844 (N_5844,N_4817,N_4076);
nor U5845 (N_5845,N_4294,N_4828);
xor U5846 (N_5846,N_4027,N_4562);
or U5847 (N_5847,N_4826,N_4401);
or U5848 (N_5848,N_4368,N_4040);
nand U5849 (N_5849,N_4960,N_4954);
and U5850 (N_5850,N_4283,N_4628);
and U5851 (N_5851,N_4672,N_4762);
nand U5852 (N_5852,N_4620,N_4752);
or U5853 (N_5853,N_4396,N_4850);
nand U5854 (N_5854,N_4116,N_4300);
nor U5855 (N_5855,N_4527,N_4627);
nand U5856 (N_5856,N_4936,N_4186);
and U5857 (N_5857,N_4947,N_4631);
and U5858 (N_5858,N_4360,N_4993);
and U5859 (N_5859,N_4576,N_4250);
nand U5860 (N_5860,N_4697,N_4554);
nor U5861 (N_5861,N_4250,N_4235);
nand U5862 (N_5862,N_4127,N_4644);
and U5863 (N_5863,N_4906,N_4755);
nand U5864 (N_5864,N_4275,N_4824);
nor U5865 (N_5865,N_4285,N_4341);
nor U5866 (N_5866,N_4763,N_4752);
and U5867 (N_5867,N_4221,N_4238);
nand U5868 (N_5868,N_4342,N_4419);
and U5869 (N_5869,N_4010,N_4230);
nor U5870 (N_5870,N_4480,N_4136);
nand U5871 (N_5871,N_4618,N_4614);
or U5872 (N_5872,N_4492,N_4594);
and U5873 (N_5873,N_4421,N_4560);
nor U5874 (N_5874,N_4249,N_4079);
nand U5875 (N_5875,N_4474,N_4334);
nand U5876 (N_5876,N_4197,N_4660);
nor U5877 (N_5877,N_4443,N_4826);
and U5878 (N_5878,N_4978,N_4923);
or U5879 (N_5879,N_4642,N_4284);
and U5880 (N_5880,N_4426,N_4472);
or U5881 (N_5881,N_4330,N_4494);
nand U5882 (N_5882,N_4823,N_4538);
nand U5883 (N_5883,N_4773,N_4394);
nor U5884 (N_5884,N_4760,N_4316);
nor U5885 (N_5885,N_4260,N_4054);
or U5886 (N_5886,N_4615,N_4090);
and U5887 (N_5887,N_4831,N_4783);
and U5888 (N_5888,N_4031,N_4839);
nand U5889 (N_5889,N_4051,N_4388);
nor U5890 (N_5890,N_4614,N_4498);
xnor U5891 (N_5891,N_4546,N_4847);
nand U5892 (N_5892,N_4743,N_4250);
or U5893 (N_5893,N_4781,N_4224);
nand U5894 (N_5894,N_4403,N_4901);
nor U5895 (N_5895,N_4514,N_4871);
nand U5896 (N_5896,N_4942,N_4534);
and U5897 (N_5897,N_4293,N_4471);
nand U5898 (N_5898,N_4321,N_4064);
nor U5899 (N_5899,N_4823,N_4950);
nor U5900 (N_5900,N_4832,N_4601);
and U5901 (N_5901,N_4516,N_4193);
or U5902 (N_5902,N_4495,N_4349);
or U5903 (N_5903,N_4643,N_4907);
nand U5904 (N_5904,N_4300,N_4363);
nand U5905 (N_5905,N_4456,N_4585);
nand U5906 (N_5906,N_4995,N_4272);
nor U5907 (N_5907,N_4006,N_4716);
xnor U5908 (N_5908,N_4173,N_4965);
nor U5909 (N_5909,N_4669,N_4997);
and U5910 (N_5910,N_4608,N_4774);
nand U5911 (N_5911,N_4208,N_4209);
or U5912 (N_5912,N_4059,N_4868);
and U5913 (N_5913,N_4641,N_4186);
nand U5914 (N_5914,N_4774,N_4351);
nand U5915 (N_5915,N_4960,N_4033);
or U5916 (N_5916,N_4936,N_4629);
nor U5917 (N_5917,N_4800,N_4836);
nand U5918 (N_5918,N_4424,N_4426);
nor U5919 (N_5919,N_4945,N_4279);
nand U5920 (N_5920,N_4901,N_4355);
xor U5921 (N_5921,N_4438,N_4820);
or U5922 (N_5922,N_4112,N_4686);
nand U5923 (N_5923,N_4424,N_4626);
and U5924 (N_5924,N_4316,N_4370);
nor U5925 (N_5925,N_4239,N_4372);
or U5926 (N_5926,N_4132,N_4466);
or U5927 (N_5927,N_4810,N_4582);
and U5928 (N_5928,N_4423,N_4496);
or U5929 (N_5929,N_4695,N_4070);
and U5930 (N_5930,N_4237,N_4067);
or U5931 (N_5931,N_4137,N_4325);
nor U5932 (N_5932,N_4439,N_4757);
nand U5933 (N_5933,N_4694,N_4243);
and U5934 (N_5934,N_4675,N_4978);
xor U5935 (N_5935,N_4618,N_4991);
and U5936 (N_5936,N_4918,N_4917);
or U5937 (N_5937,N_4582,N_4289);
or U5938 (N_5938,N_4664,N_4342);
and U5939 (N_5939,N_4661,N_4118);
xnor U5940 (N_5940,N_4402,N_4870);
or U5941 (N_5941,N_4298,N_4447);
and U5942 (N_5942,N_4728,N_4565);
nor U5943 (N_5943,N_4724,N_4766);
xor U5944 (N_5944,N_4063,N_4523);
nand U5945 (N_5945,N_4046,N_4433);
nand U5946 (N_5946,N_4089,N_4174);
nor U5947 (N_5947,N_4611,N_4140);
nor U5948 (N_5948,N_4051,N_4308);
and U5949 (N_5949,N_4975,N_4169);
nor U5950 (N_5950,N_4477,N_4251);
nor U5951 (N_5951,N_4947,N_4416);
or U5952 (N_5952,N_4393,N_4824);
nand U5953 (N_5953,N_4309,N_4425);
or U5954 (N_5954,N_4923,N_4576);
nand U5955 (N_5955,N_4477,N_4851);
nand U5956 (N_5956,N_4842,N_4268);
nor U5957 (N_5957,N_4102,N_4552);
nor U5958 (N_5958,N_4351,N_4387);
nor U5959 (N_5959,N_4769,N_4097);
nor U5960 (N_5960,N_4795,N_4494);
nand U5961 (N_5961,N_4348,N_4556);
and U5962 (N_5962,N_4970,N_4308);
and U5963 (N_5963,N_4319,N_4160);
nand U5964 (N_5964,N_4786,N_4729);
nand U5965 (N_5965,N_4788,N_4165);
nand U5966 (N_5966,N_4420,N_4430);
nor U5967 (N_5967,N_4082,N_4803);
or U5968 (N_5968,N_4535,N_4538);
nand U5969 (N_5969,N_4204,N_4259);
and U5970 (N_5970,N_4201,N_4834);
or U5971 (N_5971,N_4291,N_4872);
nor U5972 (N_5972,N_4748,N_4887);
and U5973 (N_5973,N_4902,N_4514);
nor U5974 (N_5974,N_4377,N_4670);
nor U5975 (N_5975,N_4552,N_4995);
or U5976 (N_5976,N_4375,N_4315);
nor U5977 (N_5977,N_4696,N_4486);
and U5978 (N_5978,N_4263,N_4743);
nor U5979 (N_5979,N_4670,N_4331);
or U5980 (N_5980,N_4244,N_4958);
xnor U5981 (N_5981,N_4621,N_4132);
and U5982 (N_5982,N_4501,N_4715);
xnor U5983 (N_5983,N_4150,N_4135);
or U5984 (N_5984,N_4055,N_4384);
nor U5985 (N_5985,N_4508,N_4795);
and U5986 (N_5986,N_4933,N_4643);
and U5987 (N_5987,N_4172,N_4940);
nand U5988 (N_5988,N_4977,N_4396);
and U5989 (N_5989,N_4112,N_4253);
or U5990 (N_5990,N_4380,N_4552);
and U5991 (N_5991,N_4088,N_4793);
nor U5992 (N_5992,N_4401,N_4681);
or U5993 (N_5993,N_4236,N_4675);
nand U5994 (N_5994,N_4595,N_4088);
or U5995 (N_5995,N_4767,N_4108);
xnor U5996 (N_5996,N_4799,N_4503);
nor U5997 (N_5997,N_4503,N_4379);
nor U5998 (N_5998,N_4876,N_4406);
and U5999 (N_5999,N_4067,N_4937);
nand U6000 (N_6000,N_5343,N_5027);
and U6001 (N_6001,N_5624,N_5352);
xor U6002 (N_6002,N_5065,N_5867);
xnor U6003 (N_6003,N_5994,N_5266);
or U6004 (N_6004,N_5497,N_5091);
nor U6005 (N_6005,N_5413,N_5913);
or U6006 (N_6006,N_5835,N_5766);
or U6007 (N_6007,N_5345,N_5322);
nand U6008 (N_6008,N_5415,N_5968);
xor U6009 (N_6009,N_5038,N_5315);
and U6010 (N_6010,N_5879,N_5326);
nand U6011 (N_6011,N_5708,N_5269);
nor U6012 (N_6012,N_5148,N_5334);
and U6013 (N_6013,N_5432,N_5995);
xor U6014 (N_6014,N_5061,N_5122);
and U6015 (N_6015,N_5627,N_5874);
or U6016 (N_6016,N_5872,N_5064);
nand U6017 (N_6017,N_5816,N_5156);
nor U6018 (N_6018,N_5933,N_5980);
and U6019 (N_6019,N_5438,N_5882);
nand U6020 (N_6020,N_5519,N_5821);
and U6021 (N_6021,N_5753,N_5226);
nand U6022 (N_6022,N_5107,N_5136);
and U6023 (N_6023,N_5443,N_5414);
nand U6024 (N_6024,N_5394,N_5167);
and U6025 (N_6025,N_5999,N_5244);
nand U6026 (N_6026,N_5965,N_5647);
nand U6027 (N_6027,N_5839,N_5837);
nor U6028 (N_6028,N_5364,N_5298);
nand U6029 (N_6029,N_5392,N_5197);
nand U6030 (N_6030,N_5609,N_5255);
nor U6031 (N_6031,N_5342,N_5640);
nor U6032 (N_6032,N_5823,N_5188);
and U6033 (N_6033,N_5140,N_5769);
or U6034 (N_6034,N_5370,N_5304);
nand U6035 (N_6035,N_5387,N_5530);
nand U6036 (N_6036,N_5799,N_5112);
and U6037 (N_6037,N_5551,N_5806);
xor U6038 (N_6038,N_5259,N_5291);
nand U6039 (N_6039,N_5317,N_5512);
or U6040 (N_6040,N_5402,N_5025);
nor U6041 (N_6041,N_5373,N_5355);
nor U6042 (N_6042,N_5272,N_5040);
and U6043 (N_6043,N_5274,N_5755);
nor U6044 (N_6044,N_5516,N_5729);
nand U6045 (N_6045,N_5446,N_5023);
or U6046 (N_6046,N_5719,N_5316);
nand U6047 (N_6047,N_5804,N_5570);
or U6048 (N_6048,N_5578,N_5477);
nand U6049 (N_6049,N_5553,N_5840);
xnor U6050 (N_6050,N_5212,N_5846);
and U6051 (N_6051,N_5299,N_5233);
nor U6052 (N_6052,N_5044,N_5421);
or U6053 (N_6053,N_5383,N_5526);
or U6054 (N_6054,N_5412,N_5854);
nand U6055 (N_6055,N_5836,N_5542);
or U6056 (N_6056,N_5959,N_5697);
and U6057 (N_6057,N_5945,N_5779);
or U6058 (N_6058,N_5007,N_5734);
or U6059 (N_6059,N_5435,N_5032);
and U6060 (N_6060,N_5470,N_5374);
nand U6061 (N_6061,N_5514,N_5369);
nand U6062 (N_6062,N_5715,N_5720);
and U6063 (N_6063,N_5922,N_5689);
and U6064 (N_6064,N_5240,N_5456);
or U6065 (N_6065,N_5711,N_5631);
xor U6066 (N_6066,N_5458,N_5002);
xor U6067 (N_6067,N_5507,N_5622);
and U6068 (N_6068,N_5654,N_5740);
nand U6069 (N_6069,N_5360,N_5498);
nor U6070 (N_6070,N_5775,N_5273);
nand U6071 (N_6071,N_5560,N_5353);
or U6072 (N_6072,N_5971,N_5312);
nor U6073 (N_6073,N_5379,N_5961);
nand U6074 (N_6074,N_5749,N_5489);
and U6075 (N_6075,N_5218,N_5311);
nor U6076 (N_6076,N_5985,N_5518);
nand U6077 (N_6077,N_5955,N_5651);
nand U6078 (N_6078,N_5663,N_5024);
xnor U6079 (N_6079,N_5983,N_5359);
and U6080 (N_6080,N_5405,N_5289);
and U6081 (N_6081,N_5847,N_5501);
and U6082 (N_6082,N_5488,N_5324);
nor U6083 (N_6083,N_5664,N_5826);
nand U6084 (N_6084,N_5871,N_5898);
xnor U6085 (N_6085,N_5565,N_5531);
and U6086 (N_6086,N_5855,N_5868);
or U6087 (N_6087,N_5468,N_5280);
or U6088 (N_6088,N_5060,N_5659);
and U6089 (N_6089,N_5653,N_5419);
nand U6090 (N_6090,N_5595,N_5260);
and U6091 (N_6091,N_5891,N_5957);
or U6092 (N_6092,N_5461,N_5935);
and U6093 (N_6093,N_5884,N_5680);
or U6094 (N_6094,N_5340,N_5712);
xor U6095 (N_6095,N_5811,N_5439);
or U6096 (N_6096,N_5161,N_5887);
xnor U6097 (N_6097,N_5330,N_5086);
and U6098 (N_6098,N_5250,N_5802);
nand U6099 (N_6099,N_5908,N_5704);
nor U6100 (N_6100,N_5739,N_5011);
or U6101 (N_6101,N_5440,N_5256);
and U6102 (N_6102,N_5285,N_5016);
nor U6103 (N_6103,N_5617,N_5213);
nor U6104 (N_6104,N_5964,N_5988);
and U6105 (N_6105,N_5251,N_5454);
nor U6106 (N_6106,N_5937,N_5183);
nand U6107 (N_6107,N_5248,N_5376);
nor U6108 (N_6108,N_5385,N_5911);
or U6109 (N_6109,N_5730,N_5431);
nor U6110 (N_6110,N_5276,N_5841);
and U6111 (N_6111,N_5869,N_5277);
nor U6112 (N_6112,N_5181,N_5987);
nand U6113 (N_6113,N_5574,N_5339);
nand U6114 (N_6114,N_5880,N_5114);
nor U6115 (N_6115,N_5752,N_5203);
nor U6116 (N_6116,N_5490,N_5134);
and U6117 (N_6117,N_5155,N_5579);
nor U6118 (N_6118,N_5099,N_5046);
nor U6119 (N_6119,N_5917,N_5862);
nor U6120 (N_6120,N_5106,N_5423);
and U6121 (N_6121,N_5144,N_5620);
or U6122 (N_6122,N_5978,N_5030);
nand U6123 (N_6123,N_5628,N_5282);
xor U6124 (N_6124,N_5157,N_5162);
nand U6125 (N_6125,N_5619,N_5363);
or U6126 (N_6126,N_5104,N_5142);
nand U6127 (N_6127,N_5794,N_5537);
nor U6128 (N_6128,N_5052,N_5235);
nor U6129 (N_6129,N_5783,N_5618);
or U6130 (N_6130,N_5050,N_5652);
or U6131 (N_6131,N_5418,N_5265);
nand U6132 (N_6132,N_5870,N_5688);
nand U6133 (N_6133,N_5604,N_5528);
or U6134 (N_6134,N_5223,N_5329);
nor U6135 (N_6135,N_5207,N_5337);
nor U6136 (N_6136,N_5706,N_5215);
and U6137 (N_6137,N_5566,N_5686);
and U6138 (N_6138,N_5372,N_5529);
and U6139 (N_6139,N_5453,N_5168);
nor U6140 (N_6140,N_5100,N_5781);
or U6141 (N_6141,N_5015,N_5436);
nand U6142 (N_6142,N_5028,N_5287);
and U6143 (N_6143,N_5926,N_5150);
nand U6144 (N_6144,N_5208,N_5843);
nor U6145 (N_6145,N_5877,N_5726);
nand U6146 (N_6146,N_5138,N_5696);
nand U6147 (N_6147,N_5724,N_5818);
nor U6148 (N_6148,N_5309,N_5448);
nand U6149 (N_6149,N_5656,N_5533);
and U6150 (N_6150,N_5725,N_5239);
or U6151 (N_6151,N_5261,N_5123);
nor U6152 (N_6152,N_5314,N_5262);
nor U6153 (N_6153,N_5644,N_5723);
nand U6154 (N_6154,N_5327,N_5648);
or U6155 (N_6155,N_5377,N_5069);
xnor U6156 (N_6156,N_5780,N_5705);
nand U6157 (N_6157,N_5388,N_5476);
or U6158 (N_6158,N_5117,N_5001);
xnor U6159 (N_6159,N_5613,N_5853);
nor U6160 (N_6160,N_5286,N_5119);
and U6161 (N_6161,N_5930,N_5420);
and U6162 (N_6162,N_5710,N_5083);
nand U6163 (N_6163,N_5834,N_5576);
nor U6164 (N_6164,N_5474,N_5743);
nand U6165 (N_6165,N_5568,N_5320);
and U6166 (N_6166,N_5792,N_5059);
nor U6167 (N_6167,N_5756,N_5022);
xnor U6168 (N_6168,N_5630,N_5236);
nand U6169 (N_6169,N_5916,N_5176);
nor U6170 (N_6170,N_5247,N_5778);
nand U6171 (N_6171,N_5447,N_5805);
or U6172 (N_6172,N_5808,N_5857);
nand U6173 (N_6173,N_5234,N_5881);
nand U6174 (N_6174,N_5791,N_5062);
or U6175 (N_6175,N_5534,N_5094);
xnor U6176 (N_6176,N_5469,N_5850);
xnor U6177 (N_6177,N_5058,N_5270);
and U6178 (N_6178,N_5545,N_5184);
and U6179 (N_6179,N_5829,N_5747);
nand U6180 (N_6180,N_5758,N_5169);
nor U6181 (N_6181,N_5938,N_5034);
and U6182 (N_6182,N_5400,N_5429);
xor U6183 (N_6183,N_5192,N_5583);
nand U6184 (N_6184,N_5949,N_5396);
nor U6185 (N_6185,N_5481,N_5559);
or U6186 (N_6186,N_5548,N_5641);
or U6187 (N_6187,N_5278,N_5722);
nor U6188 (N_6188,N_5198,N_5737);
xnor U6189 (N_6189,N_5092,N_5744);
xor U6190 (N_6190,N_5543,N_5249);
nand U6191 (N_6191,N_5691,N_5655);
xor U6192 (N_6192,N_5675,N_5152);
nor U6193 (N_6193,N_5075,N_5467);
or U6194 (N_6194,N_5367,N_5328);
or U6195 (N_6195,N_5500,N_5635);
xnor U6196 (N_6196,N_5056,N_5407);
nand U6197 (N_6197,N_5495,N_5389);
or U6198 (N_6198,N_5253,N_5033);
xnor U6199 (N_6199,N_5159,N_5095);
nand U6200 (N_6200,N_5931,N_5606);
nand U6201 (N_6201,N_5252,N_5943);
nand U6202 (N_6202,N_5844,N_5731);
xnor U6203 (N_6203,N_5515,N_5153);
nand U6204 (N_6204,N_5300,N_5845);
nand U6205 (N_6205,N_5129,N_5577);
nand U6206 (N_6206,N_5906,N_5079);
xor U6207 (N_6207,N_5386,N_5430);
nand U6208 (N_6208,N_5581,N_5410);
or U6209 (N_6209,N_5940,N_5896);
and U6210 (N_6210,N_5510,N_5698);
nand U6211 (N_6211,N_5685,N_5827);
and U6212 (N_6212,N_5464,N_5217);
and U6213 (N_6213,N_5546,N_5170);
nand U6214 (N_6214,N_5903,N_5325);
xor U6215 (N_6215,N_5257,N_5174);
or U6216 (N_6216,N_5625,N_5206);
nand U6217 (N_6217,N_5308,N_5102);
or U6218 (N_6218,N_5371,N_5591);
or U6219 (N_6219,N_5953,N_5848);
nand U6220 (N_6220,N_5975,N_5404);
nand U6221 (N_6221,N_5989,N_5504);
xor U6222 (N_6222,N_5358,N_5864);
nor U6223 (N_6223,N_5074,N_5541);
or U6224 (N_6224,N_5762,N_5384);
nor U6225 (N_6225,N_5146,N_5084);
nor U6226 (N_6226,N_5962,N_5788);
and U6227 (N_6227,N_5361,N_5878);
nor U6228 (N_6228,N_5090,N_5670);
or U6229 (N_6229,N_5825,N_5113);
xor U6230 (N_6230,N_5571,N_5115);
or U6231 (N_6231,N_5313,N_5970);
and U6232 (N_6232,N_5424,N_5736);
or U6233 (N_6233,N_5886,N_5876);
or U6234 (N_6234,N_5346,N_5082);
nand U6235 (N_6235,N_5411,N_5761);
nor U6236 (N_6236,N_5268,N_5661);
nor U6237 (N_6237,N_5126,N_5558);
nor U6238 (N_6238,N_5201,N_5795);
or U6239 (N_6239,N_5450,N_5671);
or U6240 (N_6240,N_5612,N_5600);
nand U6241 (N_6241,N_5171,N_5632);
nand U6242 (N_6242,N_5810,N_5919);
xnor U6243 (N_6243,N_5900,N_5323);
nor U6244 (N_6244,N_5147,N_5131);
or U6245 (N_6245,N_5101,N_5036);
and U6246 (N_6246,N_5175,N_5381);
and U6247 (N_6247,N_5139,N_5229);
or U6248 (N_6248,N_5378,N_5824);
nor U6249 (N_6249,N_5941,N_5141);
or U6250 (N_6250,N_5505,N_5746);
xor U6251 (N_6251,N_5772,N_5293);
xnor U6252 (N_6252,N_5520,N_5427);
nand U6253 (N_6253,N_5787,N_5582);
nor U6254 (N_6254,N_5899,N_5426);
nor U6255 (N_6255,N_5773,N_5770);
nor U6256 (N_6256,N_5057,N_5365);
or U6257 (N_6257,N_5748,N_5089);
or U6258 (N_6258,N_5416,N_5539);
or U6259 (N_6259,N_5110,N_5425);
or U6260 (N_6260,N_5944,N_5191);
and U6261 (N_6261,N_5692,N_5986);
and U6262 (N_6262,N_5465,N_5484);
or U6263 (N_6263,N_5925,N_5398);
nand U6264 (N_6264,N_5584,N_5290);
and U6265 (N_6265,N_5822,N_5567);
or U6266 (N_6266,N_5535,N_5759);
and U6267 (N_6267,N_5682,N_5105);
nor U6268 (N_6268,N_5194,N_5301);
or U6269 (N_6269,N_5662,N_5133);
nor U6270 (N_6270,N_5124,N_5354);
or U6271 (N_6271,N_5765,N_5803);
and U6272 (N_6272,N_5014,N_5966);
or U6273 (N_6273,N_5849,N_5634);
and U6274 (N_6274,N_5222,N_5264);
nand U6275 (N_6275,N_5564,N_5633);
xor U6276 (N_6276,N_5667,N_5511);
nor U6277 (N_6277,N_5895,N_5524);
and U6278 (N_6278,N_5590,N_5041);
or U6279 (N_6279,N_5132,N_5993);
or U6280 (N_6280,N_5160,N_5552);
nand U6281 (N_6281,N_5375,N_5972);
nand U6282 (N_6282,N_5031,N_5596);
or U6283 (N_6283,N_5592,N_5650);
nor U6284 (N_6284,N_5523,N_5910);
nor U6285 (N_6285,N_5245,N_5199);
and U6286 (N_6286,N_5563,N_5833);
nand U6287 (N_6287,N_5767,N_5401);
and U6288 (N_6288,N_5294,N_5709);
nor U6289 (N_6289,N_5555,N_5096);
and U6290 (N_6290,N_5852,N_5406);
or U6291 (N_6291,N_5382,N_5996);
nand U6292 (N_6292,N_5679,N_5391);
nor U6293 (N_6293,N_5356,N_5754);
or U6294 (N_6294,N_5066,N_5077);
and U6295 (N_6295,N_5693,N_5085);
or U6296 (N_6296,N_5888,N_5660);
and U6297 (N_6297,N_5776,N_5281);
xor U6298 (N_6298,N_5051,N_5665);
xor U6299 (N_6299,N_5437,N_5923);
and U6300 (N_6300,N_5946,N_5054);
and U6301 (N_6301,N_5399,N_5915);
and U6302 (N_6302,N_5861,N_5284);
nand U6303 (N_6303,N_5196,N_5390);
and U6304 (N_6304,N_5462,N_5936);
nand U6305 (N_6305,N_5296,N_5977);
nor U6306 (N_6306,N_5459,N_5587);
nand U6307 (N_6307,N_5485,N_5063);
or U6308 (N_6308,N_5279,N_5502);
xnor U6309 (N_6309,N_5639,N_5177);
nand U6310 (N_6310,N_5601,N_5037);
xnor U6311 (N_6311,N_5513,N_5263);
nand U6312 (N_6312,N_5602,N_5554);
or U6313 (N_6313,N_5777,N_5597);
nor U6314 (N_6314,N_5288,N_5080);
nand U6315 (N_6315,N_5081,N_5540);
xnor U6316 (N_6316,N_5594,N_5814);
and U6317 (N_6317,N_5145,N_5109);
or U6318 (N_6318,N_5669,N_5295);
nor U6319 (N_6319,N_5026,N_5344);
nand U6320 (N_6320,N_5863,N_5246);
nor U6321 (N_6321,N_5856,N_5924);
and U6322 (N_6322,N_5687,N_5678);
or U6323 (N_6323,N_5178,N_5486);
nand U6324 (N_6324,N_5463,N_5307);
nor U6325 (N_6325,N_5395,N_5842);
nor U6326 (N_6326,N_5202,N_5521);
nor U6327 (N_6327,N_5179,N_5657);
xor U6328 (N_6328,N_5434,N_5380);
nand U6329 (N_6329,N_5610,N_5956);
nand U6330 (N_6330,N_5883,N_5642);
and U6331 (N_6331,N_5681,N_5195);
nor U6332 (N_6332,N_5128,N_5478);
or U6333 (N_6333,N_5889,N_5087);
nor U6334 (N_6334,N_5433,N_5258);
and U6335 (N_6335,N_5237,N_5738);
and U6336 (N_6336,N_5333,N_5499);
nand U6337 (N_6337,N_5817,N_5154);
and U6338 (N_6338,N_5831,N_5455);
nand U6339 (N_6339,N_5366,N_5283);
and U6340 (N_6340,N_5991,N_5035);
nor U6341 (N_6341,N_5496,N_5958);
and U6342 (N_6342,N_5422,N_5690);
nand U6343 (N_6343,N_5442,N_5475);
xnor U6344 (N_6344,N_5303,N_5004);
nor U6345 (N_6345,N_5611,N_5727);
or U6346 (N_6346,N_5703,N_5733);
and U6347 (N_6347,N_5866,N_5626);
nand U6348 (N_6348,N_5585,N_5460);
or U6349 (N_6349,N_5070,N_5873);
nor U6350 (N_6350,N_5043,N_5683);
and U6351 (N_6351,N_5021,N_5047);
and U6352 (N_6352,N_5774,N_5580);
or U6353 (N_6353,N_5143,N_5045);
nand U6354 (N_6354,N_5984,N_5127);
nand U6355 (N_6355,N_5934,N_5668);
nor U6356 (N_6356,N_5221,N_5186);
xnor U6357 (N_6357,N_5947,N_5073);
and U6358 (N_6358,N_5098,N_5292);
nand U6359 (N_6359,N_5549,N_5950);
xnor U6360 (N_6360,N_5598,N_5672);
xnor U6361 (N_6361,N_5556,N_5029);
nand U6362 (N_6362,N_5714,N_5607);
and U6363 (N_6363,N_5997,N_5172);
or U6364 (N_6364,N_5932,N_5006);
and U6365 (N_6365,N_5764,N_5960);
nor U6366 (N_6366,N_5973,N_5789);
or U6367 (N_6367,N_5393,N_5562);
and U6368 (N_6368,N_5241,N_5875);
and U6369 (N_6369,N_5901,N_5321);
nor U6370 (N_6370,N_5828,N_5163);
or U6371 (N_6371,N_5479,N_5243);
nor U6372 (N_6372,N_5267,N_5674);
nand U6373 (N_6373,N_5800,N_5905);
xor U6374 (N_6374,N_5350,N_5603);
nor U6375 (N_6375,N_5527,N_5242);
nand U6376 (N_6376,N_5569,N_5232);
and U6377 (N_6377,N_5942,N_5210);
or U6378 (N_6378,N_5494,N_5649);
nand U6379 (N_6379,N_5939,N_5003);
xor U6380 (N_6380,N_5525,N_5116);
nand U6381 (N_6381,N_5111,N_5820);
or U6382 (N_6382,N_5982,N_5716);
nand U6383 (N_6383,N_5362,N_5205);
xor U6384 (N_6384,N_5677,N_5797);
and U6385 (N_6385,N_5219,N_5227);
or U6386 (N_6386,N_5979,N_5149);
nand U6387 (N_6387,N_5928,N_5165);
or U6388 (N_6388,N_5297,N_5166);
nor U6389 (N_6389,N_5801,N_5717);
or U6390 (N_6390,N_5918,N_5068);
and U6391 (N_6391,N_5491,N_5271);
nand U6392 (N_6392,N_5185,N_5676);
or U6393 (N_6393,N_5189,N_5492);
or U6394 (N_6394,N_5008,N_5684);
xor U6395 (N_6395,N_5441,N_5561);
nor U6396 (N_6396,N_5621,N_5049);
xnor U6397 (N_6397,N_5137,N_5397);
and U6398 (N_6398,N_5214,N_5990);
or U6399 (N_6399,N_5230,N_5819);
xor U6400 (N_6400,N_5713,N_5623);
and U6401 (N_6401,N_5302,N_5506);
or U6402 (N_6402,N_5575,N_5451);
and U6403 (N_6403,N_5813,N_5637);
and U6404 (N_6404,N_5417,N_5638);
nor U6405 (N_6405,N_5865,N_5190);
or U6406 (N_6406,N_5509,N_5483);
nor U6407 (N_6407,N_5912,N_5053);
nand U6408 (N_6408,N_5076,N_5216);
or U6409 (N_6409,N_5702,N_5331);
or U6410 (N_6410,N_5885,N_5586);
xnor U6411 (N_6411,N_5589,N_5547);
nor U6412 (N_6412,N_5929,N_5048);
nand U6413 (N_6413,N_5976,N_5009);
and U6414 (N_6414,N_5832,N_5643);
xnor U6415 (N_6415,N_5909,N_5793);
or U6416 (N_6416,N_5466,N_5658);
or U6417 (N_6417,N_5550,N_5005);
or U6418 (N_6418,N_5859,N_5408);
nand U6419 (N_6419,N_5254,N_5522);
xor U6420 (N_6420,N_5103,N_5851);
nand U6421 (N_6421,N_5593,N_5010);
or U6422 (N_6422,N_5967,N_5078);
nor U6423 (N_6423,N_5335,N_5457);
and U6424 (N_6424,N_5981,N_5538);
nand U6425 (N_6425,N_5645,N_5508);
nand U6426 (N_6426,N_5351,N_5088);
xnor U6427 (N_6427,N_5349,N_5220);
nand U6428 (N_6428,N_5735,N_5517);
or U6429 (N_6429,N_5125,N_5338);
nand U6430 (N_6430,N_5072,N_5615);
or U6431 (N_6431,N_5093,N_5480);
nand U6432 (N_6432,N_5636,N_5487);
nor U6433 (N_6433,N_5969,N_5409);
nand U6434 (N_6434,N_5310,N_5403);
and U6435 (N_6435,N_5536,N_5588);
nand U6436 (N_6436,N_5319,N_5721);
or U6437 (N_6437,N_5445,N_5347);
nor U6438 (N_6438,N_5557,N_5042);
nand U6439 (N_6439,N_5920,N_5471);
xnor U6440 (N_6440,N_5209,N_5763);
nor U6441 (N_6441,N_5118,N_5019);
or U6442 (N_6442,N_5605,N_5897);
nand U6443 (N_6443,N_5760,N_5182);
nor U6444 (N_6444,N_5750,N_5173);
nand U6445 (N_6445,N_5921,N_5629);
nor U6446 (N_6446,N_5097,N_5224);
or U6447 (N_6447,N_5732,N_5860);
or U6448 (N_6448,N_5666,N_5444);
and U6449 (N_6449,N_5472,N_5193);
or U6450 (N_6450,N_5812,N_5728);
and U6451 (N_6451,N_5948,N_5914);
nand U6452 (N_6452,N_5200,N_5452);
nor U6453 (N_6453,N_5306,N_5902);
and U6454 (N_6454,N_5018,N_5771);
and U6455 (N_6455,N_5482,N_5718);
nor U6456 (N_6456,N_5204,N_5893);
xnor U6457 (N_6457,N_5695,N_5020);
nand U6458 (N_6458,N_5275,N_5336);
xor U6459 (N_6459,N_5798,N_5838);
nor U6460 (N_6460,N_5238,N_5573);
nand U6461 (N_6461,N_5741,N_5786);
and U6462 (N_6462,N_5158,N_5121);
and U6463 (N_6463,N_5751,N_5784);
or U6464 (N_6464,N_5357,N_5790);
nor U6465 (N_6465,N_5503,N_5228);
nand U6466 (N_6466,N_5809,N_5120);
nor U6467 (N_6467,N_5785,N_5108);
or U6468 (N_6468,N_5348,N_5768);
and U6469 (N_6469,N_5428,N_5892);
nor U6470 (N_6470,N_5927,N_5572);
xor U6471 (N_6471,N_5700,N_5231);
and U6472 (N_6472,N_5890,N_5742);
and U6473 (N_6473,N_5616,N_5368);
nand U6474 (N_6474,N_5532,N_5694);
or U6475 (N_6475,N_5904,N_5614);
nor U6476 (N_6476,N_5013,N_5701);
or U6477 (N_6477,N_5012,N_5493);
or U6478 (N_6478,N_5305,N_5187);
nor U6479 (N_6479,N_5992,N_5544);
nand U6480 (N_6480,N_5599,N_5807);
nand U6481 (N_6481,N_5071,N_5830);
and U6482 (N_6482,N_5782,N_5707);
nand U6483 (N_6483,N_5699,N_5815);
and U6484 (N_6484,N_5796,N_5745);
nand U6485 (N_6485,N_5000,N_5318);
nor U6486 (N_6486,N_5473,N_5954);
or U6487 (N_6487,N_5039,N_5894);
xnor U6488 (N_6488,N_5164,N_5907);
or U6489 (N_6489,N_5449,N_5211);
or U6490 (N_6490,N_5646,N_5180);
xnor U6491 (N_6491,N_5608,N_5135);
and U6492 (N_6492,N_5673,N_5225);
xor U6493 (N_6493,N_5151,N_5951);
nand U6494 (N_6494,N_5130,N_5067);
xnor U6495 (N_6495,N_5974,N_5017);
and U6496 (N_6496,N_5757,N_5963);
nand U6497 (N_6497,N_5055,N_5858);
or U6498 (N_6498,N_5998,N_5341);
and U6499 (N_6499,N_5332,N_5952);
and U6500 (N_6500,N_5948,N_5889);
nor U6501 (N_6501,N_5101,N_5441);
or U6502 (N_6502,N_5665,N_5027);
nor U6503 (N_6503,N_5468,N_5273);
or U6504 (N_6504,N_5971,N_5361);
xnor U6505 (N_6505,N_5536,N_5673);
or U6506 (N_6506,N_5365,N_5454);
or U6507 (N_6507,N_5716,N_5230);
nor U6508 (N_6508,N_5636,N_5150);
or U6509 (N_6509,N_5899,N_5441);
nor U6510 (N_6510,N_5686,N_5320);
nand U6511 (N_6511,N_5454,N_5407);
and U6512 (N_6512,N_5849,N_5570);
and U6513 (N_6513,N_5096,N_5085);
nand U6514 (N_6514,N_5676,N_5624);
nor U6515 (N_6515,N_5996,N_5219);
nor U6516 (N_6516,N_5692,N_5894);
or U6517 (N_6517,N_5264,N_5853);
and U6518 (N_6518,N_5240,N_5719);
or U6519 (N_6519,N_5529,N_5146);
nor U6520 (N_6520,N_5366,N_5217);
or U6521 (N_6521,N_5185,N_5779);
nand U6522 (N_6522,N_5253,N_5461);
nand U6523 (N_6523,N_5696,N_5951);
nor U6524 (N_6524,N_5437,N_5587);
nor U6525 (N_6525,N_5819,N_5646);
xnor U6526 (N_6526,N_5494,N_5446);
nand U6527 (N_6527,N_5033,N_5408);
nand U6528 (N_6528,N_5306,N_5171);
and U6529 (N_6529,N_5379,N_5438);
nor U6530 (N_6530,N_5322,N_5976);
or U6531 (N_6531,N_5224,N_5652);
nor U6532 (N_6532,N_5286,N_5905);
and U6533 (N_6533,N_5348,N_5635);
and U6534 (N_6534,N_5120,N_5995);
and U6535 (N_6535,N_5517,N_5444);
and U6536 (N_6536,N_5077,N_5502);
nand U6537 (N_6537,N_5641,N_5892);
or U6538 (N_6538,N_5918,N_5789);
nand U6539 (N_6539,N_5226,N_5265);
nor U6540 (N_6540,N_5615,N_5723);
nor U6541 (N_6541,N_5525,N_5065);
nor U6542 (N_6542,N_5107,N_5637);
and U6543 (N_6543,N_5955,N_5922);
or U6544 (N_6544,N_5103,N_5074);
or U6545 (N_6545,N_5791,N_5060);
nand U6546 (N_6546,N_5760,N_5290);
nand U6547 (N_6547,N_5089,N_5690);
and U6548 (N_6548,N_5157,N_5008);
and U6549 (N_6549,N_5128,N_5361);
or U6550 (N_6550,N_5046,N_5291);
or U6551 (N_6551,N_5571,N_5336);
and U6552 (N_6552,N_5841,N_5580);
nand U6553 (N_6553,N_5016,N_5803);
nand U6554 (N_6554,N_5204,N_5390);
nand U6555 (N_6555,N_5979,N_5181);
nor U6556 (N_6556,N_5442,N_5381);
nand U6557 (N_6557,N_5196,N_5893);
and U6558 (N_6558,N_5471,N_5118);
nor U6559 (N_6559,N_5374,N_5747);
nor U6560 (N_6560,N_5419,N_5866);
and U6561 (N_6561,N_5753,N_5452);
nand U6562 (N_6562,N_5483,N_5806);
nor U6563 (N_6563,N_5710,N_5636);
nand U6564 (N_6564,N_5698,N_5541);
nand U6565 (N_6565,N_5395,N_5770);
or U6566 (N_6566,N_5966,N_5129);
or U6567 (N_6567,N_5843,N_5296);
or U6568 (N_6568,N_5716,N_5400);
or U6569 (N_6569,N_5579,N_5515);
nand U6570 (N_6570,N_5689,N_5223);
and U6571 (N_6571,N_5325,N_5245);
nand U6572 (N_6572,N_5830,N_5262);
or U6573 (N_6573,N_5819,N_5727);
nand U6574 (N_6574,N_5081,N_5663);
nand U6575 (N_6575,N_5602,N_5520);
or U6576 (N_6576,N_5818,N_5549);
and U6577 (N_6577,N_5609,N_5049);
nor U6578 (N_6578,N_5422,N_5804);
and U6579 (N_6579,N_5081,N_5140);
or U6580 (N_6580,N_5022,N_5918);
xnor U6581 (N_6581,N_5644,N_5342);
nor U6582 (N_6582,N_5058,N_5703);
nor U6583 (N_6583,N_5197,N_5628);
or U6584 (N_6584,N_5657,N_5761);
nor U6585 (N_6585,N_5653,N_5633);
nor U6586 (N_6586,N_5147,N_5032);
nor U6587 (N_6587,N_5435,N_5803);
and U6588 (N_6588,N_5946,N_5230);
and U6589 (N_6589,N_5001,N_5051);
nor U6590 (N_6590,N_5776,N_5906);
nor U6591 (N_6591,N_5147,N_5690);
nor U6592 (N_6592,N_5195,N_5496);
or U6593 (N_6593,N_5027,N_5899);
nor U6594 (N_6594,N_5840,N_5844);
xor U6595 (N_6595,N_5780,N_5074);
nand U6596 (N_6596,N_5227,N_5210);
nand U6597 (N_6597,N_5790,N_5440);
nand U6598 (N_6598,N_5803,N_5224);
nor U6599 (N_6599,N_5582,N_5294);
nor U6600 (N_6600,N_5393,N_5846);
and U6601 (N_6601,N_5574,N_5270);
nor U6602 (N_6602,N_5726,N_5263);
nand U6603 (N_6603,N_5780,N_5579);
or U6604 (N_6604,N_5998,N_5167);
and U6605 (N_6605,N_5814,N_5476);
and U6606 (N_6606,N_5939,N_5704);
or U6607 (N_6607,N_5596,N_5883);
nor U6608 (N_6608,N_5254,N_5564);
xnor U6609 (N_6609,N_5500,N_5011);
and U6610 (N_6610,N_5688,N_5228);
nor U6611 (N_6611,N_5293,N_5946);
xnor U6612 (N_6612,N_5847,N_5228);
nor U6613 (N_6613,N_5689,N_5226);
or U6614 (N_6614,N_5820,N_5823);
nor U6615 (N_6615,N_5931,N_5926);
xor U6616 (N_6616,N_5320,N_5206);
xnor U6617 (N_6617,N_5256,N_5702);
nand U6618 (N_6618,N_5381,N_5300);
and U6619 (N_6619,N_5214,N_5494);
nor U6620 (N_6620,N_5458,N_5267);
and U6621 (N_6621,N_5957,N_5455);
nand U6622 (N_6622,N_5517,N_5151);
or U6623 (N_6623,N_5148,N_5401);
xor U6624 (N_6624,N_5864,N_5731);
and U6625 (N_6625,N_5633,N_5972);
or U6626 (N_6626,N_5044,N_5721);
nand U6627 (N_6627,N_5459,N_5348);
or U6628 (N_6628,N_5040,N_5846);
nor U6629 (N_6629,N_5445,N_5569);
or U6630 (N_6630,N_5784,N_5330);
and U6631 (N_6631,N_5143,N_5933);
or U6632 (N_6632,N_5083,N_5688);
or U6633 (N_6633,N_5435,N_5275);
or U6634 (N_6634,N_5798,N_5712);
or U6635 (N_6635,N_5804,N_5715);
nor U6636 (N_6636,N_5911,N_5784);
nor U6637 (N_6637,N_5605,N_5180);
or U6638 (N_6638,N_5656,N_5428);
nor U6639 (N_6639,N_5138,N_5004);
or U6640 (N_6640,N_5316,N_5646);
or U6641 (N_6641,N_5450,N_5676);
nand U6642 (N_6642,N_5747,N_5077);
and U6643 (N_6643,N_5943,N_5534);
nand U6644 (N_6644,N_5786,N_5399);
nor U6645 (N_6645,N_5640,N_5043);
and U6646 (N_6646,N_5553,N_5546);
nand U6647 (N_6647,N_5438,N_5932);
and U6648 (N_6648,N_5115,N_5046);
or U6649 (N_6649,N_5053,N_5130);
and U6650 (N_6650,N_5315,N_5264);
nor U6651 (N_6651,N_5062,N_5776);
and U6652 (N_6652,N_5691,N_5062);
or U6653 (N_6653,N_5867,N_5542);
nand U6654 (N_6654,N_5581,N_5580);
nand U6655 (N_6655,N_5624,N_5537);
and U6656 (N_6656,N_5269,N_5784);
and U6657 (N_6657,N_5493,N_5527);
nand U6658 (N_6658,N_5053,N_5886);
or U6659 (N_6659,N_5221,N_5708);
or U6660 (N_6660,N_5839,N_5100);
nand U6661 (N_6661,N_5530,N_5668);
or U6662 (N_6662,N_5978,N_5305);
or U6663 (N_6663,N_5128,N_5155);
or U6664 (N_6664,N_5644,N_5276);
xnor U6665 (N_6665,N_5027,N_5672);
nor U6666 (N_6666,N_5529,N_5200);
nand U6667 (N_6667,N_5803,N_5447);
or U6668 (N_6668,N_5189,N_5606);
and U6669 (N_6669,N_5413,N_5272);
nand U6670 (N_6670,N_5971,N_5549);
or U6671 (N_6671,N_5128,N_5730);
or U6672 (N_6672,N_5408,N_5086);
or U6673 (N_6673,N_5578,N_5795);
or U6674 (N_6674,N_5125,N_5028);
or U6675 (N_6675,N_5520,N_5072);
or U6676 (N_6676,N_5607,N_5038);
and U6677 (N_6677,N_5785,N_5914);
or U6678 (N_6678,N_5010,N_5189);
or U6679 (N_6679,N_5775,N_5620);
or U6680 (N_6680,N_5998,N_5316);
and U6681 (N_6681,N_5182,N_5259);
or U6682 (N_6682,N_5133,N_5252);
nand U6683 (N_6683,N_5897,N_5904);
nor U6684 (N_6684,N_5144,N_5896);
nor U6685 (N_6685,N_5199,N_5231);
xor U6686 (N_6686,N_5195,N_5001);
or U6687 (N_6687,N_5582,N_5061);
or U6688 (N_6688,N_5501,N_5213);
and U6689 (N_6689,N_5328,N_5080);
nor U6690 (N_6690,N_5562,N_5674);
nor U6691 (N_6691,N_5196,N_5057);
nor U6692 (N_6692,N_5176,N_5551);
nor U6693 (N_6693,N_5426,N_5691);
nand U6694 (N_6694,N_5411,N_5206);
nand U6695 (N_6695,N_5055,N_5907);
xnor U6696 (N_6696,N_5092,N_5393);
nand U6697 (N_6697,N_5080,N_5944);
nor U6698 (N_6698,N_5472,N_5521);
nor U6699 (N_6699,N_5417,N_5186);
or U6700 (N_6700,N_5153,N_5661);
nor U6701 (N_6701,N_5410,N_5961);
nor U6702 (N_6702,N_5120,N_5925);
or U6703 (N_6703,N_5302,N_5282);
or U6704 (N_6704,N_5610,N_5338);
and U6705 (N_6705,N_5416,N_5399);
nor U6706 (N_6706,N_5126,N_5697);
or U6707 (N_6707,N_5995,N_5475);
and U6708 (N_6708,N_5878,N_5133);
and U6709 (N_6709,N_5381,N_5149);
nand U6710 (N_6710,N_5815,N_5040);
or U6711 (N_6711,N_5700,N_5256);
and U6712 (N_6712,N_5194,N_5364);
and U6713 (N_6713,N_5711,N_5108);
nor U6714 (N_6714,N_5360,N_5417);
and U6715 (N_6715,N_5947,N_5889);
nor U6716 (N_6716,N_5032,N_5740);
nand U6717 (N_6717,N_5961,N_5046);
and U6718 (N_6718,N_5528,N_5606);
nor U6719 (N_6719,N_5388,N_5691);
and U6720 (N_6720,N_5059,N_5585);
nand U6721 (N_6721,N_5898,N_5381);
nor U6722 (N_6722,N_5319,N_5481);
nand U6723 (N_6723,N_5415,N_5866);
and U6724 (N_6724,N_5108,N_5115);
nand U6725 (N_6725,N_5334,N_5979);
xnor U6726 (N_6726,N_5819,N_5825);
nand U6727 (N_6727,N_5229,N_5989);
xnor U6728 (N_6728,N_5542,N_5075);
and U6729 (N_6729,N_5363,N_5750);
nor U6730 (N_6730,N_5704,N_5972);
nand U6731 (N_6731,N_5768,N_5651);
nand U6732 (N_6732,N_5540,N_5444);
and U6733 (N_6733,N_5471,N_5725);
and U6734 (N_6734,N_5675,N_5605);
or U6735 (N_6735,N_5775,N_5848);
or U6736 (N_6736,N_5777,N_5352);
and U6737 (N_6737,N_5815,N_5256);
and U6738 (N_6738,N_5116,N_5563);
and U6739 (N_6739,N_5741,N_5896);
nor U6740 (N_6740,N_5880,N_5210);
and U6741 (N_6741,N_5534,N_5328);
nand U6742 (N_6742,N_5074,N_5922);
and U6743 (N_6743,N_5131,N_5689);
or U6744 (N_6744,N_5072,N_5531);
nand U6745 (N_6745,N_5298,N_5083);
nor U6746 (N_6746,N_5611,N_5259);
or U6747 (N_6747,N_5406,N_5353);
nand U6748 (N_6748,N_5862,N_5561);
nor U6749 (N_6749,N_5564,N_5807);
nor U6750 (N_6750,N_5042,N_5755);
and U6751 (N_6751,N_5372,N_5138);
or U6752 (N_6752,N_5407,N_5513);
xnor U6753 (N_6753,N_5059,N_5452);
or U6754 (N_6754,N_5543,N_5713);
or U6755 (N_6755,N_5813,N_5109);
nor U6756 (N_6756,N_5503,N_5268);
nand U6757 (N_6757,N_5802,N_5152);
and U6758 (N_6758,N_5333,N_5948);
nor U6759 (N_6759,N_5657,N_5982);
nor U6760 (N_6760,N_5468,N_5934);
or U6761 (N_6761,N_5039,N_5924);
and U6762 (N_6762,N_5562,N_5195);
nor U6763 (N_6763,N_5149,N_5629);
nand U6764 (N_6764,N_5226,N_5268);
nand U6765 (N_6765,N_5335,N_5737);
or U6766 (N_6766,N_5836,N_5085);
and U6767 (N_6767,N_5987,N_5452);
nor U6768 (N_6768,N_5930,N_5854);
or U6769 (N_6769,N_5004,N_5353);
or U6770 (N_6770,N_5377,N_5461);
nand U6771 (N_6771,N_5357,N_5376);
nor U6772 (N_6772,N_5535,N_5758);
or U6773 (N_6773,N_5922,N_5754);
and U6774 (N_6774,N_5948,N_5883);
xnor U6775 (N_6775,N_5193,N_5249);
nor U6776 (N_6776,N_5346,N_5598);
or U6777 (N_6777,N_5382,N_5154);
or U6778 (N_6778,N_5304,N_5465);
or U6779 (N_6779,N_5859,N_5586);
nor U6780 (N_6780,N_5250,N_5744);
and U6781 (N_6781,N_5792,N_5755);
and U6782 (N_6782,N_5998,N_5511);
nand U6783 (N_6783,N_5903,N_5208);
nand U6784 (N_6784,N_5345,N_5928);
and U6785 (N_6785,N_5002,N_5952);
and U6786 (N_6786,N_5141,N_5684);
or U6787 (N_6787,N_5882,N_5578);
nand U6788 (N_6788,N_5177,N_5366);
nor U6789 (N_6789,N_5599,N_5471);
and U6790 (N_6790,N_5386,N_5708);
nand U6791 (N_6791,N_5998,N_5791);
and U6792 (N_6792,N_5254,N_5309);
or U6793 (N_6793,N_5915,N_5555);
and U6794 (N_6794,N_5695,N_5636);
and U6795 (N_6795,N_5472,N_5991);
and U6796 (N_6796,N_5676,N_5506);
or U6797 (N_6797,N_5180,N_5989);
and U6798 (N_6798,N_5294,N_5913);
or U6799 (N_6799,N_5080,N_5554);
nor U6800 (N_6800,N_5425,N_5960);
and U6801 (N_6801,N_5727,N_5953);
nand U6802 (N_6802,N_5172,N_5586);
nor U6803 (N_6803,N_5451,N_5299);
and U6804 (N_6804,N_5300,N_5319);
nor U6805 (N_6805,N_5132,N_5016);
nor U6806 (N_6806,N_5942,N_5610);
or U6807 (N_6807,N_5477,N_5289);
nor U6808 (N_6808,N_5013,N_5331);
or U6809 (N_6809,N_5078,N_5417);
nand U6810 (N_6810,N_5736,N_5366);
xnor U6811 (N_6811,N_5639,N_5940);
xnor U6812 (N_6812,N_5294,N_5902);
nand U6813 (N_6813,N_5858,N_5843);
or U6814 (N_6814,N_5323,N_5238);
nor U6815 (N_6815,N_5554,N_5295);
nand U6816 (N_6816,N_5603,N_5654);
and U6817 (N_6817,N_5321,N_5732);
and U6818 (N_6818,N_5718,N_5641);
and U6819 (N_6819,N_5166,N_5366);
nor U6820 (N_6820,N_5387,N_5963);
xor U6821 (N_6821,N_5968,N_5771);
or U6822 (N_6822,N_5481,N_5891);
nand U6823 (N_6823,N_5652,N_5087);
nor U6824 (N_6824,N_5383,N_5424);
nor U6825 (N_6825,N_5627,N_5314);
or U6826 (N_6826,N_5555,N_5126);
or U6827 (N_6827,N_5889,N_5616);
nand U6828 (N_6828,N_5015,N_5463);
nor U6829 (N_6829,N_5356,N_5742);
nand U6830 (N_6830,N_5264,N_5460);
nor U6831 (N_6831,N_5831,N_5884);
or U6832 (N_6832,N_5850,N_5285);
and U6833 (N_6833,N_5549,N_5300);
and U6834 (N_6834,N_5733,N_5588);
nor U6835 (N_6835,N_5616,N_5078);
or U6836 (N_6836,N_5701,N_5545);
or U6837 (N_6837,N_5050,N_5044);
or U6838 (N_6838,N_5291,N_5932);
or U6839 (N_6839,N_5968,N_5550);
and U6840 (N_6840,N_5593,N_5747);
xor U6841 (N_6841,N_5439,N_5010);
nand U6842 (N_6842,N_5457,N_5964);
nand U6843 (N_6843,N_5685,N_5312);
or U6844 (N_6844,N_5203,N_5090);
nor U6845 (N_6845,N_5870,N_5936);
nor U6846 (N_6846,N_5929,N_5101);
or U6847 (N_6847,N_5415,N_5956);
nand U6848 (N_6848,N_5677,N_5748);
or U6849 (N_6849,N_5211,N_5864);
nand U6850 (N_6850,N_5432,N_5040);
and U6851 (N_6851,N_5988,N_5336);
nor U6852 (N_6852,N_5226,N_5132);
nand U6853 (N_6853,N_5288,N_5310);
or U6854 (N_6854,N_5018,N_5431);
nand U6855 (N_6855,N_5276,N_5718);
nor U6856 (N_6856,N_5679,N_5633);
or U6857 (N_6857,N_5017,N_5838);
or U6858 (N_6858,N_5805,N_5285);
or U6859 (N_6859,N_5097,N_5468);
nor U6860 (N_6860,N_5722,N_5826);
nand U6861 (N_6861,N_5012,N_5525);
or U6862 (N_6862,N_5162,N_5252);
nand U6863 (N_6863,N_5433,N_5221);
and U6864 (N_6864,N_5770,N_5853);
nor U6865 (N_6865,N_5740,N_5987);
and U6866 (N_6866,N_5600,N_5692);
and U6867 (N_6867,N_5850,N_5746);
and U6868 (N_6868,N_5914,N_5251);
and U6869 (N_6869,N_5227,N_5698);
xor U6870 (N_6870,N_5509,N_5058);
nand U6871 (N_6871,N_5099,N_5439);
nor U6872 (N_6872,N_5184,N_5873);
or U6873 (N_6873,N_5579,N_5802);
or U6874 (N_6874,N_5766,N_5443);
nand U6875 (N_6875,N_5182,N_5711);
nand U6876 (N_6876,N_5824,N_5887);
nand U6877 (N_6877,N_5591,N_5316);
nor U6878 (N_6878,N_5046,N_5023);
nand U6879 (N_6879,N_5845,N_5596);
nand U6880 (N_6880,N_5118,N_5925);
or U6881 (N_6881,N_5486,N_5816);
or U6882 (N_6882,N_5172,N_5813);
xor U6883 (N_6883,N_5518,N_5751);
and U6884 (N_6884,N_5407,N_5058);
and U6885 (N_6885,N_5501,N_5090);
or U6886 (N_6886,N_5885,N_5697);
and U6887 (N_6887,N_5804,N_5677);
or U6888 (N_6888,N_5273,N_5876);
and U6889 (N_6889,N_5943,N_5553);
nand U6890 (N_6890,N_5042,N_5257);
and U6891 (N_6891,N_5094,N_5566);
xnor U6892 (N_6892,N_5287,N_5381);
nand U6893 (N_6893,N_5782,N_5399);
nand U6894 (N_6894,N_5220,N_5308);
nor U6895 (N_6895,N_5615,N_5410);
and U6896 (N_6896,N_5827,N_5215);
or U6897 (N_6897,N_5767,N_5512);
xor U6898 (N_6898,N_5678,N_5650);
or U6899 (N_6899,N_5117,N_5645);
or U6900 (N_6900,N_5531,N_5619);
nor U6901 (N_6901,N_5658,N_5990);
xor U6902 (N_6902,N_5990,N_5973);
or U6903 (N_6903,N_5459,N_5224);
and U6904 (N_6904,N_5659,N_5450);
nand U6905 (N_6905,N_5563,N_5577);
nor U6906 (N_6906,N_5302,N_5334);
and U6907 (N_6907,N_5753,N_5310);
and U6908 (N_6908,N_5327,N_5013);
and U6909 (N_6909,N_5116,N_5291);
nor U6910 (N_6910,N_5209,N_5719);
xor U6911 (N_6911,N_5051,N_5890);
or U6912 (N_6912,N_5944,N_5383);
nand U6913 (N_6913,N_5639,N_5834);
and U6914 (N_6914,N_5110,N_5716);
and U6915 (N_6915,N_5417,N_5180);
or U6916 (N_6916,N_5293,N_5622);
nand U6917 (N_6917,N_5487,N_5598);
and U6918 (N_6918,N_5384,N_5767);
nor U6919 (N_6919,N_5734,N_5597);
and U6920 (N_6920,N_5182,N_5002);
nor U6921 (N_6921,N_5239,N_5229);
nand U6922 (N_6922,N_5190,N_5580);
and U6923 (N_6923,N_5389,N_5403);
nor U6924 (N_6924,N_5194,N_5070);
or U6925 (N_6925,N_5373,N_5429);
nor U6926 (N_6926,N_5673,N_5763);
or U6927 (N_6927,N_5988,N_5724);
and U6928 (N_6928,N_5447,N_5776);
and U6929 (N_6929,N_5470,N_5928);
nand U6930 (N_6930,N_5578,N_5179);
or U6931 (N_6931,N_5795,N_5043);
or U6932 (N_6932,N_5836,N_5501);
nand U6933 (N_6933,N_5823,N_5100);
or U6934 (N_6934,N_5529,N_5461);
nand U6935 (N_6935,N_5482,N_5274);
nand U6936 (N_6936,N_5104,N_5169);
nand U6937 (N_6937,N_5213,N_5351);
nand U6938 (N_6938,N_5055,N_5208);
nand U6939 (N_6939,N_5010,N_5530);
and U6940 (N_6940,N_5768,N_5912);
and U6941 (N_6941,N_5345,N_5753);
nor U6942 (N_6942,N_5429,N_5799);
nor U6943 (N_6943,N_5148,N_5968);
nand U6944 (N_6944,N_5826,N_5379);
and U6945 (N_6945,N_5087,N_5304);
nor U6946 (N_6946,N_5962,N_5997);
and U6947 (N_6947,N_5375,N_5294);
and U6948 (N_6948,N_5240,N_5670);
or U6949 (N_6949,N_5949,N_5497);
or U6950 (N_6950,N_5939,N_5972);
and U6951 (N_6951,N_5220,N_5733);
nor U6952 (N_6952,N_5238,N_5870);
xor U6953 (N_6953,N_5110,N_5127);
and U6954 (N_6954,N_5710,N_5326);
and U6955 (N_6955,N_5207,N_5078);
or U6956 (N_6956,N_5739,N_5124);
or U6957 (N_6957,N_5516,N_5336);
and U6958 (N_6958,N_5414,N_5184);
nor U6959 (N_6959,N_5529,N_5652);
nor U6960 (N_6960,N_5282,N_5018);
or U6961 (N_6961,N_5543,N_5624);
nor U6962 (N_6962,N_5355,N_5811);
and U6963 (N_6963,N_5938,N_5104);
nand U6964 (N_6964,N_5403,N_5545);
and U6965 (N_6965,N_5570,N_5006);
nand U6966 (N_6966,N_5941,N_5324);
and U6967 (N_6967,N_5598,N_5334);
and U6968 (N_6968,N_5298,N_5245);
nor U6969 (N_6969,N_5964,N_5855);
nand U6970 (N_6970,N_5396,N_5462);
nand U6971 (N_6971,N_5997,N_5476);
or U6972 (N_6972,N_5500,N_5856);
nor U6973 (N_6973,N_5254,N_5758);
nand U6974 (N_6974,N_5448,N_5784);
and U6975 (N_6975,N_5841,N_5200);
nor U6976 (N_6976,N_5863,N_5739);
or U6977 (N_6977,N_5982,N_5183);
nand U6978 (N_6978,N_5961,N_5656);
nor U6979 (N_6979,N_5160,N_5159);
or U6980 (N_6980,N_5697,N_5148);
nor U6981 (N_6981,N_5431,N_5604);
xnor U6982 (N_6982,N_5129,N_5947);
nor U6983 (N_6983,N_5104,N_5965);
and U6984 (N_6984,N_5275,N_5287);
or U6985 (N_6985,N_5449,N_5911);
xor U6986 (N_6986,N_5080,N_5240);
nand U6987 (N_6987,N_5991,N_5128);
nand U6988 (N_6988,N_5195,N_5714);
nor U6989 (N_6989,N_5730,N_5284);
and U6990 (N_6990,N_5040,N_5509);
nand U6991 (N_6991,N_5772,N_5745);
nor U6992 (N_6992,N_5683,N_5876);
nand U6993 (N_6993,N_5379,N_5991);
nand U6994 (N_6994,N_5316,N_5094);
nor U6995 (N_6995,N_5618,N_5752);
and U6996 (N_6996,N_5178,N_5122);
and U6997 (N_6997,N_5160,N_5134);
and U6998 (N_6998,N_5809,N_5216);
nor U6999 (N_6999,N_5609,N_5261);
nor U7000 (N_7000,N_6271,N_6452);
nor U7001 (N_7001,N_6165,N_6614);
nor U7002 (N_7002,N_6529,N_6528);
and U7003 (N_7003,N_6938,N_6622);
nor U7004 (N_7004,N_6579,N_6182);
nand U7005 (N_7005,N_6803,N_6988);
or U7006 (N_7006,N_6467,N_6204);
nand U7007 (N_7007,N_6892,N_6355);
or U7008 (N_7008,N_6687,N_6127);
nor U7009 (N_7009,N_6461,N_6694);
nand U7010 (N_7010,N_6998,N_6218);
nor U7011 (N_7011,N_6755,N_6542);
nor U7012 (N_7012,N_6214,N_6714);
or U7013 (N_7013,N_6370,N_6860);
and U7014 (N_7014,N_6728,N_6399);
nand U7015 (N_7015,N_6572,N_6541);
nor U7016 (N_7016,N_6293,N_6014);
xnor U7017 (N_7017,N_6865,N_6914);
nor U7018 (N_7018,N_6908,N_6979);
xor U7019 (N_7019,N_6893,N_6309);
and U7020 (N_7020,N_6828,N_6344);
xor U7021 (N_7021,N_6487,N_6325);
nand U7022 (N_7022,N_6782,N_6466);
or U7023 (N_7023,N_6683,N_6984);
and U7024 (N_7024,N_6665,N_6959);
nand U7025 (N_7025,N_6157,N_6815);
nand U7026 (N_7026,N_6718,N_6457);
nor U7027 (N_7027,N_6776,N_6381);
and U7028 (N_7028,N_6846,N_6662);
nor U7029 (N_7029,N_6795,N_6703);
xnor U7030 (N_7030,N_6653,N_6296);
and U7031 (N_7031,N_6400,N_6544);
nand U7032 (N_7032,N_6581,N_6512);
and U7033 (N_7033,N_6352,N_6336);
and U7034 (N_7034,N_6033,N_6645);
and U7035 (N_7035,N_6748,N_6739);
nor U7036 (N_7036,N_6882,N_6143);
and U7037 (N_7037,N_6267,N_6691);
nand U7038 (N_7038,N_6227,N_6517);
nand U7039 (N_7039,N_6875,N_6798);
or U7040 (N_7040,N_6811,N_6278);
nor U7041 (N_7041,N_6616,N_6767);
xor U7042 (N_7042,N_6639,N_6485);
and U7043 (N_7043,N_6423,N_6345);
nor U7044 (N_7044,N_6580,N_6774);
and U7045 (N_7045,N_6824,N_6950);
or U7046 (N_7046,N_6629,N_6174);
nor U7047 (N_7047,N_6747,N_6299);
nand U7048 (N_7048,N_6900,N_6577);
and U7049 (N_7049,N_6112,N_6785);
and U7050 (N_7050,N_6131,N_6801);
and U7051 (N_7051,N_6744,N_6997);
nor U7052 (N_7052,N_6499,N_6954);
or U7053 (N_7053,N_6040,N_6897);
or U7054 (N_7054,N_6178,N_6496);
xor U7055 (N_7055,N_6362,N_6823);
or U7056 (N_7056,N_6389,N_6842);
nor U7057 (N_7057,N_6809,N_6085);
or U7058 (N_7058,N_6519,N_6151);
nand U7059 (N_7059,N_6546,N_6834);
nor U7060 (N_7060,N_6090,N_6409);
nor U7061 (N_7061,N_6565,N_6732);
nor U7062 (N_7062,N_6027,N_6664);
nor U7063 (N_7063,N_6859,N_6552);
nand U7064 (N_7064,N_6913,N_6265);
and U7065 (N_7065,N_6074,N_6205);
xnor U7066 (N_7066,N_6943,N_6874);
nand U7067 (N_7067,N_6831,N_6696);
and U7068 (N_7068,N_6030,N_6435);
nor U7069 (N_7069,N_6289,N_6987);
and U7070 (N_7070,N_6634,N_6353);
nand U7071 (N_7071,N_6092,N_6044);
and U7072 (N_7072,N_6240,N_6887);
and U7073 (N_7073,N_6695,N_6500);
or U7074 (N_7074,N_6198,N_6327);
nand U7075 (N_7075,N_6641,N_6012);
nand U7076 (N_7076,N_6369,N_6656);
nor U7077 (N_7077,N_6720,N_6920);
nand U7078 (N_7078,N_6889,N_6956);
or U7079 (N_7079,N_6319,N_6197);
and U7080 (N_7080,N_6642,N_6091);
xnor U7081 (N_7081,N_6762,N_6212);
nor U7082 (N_7082,N_6032,N_6225);
nor U7083 (N_7083,N_6095,N_6488);
and U7084 (N_7084,N_6245,N_6510);
and U7085 (N_7085,N_6312,N_6392);
and U7086 (N_7086,N_6324,N_6383);
and U7087 (N_7087,N_6810,N_6279);
and U7088 (N_7088,N_6428,N_6813);
nor U7089 (N_7089,N_6072,N_6415);
nand U7090 (N_7090,N_6193,N_6141);
and U7091 (N_7091,N_6602,N_6967);
and U7092 (N_7092,N_6019,N_6323);
nor U7093 (N_7093,N_6338,N_6612);
nor U7094 (N_7094,N_6083,N_6166);
or U7095 (N_7095,N_6374,N_6591);
and U7096 (N_7096,N_6890,N_6121);
or U7097 (N_7097,N_6560,N_6231);
or U7098 (N_7098,N_6805,N_6340);
nand U7099 (N_7099,N_6727,N_6358);
xor U7100 (N_7100,N_6750,N_6526);
and U7101 (N_7101,N_6063,N_6416);
nor U7102 (N_7102,N_6631,N_6723);
and U7103 (N_7103,N_6636,N_6162);
nor U7104 (N_7104,N_6548,N_6253);
and U7105 (N_7105,N_6351,N_6427);
nand U7106 (N_7106,N_6125,N_6754);
nand U7107 (N_7107,N_6071,N_6130);
nand U7108 (N_7108,N_6717,N_6001);
nor U7109 (N_7109,N_6903,N_6186);
xnor U7110 (N_7110,N_6497,N_6827);
xnor U7111 (N_7111,N_6473,N_6521);
nor U7112 (N_7112,N_6486,N_6758);
nand U7113 (N_7113,N_6632,N_6835);
nand U7114 (N_7114,N_6649,N_6054);
nand U7115 (N_7115,N_6465,N_6413);
or U7116 (N_7116,N_6849,N_6742);
or U7117 (N_7117,N_6094,N_6724);
nor U7118 (N_7118,N_6609,N_6244);
xor U7119 (N_7119,N_6567,N_6421);
nand U7120 (N_7120,N_6833,N_6295);
nand U7121 (N_7121,N_6553,N_6183);
nand U7122 (N_7122,N_6264,N_6707);
nor U7123 (N_7123,N_6149,N_6238);
nand U7124 (N_7124,N_6064,N_6284);
nor U7125 (N_7125,N_6224,N_6390);
and U7126 (N_7126,N_6177,N_6441);
nor U7127 (N_7127,N_6363,N_6442);
nor U7128 (N_7128,N_6453,N_6053);
and U7129 (N_7129,N_6132,N_6504);
nor U7130 (N_7130,N_6573,N_6733);
nor U7131 (N_7131,N_6076,N_6912);
and U7132 (N_7132,N_6059,N_6230);
nand U7133 (N_7133,N_6443,N_6626);
and U7134 (N_7134,N_6305,N_6765);
xor U7135 (N_7135,N_6719,N_6412);
nand U7136 (N_7136,N_6145,N_6582);
xnor U7137 (N_7137,N_6839,N_6438);
nand U7138 (N_7138,N_6450,N_6667);
nand U7139 (N_7139,N_6456,N_6140);
xor U7140 (N_7140,N_6909,N_6037);
nor U7141 (N_7141,N_6003,N_6070);
nor U7142 (N_7142,N_6069,N_6316);
or U7143 (N_7143,N_6471,N_6856);
and U7144 (N_7144,N_6304,N_6734);
xnor U7145 (N_7145,N_6953,N_6995);
nor U7146 (N_7146,N_6256,N_6712);
or U7147 (N_7147,N_6259,N_6373);
nand U7148 (N_7148,N_6797,N_6819);
and U7149 (N_7149,N_6035,N_6671);
nor U7150 (N_7150,N_6670,N_6168);
or U7151 (N_7151,N_6368,N_6966);
or U7152 (N_7152,N_6655,N_6233);
nand U7153 (N_7153,N_6398,N_6502);
nor U7154 (N_7154,N_6376,N_6922);
and U7155 (N_7155,N_6490,N_6977);
nor U7156 (N_7156,N_6690,N_6867);
nand U7157 (N_7157,N_6756,N_6692);
nand U7158 (N_7158,N_6148,N_6152);
nand U7159 (N_7159,N_6885,N_6300);
nor U7160 (N_7160,N_6679,N_6223);
xor U7161 (N_7161,N_6899,N_6705);
nor U7162 (N_7162,N_6559,N_6396);
or U7163 (N_7163,N_6023,N_6406);
nor U7164 (N_7164,N_6258,N_6713);
or U7165 (N_7165,N_6605,N_6992);
or U7166 (N_7166,N_6458,N_6429);
nor U7167 (N_7167,N_6317,N_6688);
and U7168 (N_7168,N_6120,N_6949);
xnor U7169 (N_7169,N_6587,N_6419);
nor U7170 (N_7170,N_6737,N_6968);
nor U7171 (N_7171,N_6078,N_6888);
and U7172 (N_7172,N_6270,N_6154);
and U7173 (N_7173,N_6176,N_6930);
nor U7174 (N_7174,N_6026,N_6530);
nor U7175 (N_7175,N_6880,N_6836);
xor U7176 (N_7176,N_6848,N_6958);
nor U7177 (N_7177,N_6437,N_6476);
nand U7178 (N_7178,N_6318,N_6170);
and U7179 (N_7179,N_6523,N_6247);
nand U7180 (N_7180,N_6185,N_6661);
or U7181 (N_7181,N_6303,N_6096);
xnor U7182 (N_7182,N_6901,N_6829);
nor U7183 (N_7183,N_6055,N_6147);
xnor U7184 (N_7184,N_6232,N_6320);
or U7185 (N_7185,N_6146,N_6425);
and U7186 (N_7186,N_6210,N_6886);
and U7187 (N_7187,N_6804,N_6764);
and U7188 (N_7188,N_6630,N_6161);
nor U7189 (N_7189,N_6643,N_6648);
and U7190 (N_7190,N_6098,N_6025);
and U7191 (N_7191,N_6633,N_6217);
or U7192 (N_7192,N_6432,N_6159);
nor U7193 (N_7193,N_6535,N_6329);
and U7194 (N_7194,N_6857,N_6934);
and U7195 (N_7195,N_6382,N_6640);
nor U7196 (N_7196,N_6556,N_6980);
xor U7197 (N_7197,N_6674,N_6678);
and U7198 (N_7198,N_6343,N_6547);
or U7199 (N_7199,N_6749,N_6153);
nand U7200 (N_7200,N_6575,N_6878);
xor U7201 (N_7201,N_6192,N_6701);
nand U7202 (N_7202,N_6104,N_6221);
nor U7203 (N_7203,N_6203,N_6783);
and U7204 (N_7204,N_6150,N_6771);
xnor U7205 (N_7205,N_6851,N_6472);
and U7206 (N_7206,N_6925,N_6698);
or U7207 (N_7207,N_6013,N_6468);
nand U7208 (N_7208,N_6790,N_6781);
nor U7209 (N_7209,N_6464,N_6761);
or U7210 (N_7210,N_6113,N_6326);
nor U7211 (N_7211,N_6584,N_6711);
nor U7212 (N_7212,N_6501,N_6211);
and U7213 (N_7213,N_6016,N_6593);
nand U7214 (N_7214,N_6179,N_6778);
xnor U7215 (N_7215,N_6847,N_6672);
nand U7216 (N_7216,N_6024,N_6613);
xnor U7217 (N_7217,N_6226,N_6481);
nand U7218 (N_7218,N_6566,N_6290);
and U7219 (N_7219,N_6955,N_6298);
or U7220 (N_7220,N_6377,N_6974);
and U7221 (N_7221,N_6628,N_6163);
nor U7222 (N_7222,N_6236,N_6272);
or U7223 (N_7223,N_6422,N_6619);
nand U7224 (N_7224,N_6917,N_6963);
and U7225 (N_7225,N_6038,N_6763);
or U7226 (N_7226,N_6511,N_6136);
and U7227 (N_7227,N_6855,N_6638);
and U7228 (N_7228,N_6342,N_6050);
nor U7229 (N_7229,N_6410,N_6248);
and U7230 (N_7230,N_6215,N_6015);
nand U7231 (N_7231,N_6283,N_6460);
nor U7232 (N_7232,N_6818,N_6328);
or U7233 (N_7233,N_6424,N_6492);
and U7234 (N_7234,N_6905,N_6172);
nor U7235 (N_7235,N_6725,N_6589);
and U7236 (N_7236,N_6624,N_6077);
and U7237 (N_7237,N_6650,N_6620);
and U7238 (N_7238,N_6503,N_6550);
or U7239 (N_7239,N_6845,N_6594);
or U7240 (N_7240,N_6516,N_6455);
nand U7241 (N_7241,N_6266,N_6364);
and U7242 (N_7242,N_6869,N_6598);
nand U7243 (N_7243,N_6787,N_6658);
xor U7244 (N_7244,N_6103,N_6046);
and U7245 (N_7245,N_6757,N_6005);
or U7246 (N_7246,N_6056,N_6234);
and U7247 (N_7247,N_6135,N_6359);
nand U7248 (N_7248,N_6534,N_6447);
or U7249 (N_7249,N_6983,N_6099);
and U7250 (N_7250,N_6181,N_6647);
nor U7251 (N_7251,N_6796,N_6372);
and U7252 (N_7252,N_6506,N_6693);
nand U7253 (N_7253,N_6902,N_6876);
nand U7254 (N_7254,N_6538,N_6107);
nor U7255 (N_7255,N_6375,N_6404);
nand U7256 (N_7256,N_6208,N_6000);
or U7257 (N_7257,N_6239,N_6669);
or U7258 (N_7258,N_6576,N_6307);
and U7259 (N_7259,N_6898,N_6254);
or U7260 (N_7260,N_6514,N_6426);
xor U7261 (N_7261,N_6607,N_6479);
and U7262 (N_7262,N_6606,N_6866);
nand U7263 (N_7263,N_6923,N_6268);
nor U7264 (N_7264,N_6926,N_6101);
or U7265 (N_7265,N_6011,N_6568);
or U7266 (N_7266,N_6525,N_6219);
nor U7267 (N_7267,N_6405,N_6189);
nor U7268 (N_7268,N_6387,N_6929);
nor U7269 (N_7269,N_6445,N_6483);
nand U7270 (N_7270,N_6508,N_6142);
nand U7271 (N_7271,N_6623,N_6513);
nor U7272 (N_7272,N_6228,N_6291);
xor U7273 (N_7273,N_6985,N_6021);
nand U7274 (N_7274,N_6518,N_6562);
nand U7275 (N_7275,N_6947,N_6816);
or U7276 (N_7276,N_6944,N_6989);
and U7277 (N_7277,N_6388,N_6158);
and U7278 (N_7278,N_6294,N_6574);
or U7279 (N_7279,N_6052,N_6666);
and U7280 (N_7280,N_6333,N_6608);
nand U7281 (N_7281,N_6615,N_6675);
and U7282 (N_7282,N_6039,N_6124);
nand U7283 (N_7283,N_6596,N_6561);
xor U7284 (N_7284,N_6524,N_6741);
nand U7285 (N_7285,N_6451,N_6600);
nand U7286 (N_7286,N_6117,N_6792);
xnor U7287 (N_7287,N_6332,N_6420);
nor U7288 (N_7288,N_6459,N_6814);
nand U7289 (N_7289,N_6837,N_6079);
nor U7290 (N_7290,N_6306,N_6663);
nor U7291 (N_7291,N_6180,N_6122);
nand U7292 (N_7292,N_6269,N_6048);
xnor U7293 (N_7293,N_6433,N_6945);
nor U7294 (N_7294,N_6061,N_6031);
nor U7295 (N_7295,N_6872,N_6206);
and U7296 (N_7296,N_6682,N_6277);
nor U7297 (N_7297,N_6430,N_6708);
and U7298 (N_7298,N_6769,N_6060);
xnor U7299 (N_7299,N_6993,N_6106);
and U7300 (N_7300,N_6273,N_6991);
or U7301 (N_7301,N_6007,N_6788);
and U7302 (N_7302,N_6540,N_6474);
and U7303 (N_7303,N_6794,N_6111);
or U7304 (N_7304,N_6262,N_6209);
nor U7305 (N_7305,N_6196,N_6093);
nor U7306 (N_7306,N_6173,N_6604);
or U7307 (N_7307,N_6384,N_6380);
and U7308 (N_7308,N_6557,N_6895);
nor U7309 (N_7309,N_6082,N_6928);
and U7310 (N_7310,N_6285,N_6951);
or U7311 (N_7311,N_6924,N_6042);
and U7312 (N_7312,N_6004,N_6644);
or U7313 (N_7313,N_6578,N_6617);
xor U7314 (N_7314,N_6393,N_6799);
nor U7315 (N_7315,N_6652,N_6213);
xnor U7316 (N_7316,N_6657,N_6469);
nand U7317 (N_7317,N_6558,N_6873);
xnor U7318 (N_7318,N_6356,N_6879);
nor U7319 (N_7319,N_6462,N_6709);
nor U7320 (N_7320,N_6041,N_6097);
or U7321 (N_7321,N_6759,N_6454);
nand U7322 (N_7322,N_6791,N_6896);
nand U7323 (N_7323,N_6821,N_6676);
xnor U7324 (N_7324,N_6417,N_6569);
nor U7325 (N_7325,N_6721,N_6366);
or U7326 (N_7326,N_6302,N_6864);
nand U7327 (N_7327,N_6118,N_6049);
xor U7328 (N_7328,N_6108,N_6337);
or U7329 (N_7329,N_6301,N_6706);
nand U7330 (N_7330,N_6965,N_6820);
nand U7331 (N_7331,N_6841,N_6123);
and U7332 (N_7332,N_6697,N_6745);
nand U7333 (N_7333,N_6507,N_6618);
or U7334 (N_7334,N_6736,N_6017);
or U7335 (N_7335,N_6137,N_6431);
nand U7336 (N_7336,N_6981,N_6806);
nor U7337 (N_7337,N_6884,N_6844);
and U7338 (N_7338,N_6116,N_6347);
and U7339 (N_7339,N_6308,N_6190);
nor U7340 (N_7340,N_6766,N_6590);
nand U7341 (N_7341,N_6365,N_6686);
nand U7342 (N_7342,N_6493,N_6971);
or U7343 (N_7343,N_6463,N_6635);
nor U7344 (N_7344,N_6379,N_6952);
and U7345 (N_7345,N_6187,N_6539);
nand U7346 (N_7346,N_6537,N_6045);
nor U7347 (N_7347,N_6020,N_6843);
and U7348 (N_7348,N_6029,N_6969);
nor U7349 (N_7349,N_6793,N_6065);
and U7350 (N_7350,N_6401,N_6200);
nor U7351 (N_7351,N_6941,N_6339);
nor U7352 (N_7352,N_6034,N_6036);
nand U7353 (N_7353,N_6109,N_6348);
and U7354 (N_7354,N_6659,N_6222);
nor U7355 (N_7355,N_6910,N_6704);
or U7356 (N_7356,N_6940,N_6973);
and U7357 (N_7357,N_6354,N_6982);
nand U7358 (N_7358,N_6868,N_6533);
nand U7359 (N_7359,N_6395,N_6436);
nor U7360 (N_7360,N_6391,N_6440);
or U7361 (N_7361,N_6194,N_6775);
or U7362 (N_7362,N_6660,N_6861);
nor U7363 (N_7363,N_6449,N_6826);
and U7364 (N_7364,N_6780,N_6891);
nor U7365 (N_7365,N_6768,N_6164);
or U7366 (N_7366,N_6066,N_6853);
and U7367 (N_7367,N_6532,N_6681);
xnor U7368 (N_7368,N_6087,N_6047);
and U7369 (N_7369,N_6509,N_6838);
and U7370 (N_7370,N_6010,N_6314);
nor U7371 (N_7371,N_6946,N_6731);
nand U7372 (N_7372,N_6084,N_6018);
nand U7373 (N_7373,N_6119,N_6904);
nor U7374 (N_7374,N_6520,N_6330);
nand U7375 (N_7375,N_6089,N_6331);
nand U7376 (N_7376,N_6832,N_6994);
nor U7377 (N_7377,N_6716,N_6760);
nor U7378 (N_7378,N_6321,N_6505);
nand U7379 (N_7379,N_6729,N_6478);
or U7380 (N_7380,N_6522,N_6699);
or U7381 (N_7381,N_6184,N_6482);
or U7382 (N_7382,N_6752,N_6877);
nand U7383 (N_7383,N_6102,N_6543);
nor U7384 (N_7384,N_6651,N_6527);
nand U7385 (N_7385,N_6397,N_6073);
nand U7386 (N_7386,N_6175,N_6939);
nand U7387 (N_7387,N_6009,N_6646);
nor U7388 (N_7388,N_6545,N_6188);
and U7389 (N_7389,N_6075,N_6942);
or U7390 (N_7390,N_6583,N_6255);
nand U7391 (N_7391,N_6601,N_6536);
xor U7392 (N_7392,N_6549,N_6281);
nand U7393 (N_7393,N_6160,N_6571);
nor U7394 (N_7394,N_6680,N_6685);
or U7395 (N_7395,N_6080,N_6414);
or U7396 (N_7396,N_6260,N_6726);
nand U7397 (N_7397,N_6110,N_6779);
and U7398 (N_7398,N_6126,N_6241);
or U7399 (N_7399,N_6207,N_6371);
nor U7400 (N_7400,N_6385,N_6555);
xor U7401 (N_7401,N_6246,N_6280);
or U7402 (N_7402,N_6439,N_6274);
and U7403 (N_7403,N_6134,N_6169);
or U7404 (N_7404,N_6297,N_6250);
or U7405 (N_7405,N_6057,N_6599);
nor U7406 (N_7406,N_6022,N_6006);
and U7407 (N_7407,N_6933,N_6677);
nor U7408 (N_7408,N_6961,N_6751);
nand U7409 (N_7409,N_6144,N_6216);
nand U7410 (N_7410,N_6081,N_6171);
nand U7411 (N_7411,N_6100,N_6770);
nand U7412 (N_7412,N_6287,N_6883);
and U7413 (N_7413,N_6715,N_6588);
or U7414 (N_7414,N_6852,N_6251);
or U7415 (N_7415,N_6315,N_6911);
nand U7416 (N_7416,N_6915,N_6585);
or U7417 (N_7417,N_6722,N_6978);
nand U7418 (N_7418,N_6480,N_6043);
nand U7419 (N_7419,N_6777,N_6288);
or U7420 (N_7420,N_6921,N_6341);
and U7421 (N_7421,N_6964,N_6361);
nand U7422 (N_7422,N_6700,N_6403);
nor U7423 (N_7423,N_6554,N_6970);
nand U7424 (N_7424,N_6948,N_6346);
nor U7425 (N_7425,N_6531,N_6470);
nand U7426 (N_7426,N_6411,N_6444);
nor U7427 (N_7427,N_6935,N_6062);
nor U7428 (N_7428,N_6962,N_6475);
and U7429 (N_7429,N_6282,N_6802);
or U7430 (N_7430,N_6907,N_6067);
nor U7431 (N_7431,N_6990,N_6916);
nor U7432 (N_7432,N_6932,N_6199);
and U7433 (N_7433,N_6275,N_6919);
nand U7434 (N_7434,N_6972,N_6495);
or U7435 (N_7435,N_6394,N_6261);
nand U7436 (N_7436,N_6105,N_6570);
nor U7437 (N_7437,N_6863,N_6220);
nor U7438 (N_7438,N_6386,N_6367);
and U7439 (N_7439,N_6957,N_6931);
nand U7440 (N_7440,N_6894,N_6051);
nand U7441 (N_7441,N_6237,N_6133);
and U7442 (N_7442,N_6322,N_6229);
nand U7443 (N_7443,N_6310,N_6286);
nand U7444 (N_7444,N_6800,N_6592);
nand U7445 (N_7445,N_6689,N_6918);
nor U7446 (N_7446,N_6292,N_6746);
and U7447 (N_7447,N_6871,N_6937);
nand U7448 (N_7448,N_6668,N_6448);
nor U7449 (N_7449,N_6128,N_6350);
and U7450 (N_7450,N_6378,N_6881);
nand U7451 (N_7451,N_6335,N_6976);
or U7452 (N_7452,N_6595,N_6167);
nand U7453 (N_7453,N_6975,N_6515);
nand U7454 (N_7454,N_6654,N_6418);
nand U7455 (N_7455,N_6434,N_6008);
nor U7456 (N_7456,N_6407,N_6563);
and U7457 (N_7457,N_6202,N_6743);
nor U7458 (N_7458,N_6586,N_6195);
or U7459 (N_7459,N_6738,N_6772);
and U7460 (N_7460,N_6673,N_6812);
nand U7461 (N_7461,N_6597,N_6357);
nor U7462 (N_7462,N_6817,N_6242);
xor U7463 (N_7463,N_6002,N_6627);
and U7464 (N_7464,N_6276,N_6927);
or U7465 (N_7465,N_6408,N_6201);
nor U7466 (N_7466,N_6784,N_6257);
and U7467 (N_7467,N_6611,N_6960);
nand U7468 (N_7468,N_6789,N_6730);
or U7469 (N_7469,N_6807,N_6625);
and U7470 (N_7470,N_6491,N_6786);
nand U7471 (N_7471,N_6610,N_6138);
or U7472 (N_7472,N_6773,N_6360);
nand U7473 (N_7473,N_6477,N_6735);
or U7474 (N_7474,N_6058,N_6139);
or U7475 (N_7475,N_6621,N_6252);
nor U7476 (N_7476,N_6740,N_6999);
or U7477 (N_7477,N_6936,N_6840);
nor U7478 (N_7478,N_6822,N_6808);
and U7479 (N_7479,N_6484,N_6862);
nor U7480 (N_7480,N_6446,N_6068);
or U7481 (N_7481,N_6086,N_6996);
and U7482 (N_7482,N_6710,N_6830);
nand U7483 (N_7483,N_6854,N_6129);
xor U7484 (N_7484,N_6564,N_6603);
or U7485 (N_7485,N_6191,N_6088);
xnor U7486 (N_7486,N_6156,N_6551);
nor U7487 (N_7487,N_6235,N_6334);
or U7488 (N_7488,N_6311,N_6313);
xnor U7489 (N_7489,N_6115,N_6243);
xnor U7490 (N_7490,N_6858,N_6263);
nand U7491 (N_7491,N_6249,N_6702);
nor U7492 (N_7492,N_6870,N_6825);
and U7493 (N_7493,N_6114,N_6494);
nor U7494 (N_7494,N_6637,N_6349);
nor U7495 (N_7495,N_6489,N_6986);
and U7496 (N_7496,N_6906,N_6498);
nand U7497 (N_7497,N_6850,N_6402);
and U7498 (N_7498,N_6753,N_6028);
or U7499 (N_7499,N_6155,N_6684);
nand U7500 (N_7500,N_6110,N_6212);
or U7501 (N_7501,N_6759,N_6090);
nand U7502 (N_7502,N_6597,N_6322);
nor U7503 (N_7503,N_6316,N_6999);
nand U7504 (N_7504,N_6273,N_6376);
and U7505 (N_7505,N_6639,N_6575);
and U7506 (N_7506,N_6191,N_6764);
or U7507 (N_7507,N_6671,N_6408);
nand U7508 (N_7508,N_6146,N_6610);
nor U7509 (N_7509,N_6663,N_6987);
nand U7510 (N_7510,N_6381,N_6575);
nand U7511 (N_7511,N_6964,N_6241);
nor U7512 (N_7512,N_6815,N_6666);
or U7513 (N_7513,N_6099,N_6003);
and U7514 (N_7514,N_6260,N_6155);
or U7515 (N_7515,N_6647,N_6624);
xnor U7516 (N_7516,N_6460,N_6007);
nand U7517 (N_7517,N_6784,N_6873);
xnor U7518 (N_7518,N_6684,N_6611);
xnor U7519 (N_7519,N_6558,N_6470);
nand U7520 (N_7520,N_6503,N_6038);
nand U7521 (N_7521,N_6863,N_6159);
xnor U7522 (N_7522,N_6741,N_6645);
and U7523 (N_7523,N_6077,N_6849);
or U7524 (N_7524,N_6102,N_6729);
nand U7525 (N_7525,N_6996,N_6071);
and U7526 (N_7526,N_6445,N_6472);
or U7527 (N_7527,N_6622,N_6731);
and U7528 (N_7528,N_6291,N_6264);
nor U7529 (N_7529,N_6753,N_6872);
or U7530 (N_7530,N_6671,N_6833);
and U7531 (N_7531,N_6975,N_6891);
or U7532 (N_7532,N_6386,N_6555);
nor U7533 (N_7533,N_6021,N_6214);
or U7534 (N_7534,N_6695,N_6918);
nor U7535 (N_7535,N_6468,N_6481);
nor U7536 (N_7536,N_6534,N_6307);
nand U7537 (N_7537,N_6098,N_6791);
or U7538 (N_7538,N_6991,N_6740);
and U7539 (N_7539,N_6697,N_6533);
and U7540 (N_7540,N_6770,N_6182);
and U7541 (N_7541,N_6175,N_6316);
or U7542 (N_7542,N_6137,N_6539);
and U7543 (N_7543,N_6007,N_6223);
and U7544 (N_7544,N_6443,N_6387);
or U7545 (N_7545,N_6885,N_6535);
nand U7546 (N_7546,N_6194,N_6542);
or U7547 (N_7547,N_6058,N_6264);
nor U7548 (N_7548,N_6617,N_6293);
or U7549 (N_7549,N_6014,N_6004);
nand U7550 (N_7550,N_6406,N_6072);
nand U7551 (N_7551,N_6619,N_6755);
nor U7552 (N_7552,N_6026,N_6985);
and U7553 (N_7553,N_6041,N_6603);
nand U7554 (N_7554,N_6284,N_6565);
nor U7555 (N_7555,N_6052,N_6132);
nand U7556 (N_7556,N_6514,N_6435);
nor U7557 (N_7557,N_6198,N_6069);
nor U7558 (N_7558,N_6384,N_6863);
nand U7559 (N_7559,N_6838,N_6548);
nor U7560 (N_7560,N_6737,N_6498);
nor U7561 (N_7561,N_6477,N_6856);
nand U7562 (N_7562,N_6486,N_6291);
nor U7563 (N_7563,N_6016,N_6840);
or U7564 (N_7564,N_6821,N_6948);
nand U7565 (N_7565,N_6601,N_6458);
or U7566 (N_7566,N_6556,N_6965);
and U7567 (N_7567,N_6317,N_6048);
nand U7568 (N_7568,N_6335,N_6449);
and U7569 (N_7569,N_6999,N_6800);
nor U7570 (N_7570,N_6033,N_6854);
and U7571 (N_7571,N_6734,N_6709);
nand U7572 (N_7572,N_6863,N_6083);
and U7573 (N_7573,N_6700,N_6852);
nand U7574 (N_7574,N_6096,N_6228);
nand U7575 (N_7575,N_6523,N_6646);
xor U7576 (N_7576,N_6906,N_6307);
and U7577 (N_7577,N_6837,N_6033);
or U7578 (N_7578,N_6965,N_6423);
or U7579 (N_7579,N_6017,N_6621);
or U7580 (N_7580,N_6918,N_6917);
and U7581 (N_7581,N_6688,N_6906);
nor U7582 (N_7582,N_6917,N_6870);
nand U7583 (N_7583,N_6365,N_6079);
nand U7584 (N_7584,N_6731,N_6113);
and U7585 (N_7585,N_6949,N_6191);
or U7586 (N_7586,N_6135,N_6410);
or U7587 (N_7587,N_6485,N_6504);
nand U7588 (N_7588,N_6553,N_6800);
nor U7589 (N_7589,N_6167,N_6438);
and U7590 (N_7590,N_6464,N_6406);
nand U7591 (N_7591,N_6207,N_6307);
nand U7592 (N_7592,N_6783,N_6189);
nor U7593 (N_7593,N_6423,N_6638);
nor U7594 (N_7594,N_6597,N_6027);
and U7595 (N_7595,N_6968,N_6388);
nor U7596 (N_7596,N_6114,N_6587);
nand U7597 (N_7597,N_6523,N_6593);
nand U7598 (N_7598,N_6201,N_6951);
and U7599 (N_7599,N_6990,N_6533);
xor U7600 (N_7600,N_6771,N_6938);
or U7601 (N_7601,N_6509,N_6791);
and U7602 (N_7602,N_6132,N_6491);
nand U7603 (N_7603,N_6329,N_6352);
and U7604 (N_7604,N_6193,N_6948);
nand U7605 (N_7605,N_6986,N_6494);
nor U7606 (N_7606,N_6540,N_6558);
nor U7607 (N_7607,N_6125,N_6359);
nor U7608 (N_7608,N_6050,N_6652);
xnor U7609 (N_7609,N_6446,N_6733);
and U7610 (N_7610,N_6271,N_6900);
nand U7611 (N_7611,N_6428,N_6729);
and U7612 (N_7612,N_6097,N_6083);
nor U7613 (N_7613,N_6118,N_6900);
nand U7614 (N_7614,N_6062,N_6401);
and U7615 (N_7615,N_6486,N_6557);
nand U7616 (N_7616,N_6779,N_6365);
and U7617 (N_7617,N_6035,N_6362);
and U7618 (N_7618,N_6058,N_6861);
nand U7619 (N_7619,N_6685,N_6290);
and U7620 (N_7620,N_6365,N_6880);
and U7621 (N_7621,N_6540,N_6054);
and U7622 (N_7622,N_6252,N_6985);
nand U7623 (N_7623,N_6997,N_6884);
and U7624 (N_7624,N_6066,N_6700);
nand U7625 (N_7625,N_6798,N_6707);
and U7626 (N_7626,N_6008,N_6592);
xnor U7627 (N_7627,N_6811,N_6975);
or U7628 (N_7628,N_6343,N_6749);
or U7629 (N_7629,N_6813,N_6006);
or U7630 (N_7630,N_6433,N_6999);
or U7631 (N_7631,N_6809,N_6652);
xor U7632 (N_7632,N_6609,N_6527);
and U7633 (N_7633,N_6843,N_6996);
nand U7634 (N_7634,N_6863,N_6826);
nand U7635 (N_7635,N_6815,N_6550);
and U7636 (N_7636,N_6921,N_6335);
nor U7637 (N_7637,N_6970,N_6226);
nor U7638 (N_7638,N_6327,N_6834);
or U7639 (N_7639,N_6002,N_6217);
nand U7640 (N_7640,N_6960,N_6883);
or U7641 (N_7641,N_6974,N_6975);
or U7642 (N_7642,N_6873,N_6928);
and U7643 (N_7643,N_6155,N_6821);
nand U7644 (N_7644,N_6688,N_6024);
nor U7645 (N_7645,N_6026,N_6148);
xor U7646 (N_7646,N_6818,N_6816);
nand U7647 (N_7647,N_6751,N_6502);
nor U7648 (N_7648,N_6696,N_6903);
nor U7649 (N_7649,N_6004,N_6655);
and U7650 (N_7650,N_6328,N_6693);
nand U7651 (N_7651,N_6790,N_6697);
or U7652 (N_7652,N_6644,N_6380);
xor U7653 (N_7653,N_6116,N_6639);
xor U7654 (N_7654,N_6100,N_6211);
nor U7655 (N_7655,N_6439,N_6401);
and U7656 (N_7656,N_6175,N_6686);
nor U7657 (N_7657,N_6032,N_6643);
nand U7658 (N_7658,N_6602,N_6043);
and U7659 (N_7659,N_6573,N_6980);
and U7660 (N_7660,N_6451,N_6739);
nor U7661 (N_7661,N_6897,N_6143);
and U7662 (N_7662,N_6979,N_6404);
nor U7663 (N_7663,N_6880,N_6386);
nand U7664 (N_7664,N_6006,N_6161);
and U7665 (N_7665,N_6146,N_6668);
nor U7666 (N_7666,N_6552,N_6212);
and U7667 (N_7667,N_6009,N_6353);
or U7668 (N_7668,N_6615,N_6673);
nand U7669 (N_7669,N_6216,N_6801);
or U7670 (N_7670,N_6326,N_6156);
nor U7671 (N_7671,N_6500,N_6429);
nor U7672 (N_7672,N_6586,N_6423);
nor U7673 (N_7673,N_6564,N_6360);
and U7674 (N_7674,N_6413,N_6837);
nand U7675 (N_7675,N_6843,N_6679);
and U7676 (N_7676,N_6812,N_6575);
nand U7677 (N_7677,N_6903,N_6796);
nor U7678 (N_7678,N_6255,N_6990);
xor U7679 (N_7679,N_6508,N_6758);
nand U7680 (N_7680,N_6338,N_6839);
nor U7681 (N_7681,N_6115,N_6502);
and U7682 (N_7682,N_6035,N_6796);
nor U7683 (N_7683,N_6058,N_6527);
or U7684 (N_7684,N_6703,N_6884);
nor U7685 (N_7685,N_6658,N_6156);
nor U7686 (N_7686,N_6641,N_6851);
and U7687 (N_7687,N_6210,N_6509);
or U7688 (N_7688,N_6511,N_6480);
xnor U7689 (N_7689,N_6992,N_6878);
or U7690 (N_7690,N_6633,N_6109);
and U7691 (N_7691,N_6804,N_6119);
or U7692 (N_7692,N_6150,N_6684);
or U7693 (N_7693,N_6387,N_6432);
nand U7694 (N_7694,N_6131,N_6959);
nand U7695 (N_7695,N_6059,N_6767);
nand U7696 (N_7696,N_6985,N_6343);
xor U7697 (N_7697,N_6264,N_6279);
or U7698 (N_7698,N_6708,N_6775);
or U7699 (N_7699,N_6634,N_6942);
nand U7700 (N_7700,N_6108,N_6186);
and U7701 (N_7701,N_6041,N_6486);
and U7702 (N_7702,N_6601,N_6790);
xor U7703 (N_7703,N_6709,N_6507);
nand U7704 (N_7704,N_6655,N_6574);
or U7705 (N_7705,N_6278,N_6876);
nand U7706 (N_7706,N_6683,N_6864);
nand U7707 (N_7707,N_6316,N_6500);
or U7708 (N_7708,N_6559,N_6737);
or U7709 (N_7709,N_6944,N_6353);
nor U7710 (N_7710,N_6234,N_6646);
nor U7711 (N_7711,N_6849,N_6555);
or U7712 (N_7712,N_6455,N_6242);
and U7713 (N_7713,N_6294,N_6073);
nor U7714 (N_7714,N_6412,N_6919);
or U7715 (N_7715,N_6367,N_6646);
nor U7716 (N_7716,N_6518,N_6204);
and U7717 (N_7717,N_6534,N_6484);
or U7718 (N_7718,N_6463,N_6273);
and U7719 (N_7719,N_6236,N_6313);
xor U7720 (N_7720,N_6776,N_6648);
xnor U7721 (N_7721,N_6494,N_6048);
or U7722 (N_7722,N_6411,N_6718);
nand U7723 (N_7723,N_6153,N_6824);
or U7724 (N_7724,N_6893,N_6239);
xor U7725 (N_7725,N_6533,N_6407);
and U7726 (N_7726,N_6190,N_6861);
nor U7727 (N_7727,N_6036,N_6829);
nand U7728 (N_7728,N_6556,N_6271);
xnor U7729 (N_7729,N_6106,N_6823);
and U7730 (N_7730,N_6043,N_6346);
nand U7731 (N_7731,N_6785,N_6683);
nand U7732 (N_7732,N_6152,N_6605);
nand U7733 (N_7733,N_6297,N_6452);
nor U7734 (N_7734,N_6522,N_6348);
nor U7735 (N_7735,N_6150,N_6820);
nand U7736 (N_7736,N_6530,N_6615);
nor U7737 (N_7737,N_6780,N_6145);
nand U7738 (N_7738,N_6819,N_6332);
nor U7739 (N_7739,N_6477,N_6375);
and U7740 (N_7740,N_6998,N_6470);
xnor U7741 (N_7741,N_6399,N_6145);
xnor U7742 (N_7742,N_6979,N_6249);
xor U7743 (N_7743,N_6266,N_6057);
and U7744 (N_7744,N_6347,N_6613);
or U7745 (N_7745,N_6159,N_6219);
nor U7746 (N_7746,N_6842,N_6194);
nand U7747 (N_7747,N_6123,N_6896);
nor U7748 (N_7748,N_6980,N_6371);
nor U7749 (N_7749,N_6379,N_6617);
and U7750 (N_7750,N_6943,N_6801);
nand U7751 (N_7751,N_6614,N_6673);
nor U7752 (N_7752,N_6416,N_6445);
nor U7753 (N_7753,N_6967,N_6834);
and U7754 (N_7754,N_6921,N_6725);
nand U7755 (N_7755,N_6008,N_6802);
or U7756 (N_7756,N_6759,N_6224);
nor U7757 (N_7757,N_6165,N_6785);
nand U7758 (N_7758,N_6373,N_6822);
nand U7759 (N_7759,N_6530,N_6434);
xor U7760 (N_7760,N_6290,N_6472);
nand U7761 (N_7761,N_6253,N_6709);
nand U7762 (N_7762,N_6979,N_6347);
nor U7763 (N_7763,N_6830,N_6199);
or U7764 (N_7764,N_6339,N_6277);
xnor U7765 (N_7765,N_6944,N_6186);
nor U7766 (N_7766,N_6308,N_6309);
nand U7767 (N_7767,N_6023,N_6352);
nand U7768 (N_7768,N_6240,N_6493);
nor U7769 (N_7769,N_6182,N_6265);
nor U7770 (N_7770,N_6089,N_6045);
nand U7771 (N_7771,N_6946,N_6600);
nor U7772 (N_7772,N_6622,N_6226);
nand U7773 (N_7773,N_6624,N_6178);
nand U7774 (N_7774,N_6069,N_6835);
and U7775 (N_7775,N_6564,N_6151);
nor U7776 (N_7776,N_6542,N_6802);
and U7777 (N_7777,N_6271,N_6703);
or U7778 (N_7778,N_6540,N_6467);
nor U7779 (N_7779,N_6414,N_6945);
and U7780 (N_7780,N_6909,N_6255);
xnor U7781 (N_7781,N_6917,N_6885);
xor U7782 (N_7782,N_6489,N_6996);
or U7783 (N_7783,N_6691,N_6855);
nor U7784 (N_7784,N_6517,N_6963);
and U7785 (N_7785,N_6047,N_6615);
and U7786 (N_7786,N_6462,N_6602);
nor U7787 (N_7787,N_6595,N_6726);
or U7788 (N_7788,N_6943,N_6490);
nand U7789 (N_7789,N_6065,N_6708);
and U7790 (N_7790,N_6441,N_6325);
xor U7791 (N_7791,N_6049,N_6715);
or U7792 (N_7792,N_6685,N_6164);
or U7793 (N_7793,N_6618,N_6547);
or U7794 (N_7794,N_6121,N_6760);
nand U7795 (N_7795,N_6458,N_6702);
nor U7796 (N_7796,N_6412,N_6334);
nand U7797 (N_7797,N_6549,N_6914);
nor U7798 (N_7798,N_6105,N_6125);
nand U7799 (N_7799,N_6039,N_6791);
nor U7800 (N_7800,N_6268,N_6935);
nand U7801 (N_7801,N_6801,N_6008);
and U7802 (N_7802,N_6006,N_6636);
nor U7803 (N_7803,N_6124,N_6943);
nor U7804 (N_7804,N_6808,N_6825);
and U7805 (N_7805,N_6775,N_6374);
nand U7806 (N_7806,N_6450,N_6211);
nand U7807 (N_7807,N_6781,N_6082);
or U7808 (N_7808,N_6163,N_6269);
nor U7809 (N_7809,N_6637,N_6776);
nand U7810 (N_7810,N_6056,N_6426);
and U7811 (N_7811,N_6526,N_6712);
nor U7812 (N_7812,N_6738,N_6538);
and U7813 (N_7813,N_6622,N_6503);
or U7814 (N_7814,N_6660,N_6894);
nand U7815 (N_7815,N_6255,N_6219);
and U7816 (N_7816,N_6714,N_6968);
and U7817 (N_7817,N_6522,N_6184);
and U7818 (N_7818,N_6029,N_6276);
or U7819 (N_7819,N_6710,N_6875);
nor U7820 (N_7820,N_6224,N_6988);
nor U7821 (N_7821,N_6999,N_6271);
nor U7822 (N_7822,N_6685,N_6923);
nor U7823 (N_7823,N_6306,N_6033);
nand U7824 (N_7824,N_6434,N_6754);
and U7825 (N_7825,N_6921,N_6710);
nor U7826 (N_7826,N_6248,N_6368);
and U7827 (N_7827,N_6536,N_6426);
or U7828 (N_7828,N_6152,N_6374);
and U7829 (N_7829,N_6304,N_6851);
nand U7830 (N_7830,N_6240,N_6271);
and U7831 (N_7831,N_6010,N_6272);
and U7832 (N_7832,N_6832,N_6027);
or U7833 (N_7833,N_6404,N_6275);
nand U7834 (N_7834,N_6974,N_6684);
or U7835 (N_7835,N_6405,N_6667);
nand U7836 (N_7836,N_6116,N_6925);
or U7837 (N_7837,N_6877,N_6443);
and U7838 (N_7838,N_6823,N_6847);
and U7839 (N_7839,N_6776,N_6874);
and U7840 (N_7840,N_6573,N_6299);
or U7841 (N_7841,N_6242,N_6449);
and U7842 (N_7842,N_6291,N_6950);
nand U7843 (N_7843,N_6428,N_6563);
nor U7844 (N_7844,N_6869,N_6516);
and U7845 (N_7845,N_6503,N_6991);
or U7846 (N_7846,N_6980,N_6636);
nand U7847 (N_7847,N_6083,N_6215);
nand U7848 (N_7848,N_6130,N_6769);
or U7849 (N_7849,N_6233,N_6148);
and U7850 (N_7850,N_6561,N_6120);
or U7851 (N_7851,N_6737,N_6007);
or U7852 (N_7852,N_6539,N_6085);
nand U7853 (N_7853,N_6762,N_6797);
and U7854 (N_7854,N_6500,N_6990);
nor U7855 (N_7855,N_6387,N_6225);
nand U7856 (N_7856,N_6768,N_6890);
or U7857 (N_7857,N_6188,N_6670);
nor U7858 (N_7858,N_6852,N_6711);
and U7859 (N_7859,N_6971,N_6912);
nand U7860 (N_7860,N_6596,N_6872);
nand U7861 (N_7861,N_6471,N_6937);
nor U7862 (N_7862,N_6596,N_6369);
nand U7863 (N_7863,N_6172,N_6731);
nand U7864 (N_7864,N_6716,N_6330);
xnor U7865 (N_7865,N_6338,N_6103);
and U7866 (N_7866,N_6322,N_6214);
or U7867 (N_7867,N_6581,N_6396);
nor U7868 (N_7868,N_6921,N_6212);
and U7869 (N_7869,N_6924,N_6216);
nor U7870 (N_7870,N_6345,N_6598);
nand U7871 (N_7871,N_6360,N_6314);
nand U7872 (N_7872,N_6971,N_6856);
or U7873 (N_7873,N_6527,N_6213);
nor U7874 (N_7874,N_6379,N_6183);
nor U7875 (N_7875,N_6404,N_6830);
and U7876 (N_7876,N_6561,N_6348);
nor U7877 (N_7877,N_6652,N_6695);
or U7878 (N_7878,N_6824,N_6861);
nand U7879 (N_7879,N_6570,N_6163);
nor U7880 (N_7880,N_6827,N_6756);
nor U7881 (N_7881,N_6841,N_6101);
nand U7882 (N_7882,N_6144,N_6095);
and U7883 (N_7883,N_6543,N_6219);
or U7884 (N_7884,N_6937,N_6553);
nor U7885 (N_7885,N_6650,N_6081);
nor U7886 (N_7886,N_6024,N_6267);
and U7887 (N_7887,N_6805,N_6342);
nand U7888 (N_7888,N_6170,N_6247);
and U7889 (N_7889,N_6304,N_6932);
and U7890 (N_7890,N_6592,N_6323);
and U7891 (N_7891,N_6837,N_6507);
or U7892 (N_7892,N_6571,N_6329);
xor U7893 (N_7893,N_6514,N_6319);
nand U7894 (N_7894,N_6907,N_6557);
nor U7895 (N_7895,N_6369,N_6626);
or U7896 (N_7896,N_6001,N_6037);
and U7897 (N_7897,N_6171,N_6832);
or U7898 (N_7898,N_6857,N_6852);
and U7899 (N_7899,N_6611,N_6073);
nor U7900 (N_7900,N_6281,N_6475);
and U7901 (N_7901,N_6030,N_6596);
and U7902 (N_7902,N_6068,N_6145);
or U7903 (N_7903,N_6444,N_6161);
nor U7904 (N_7904,N_6296,N_6075);
nand U7905 (N_7905,N_6409,N_6162);
or U7906 (N_7906,N_6929,N_6001);
or U7907 (N_7907,N_6243,N_6300);
nor U7908 (N_7908,N_6687,N_6165);
xnor U7909 (N_7909,N_6771,N_6819);
xor U7910 (N_7910,N_6285,N_6909);
or U7911 (N_7911,N_6854,N_6916);
or U7912 (N_7912,N_6289,N_6386);
xnor U7913 (N_7913,N_6496,N_6726);
and U7914 (N_7914,N_6270,N_6813);
and U7915 (N_7915,N_6076,N_6527);
and U7916 (N_7916,N_6312,N_6820);
or U7917 (N_7917,N_6555,N_6654);
nor U7918 (N_7918,N_6221,N_6694);
and U7919 (N_7919,N_6532,N_6030);
nor U7920 (N_7920,N_6495,N_6568);
and U7921 (N_7921,N_6780,N_6366);
and U7922 (N_7922,N_6394,N_6974);
nand U7923 (N_7923,N_6040,N_6496);
or U7924 (N_7924,N_6007,N_6012);
nor U7925 (N_7925,N_6361,N_6893);
or U7926 (N_7926,N_6088,N_6344);
xor U7927 (N_7927,N_6289,N_6449);
and U7928 (N_7928,N_6226,N_6081);
nand U7929 (N_7929,N_6234,N_6180);
nor U7930 (N_7930,N_6811,N_6893);
xnor U7931 (N_7931,N_6322,N_6351);
nand U7932 (N_7932,N_6093,N_6532);
nand U7933 (N_7933,N_6826,N_6977);
nor U7934 (N_7934,N_6939,N_6970);
nor U7935 (N_7935,N_6582,N_6782);
or U7936 (N_7936,N_6927,N_6488);
or U7937 (N_7937,N_6204,N_6365);
and U7938 (N_7938,N_6253,N_6038);
xor U7939 (N_7939,N_6612,N_6461);
nor U7940 (N_7940,N_6552,N_6477);
nand U7941 (N_7941,N_6851,N_6467);
nand U7942 (N_7942,N_6861,N_6562);
nor U7943 (N_7943,N_6013,N_6855);
nor U7944 (N_7944,N_6156,N_6707);
and U7945 (N_7945,N_6423,N_6775);
or U7946 (N_7946,N_6527,N_6758);
and U7947 (N_7947,N_6362,N_6279);
xnor U7948 (N_7948,N_6375,N_6387);
and U7949 (N_7949,N_6624,N_6910);
nand U7950 (N_7950,N_6388,N_6360);
nor U7951 (N_7951,N_6945,N_6636);
nor U7952 (N_7952,N_6860,N_6531);
nand U7953 (N_7953,N_6762,N_6908);
nand U7954 (N_7954,N_6008,N_6464);
or U7955 (N_7955,N_6290,N_6240);
xnor U7956 (N_7956,N_6676,N_6161);
nand U7957 (N_7957,N_6547,N_6234);
nor U7958 (N_7958,N_6574,N_6319);
nand U7959 (N_7959,N_6831,N_6973);
nor U7960 (N_7960,N_6529,N_6554);
and U7961 (N_7961,N_6317,N_6535);
xor U7962 (N_7962,N_6614,N_6651);
nand U7963 (N_7963,N_6770,N_6547);
and U7964 (N_7964,N_6964,N_6953);
nand U7965 (N_7965,N_6888,N_6567);
nand U7966 (N_7966,N_6674,N_6017);
nor U7967 (N_7967,N_6868,N_6176);
xor U7968 (N_7968,N_6712,N_6272);
nor U7969 (N_7969,N_6024,N_6420);
and U7970 (N_7970,N_6943,N_6868);
nor U7971 (N_7971,N_6262,N_6154);
xor U7972 (N_7972,N_6696,N_6552);
or U7973 (N_7973,N_6506,N_6565);
or U7974 (N_7974,N_6481,N_6171);
or U7975 (N_7975,N_6494,N_6513);
nand U7976 (N_7976,N_6013,N_6085);
nor U7977 (N_7977,N_6093,N_6750);
nand U7978 (N_7978,N_6565,N_6941);
or U7979 (N_7979,N_6093,N_6807);
xor U7980 (N_7980,N_6890,N_6629);
nor U7981 (N_7981,N_6825,N_6329);
nor U7982 (N_7982,N_6438,N_6395);
nor U7983 (N_7983,N_6754,N_6816);
and U7984 (N_7984,N_6580,N_6493);
nand U7985 (N_7985,N_6422,N_6547);
or U7986 (N_7986,N_6071,N_6002);
nand U7987 (N_7987,N_6630,N_6998);
and U7988 (N_7988,N_6149,N_6394);
and U7989 (N_7989,N_6482,N_6721);
nor U7990 (N_7990,N_6758,N_6229);
and U7991 (N_7991,N_6185,N_6644);
nand U7992 (N_7992,N_6261,N_6717);
and U7993 (N_7993,N_6015,N_6348);
and U7994 (N_7994,N_6795,N_6354);
xor U7995 (N_7995,N_6837,N_6349);
nor U7996 (N_7996,N_6238,N_6947);
nor U7997 (N_7997,N_6273,N_6016);
or U7998 (N_7998,N_6006,N_6429);
or U7999 (N_7999,N_6676,N_6384);
nor U8000 (N_8000,N_7017,N_7007);
or U8001 (N_8001,N_7078,N_7195);
and U8002 (N_8002,N_7056,N_7767);
nor U8003 (N_8003,N_7457,N_7994);
nor U8004 (N_8004,N_7582,N_7507);
nor U8005 (N_8005,N_7100,N_7104);
nand U8006 (N_8006,N_7051,N_7879);
and U8007 (N_8007,N_7283,N_7090);
or U8008 (N_8008,N_7167,N_7103);
and U8009 (N_8009,N_7781,N_7539);
and U8010 (N_8010,N_7757,N_7267);
or U8011 (N_8011,N_7536,N_7926);
nor U8012 (N_8012,N_7293,N_7228);
nor U8013 (N_8013,N_7262,N_7111);
xor U8014 (N_8014,N_7600,N_7787);
nor U8015 (N_8015,N_7406,N_7303);
nor U8016 (N_8016,N_7191,N_7619);
or U8017 (N_8017,N_7128,N_7834);
nor U8018 (N_8018,N_7363,N_7851);
or U8019 (N_8019,N_7647,N_7748);
nand U8020 (N_8020,N_7273,N_7416);
and U8021 (N_8021,N_7384,N_7339);
nand U8022 (N_8022,N_7469,N_7255);
nand U8023 (N_8023,N_7999,N_7265);
or U8024 (N_8024,N_7620,N_7798);
nor U8025 (N_8025,N_7183,N_7014);
nand U8026 (N_8026,N_7541,N_7625);
and U8027 (N_8027,N_7478,N_7066);
or U8028 (N_8028,N_7525,N_7743);
nand U8029 (N_8029,N_7744,N_7681);
nor U8030 (N_8030,N_7233,N_7586);
nand U8031 (N_8031,N_7797,N_7423);
or U8032 (N_8032,N_7370,N_7943);
or U8033 (N_8033,N_7706,N_7520);
or U8034 (N_8034,N_7872,N_7122);
or U8035 (N_8035,N_7626,N_7421);
nor U8036 (N_8036,N_7947,N_7962);
and U8037 (N_8037,N_7613,N_7717);
xnor U8038 (N_8038,N_7393,N_7063);
or U8039 (N_8039,N_7208,N_7048);
nand U8040 (N_8040,N_7544,N_7018);
nand U8041 (N_8041,N_7952,N_7455);
or U8042 (N_8042,N_7115,N_7969);
or U8043 (N_8043,N_7269,N_7519);
or U8044 (N_8044,N_7139,N_7082);
nand U8045 (N_8045,N_7538,N_7832);
and U8046 (N_8046,N_7511,N_7383);
nor U8047 (N_8047,N_7243,N_7719);
nor U8048 (N_8048,N_7428,N_7808);
and U8049 (N_8049,N_7418,N_7098);
nand U8050 (N_8050,N_7465,N_7321);
and U8051 (N_8051,N_7502,N_7861);
or U8052 (N_8052,N_7693,N_7144);
or U8053 (N_8053,N_7915,N_7229);
nand U8054 (N_8054,N_7803,N_7891);
and U8055 (N_8055,N_7415,N_7445);
and U8056 (N_8056,N_7985,N_7386);
xnor U8057 (N_8057,N_7825,N_7942);
nor U8058 (N_8058,N_7594,N_7147);
or U8059 (N_8059,N_7483,N_7252);
nor U8060 (N_8060,N_7816,N_7932);
nor U8061 (N_8061,N_7577,N_7146);
or U8062 (N_8062,N_7157,N_7186);
or U8063 (N_8063,N_7019,N_7093);
nor U8064 (N_8064,N_7648,N_7737);
and U8065 (N_8065,N_7106,N_7112);
nor U8066 (N_8066,N_7896,N_7012);
nor U8067 (N_8067,N_7306,N_7351);
and U8068 (N_8068,N_7836,N_7599);
nor U8069 (N_8069,N_7721,N_7881);
xor U8070 (N_8070,N_7123,N_7953);
nor U8071 (N_8071,N_7704,N_7451);
nand U8072 (N_8072,N_7134,N_7855);
and U8073 (N_8073,N_7535,N_7518);
and U8074 (N_8074,N_7378,N_7500);
nor U8075 (N_8075,N_7324,N_7608);
and U8076 (N_8076,N_7564,N_7125);
or U8077 (N_8077,N_7245,N_7226);
xor U8078 (N_8078,N_7189,N_7772);
nand U8079 (N_8079,N_7910,N_7687);
or U8080 (N_8080,N_7764,N_7472);
nand U8081 (N_8081,N_7005,N_7231);
or U8082 (N_8082,N_7227,N_7715);
nand U8083 (N_8083,N_7391,N_7169);
or U8084 (N_8084,N_7081,N_7568);
or U8085 (N_8085,N_7176,N_7927);
or U8086 (N_8086,N_7662,N_7101);
and U8087 (N_8087,N_7549,N_7546);
nand U8088 (N_8088,N_7686,N_7411);
nor U8089 (N_8089,N_7184,N_7041);
nor U8090 (N_8090,N_7340,N_7034);
and U8091 (N_8091,N_7460,N_7946);
xor U8092 (N_8092,N_7348,N_7792);
and U8093 (N_8093,N_7300,N_7848);
and U8094 (N_8094,N_7712,N_7897);
nand U8095 (N_8095,N_7641,N_7033);
or U8096 (N_8096,N_7268,N_7696);
nor U8097 (N_8097,N_7220,N_7408);
xor U8098 (N_8098,N_7410,N_7130);
nor U8099 (N_8099,N_7554,N_7360);
or U8100 (N_8100,N_7863,N_7288);
nand U8101 (N_8101,N_7447,N_7672);
nor U8102 (N_8102,N_7677,N_7930);
xor U8103 (N_8103,N_7609,N_7674);
nor U8104 (N_8104,N_7552,N_7563);
nand U8105 (N_8105,N_7742,N_7659);
or U8106 (N_8106,N_7016,N_7811);
xnor U8107 (N_8107,N_7371,N_7565);
or U8108 (N_8108,N_7020,N_7357);
or U8109 (N_8109,N_7660,N_7368);
nand U8110 (N_8110,N_7069,N_7889);
nor U8111 (N_8111,N_7289,N_7774);
nand U8112 (N_8112,N_7933,N_7598);
nand U8113 (N_8113,N_7023,N_7367);
nand U8114 (N_8114,N_7601,N_7562);
and U8115 (N_8115,N_7871,N_7485);
and U8116 (N_8116,N_7860,N_7072);
nor U8117 (N_8117,N_7459,N_7917);
nor U8118 (N_8118,N_7603,N_7334);
nand U8119 (N_8119,N_7387,N_7096);
or U8120 (N_8120,N_7655,N_7344);
nor U8121 (N_8121,N_7777,N_7403);
and U8122 (N_8122,N_7276,N_7595);
xor U8123 (N_8123,N_7119,N_7888);
nor U8124 (N_8124,N_7008,N_7296);
nand U8125 (N_8125,N_7205,N_7701);
nand U8126 (N_8126,N_7318,N_7958);
or U8127 (N_8127,N_7622,N_7993);
xor U8128 (N_8128,N_7558,N_7473);
xnor U8129 (N_8129,N_7352,N_7467);
nand U8130 (N_8130,N_7264,N_7250);
and U8131 (N_8131,N_7867,N_7928);
or U8132 (N_8132,N_7165,N_7761);
nand U8133 (N_8133,N_7698,N_7295);
or U8134 (N_8134,N_7050,N_7105);
nand U8135 (N_8135,N_7692,N_7510);
xor U8136 (N_8136,N_7124,N_7437);
xor U8137 (N_8137,N_7854,N_7089);
or U8138 (N_8138,N_7644,N_7611);
or U8139 (N_8139,N_7079,N_7301);
nor U8140 (N_8140,N_7905,N_7976);
xor U8141 (N_8141,N_7364,N_7548);
or U8142 (N_8142,N_7446,N_7290);
nand U8143 (N_8143,N_7336,N_7901);
or U8144 (N_8144,N_7136,N_7874);
or U8145 (N_8145,N_7013,N_7211);
and U8146 (N_8146,N_7326,N_7738);
nor U8147 (N_8147,N_7085,N_7653);
and U8148 (N_8148,N_7214,N_7244);
or U8149 (N_8149,N_7920,N_7924);
and U8150 (N_8150,N_7990,N_7657);
or U8151 (N_8151,N_7037,N_7236);
nand U8152 (N_8152,N_7617,N_7057);
nand U8153 (N_8153,N_7941,N_7570);
xor U8154 (N_8154,N_7054,N_7576);
nor U8155 (N_8155,N_7964,N_7802);
or U8156 (N_8156,N_7097,N_7652);
nand U8157 (N_8157,N_7064,N_7199);
or U8158 (N_8158,N_7398,N_7751);
nor U8159 (N_8159,N_7382,N_7271);
nor U8160 (N_8160,N_7088,N_7419);
nand U8161 (N_8161,N_7249,N_7579);
nor U8162 (N_8162,N_7639,N_7936);
xor U8163 (N_8163,N_7480,N_7261);
and U8164 (N_8164,N_7476,N_7673);
or U8165 (N_8165,N_7397,N_7656);
nor U8166 (N_8166,N_7893,N_7602);
nor U8167 (N_8167,N_7060,N_7996);
nand U8168 (N_8168,N_7151,N_7708);
or U8169 (N_8169,N_7722,N_7818);
nand U8170 (N_8170,N_7522,N_7335);
and U8171 (N_8171,N_7468,N_7389);
nor U8172 (N_8172,N_7845,N_7281);
or U8173 (N_8173,N_7831,N_7346);
nand U8174 (N_8174,N_7730,N_7192);
nor U8175 (N_8175,N_7799,N_7443);
nor U8176 (N_8176,N_7177,N_7373);
xor U8177 (N_8177,N_7052,N_7666);
nand U8178 (N_8178,N_7040,N_7745);
nand U8179 (N_8179,N_7175,N_7689);
and U8180 (N_8180,N_7275,N_7330);
nor U8181 (N_8181,N_7804,N_7618);
or U8182 (N_8182,N_7606,N_7203);
nand U8183 (N_8183,N_7667,N_7463);
and U8184 (N_8184,N_7883,N_7945);
nand U8185 (N_8185,N_7207,N_7172);
and U8186 (N_8186,N_7381,N_7530);
and U8187 (N_8187,N_7545,N_7297);
or U8188 (N_8188,N_7746,N_7524);
or U8189 (N_8189,N_7669,N_7982);
nor U8190 (N_8190,N_7833,N_7705);
xnor U8191 (N_8191,N_7102,N_7237);
xnor U8192 (N_8192,N_7430,N_7484);
xnor U8193 (N_8193,N_7028,N_7826);
nand U8194 (N_8194,N_7940,N_7957);
nor U8195 (N_8195,N_7315,N_7076);
xor U8196 (N_8196,N_7880,N_7849);
or U8197 (N_8197,N_7286,N_7670);
nand U8198 (N_8198,N_7453,N_7212);
nand U8199 (N_8199,N_7140,N_7375);
or U8200 (N_8200,N_7747,N_7458);
nor U8201 (N_8201,N_7328,N_7526);
xor U8202 (N_8202,N_7004,N_7316);
or U8203 (N_8203,N_7338,N_7278);
nor U8204 (N_8204,N_7790,N_7534);
and U8205 (N_8205,N_7068,N_7827);
nor U8206 (N_8206,N_7835,N_7841);
nor U8207 (N_8207,N_7966,N_7059);
and U8208 (N_8208,N_7651,N_7163);
or U8209 (N_8209,N_7995,N_7187);
and U8210 (N_8210,N_7537,N_7137);
and U8211 (N_8211,N_7200,N_7912);
and U8212 (N_8212,N_7080,N_7560);
or U8213 (N_8213,N_7980,N_7168);
xnor U8214 (N_8214,N_7215,N_7970);
nand U8215 (N_8215,N_7780,N_7197);
or U8216 (N_8216,N_7094,N_7160);
and U8217 (N_8217,N_7353,N_7809);
or U8218 (N_8218,N_7760,N_7035);
nand U8219 (N_8219,N_7204,N_7110);
and U8220 (N_8220,N_7314,N_7770);
nor U8221 (N_8221,N_7796,N_7311);
nor U8222 (N_8222,N_7319,N_7002);
and U8223 (N_8223,N_7876,N_7989);
nor U8224 (N_8224,N_7141,N_7143);
xor U8225 (N_8225,N_7120,N_7634);
and U8226 (N_8226,N_7025,N_7277);
and U8227 (N_8227,N_7046,N_7934);
nand U8228 (N_8228,N_7417,N_7263);
or U8229 (N_8229,N_7873,N_7911);
or U8230 (N_8230,N_7426,N_7532);
xor U8231 (N_8231,N_7894,N_7327);
nand U8232 (N_8232,N_7840,N_7355);
nor U8233 (N_8233,N_7640,N_7773);
nor U8234 (N_8234,N_7182,N_7179);
nor U8235 (N_8235,N_7067,N_7358);
and U8236 (N_8236,N_7971,N_7939);
nor U8237 (N_8237,N_7758,N_7566);
and U8238 (N_8238,N_7492,N_7438);
or U8239 (N_8239,N_7178,N_7127);
xor U8240 (N_8240,N_7892,N_7516);
nor U8241 (N_8241,N_7793,N_7533);
and U8242 (N_8242,N_7983,N_7540);
nand U8243 (N_8243,N_7728,N_7006);
xor U8244 (N_8244,N_7107,N_7736);
and U8245 (N_8245,N_7095,N_7049);
nor U8246 (N_8246,N_7741,N_7223);
nor U8247 (N_8247,N_7762,N_7332);
nand U8248 (N_8248,N_7258,N_7272);
and U8249 (N_8249,N_7714,N_7077);
nor U8250 (N_8250,N_7400,N_7190);
and U8251 (N_8251,N_7694,N_7691);
and U8252 (N_8252,N_7788,N_7061);
xnor U8253 (N_8253,N_7528,N_7663);
or U8254 (N_8254,N_7282,N_7477);
nor U8255 (N_8255,N_7441,N_7612);
nor U8256 (N_8256,N_7439,N_7753);
nor U8257 (N_8257,N_7242,N_7654);
nor U8258 (N_8258,N_7045,N_7495);
and U8259 (N_8259,N_7481,N_7631);
and U8260 (N_8260,N_7664,N_7645);
or U8261 (N_8261,N_7022,N_7531);
nor U8262 (N_8262,N_7853,N_7359);
nor U8263 (N_8263,N_7716,N_7404);
or U8264 (N_8264,N_7345,N_7369);
or U8265 (N_8265,N_7121,N_7521);
and U8266 (N_8266,N_7009,N_7444);
nor U8267 (N_8267,N_7188,N_7610);
or U8268 (N_8268,N_7320,N_7587);
nand U8269 (N_8269,N_7253,N_7350);
or U8270 (N_8270,N_7882,N_7193);
and U8271 (N_8271,N_7752,N_7877);
nor U8272 (N_8272,N_7150,N_7968);
nand U8273 (N_8273,N_7887,N_7232);
nor U8274 (N_8274,N_7550,N_7209);
and U8275 (N_8275,N_7471,N_7024);
and U8276 (N_8276,N_7260,N_7794);
nand U8277 (N_8277,N_7201,N_7431);
nor U8278 (N_8278,N_7828,N_7815);
nand U8279 (N_8279,N_7279,N_7731);
nand U8280 (N_8280,N_7585,N_7432);
or U8281 (N_8281,N_7739,N_7702);
nor U8282 (N_8282,N_7365,N_7711);
nand U8283 (N_8283,N_7856,N_7087);
nor U8284 (N_8284,N_7109,N_7908);
and U8285 (N_8285,N_7294,N_7394);
or U8286 (N_8286,N_7557,N_7914);
or U8287 (N_8287,N_7091,N_7196);
or U8288 (N_8288,N_7073,N_7749);
and U8289 (N_8289,N_7699,N_7623);
or U8290 (N_8290,N_7593,N_7847);
nand U8291 (N_8291,N_7627,N_7885);
and U8292 (N_8292,N_7629,N_7824);
nand U8293 (N_8293,N_7489,N_7043);
nand U8294 (N_8294,N_7361,N_7784);
nand U8295 (N_8295,N_7700,N_7956);
nor U8296 (N_8296,N_7668,N_7292);
and U8297 (N_8297,N_7895,N_7735);
nand U8298 (N_8298,N_7723,N_7161);
and U8299 (N_8299,N_7450,N_7392);
nand U8300 (N_8300,N_7807,N_7578);
or U8301 (N_8301,N_7454,N_7597);
and U8302 (N_8302,N_7981,N_7356);
and U8303 (N_8303,N_7857,N_7331);
and U8304 (N_8304,N_7021,N_7813);
or U8305 (N_8305,N_7114,N_7274);
nor U8306 (N_8306,N_7084,N_7224);
or U8307 (N_8307,N_7075,N_7218);
nand U8308 (N_8308,N_7513,N_7581);
nand U8309 (N_8309,N_7395,N_7000);
nand U8310 (N_8310,N_7961,N_7198);
nor U8311 (N_8311,N_7304,N_7142);
nor U8312 (N_8312,N_7763,N_7750);
or U8313 (N_8313,N_7221,N_7222);
and U8314 (N_8314,N_7624,N_7820);
and U8315 (N_8315,N_7173,N_7616);
xor U8316 (N_8316,N_7703,N_7030);
nor U8317 (N_8317,N_7442,N_7771);
nand U8318 (N_8318,N_7680,N_7814);
and U8319 (N_8319,N_7026,N_7592);
xnor U8320 (N_8320,N_7907,N_7377);
and U8321 (N_8321,N_7427,N_7514);
nand U8322 (N_8322,N_7074,N_7789);
and U8323 (N_8323,N_7174,N_7153);
xor U8324 (N_8324,N_7979,N_7129);
and U8325 (N_8325,N_7571,N_7974);
nor U8326 (N_8326,N_7366,N_7003);
or U8327 (N_8327,N_7607,N_7402);
and U8328 (N_8328,N_7806,N_7862);
nand U8329 (N_8329,N_7247,N_7036);
or U8330 (N_8330,N_7829,N_7527);
or U8331 (N_8331,N_7935,N_7695);
nor U8332 (N_8332,N_7372,N_7919);
nand U8333 (N_8333,N_7342,N_7291);
nand U8334 (N_8334,N_7376,N_7878);
or U8335 (N_8335,N_7733,N_7852);
nor U8336 (N_8336,N_7117,N_7671);
nand U8337 (N_8337,N_7474,N_7230);
nor U8338 (N_8338,N_7775,N_7967);
nand U8339 (N_8339,N_7734,N_7709);
nor U8340 (N_8340,N_7621,N_7317);
xnor U8341 (N_8341,N_7171,N_7062);
and U8342 (N_8342,N_7194,N_7429);
nor U8343 (N_8343,N_7108,N_7452);
nor U8344 (N_8344,N_7913,N_7333);
xor U8345 (N_8345,N_7584,N_7843);
or U8346 (N_8346,N_7032,N_7313);
or U8347 (N_8347,N_7869,N_7424);
and U8348 (N_8348,N_7152,N_7949);
and U8349 (N_8349,N_7678,N_7512);
nor U8350 (N_8350,N_7440,N_7523);
nor U8351 (N_8351,N_7099,N_7238);
or U8352 (N_8352,N_7162,N_7690);
and U8353 (N_8353,N_7396,N_7844);
and U8354 (N_8354,N_7042,N_7219);
or U8355 (N_8355,N_7713,N_7065);
nor U8356 (N_8356,N_7838,N_7633);
and U8357 (N_8357,N_7707,N_7148);
and U8358 (N_8358,N_7984,N_7234);
nand U8359 (N_8359,N_7116,N_7149);
xor U8360 (N_8360,N_7322,N_7011);
nand U8361 (N_8361,N_7490,N_7185);
and U8362 (N_8362,N_7070,N_7795);
or U8363 (N_8363,N_7786,N_7944);
and U8364 (N_8364,N_7676,N_7055);
or U8365 (N_8365,N_7284,N_7092);
nor U8366 (N_8366,N_7859,N_7015);
or U8367 (N_8367,N_7414,N_7422);
or U8368 (N_8368,N_7323,N_7886);
and U8369 (N_8369,N_7380,N_7710);
and U8370 (N_8370,N_7823,N_7213);
or U8371 (N_8371,N_7925,N_7462);
nand U8372 (N_8372,N_7665,N_7503);
and U8373 (N_8373,N_7217,N_7001);
and U8374 (N_8374,N_7254,N_7280);
nor U8375 (N_8375,N_7158,N_7922);
and U8376 (N_8376,N_7246,N_7409);
nand U8377 (N_8377,N_7636,N_7684);
and U8378 (N_8378,N_7769,N_7504);
or U8379 (N_8379,N_7170,N_7044);
nand U8380 (N_8380,N_7858,N_7482);
and U8381 (N_8381,N_7567,N_7010);
and U8382 (N_8382,N_7569,N_7965);
nand U8383 (N_8383,N_7830,N_7766);
or U8384 (N_8384,N_7805,N_7488);
or U8385 (N_8385,N_7385,N_7909);
nor U8386 (N_8386,N_7866,N_7181);
or U8387 (N_8387,N_7259,N_7850);
and U8388 (N_8388,N_7257,N_7029);
nor U8389 (N_8389,N_7632,N_7456);
nand U8390 (N_8390,N_7812,N_7225);
or U8391 (N_8391,N_7135,N_7498);
nor U8392 (N_8392,N_7058,N_7954);
or U8393 (N_8393,N_7515,N_7337);
nor U8394 (N_8394,N_7325,N_7251);
nor U8395 (N_8395,N_7642,N_7658);
and U8396 (N_8396,N_7782,N_7759);
or U8397 (N_8397,N_7591,N_7487);
and U8398 (N_8398,N_7596,N_7697);
or U8399 (N_8399,N_7837,N_7497);
and U8400 (N_8400,N_7166,N_7675);
nor U8401 (N_8401,N_7991,N_7461);
nor U8402 (N_8402,N_7561,N_7499);
and U8403 (N_8403,N_7755,N_7987);
xnor U8404 (N_8404,N_7902,N_7494);
or U8405 (N_8405,N_7951,N_7756);
and U8406 (N_8406,N_7630,N_7683);
xor U8407 (N_8407,N_7923,N_7720);
or U8408 (N_8408,N_7401,N_7972);
and U8409 (N_8409,N_7615,N_7343);
or U8410 (N_8410,N_7038,N_7349);
nor U8411 (N_8411,N_7180,N_7638);
xor U8412 (N_8412,N_7138,N_7464);
or U8413 (N_8413,N_7682,N_7420);
nor U8414 (N_8414,N_7154,N_7312);
nand U8415 (N_8415,N_7978,N_7580);
nor U8416 (N_8416,N_7839,N_7407);
nand U8417 (N_8417,N_7216,N_7308);
xnor U8418 (N_8418,N_7959,N_7899);
or U8419 (N_8419,N_7846,N_7575);
or U8420 (N_8420,N_7998,N_7133);
nor U8421 (N_8421,N_7132,N_7725);
nand U8422 (N_8422,N_7310,N_7727);
or U8423 (N_8423,N_7950,N_7031);
and U8424 (N_8424,N_7307,N_7573);
nor U8425 (N_8425,N_7604,N_7754);
nor U8426 (N_8426,N_7302,N_7449);
nand U8427 (N_8427,N_7239,N_7685);
nand U8428 (N_8428,N_7486,N_7235);
nor U8429 (N_8429,N_7551,N_7543);
xor U8430 (N_8430,N_7362,N_7379);
nand U8431 (N_8431,N_7821,N_7810);
xnor U8432 (N_8432,N_7875,N_7864);
xor U8433 (N_8433,N_7776,N_7791);
or U8434 (N_8434,N_7156,N_7590);
xnor U8435 (N_8435,N_7206,N_7027);
xnor U8436 (N_8436,N_7131,N_7555);
and U8437 (N_8437,N_7501,N_7955);
nor U8438 (N_8438,N_7083,N_7768);
or U8439 (N_8439,N_7868,N_7817);
xor U8440 (N_8440,N_7433,N_7491);
xor U8441 (N_8441,N_7210,N_7405);
and U8442 (N_8442,N_7053,N_7509);
nand U8443 (N_8443,N_7884,N_7574);
and U8444 (N_8444,N_7679,N_7783);
and U8445 (N_8445,N_7412,N_7298);
or U8446 (N_8446,N_7299,N_7724);
or U8447 (N_8447,N_7938,N_7778);
nand U8448 (N_8448,N_7740,N_7649);
nor U8449 (N_8449,N_7466,N_7992);
xor U8450 (N_8450,N_7475,N_7256);
nor U8451 (N_8451,N_7605,N_7635);
nand U8452 (N_8452,N_7270,N_7496);
and U8453 (N_8453,N_7448,N_7086);
xnor U8454 (N_8454,N_7588,N_7388);
or U8455 (N_8455,N_7118,N_7434);
and U8456 (N_8456,N_7155,N_7559);
nor U8457 (N_8457,N_7240,N_7159);
xnor U8458 (N_8458,N_7732,N_7918);
or U8459 (N_8459,N_7202,N_7542);
nand U8460 (N_8460,N_7800,N_7929);
or U8461 (N_8461,N_7493,N_7329);
or U8462 (N_8462,N_7517,N_7801);
and U8463 (N_8463,N_7948,N_7986);
and U8464 (N_8464,N_7583,N_7047);
nor U8465 (N_8465,N_7071,N_7973);
or U8466 (N_8466,N_7646,N_7505);
and U8467 (N_8467,N_7113,N_7988);
nor U8468 (N_8468,N_7765,N_7425);
nand U8469 (N_8469,N_7399,N_7164);
nand U8470 (N_8470,N_7903,N_7650);
or U8471 (N_8471,N_7553,N_7637);
xor U8472 (N_8472,N_7354,N_7900);
or U8473 (N_8473,N_7309,N_7785);
nor U8474 (N_8474,N_7937,N_7718);
nand U8475 (N_8475,N_7413,N_7390);
and U8476 (N_8476,N_7285,N_7865);
nand U8477 (N_8477,N_7508,N_7726);
nand U8478 (N_8478,N_7931,N_7305);
or U8479 (N_8479,N_7556,N_7506);
nand U8480 (N_8480,N_7039,N_7977);
xor U8481 (N_8481,N_7729,N_7779);
or U8482 (N_8482,N_7688,N_7819);
nand U8483 (N_8483,N_7341,N_7479);
and U8484 (N_8484,N_7126,N_7266);
nor U8485 (N_8485,N_7628,N_7963);
and U8486 (N_8486,N_7248,N_7547);
nand U8487 (N_8487,N_7287,N_7870);
nand U8488 (N_8488,N_7145,N_7241);
xnor U8489 (N_8489,N_7906,N_7890);
or U8490 (N_8490,N_7822,N_7904);
nand U8491 (N_8491,N_7661,N_7898);
and U8492 (N_8492,N_7347,N_7842);
or U8493 (N_8493,N_7997,N_7572);
or U8494 (N_8494,N_7470,N_7916);
nand U8495 (N_8495,N_7975,N_7374);
nand U8496 (N_8496,N_7436,N_7529);
xor U8497 (N_8497,N_7960,N_7921);
nand U8498 (N_8498,N_7435,N_7643);
and U8499 (N_8499,N_7614,N_7589);
nor U8500 (N_8500,N_7084,N_7062);
xor U8501 (N_8501,N_7771,N_7497);
and U8502 (N_8502,N_7642,N_7015);
nand U8503 (N_8503,N_7016,N_7610);
xnor U8504 (N_8504,N_7393,N_7032);
nand U8505 (N_8505,N_7880,N_7931);
or U8506 (N_8506,N_7507,N_7744);
and U8507 (N_8507,N_7790,N_7522);
and U8508 (N_8508,N_7747,N_7502);
and U8509 (N_8509,N_7858,N_7683);
nand U8510 (N_8510,N_7127,N_7079);
nor U8511 (N_8511,N_7030,N_7468);
nand U8512 (N_8512,N_7658,N_7115);
xor U8513 (N_8513,N_7980,N_7186);
or U8514 (N_8514,N_7908,N_7102);
or U8515 (N_8515,N_7975,N_7576);
nand U8516 (N_8516,N_7112,N_7833);
and U8517 (N_8517,N_7986,N_7386);
or U8518 (N_8518,N_7827,N_7605);
and U8519 (N_8519,N_7941,N_7715);
and U8520 (N_8520,N_7811,N_7640);
nand U8521 (N_8521,N_7808,N_7843);
nor U8522 (N_8522,N_7750,N_7882);
or U8523 (N_8523,N_7921,N_7367);
nand U8524 (N_8524,N_7221,N_7949);
or U8525 (N_8525,N_7786,N_7184);
and U8526 (N_8526,N_7371,N_7059);
nand U8527 (N_8527,N_7423,N_7541);
and U8528 (N_8528,N_7426,N_7080);
and U8529 (N_8529,N_7022,N_7124);
nor U8530 (N_8530,N_7190,N_7417);
nor U8531 (N_8531,N_7847,N_7175);
nand U8532 (N_8532,N_7417,N_7456);
and U8533 (N_8533,N_7095,N_7396);
nand U8534 (N_8534,N_7515,N_7822);
nand U8535 (N_8535,N_7898,N_7200);
and U8536 (N_8536,N_7987,N_7244);
xnor U8537 (N_8537,N_7586,N_7884);
nor U8538 (N_8538,N_7149,N_7411);
xnor U8539 (N_8539,N_7657,N_7702);
or U8540 (N_8540,N_7435,N_7797);
xnor U8541 (N_8541,N_7306,N_7333);
xor U8542 (N_8542,N_7434,N_7845);
and U8543 (N_8543,N_7502,N_7424);
or U8544 (N_8544,N_7605,N_7283);
xor U8545 (N_8545,N_7681,N_7123);
or U8546 (N_8546,N_7883,N_7143);
nand U8547 (N_8547,N_7781,N_7140);
xnor U8548 (N_8548,N_7462,N_7105);
nor U8549 (N_8549,N_7864,N_7492);
xor U8550 (N_8550,N_7084,N_7445);
nand U8551 (N_8551,N_7377,N_7896);
or U8552 (N_8552,N_7942,N_7656);
and U8553 (N_8553,N_7477,N_7849);
nor U8554 (N_8554,N_7377,N_7567);
and U8555 (N_8555,N_7486,N_7488);
and U8556 (N_8556,N_7740,N_7484);
nor U8557 (N_8557,N_7029,N_7306);
nor U8558 (N_8558,N_7247,N_7885);
nand U8559 (N_8559,N_7935,N_7767);
and U8560 (N_8560,N_7284,N_7208);
and U8561 (N_8561,N_7576,N_7719);
xor U8562 (N_8562,N_7373,N_7895);
and U8563 (N_8563,N_7325,N_7165);
nor U8564 (N_8564,N_7790,N_7138);
and U8565 (N_8565,N_7587,N_7883);
or U8566 (N_8566,N_7783,N_7502);
nand U8567 (N_8567,N_7385,N_7347);
and U8568 (N_8568,N_7363,N_7840);
nand U8569 (N_8569,N_7216,N_7903);
nor U8570 (N_8570,N_7719,N_7499);
or U8571 (N_8571,N_7468,N_7483);
or U8572 (N_8572,N_7902,N_7750);
nor U8573 (N_8573,N_7439,N_7733);
or U8574 (N_8574,N_7446,N_7919);
nor U8575 (N_8575,N_7625,N_7395);
nor U8576 (N_8576,N_7631,N_7365);
xor U8577 (N_8577,N_7879,N_7617);
nor U8578 (N_8578,N_7496,N_7870);
and U8579 (N_8579,N_7826,N_7547);
and U8580 (N_8580,N_7812,N_7800);
or U8581 (N_8581,N_7795,N_7059);
nor U8582 (N_8582,N_7101,N_7872);
or U8583 (N_8583,N_7371,N_7493);
and U8584 (N_8584,N_7464,N_7053);
and U8585 (N_8585,N_7656,N_7927);
or U8586 (N_8586,N_7574,N_7152);
nor U8587 (N_8587,N_7013,N_7136);
or U8588 (N_8588,N_7625,N_7680);
nor U8589 (N_8589,N_7036,N_7668);
and U8590 (N_8590,N_7700,N_7568);
or U8591 (N_8591,N_7470,N_7994);
xor U8592 (N_8592,N_7942,N_7804);
nor U8593 (N_8593,N_7824,N_7236);
and U8594 (N_8594,N_7584,N_7158);
nand U8595 (N_8595,N_7605,N_7885);
and U8596 (N_8596,N_7579,N_7900);
or U8597 (N_8597,N_7275,N_7288);
and U8598 (N_8598,N_7691,N_7651);
and U8599 (N_8599,N_7478,N_7361);
xor U8600 (N_8600,N_7609,N_7048);
or U8601 (N_8601,N_7151,N_7145);
or U8602 (N_8602,N_7331,N_7728);
xor U8603 (N_8603,N_7996,N_7262);
or U8604 (N_8604,N_7558,N_7604);
nand U8605 (N_8605,N_7922,N_7479);
nand U8606 (N_8606,N_7046,N_7580);
or U8607 (N_8607,N_7488,N_7881);
nand U8608 (N_8608,N_7036,N_7042);
or U8609 (N_8609,N_7662,N_7445);
or U8610 (N_8610,N_7888,N_7615);
and U8611 (N_8611,N_7270,N_7223);
nand U8612 (N_8612,N_7798,N_7507);
or U8613 (N_8613,N_7157,N_7651);
xnor U8614 (N_8614,N_7122,N_7540);
and U8615 (N_8615,N_7300,N_7568);
nand U8616 (N_8616,N_7271,N_7917);
nor U8617 (N_8617,N_7394,N_7742);
and U8618 (N_8618,N_7471,N_7467);
nand U8619 (N_8619,N_7819,N_7698);
nor U8620 (N_8620,N_7392,N_7429);
nor U8621 (N_8621,N_7090,N_7546);
nor U8622 (N_8622,N_7683,N_7123);
nand U8623 (N_8623,N_7831,N_7501);
nor U8624 (N_8624,N_7261,N_7796);
and U8625 (N_8625,N_7230,N_7573);
and U8626 (N_8626,N_7395,N_7298);
or U8627 (N_8627,N_7664,N_7575);
xor U8628 (N_8628,N_7459,N_7096);
and U8629 (N_8629,N_7176,N_7252);
nand U8630 (N_8630,N_7986,N_7720);
nand U8631 (N_8631,N_7282,N_7085);
and U8632 (N_8632,N_7502,N_7932);
or U8633 (N_8633,N_7344,N_7923);
xnor U8634 (N_8634,N_7974,N_7452);
nand U8635 (N_8635,N_7990,N_7550);
and U8636 (N_8636,N_7854,N_7262);
and U8637 (N_8637,N_7643,N_7679);
and U8638 (N_8638,N_7691,N_7968);
or U8639 (N_8639,N_7152,N_7051);
or U8640 (N_8640,N_7120,N_7130);
nor U8641 (N_8641,N_7002,N_7536);
and U8642 (N_8642,N_7711,N_7750);
nand U8643 (N_8643,N_7562,N_7261);
and U8644 (N_8644,N_7444,N_7241);
or U8645 (N_8645,N_7603,N_7271);
nand U8646 (N_8646,N_7415,N_7331);
xor U8647 (N_8647,N_7212,N_7094);
and U8648 (N_8648,N_7041,N_7231);
nor U8649 (N_8649,N_7724,N_7661);
or U8650 (N_8650,N_7715,N_7831);
nor U8651 (N_8651,N_7166,N_7219);
xnor U8652 (N_8652,N_7957,N_7490);
nand U8653 (N_8653,N_7481,N_7246);
and U8654 (N_8654,N_7144,N_7322);
and U8655 (N_8655,N_7418,N_7528);
nand U8656 (N_8656,N_7703,N_7842);
and U8657 (N_8657,N_7295,N_7904);
or U8658 (N_8658,N_7946,N_7645);
nor U8659 (N_8659,N_7216,N_7054);
or U8660 (N_8660,N_7795,N_7656);
and U8661 (N_8661,N_7730,N_7006);
nor U8662 (N_8662,N_7809,N_7262);
or U8663 (N_8663,N_7916,N_7089);
or U8664 (N_8664,N_7561,N_7856);
xor U8665 (N_8665,N_7044,N_7715);
xor U8666 (N_8666,N_7119,N_7078);
or U8667 (N_8667,N_7568,N_7212);
nor U8668 (N_8668,N_7992,N_7916);
xnor U8669 (N_8669,N_7376,N_7392);
nand U8670 (N_8670,N_7476,N_7202);
or U8671 (N_8671,N_7695,N_7153);
xnor U8672 (N_8672,N_7501,N_7885);
and U8673 (N_8673,N_7784,N_7212);
and U8674 (N_8674,N_7587,N_7659);
or U8675 (N_8675,N_7062,N_7987);
nor U8676 (N_8676,N_7711,N_7699);
nand U8677 (N_8677,N_7991,N_7271);
nand U8678 (N_8678,N_7870,N_7709);
and U8679 (N_8679,N_7211,N_7931);
nand U8680 (N_8680,N_7886,N_7666);
and U8681 (N_8681,N_7056,N_7683);
and U8682 (N_8682,N_7957,N_7431);
and U8683 (N_8683,N_7233,N_7602);
nor U8684 (N_8684,N_7578,N_7873);
nand U8685 (N_8685,N_7501,N_7276);
and U8686 (N_8686,N_7083,N_7271);
nor U8687 (N_8687,N_7742,N_7269);
or U8688 (N_8688,N_7550,N_7988);
or U8689 (N_8689,N_7140,N_7308);
xor U8690 (N_8690,N_7583,N_7466);
and U8691 (N_8691,N_7260,N_7319);
xor U8692 (N_8692,N_7045,N_7002);
and U8693 (N_8693,N_7105,N_7696);
nand U8694 (N_8694,N_7403,N_7954);
xor U8695 (N_8695,N_7308,N_7703);
nand U8696 (N_8696,N_7844,N_7045);
or U8697 (N_8697,N_7296,N_7507);
or U8698 (N_8698,N_7980,N_7573);
nand U8699 (N_8699,N_7560,N_7742);
or U8700 (N_8700,N_7484,N_7966);
or U8701 (N_8701,N_7394,N_7378);
and U8702 (N_8702,N_7283,N_7471);
and U8703 (N_8703,N_7936,N_7935);
nor U8704 (N_8704,N_7925,N_7899);
and U8705 (N_8705,N_7803,N_7241);
nor U8706 (N_8706,N_7172,N_7458);
nand U8707 (N_8707,N_7123,N_7940);
and U8708 (N_8708,N_7205,N_7260);
or U8709 (N_8709,N_7967,N_7033);
or U8710 (N_8710,N_7951,N_7075);
and U8711 (N_8711,N_7169,N_7201);
nor U8712 (N_8712,N_7653,N_7855);
nor U8713 (N_8713,N_7960,N_7633);
nand U8714 (N_8714,N_7103,N_7902);
and U8715 (N_8715,N_7340,N_7391);
nor U8716 (N_8716,N_7635,N_7657);
nor U8717 (N_8717,N_7094,N_7699);
nor U8718 (N_8718,N_7389,N_7223);
nand U8719 (N_8719,N_7025,N_7056);
nand U8720 (N_8720,N_7397,N_7914);
and U8721 (N_8721,N_7795,N_7419);
or U8722 (N_8722,N_7226,N_7147);
nor U8723 (N_8723,N_7471,N_7120);
or U8724 (N_8724,N_7215,N_7839);
nor U8725 (N_8725,N_7105,N_7312);
and U8726 (N_8726,N_7533,N_7846);
or U8727 (N_8727,N_7097,N_7155);
nand U8728 (N_8728,N_7976,N_7761);
and U8729 (N_8729,N_7003,N_7659);
nand U8730 (N_8730,N_7497,N_7982);
nand U8731 (N_8731,N_7468,N_7512);
and U8732 (N_8732,N_7944,N_7698);
nor U8733 (N_8733,N_7664,N_7328);
and U8734 (N_8734,N_7303,N_7735);
and U8735 (N_8735,N_7800,N_7241);
xor U8736 (N_8736,N_7988,N_7634);
and U8737 (N_8737,N_7863,N_7181);
nand U8738 (N_8738,N_7019,N_7919);
or U8739 (N_8739,N_7743,N_7632);
and U8740 (N_8740,N_7104,N_7648);
or U8741 (N_8741,N_7543,N_7440);
nor U8742 (N_8742,N_7028,N_7114);
or U8743 (N_8743,N_7261,N_7297);
xor U8744 (N_8744,N_7488,N_7894);
and U8745 (N_8745,N_7402,N_7251);
and U8746 (N_8746,N_7021,N_7361);
and U8747 (N_8747,N_7905,N_7346);
nand U8748 (N_8748,N_7187,N_7764);
xor U8749 (N_8749,N_7847,N_7681);
nor U8750 (N_8750,N_7271,N_7459);
nand U8751 (N_8751,N_7571,N_7693);
or U8752 (N_8752,N_7742,N_7246);
nand U8753 (N_8753,N_7858,N_7300);
nand U8754 (N_8754,N_7629,N_7244);
and U8755 (N_8755,N_7344,N_7435);
nand U8756 (N_8756,N_7611,N_7682);
or U8757 (N_8757,N_7446,N_7691);
or U8758 (N_8758,N_7731,N_7615);
nand U8759 (N_8759,N_7615,N_7056);
or U8760 (N_8760,N_7587,N_7318);
nand U8761 (N_8761,N_7323,N_7569);
and U8762 (N_8762,N_7316,N_7190);
nand U8763 (N_8763,N_7617,N_7073);
nand U8764 (N_8764,N_7254,N_7671);
nand U8765 (N_8765,N_7480,N_7922);
nor U8766 (N_8766,N_7766,N_7768);
or U8767 (N_8767,N_7664,N_7896);
nand U8768 (N_8768,N_7087,N_7722);
and U8769 (N_8769,N_7539,N_7311);
nand U8770 (N_8770,N_7748,N_7417);
nand U8771 (N_8771,N_7080,N_7895);
or U8772 (N_8772,N_7778,N_7223);
nand U8773 (N_8773,N_7366,N_7299);
and U8774 (N_8774,N_7102,N_7743);
nor U8775 (N_8775,N_7262,N_7340);
or U8776 (N_8776,N_7080,N_7599);
and U8777 (N_8777,N_7439,N_7891);
nand U8778 (N_8778,N_7232,N_7845);
nand U8779 (N_8779,N_7571,N_7623);
or U8780 (N_8780,N_7724,N_7326);
nand U8781 (N_8781,N_7185,N_7257);
or U8782 (N_8782,N_7189,N_7718);
and U8783 (N_8783,N_7052,N_7643);
nor U8784 (N_8784,N_7060,N_7735);
and U8785 (N_8785,N_7179,N_7045);
or U8786 (N_8786,N_7063,N_7656);
nor U8787 (N_8787,N_7027,N_7065);
and U8788 (N_8788,N_7859,N_7530);
xor U8789 (N_8789,N_7510,N_7967);
nand U8790 (N_8790,N_7254,N_7814);
xnor U8791 (N_8791,N_7625,N_7935);
or U8792 (N_8792,N_7441,N_7726);
xor U8793 (N_8793,N_7443,N_7805);
and U8794 (N_8794,N_7380,N_7270);
and U8795 (N_8795,N_7659,N_7432);
or U8796 (N_8796,N_7250,N_7678);
and U8797 (N_8797,N_7304,N_7756);
or U8798 (N_8798,N_7382,N_7158);
nor U8799 (N_8799,N_7182,N_7490);
nor U8800 (N_8800,N_7301,N_7477);
nand U8801 (N_8801,N_7636,N_7996);
or U8802 (N_8802,N_7144,N_7796);
xor U8803 (N_8803,N_7811,N_7859);
nand U8804 (N_8804,N_7423,N_7168);
nand U8805 (N_8805,N_7073,N_7956);
xor U8806 (N_8806,N_7365,N_7012);
or U8807 (N_8807,N_7409,N_7561);
nor U8808 (N_8808,N_7425,N_7893);
or U8809 (N_8809,N_7219,N_7561);
or U8810 (N_8810,N_7569,N_7947);
or U8811 (N_8811,N_7970,N_7149);
and U8812 (N_8812,N_7054,N_7338);
and U8813 (N_8813,N_7627,N_7598);
nand U8814 (N_8814,N_7153,N_7321);
nand U8815 (N_8815,N_7099,N_7713);
nand U8816 (N_8816,N_7090,N_7056);
xor U8817 (N_8817,N_7654,N_7896);
nand U8818 (N_8818,N_7427,N_7036);
nand U8819 (N_8819,N_7102,N_7660);
xnor U8820 (N_8820,N_7720,N_7364);
nand U8821 (N_8821,N_7132,N_7049);
and U8822 (N_8822,N_7413,N_7411);
and U8823 (N_8823,N_7118,N_7501);
nor U8824 (N_8824,N_7506,N_7922);
or U8825 (N_8825,N_7198,N_7748);
nand U8826 (N_8826,N_7937,N_7467);
xor U8827 (N_8827,N_7379,N_7462);
and U8828 (N_8828,N_7350,N_7704);
or U8829 (N_8829,N_7213,N_7944);
and U8830 (N_8830,N_7343,N_7581);
nor U8831 (N_8831,N_7061,N_7996);
nor U8832 (N_8832,N_7509,N_7883);
and U8833 (N_8833,N_7392,N_7152);
or U8834 (N_8834,N_7392,N_7421);
nand U8835 (N_8835,N_7852,N_7104);
nand U8836 (N_8836,N_7504,N_7205);
nor U8837 (N_8837,N_7603,N_7004);
nand U8838 (N_8838,N_7870,N_7286);
and U8839 (N_8839,N_7654,N_7444);
or U8840 (N_8840,N_7702,N_7079);
nand U8841 (N_8841,N_7990,N_7781);
xnor U8842 (N_8842,N_7914,N_7358);
or U8843 (N_8843,N_7151,N_7158);
and U8844 (N_8844,N_7479,N_7024);
and U8845 (N_8845,N_7272,N_7907);
or U8846 (N_8846,N_7346,N_7545);
and U8847 (N_8847,N_7021,N_7126);
xnor U8848 (N_8848,N_7855,N_7523);
nand U8849 (N_8849,N_7376,N_7615);
and U8850 (N_8850,N_7930,N_7855);
nor U8851 (N_8851,N_7481,N_7442);
nor U8852 (N_8852,N_7104,N_7165);
nor U8853 (N_8853,N_7259,N_7895);
and U8854 (N_8854,N_7844,N_7198);
and U8855 (N_8855,N_7920,N_7443);
nor U8856 (N_8856,N_7609,N_7157);
or U8857 (N_8857,N_7286,N_7925);
nand U8858 (N_8858,N_7358,N_7944);
nand U8859 (N_8859,N_7895,N_7750);
and U8860 (N_8860,N_7506,N_7759);
xnor U8861 (N_8861,N_7298,N_7965);
or U8862 (N_8862,N_7195,N_7891);
nand U8863 (N_8863,N_7126,N_7075);
nor U8864 (N_8864,N_7422,N_7261);
xnor U8865 (N_8865,N_7640,N_7958);
and U8866 (N_8866,N_7647,N_7774);
or U8867 (N_8867,N_7037,N_7008);
nand U8868 (N_8868,N_7214,N_7298);
nor U8869 (N_8869,N_7281,N_7781);
nor U8870 (N_8870,N_7307,N_7437);
nand U8871 (N_8871,N_7139,N_7651);
nand U8872 (N_8872,N_7455,N_7541);
nand U8873 (N_8873,N_7393,N_7003);
nand U8874 (N_8874,N_7244,N_7551);
and U8875 (N_8875,N_7372,N_7022);
or U8876 (N_8876,N_7885,N_7479);
nand U8877 (N_8877,N_7007,N_7381);
and U8878 (N_8878,N_7967,N_7260);
nor U8879 (N_8879,N_7957,N_7907);
and U8880 (N_8880,N_7650,N_7077);
or U8881 (N_8881,N_7021,N_7934);
or U8882 (N_8882,N_7637,N_7500);
or U8883 (N_8883,N_7720,N_7795);
nor U8884 (N_8884,N_7925,N_7893);
and U8885 (N_8885,N_7269,N_7917);
nor U8886 (N_8886,N_7997,N_7385);
nor U8887 (N_8887,N_7189,N_7496);
or U8888 (N_8888,N_7343,N_7346);
nor U8889 (N_8889,N_7999,N_7142);
xor U8890 (N_8890,N_7698,N_7179);
nand U8891 (N_8891,N_7010,N_7919);
nand U8892 (N_8892,N_7109,N_7588);
nor U8893 (N_8893,N_7983,N_7176);
nand U8894 (N_8894,N_7575,N_7494);
nand U8895 (N_8895,N_7054,N_7995);
nand U8896 (N_8896,N_7975,N_7455);
nand U8897 (N_8897,N_7927,N_7376);
nor U8898 (N_8898,N_7885,N_7985);
nor U8899 (N_8899,N_7412,N_7407);
xor U8900 (N_8900,N_7487,N_7510);
nor U8901 (N_8901,N_7489,N_7931);
and U8902 (N_8902,N_7970,N_7954);
xnor U8903 (N_8903,N_7539,N_7645);
and U8904 (N_8904,N_7003,N_7424);
xor U8905 (N_8905,N_7670,N_7373);
nor U8906 (N_8906,N_7485,N_7741);
xnor U8907 (N_8907,N_7534,N_7497);
and U8908 (N_8908,N_7741,N_7314);
nor U8909 (N_8909,N_7294,N_7426);
nand U8910 (N_8910,N_7035,N_7282);
nor U8911 (N_8911,N_7123,N_7235);
nand U8912 (N_8912,N_7707,N_7584);
and U8913 (N_8913,N_7992,N_7352);
nor U8914 (N_8914,N_7571,N_7883);
nand U8915 (N_8915,N_7110,N_7999);
nand U8916 (N_8916,N_7330,N_7138);
xnor U8917 (N_8917,N_7981,N_7295);
nor U8918 (N_8918,N_7264,N_7615);
xnor U8919 (N_8919,N_7540,N_7215);
or U8920 (N_8920,N_7680,N_7315);
or U8921 (N_8921,N_7821,N_7964);
and U8922 (N_8922,N_7433,N_7959);
nor U8923 (N_8923,N_7588,N_7695);
nor U8924 (N_8924,N_7177,N_7675);
nand U8925 (N_8925,N_7374,N_7488);
and U8926 (N_8926,N_7539,N_7649);
nor U8927 (N_8927,N_7793,N_7881);
nand U8928 (N_8928,N_7540,N_7037);
nor U8929 (N_8929,N_7913,N_7160);
nor U8930 (N_8930,N_7032,N_7425);
and U8931 (N_8931,N_7147,N_7655);
and U8932 (N_8932,N_7932,N_7985);
nand U8933 (N_8933,N_7363,N_7890);
nand U8934 (N_8934,N_7785,N_7979);
or U8935 (N_8935,N_7902,N_7674);
or U8936 (N_8936,N_7373,N_7757);
nor U8937 (N_8937,N_7796,N_7975);
nor U8938 (N_8938,N_7928,N_7451);
nor U8939 (N_8939,N_7993,N_7915);
or U8940 (N_8940,N_7955,N_7492);
nor U8941 (N_8941,N_7274,N_7812);
nor U8942 (N_8942,N_7809,N_7931);
nor U8943 (N_8943,N_7882,N_7092);
nand U8944 (N_8944,N_7974,N_7856);
nand U8945 (N_8945,N_7363,N_7073);
and U8946 (N_8946,N_7681,N_7577);
nand U8947 (N_8947,N_7583,N_7944);
nor U8948 (N_8948,N_7778,N_7281);
nand U8949 (N_8949,N_7070,N_7212);
and U8950 (N_8950,N_7383,N_7752);
and U8951 (N_8951,N_7417,N_7126);
nand U8952 (N_8952,N_7900,N_7243);
and U8953 (N_8953,N_7465,N_7962);
nand U8954 (N_8954,N_7403,N_7102);
nand U8955 (N_8955,N_7257,N_7369);
and U8956 (N_8956,N_7268,N_7156);
and U8957 (N_8957,N_7769,N_7618);
and U8958 (N_8958,N_7221,N_7919);
xnor U8959 (N_8959,N_7676,N_7637);
and U8960 (N_8960,N_7725,N_7178);
xnor U8961 (N_8961,N_7189,N_7415);
nor U8962 (N_8962,N_7115,N_7951);
and U8963 (N_8963,N_7748,N_7859);
nor U8964 (N_8964,N_7334,N_7687);
nand U8965 (N_8965,N_7059,N_7403);
nand U8966 (N_8966,N_7836,N_7732);
and U8967 (N_8967,N_7208,N_7932);
nor U8968 (N_8968,N_7803,N_7714);
nor U8969 (N_8969,N_7279,N_7622);
or U8970 (N_8970,N_7896,N_7080);
nand U8971 (N_8971,N_7022,N_7389);
and U8972 (N_8972,N_7918,N_7746);
nand U8973 (N_8973,N_7726,N_7500);
or U8974 (N_8974,N_7700,N_7833);
nor U8975 (N_8975,N_7506,N_7152);
and U8976 (N_8976,N_7151,N_7602);
and U8977 (N_8977,N_7535,N_7906);
nand U8978 (N_8978,N_7491,N_7693);
nand U8979 (N_8979,N_7366,N_7922);
xnor U8980 (N_8980,N_7194,N_7160);
xnor U8981 (N_8981,N_7368,N_7400);
nand U8982 (N_8982,N_7272,N_7223);
xor U8983 (N_8983,N_7403,N_7056);
or U8984 (N_8984,N_7654,N_7214);
nor U8985 (N_8985,N_7667,N_7453);
or U8986 (N_8986,N_7497,N_7249);
and U8987 (N_8987,N_7054,N_7333);
or U8988 (N_8988,N_7424,N_7107);
or U8989 (N_8989,N_7234,N_7909);
nor U8990 (N_8990,N_7681,N_7810);
and U8991 (N_8991,N_7564,N_7105);
nand U8992 (N_8992,N_7264,N_7771);
or U8993 (N_8993,N_7265,N_7792);
nand U8994 (N_8994,N_7364,N_7068);
nand U8995 (N_8995,N_7456,N_7118);
or U8996 (N_8996,N_7369,N_7353);
xnor U8997 (N_8997,N_7480,N_7884);
or U8998 (N_8998,N_7075,N_7480);
xnor U8999 (N_8999,N_7746,N_7670);
or U9000 (N_9000,N_8752,N_8689);
nor U9001 (N_9001,N_8928,N_8500);
nand U9002 (N_9002,N_8263,N_8360);
or U9003 (N_9003,N_8520,N_8591);
and U9004 (N_9004,N_8904,N_8207);
nand U9005 (N_9005,N_8555,N_8456);
or U9006 (N_9006,N_8477,N_8652);
nor U9007 (N_9007,N_8947,N_8473);
xor U9008 (N_9008,N_8205,N_8640);
xnor U9009 (N_9009,N_8999,N_8567);
nor U9010 (N_9010,N_8424,N_8940);
or U9011 (N_9011,N_8715,N_8796);
nand U9012 (N_9012,N_8891,N_8923);
or U9013 (N_9013,N_8043,N_8091);
nand U9014 (N_9014,N_8494,N_8980);
nor U9015 (N_9015,N_8570,N_8304);
or U9016 (N_9016,N_8387,N_8505);
xor U9017 (N_9017,N_8038,N_8259);
and U9018 (N_9018,N_8322,N_8331);
or U9019 (N_9019,N_8156,N_8006);
or U9020 (N_9020,N_8084,N_8454);
nand U9021 (N_9021,N_8265,N_8614);
nand U9022 (N_9022,N_8440,N_8499);
xor U9023 (N_9023,N_8177,N_8072);
and U9024 (N_9024,N_8585,N_8460);
nor U9025 (N_9025,N_8306,N_8189);
nand U9026 (N_9026,N_8991,N_8924);
xnor U9027 (N_9027,N_8982,N_8280);
xor U9028 (N_9028,N_8136,N_8335);
xor U9029 (N_9029,N_8654,N_8800);
and U9030 (N_9030,N_8121,N_8854);
and U9031 (N_9031,N_8708,N_8476);
nor U9032 (N_9032,N_8432,N_8817);
nor U9033 (N_9033,N_8251,N_8158);
or U9034 (N_9034,N_8168,N_8879);
or U9035 (N_9035,N_8351,N_8563);
nor U9036 (N_9036,N_8428,N_8086);
xor U9037 (N_9037,N_8639,N_8678);
nand U9038 (N_9038,N_8455,N_8436);
nand U9039 (N_9039,N_8648,N_8897);
or U9040 (N_9040,N_8378,N_8269);
or U9041 (N_9041,N_8816,N_8944);
and U9042 (N_9042,N_8707,N_8041);
and U9043 (N_9043,N_8221,N_8782);
nor U9044 (N_9044,N_8336,N_8399);
xor U9045 (N_9045,N_8303,N_8890);
nor U9046 (N_9046,N_8092,N_8178);
or U9047 (N_9047,N_8755,N_8865);
and U9048 (N_9048,N_8357,N_8425);
and U9049 (N_9049,N_8556,N_8821);
and U9050 (N_9050,N_8762,N_8324);
or U9051 (N_9051,N_8036,N_8258);
nand U9052 (N_9052,N_8135,N_8321);
nand U9053 (N_9053,N_8300,N_8709);
or U9054 (N_9054,N_8729,N_8358);
and U9055 (N_9055,N_8055,N_8483);
or U9056 (N_9056,N_8840,N_8881);
or U9057 (N_9057,N_8393,N_8549);
or U9058 (N_9058,N_8116,N_8908);
nand U9059 (N_9059,N_8400,N_8815);
xnor U9060 (N_9060,N_8554,N_8023);
xnor U9061 (N_9061,N_8594,N_8273);
or U9062 (N_9062,N_8605,N_8785);
and U9063 (N_9063,N_8231,N_8769);
xnor U9064 (N_9064,N_8284,N_8392);
nor U9065 (N_9065,N_8215,N_8370);
or U9066 (N_9066,N_8489,N_8507);
nand U9067 (N_9067,N_8958,N_8464);
nor U9068 (N_9068,N_8443,N_8623);
nand U9069 (N_9069,N_8186,N_8001);
and U9070 (N_9070,N_8046,N_8730);
and U9071 (N_9071,N_8849,N_8426);
nor U9072 (N_9072,N_8588,N_8701);
and U9073 (N_9073,N_8653,N_8169);
and U9074 (N_9074,N_8634,N_8774);
or U9075 (N_9075,N_8777,N_8248);
nor U9076 (N_9076,N_8667,N_8693);
nand U9077 (N_9077,N_8564,N_8236);
nand U9078 (N_9078,N_8801,N_8346);
and U9079 (N_9079,N_8575,N_8759);
nand U9080 (N_9080,N_8917,N_8082);
or U9081 (N_9081,N_8385,N_8820);
or U9082 (N_9082,N_8149,N_8502);
nand U9083 (N_9083,N_8617,N_8676);
nand U9084 (N_9084,N_8713,N_8872);
nor U9085 (N_9085,N_8629,N_8067);
nand U9086 (N_9086,N_8412,N_8397);
and U9087 (N_9087,N_8931,N_8766);
or U9088 (N_9088,N_8161,N_8313);
nor U9089 (N_9089,N_8990,N_8929);
nor U9090 (N_9090,N_8497,N_8240);
nand U9091 (N_9091,N_8895,N_8218);
and U9092 (N_9092,N_8568,N_8319);
nor U9093 (N_9093,N_8910,N_8139);
or U9094 (N_9094,N_8470,N_8467);
nor U9095 (N_9095,N_8475,N_8297);
nor U9096 (N_9096,N_8934,N_8655);
xor U9097 (N_9097,N_8317,N_8988);
xor U9098 (N_9098,N_8057,N_8798);
nor U9099 (N_9099,N_8033,N_8789);
and U9100 (N_9100,N_8957,N_8449);
xnor U9101 (N_9101,N_8551,N_8989);
nor U9102 (N_9102,N_8353,N_8228);
and U9103 (N_9103,N_8486,N_8187);
or U9104 (N_9104,N_8878,N_8682);
and U9105 (N_9105,N_8326,N_8492);
nand U9106 (N_9106,N_8184,N_8372);
or U9107 (N_9107,N_8018,N_8237);
or U9108 (N_9108,N_8243,N_8926);
nand U9109 (N_9109,N_8998,N_8340);
nor U9110 (N_9110,N_8000,N_8666);
nand U9111 (N_9111,N_8312,N_8584);
nand U9112 (N_9112,N_8469,N_8223);
nor U9113 (N_9113,N_8129,N_8222);
nor U9114 (N_9114,N_8814,N_8735);
nand U9115 (N_9115,N_8775,N_8674);
or U9116 (N_9116,N_8414,N_8029);
nor U9117 (N_9117,N_8242,N_8083);
or U9118 (N_9118,N_8145,N_8379);
and U9119 (N_9119,N_8946,N_8662);
and U9120 (N_9120,N_8102,N_8960);
nor U9121 (N_9121,N_8108,N_8660);
nand U9122 (N_9122,N_8636,N_8097);
xor U9123 (N_9123,N_8423,N_8528);
nand U9124 (N_9124,N_8628,N_8441);
nand U9125 (N_9125,N_8790,N_8948);
xor U9126 (N_9126,N_8277,N_8482);
nor U9127 (N_9127,N_8192,N_8085);
nand U9128 (N_9128,N_8531,N_8472);
and U9129 (N_9129,N_8155,N_8870);
nand U9130 (N_9130,N_8421,N_8573);
or U9131 (N_9131,N_8690,N_8040);
xor U9132 (N_9132,N_8495,N_8506);
xor U9133 (N_9133,N_8491,N_8056);
xor U9134 (N_9134,N_8451,N_8941);
xnor U9135 (N_9135,N_8318,N_8925);
or U9136 (N_9136,N_8874,N_8356);
xor U9137 (N_9137,N_8569,N_8389);
nor U9138 (N_9138,N_8013,N_8119);
nor U9139 (N_9139,N_8912,N_8252);
and U9140 (N_9140,N_8413,N_8856);
nor U9141 (N_9141,N_8807,N_8788);
nand U9142 (N_9142,N_8619,N_8953);
and U9143 (N_9143,N_8852,N_8268);
and U9144 (N_9144,N_8008,N_8671);
nand U9145 (N_9145,N_8808,N_8739);
and U9146 (N_9146,N_8542,N_8922);
and U9147 (N_9147,N_8576,N_8471);
nor U9148 (N_9148,N_8691,N_8921);
xnor U9149 (N_9149,N_8641,N_8011);
and U9150 (N_9150,N_8521,N_8185);
nor U9151 (N_9151,N_8118,N_8835);
xnor U9152 (N_9152,N_8409,N_8054);
and U9153 (N_9153,N_8779,N_8274);
or U9154 (N_9154,N_8203,N_8174);
and U9155 (N_9155,N_8294,N_8098);
or U9156 (N_9156,N_8992,N_8776);
and U9157 (N_9157,N_8981,N_8193);
nor U9158 (N_9158,N_8985,N_8381);
xor U9159 (N_9159,N_8883,N_8200);
xnor U9160 (N_9160,N_8532,N_8697);
or U9161 (N_9161,N_8861,N_8430);
nor U9162 (N_9162,N_8626,N_8075);
or U9163 (N_9163,N_8937,N_8442);
nand U9164 (N_9164,N_8371,N_8645);
or U9165 (N_9165,N_8996,N_8949);
nor U9166 (N_9166,N_8087,N_8490);
nand U9167 (N_9167,N_8420,N_8354);
nand U9168 (N_9168,N_8906,N_8787);
nand U9169 (N_9169,N_8819,N_8275);
nor U9170 (N_9170,N_8141,N_8638);
nor U9171 (N_9171,N_8212,N_8797);
nor U9172 (N_9172,N_8510,N_8465);
or U9173 (N_9173,N_8493,N_8952);
nor U9174 (N_9174,N_8836,N_8577);
and U9175 (N_9175,N_8703,N_8767);
or U9176 (N_9176,N_8954,N_8262);
nor U9177 (N_9177,N_8911,N_8437);
and U9178 (N_9178,N_8019,N_8106);
nand U9179 (N_9179,N_8152,N_8384);
nor U9180 (N_9180,N_8227,N_8005);
or U9181 (N_9181,N_8088,N_8809);
and U9182 (N_9182,N_8986,N_8675);
nor U9183 (N_9183,N_8403,N_8366);
and U9184 (N_9184,N_8095,N_8406);
nor U9185 (N_9185,N_8799,N_8276);
xnor U9186 (N_9186,N_8665,N_8858);
nand U9187 (N_9187,N_8344,N_8602);
nor U9188 (N_9188,N_8833,N_8289);
or U9189 (N_9189,N_8260,N_8620);
or U9190 (N_9190,N_8504,N_8191);
or U9191 (N_9191,N_8478,N_8501);
and U9192 (N_9192,N_8285,N_8452);
nor U9193 (N_9193,N_8229,N_8828);
nor U9194 (N_9194,N_8073,N_8651);
nand U9195 (N_9195,N_8672,N_8206);
xnor U9196 (N_9196,N_8182,N_8134);
nand U9197 (N_9197,N_8030,N_8624);
nor U9198 (N_9198,N_8100,N_8903);
and U9199 (N_9199,N_8927,N_8806);
and U9200 (N_9200,N_8644,N_8611);
and U9201 (N_9201,N_8810,N_8525);
and U9202 (N_9202,N_8932,N_8834);
nor U9203 (N_9203,N_8760,N_8059);
and U9204 (N_9204,N_8670,N_8310);
or U9205 (N_9205,N_8365,N_8818);
or U9206 (N_9206,N_8445,N_8338);
and U9207 (N_9207,N_8377,N_8843);
and U9208 (N_9208,N_8411,N_8435);
and U9209 (N_9209,N_8553,N_8942);
and U9210 (N_9210,N_8786,N_8388);
and U9211 (N_9211,N_8140,N_8291);
nor U9212 (N_9212,N_8320,N_8552);
nand U9213 (N_9213,N_8327,N_8349);
nor U9214 (N_9214,N_8416,N_8744);
nor U9215 (N_9215,N_8973,N_8967);
and U9216 (N_9216,N_8875,N_8714);
or U9217 (N_9217,N_8842,N_8511);
or U9218 (N_9218,N_8877,N_8721);
and U9219 (N_9219,N_8813,N_8894);
and U9220 (N_9220,N_8196,N_8802);
nor U9221 (N_9221,N_8078,N_8474);
nor U9222 (N_9222,N_8811,N_8523);
nor U9223 (N_9223,N_8664,N_8012);
and U9224 (N_9224,N_8613,N_8279);
and U9225 (N_9225,N_8914,N_8101);
nor U9226 (N_9226,N_8292,N_8188);
nor U9227 (N_9227,N_8278,N_8547);
nand U9228 (N_9228,N_8466,N_8930);
nand U9229 (N_9229,N_8658,N_8582);
nor U9230 (N_9230,N_8592,N_8603);
or U9231 (N_9231,N_8050,N_8368);
nor U9232 (N_9232,N_8719,N_8245);
and U9233 (N_9233,N_8123,N_8450);
xor U9234 (N_9234,N_8103,N_8749);
or U9235 (N_9235,N_8838,N_8299);
xor U9236 (N_9236,N_8939,N_8010);
nand U9237 (N_9237,N_8740,N_8286);
xnor U9238 (N_9238,N_8448,N_8131);
nand U9239 (N_9239,N_8604,N_8688);
nor U9240 (N_9240,N_8888,N_8021);
or U9241 (N_9241,N_8997,N_8805);
nand U9242 (N_9242,N_8247,N_8768);
and U9243 (N_9243,N_8488,N_8090);
xnor U9244 (N_9244,N_8873,N_8723);
or U9245 (N_9245,N_8042,N_8915);
and U9246 (N_9246,N_8181,N_8770);
nand U9247 (N_9247,N_8253,N_8081);
nor U9248 (N_9248,N_8052,N_8794);
or U9249 (N_9249,N_8905,N_8401);
or U9250 (N_9250,N_8147,N_8065);
nand U9251 (N_9251,N_8159,N_8516);
nor U9252 (N_9252,N_8020,N_8198);
and U9253 (N_9253,N_8481,N_8296);
and U9254 (N_9254,N_8746,N_8239);
nand U9255 (N_9255,N_8642,N_8138);
nor U9256 (N_9256,N_8938,N_8049);
nand U9257 (N_9257,N_8745,N_8431);
nor U9258 (N_9258,N_8064,N_8079);
nor U9259 (N_9259,N_8829,N_8183);
or U9260 (N_9260,N_8971,N_8876);
nand U9261 (N_9261,N_8560,N_8150);
nor U9262 (N_9262,N_8860,N_8758);
xnor U9263 (N_9263,N_8120,N_8864);
nor U9264 (N_9264,N_8541,N_8784);
nor U9265 (N_9265,N_8741,N_8831);
xnor U9266 (N_9266,N_8830,N_8711);
and U9267 (N_9267,N_8094,N_8859);
nand U9268 (N_9268,N_8071,N_8909);
nor U9269 (N_9269,N_8733,N_8060);
and U9270 (N_9270,N_8122,N_8132);
nand U9271 (N_9271,N_8956,N_8540);
nand U9272 (N_9272,N_8234,N_8783);
nor U9273 (N_9273,N_8308,N_8882);
or U9274 (N_9274,N_8208,N_8526);
and U9275 (N_9275,N_8548,N_8847);
xor U9276 (N_9276,N_8647,N_8316);
nand U9277 (N_9277,N_8061,N_8974);
nand U9278 (N_9278,N_8673,N_8561);
nor U9279 (N_9279,N_8434,N_8076);
nand U9280 (N_9280,N_8515,N_8298);
nand U9281 (N_9281,N_8302,N_8718);
and U9282 (N_9282,N_8332,N_8407);
and U9283 (N_9283,N_8750,N_8364);
nor U9284 (N_9284,N_8536,N_8621);
nor U9285 (N_9285,N_8173,N_8293);
nor U9286 (N_9286,N_8257,N_8633);
nand U9287 (N_9287,N_8069,N_8350);
or U9288 (N_9288,N_8699,N_8601);
or U9289 (N_9289,N_8722,N_8841);
and U9290 (N_9290,N_8144,N_8734);
or U9291 (N_9291,N_8680,N_8889);
nor U9292 (N_9292,N_8975,N_8677);
nor U9293 (N_9293,N_8839,N_8596);
and U9294 (N_9294,N_8405,N_8230);
or U9295 (N_9295,N_8583,N_8165);
nor U9296 (N_9296,N_8649,N_8580);
and U9297 (N_9297,N_8812,N_8727);
nand U9298 (N_9298,N_8866,N_8395);
or U9299 (N_9299,N_8402,N_8194);
nor U9300 (N_9300,N_8587,N_8111);
nand U9301 (N_9301,N_8862,N_8534);
nand U9302 (N_9302,N_8487,N_8266);
or U9303 (N_9303,N_8345,N_8117);
nand U9304 (N_9304,N_8128,N_8920);
nand U9305 (N_9305,N_8538,N_8522);
and U9306 (N_9306,N_8679,N_8375);
or U9307 (N_9307,N_8290,N_8918);
or U9308 (N_9308,N_8513,N_8537);
nor U9309 (N_9309,N_8352,N_8307);
nor U9310 (N_9310,N_8026,N_8343);
nor U9311 (N_9311,N_8512,N_8219);
nand U9312 (N_9312,N_8314,N_8885);
and U9313 (N_9313,N_8951,N_8950);
or U9314 (N_9314,N_8668,N_8706);
or U9315 (N_9315,N_8410,N_8976);
or U9316 (N_9316,N_8579,N_8398);
or U9317 (N_9317,N_8791,N_8618);
or U9318 (N_9318,N_8823,N_8685);
nand U9319 (N_9319,N_8089,N_8333);
or U9320 (N_9320,N_8943,N_8133);
and U9321 (N_9321,N_8826,N_8337);
and U9322 (N_9322,N_8979,N_8963);
nand U9323 (N_9323,N_8376,N_8978);
and U9324 (N_9324,N_8533,N_8753);
or U9325 (N_9325,N_8855,N_8382);
nand U9326 (N_9326,N_8272,N_8287);
or U9327 (N_9327,N_8822,N_8386);
and U9328 (N_9328,N_8014,N_8608);
nor U9329 (N_9329,N_8616,N_8650);
nor U9330 (N_9330,N_8545,N_8543);
nor U9331 (N_9331,N_8566,N_8226);
or U9332 (N_9332,N_8367,N_8394);
or U9333 (N_9333,N_8562,N_8362);
nand U9334 (N_9334,N_8484,N_8732);
nor U9335 (N_9335,N_8323,N_8224);
nor U9336 (N_9336,N_8028,N_8172);
nand U9337 (N_9337,N_8764,N_8438);
or U9338 (N_9338,N_8984,N_8558);
nor U9339 (N_9339,N_8748,N_8422);
nand U9340 (N_9340,N_8341,N_8105);
nand U9341 (N_9341,N_8166,N_8993);
or U9342 (N_9342,N_8305,N_8074);
nor U9343 (N_9343,N_8032,N_8039);
nor U9344 (N_9344,N_8164,N_8270);
xnor U9345 (N_9345,N_8597,N_8557);
or U9346 (N_9346,N_8824,N_8965);
nor U9347 (N_9347,N_8220,N_8970);
nor U9348 (N_9348,N_8867,N_8408);
and U9349 (N_9349,N_8295,N_8151);
nand U9350 (N_9350,N_8687,N_8480);
nor U9351 (N_9351,N_8955,N_8025);
and U9352 (N_9352,N_8574,N_8099);
xor U9353 (N_9353,N_8130,N_8209);
nand U9354 (N_9354,N_8246,N_8977);
nand U9355 (N_9355,N_8517,N_8742);
and U9356 (N_9356,N_8696,N_8459);
nor U9357 (N_9357,N_8197,N_8419);
nand U9358 (N_9358,N_8539,N_8017);
nand U9359 (N_9359,N_8485,N_8463);
or U9360 (N_9360,N_8590,N_8051);
and U9361 (N_9361,N_8850,N_8509);
xnor U9362 (N_9362,N_8329,N_8846);
or U9363 (N_9363,N_8615,N_8726);
and U9364 (N_9364,N_8004,N_8261);
or U9365 (N_9365,N_8612,N_8361);
nand U9366 (N_9366,N_8896,N_8363);
and U9367 (N_9367,N_8880,N_8593);
nor U9368 (N_9368,N_8439,N_8249);
and U9369 (N_9369,N_8109,N_8728);
nor U9370 (N_9370,N_8610,N_8646);
nor U9371 (N_9371,N_8048,N_8669);
nor U9372 (N_9372,N_8535,N_8589);
nand U9373 (N_9373,N_8383,N_8795);
nor U9374 (N_9374,N_8447,N_8162);
or U9375 (N_9375,N_8827,N_8886);
nand U9376 (N_9376,N_8832,N_8756);
nor U9377 (N_9377,N_8757,N_8496);
nand U9378 (N_9378,N_8170,N_8962);
nor U9379 (N_9379,N_8544,N_8175);
xor U9380 (N_9380,N_8235,N_8772);
xnor U9381 (N_9381,N_8034,N_8113);
or U9382 (N_9382,N_8717,N_8907);
nand U9383 (N_9383,N_8114,N_8233);
and U9384 (N_9384,N_8195,N_8288);
and U9385 (N_9385,N_8972,N_8446);
or U9386 (N_9386,N_8961,N_8180);
nand U9387 (N_9387,N_8153,N_8334);
nor U9388 (N_9388,N_8966,N_8044);
nor U9389 (N_9389,N_8063,N_8763);
xnor U9390 (N_9390,N_8933,N_8415);
or U9391 (N_9391,N_8630,N_8804);
and U9392 (N_9392,N_8869,N_8214);
or U9393 (N_9393,N_8254,N_8256);
nor U9394 (N_9394,N_8663,N_8694);
nor U9395 (N_9395,N_8916,N_8282);
nor U9396 (N_9396,N_8163,N_8007);
or U9397 (N_9397,N_8390,N_8716);
or U9398 (N_9398,N_8062,N_8204);
nand U9399 (N_9399,N_8825,N_8190);
and U9400 (N_9400,N_8142,N_8241);
nor U9401 (N_9401,N_8462,N_8712);
or U9402 (N_9402,N_8342,N_8781);
nand U9403 (N_9403,N_8373,N_8045);
xor U9404 (N_9404,N_8148,N_8154);
nor U9405 (N_9405,N_8857,N_8684);
and U9406 (N_9406,N_8632,N_8244);
or U9407 (N_9407,N_8529,N_8107);
and U9408 (N_9408,N_8035,N_8199);
nand U9409 (N_9409,N_8015,N_8609);
and U9410 (N_9410,N_8803,N_8725);
or U9411 (N_9411,N_8738,N_8112);
or U9412 (N_9412,N_8037,N_8657);
or U9413 (N_9413,N_8635,N_8778);
nor U9414 (N_9414,N_8380,N_8213);
nor U9415 (N_9415,N_8429,N_8009);
nand U9416 (N_9416,N_8625,N_8369);
or U9417 (N_9417,N_8068,N_8127);
and U9418 (N_9418,N_8751,N_8724);
and U9419 (N_9419,N_8622,N_8093);
nand U9420 (N_9420,N_8457,N_8845);
nand U9421 (N_9421,N_8704,N_8550);
nand U9422 (N_9422,N_8731,N_8264);
nor U9423 (N_9423,N_8659,N_8643);
xor U9424 (N_9424,N_8315,N_8271);
nand U9425 (N_9425,N_8255,N_8404);
or U9426 (N_9426,N_8848,N_8453);
nor U9427 (N_9427,N_8844,N_8565);
nor U9428 (N_9428,N_8524,N_8301);
nand U9429 (N_9429,N_8125,N_8935);
nor U9430 (N_9430,N_8571,N_8546);
nor U9431 (N_9431,N_8627,N_8681);
nor U9432 (N_9432,N_8994,N_8683);
nand U9433 (N_9433,N_8902,N_8016);
nand U9434 (N_9434,N_8047,N_8747);
nand U9435 (N_9435,N_8936,N_8325);
xor U9436 (N_9436,N_8656,N_8468);
or U9437 (N_9437,N_8900,N_8913);
nand U9438 (N_9438,N_8959,N_8232);
xnor U9439 (N_9439,N_8987,N_8773);
xor U9440 (N_9440,N_8899,N_8598);
nand U9441 (N_9441,N_8418,N_8743);
and U9442 (N_9442,N_8606,N_8096);
nor U9443 (N_9443,N_8868,N_8225);
nand U9444 (N_9444,N_8080,N_8710);
and U9445 (N_9445,N_8359,N_8347);
or U9446 (N_9446,N_8355,N_8143);
or U9447 (N_9447,N_8115,N_8503);
nand U9448 (N_9448,N_8027,N_8311);
nand U9449 (N_9449,N_8871,N_8146);
or U9450 (N_9450,N_8519,N_8330);
nand U9451 (N_9451,N_8964,N_8765);
nor U9452 (N_9452,N_8024,N_8901);
and U9453 (N_9453,N_8217,N_8884);
or U9454 (N_9454,N_8736,N_8461);
or U9455 (N_9455,N_8137,N_8281);
nor U9456 (N_9456,N_8720,N_8031);
and U9457 (N_9457,N_8586,N_8527);
xnor U9458 (N_9458,N_8124,N_8216);
or U9459 (N_9459,N_8238,N_8737);
or U9460 (N_9460,N_8458,N_8919);
nor U9461 (N_9461,N_8695,N_8022);
nand U9462 (N_9462,N_8698,N_8702);
nand U9463 (N_9463,N_8160,N_8968);
nor U9464 (N_9464,N_8771,N_8250);
nand U9465 (N_9465,N_8479,N_8211);
nor U9466 (N_9466,N_8077,N_8599);
and U9467 (N_9467,N_8348,N_8686);
or U9468 (N_9468,N_8863,N_8110);
nand U9469 (N_9469,N_8267,N_8058);
nand U9470 (N_9470,N_8995,N_8283);
xor U9471 (N_9471,N_8631,N_8427);
xnor U9472 (N_9472,N_8498,N_8572);
or U9473 (N_9473,N_8607,N_8595);
xor U9474 (N_9474,N_8391,N_8851);
or U9475 (N_9475,N_8126,N_8104);
nand U9476 (N_9476,N_8167,N_8581);
nor U9477 (N_9477,N_8898,N_8780);
or U9478 (N_9478,N_8692,N_8417);
nor U9479 (N_9479,N_8559,N_8070);
or U9480 (N_9480,N_8002,N_8157);
nand U9481 (N_9481,N_8600,N_8700);
and U9482 (N_9482,N_8578,N_8983);
nor U9483 (N_9483,N_8176,N_8530);
and U9484 (N_9484,N_8661,N_8705);
nor U9485 (N_9485,N_8793,N_8179);
nor U9486 (N_9486,N_8066,N_8837);
xnor U9487 (N_9487,N_8328,N_8792);
nor U9488 (N_9488,N_8754,N_8374);
or U9489 (N_9489,N_8892,N_8518);
or U9490 (N_9490,N_8202,N_8893);
nand U9491 (N_9491,N_8396,N_8339);
and U9492 (N_9492,N_8853,N_8201);
or U9493 (N_9493,N_8171,N_8508);
nor U9494 (N_9494,N_8514,N_8637);
or U9495 (N_9495,N_8053,N_8309);
and U9496 (N_9496,N_8003,N_8887);
or U9497 (N_9497,N_8761,N_8210);
nor U9498 (N_9498,N_8433,N_8945);
xor U9499 (N_9499,N_8444,N_8969);
xor U9500 (N_9500,N_8573,N_8880);
nor U9501 (N_9501,N_8689,N_8129);
nand U9502 (N_9502,N_8749,N_8342);
nor U9503 (N_9503,N_8306,N_8375);
nor U9504 (N_9504,N_8042,N_8477);
nand U9505 (N_9505,N_8708,N_8020);
and U9506 (N_9506,N_8244,N_8783);
nand U9507 (N_9507,N_8813,N_8948);
nand U9508 (N_9508,N_8453,N_8950);
nor U9509 (N_9509,N_8411,N_8182);
and U9510 (N_9510,N_8868,N_8217);
or U9511 (N_9511,N_8389,N_8743);
or U9512 (N_9512,N_8293,N_8691);
nor U9513 (N_9513,N_8296,N_8519);
xnor U9514 (N_9514,N_8130,N_8548);
xnor U9515 (N_9515,N_8015,N_8284);
or U9516 (N_9516,N_8620,N_8336);
or U9517 (N_9517,N_8765,N_8165);
xor U9518 (N_9518,N_8133,N_8542);
and U9519 (N_9519,N_8916,N_8627);
nand U9520 (N_9520,N_8973,N_8021);
or U9521 (N_9521,N_8923,N_8425);
and U9522 (N_9522,N_8337,N_8241);
and U9523 (N_9523,N_8881,N_8007);
or U9524 (N_9524,N_8939,N_8808);
nand U9525 (N_9525,N_8674,N_8305);
nand U9526 (N_9526,N_8902,N_8544);
nor U9527 (N_9527,N_8128,N_8923);
and U9528 (N_9528,N_8322,N_8157);
or U9529 (N_9529,N_8981,N_8478);
or U9530 (N_9530,N_8610,N_8334);
xor U9531 (N_9531,N_8344,N_8999);
or U9532 (N_9532,N_8921,N_8769);
and U9533 (N_9533,N_8875,N_8547);
nor U9534 (N_9534,N_8951,N_8489);
and U9535 (N_9535,N_8554,N_8257);
and U9536 (N_9536,N_8158,N_8492);
nor U9537 (N_9537,N_8538,N_8713);
nor U9538 (N_9538,N_8504,N_8764);
and U9539 (N_9539,N_8181,N_8185);
xnor U9540 (N_9540,N_8390,N_8782);
nand U9541 (N_9541,N_8640,N_8009);
or U9542 (N_9542,N_8647,N_8638);
xor U9543 (N_9543,N_8784,N_8344);
or U9544 (N_9544,N_8328,N_8998);
xnor U9545 (N_9545,N_8858,N_8181);
or U9546 (N_9546,N_8504,N_8480);
nand U9547 (N_9547,N_8182,N_8114);
nand U9548 (N_9548,N_8844,N_8174);
and U9549 (N_9549,N_8480,N_8426);
and U9550 (N_9550,N_8024,N_8717);
nor U9551 (N_9551,N_8394,N_8049);
nor U9552 (N_9552,N_8802,N_8941);
or U9553 (N_9553,N_8586,N_8496);
xor U9554 (N_9554,N_8678,N_8840);
nand U9555 (N_9555,N_8619,N_8829);
or U9556 (N_9556,N_8801,N_8939);
and U9557 (N_9557,N_8006,N_8799);
xor U9558 (N_9558,N_8185,N_8473);
nand U9559 (N_9559,N_8698,N_8511);
or U9560 (N_9560,N_8891,N_8699);
nor U9561 (N_9561,N_8088,N_8875);
or U9562 (N_9562,N_8537,N_8755);
and U9563 (N_9563,N_8207,N_8926);
nand U9564 (N_9564,N_8733,N_8081);
nand U9565 (N_9565,N_8941,N_8637);
and U9566 (N_9566,N_8494,N_8285);
nor U9567 (N_9567,N_8659,N_8793);
nor U9568 (N_9568,N_8135,N_8583);
and U9569 (N_9569,N_8211,N_8056);
xnor U9570 (N_9570,N_8851,N_8938);
nor U9571 (N_9571,N_8761,N_8485);
nor U9572 (N_9572,N_8227,N_8510);
nor U9573 (N_9573,N_8599,N_8612);
and U9574 (N_9574,N_8619,N_8538);
nor U9575 (N_9575,N_8142,N_8260);
and U9576 (N_9576,N_8808,N_8425);
nand U9577 (N_9577,N_8134,N_8480);
or U9578 (N_9578,N_8570,N_8817);
or U9579 (N_9579,N_8692,N_8320);
or U9580 (N_9580,N_8435,N_8617);
or U9581 (N_9581,N_8062,N_8408);
or U9582 (N_9582,N_8288,N_8046);
and U9583 (N_9583,N_8877,N_8817);
nor U9584 (N_9584,N_8335,N_8290);
and U9585 (N_9585,N_8754,N_8890);
or U9586 (N_9586,N_8453,N_8718);
nand U9587 (N_9587,N_8081,N_8116);
nand U9588 (N_9588,N_8345,N_8565);
and U9589 (N_9589,N_8476,N_8344);
nor U9590 (N_9590,N_8471,N_8046);
nor U9591 (N_9591,N_8578,N_8041);
xnor U9592 (N_9592,N_8086,N_8295);
nand U9593 (N_9593,N_8634,N_8129);
and U9594 (N_9594,N_8088,N_8328);
xnor U9595 (N_9595,N_8787,N_8774);
and U9596 (N_9596,N_8542,N_8755);
nor U9597 (N_9597,N_8795,N_8729);
or U9598 (N_9598,N_8887,N_8345);
and U9599 (N_9599,N_8560,N_8175);
nor U9600 (N_9600,N_8854,N_8736);
nor U9601 (N_9601,N_8970,N_8159);
nand U9602 (N_9602,N_8092,N_8825);
nor U9603 (N_9603,N_8284,N_8092);
nand U9604 (N_9604,N_8401,N_8429);
nand U9605 (N_9605,N_8163,N_8439);
and U9606 (N_9606,N_8298,N_8152);
nand U9607 (N_9607,N_8841,N_8434);
nor U9608 (N_9608,N_8826,N_8039);
or U9609 (N_9609,N_8861,N_8646);
nor U9610 (N_9610,N_8956,N_8632);
or U9611 (N_9611,N_8117,N_8754);
nand U9612 (N_9612,N_8913,N_8833);
or U9613 (N_9613,N_8398,N_8003);
nand U9614 (N_9614,N_8741,N_8923);
and U9615 (N_9615,N_8428,N_8631);
nor U9616 (N_9616,N_8051,N_8127);
and U9617 (N_9617,N_8687,N_8177);
and U9618 (N_9618,N_8403,N_8291);
or U9619 (N_9619,N_8902,N_8190);
or U9620 (N_9620,N_8112,N_8647);
nand U9621 (N_9621,N_8986,N_8373);
nor U9622 (N_9622,N_8718,N_8805);
nand U9623 (N_9623,N_8211,N_8299);
or U9624 (N_9624,N_8597,N_8140);
nand U9625 (N_9625,N_8455,N_8477);
and U9626 (N_9626,N_8004,N_8011);
and U9627 (N_9627,N_8713,N_8050);
and U9628 (N_9628,N_8935,N_8511);
nor U9629 (N_9629,N_8576,N_8469);
xnor U9630 (N_9630,N_8781,N_8855);
nand U9631 (N_9631,N_8669,N_8627);
or U9632 (N_9632,N_8607,N_8433);
nor U9633 (N_9633,N_8549,N_8602);
nand U9634 (N_9634,N_8544,N_8760);
nand U9635 (N_9635,N_8449,N_8830);
nor U9636 (N_9636,N_8886,N_8940);
or U9637 (N_9637,N_8718,N_8670);
nor U9638 (N_9638,N_8240,N_8595);
nor U9639 (N_9639,N_8322,N_8213);
and U9640 (N_9640,N_8775,N_8291);
nor U9641 (N_9641,N_8361,N_8240);
xor U9642 (N_9642,N_8015,N_8303);
and U9643 (N_9643,N_8398,N_8174);
or U9644 (N_9644,N_8310,N_8358);
nand U9645 (N_9645,N_8993,N_8386);
or U9646 (N_9646,N_8756,N_8340);
nor U9647 (N_9647,N_8062,N_8378);
xor U9648 (N_9648,N_8068,N_8217);
nand U9649 (N_9649,N_8731,N_8533);
xnor U9650 (N_9650,N_8732,N_8129);
xor U9651 (N_9651,N_8865,N_8990);
nor U9652 (N_9652,N_8117,N_8137);
and U9653 (N_9653,N_8733,N_8419);
nand U9654 (N_9654,N_8698,N_8082);
nor U9655 (N_9655,N_8756,N_8990);
or U9656 (N_9656,N_8746,N_8106);
and U9657 (N_9657,N_8139,N_8187);
or U9658 (N_9658,N_8524,N_8948);
nand U9659 (N_9659,N_8895,N_8803);
and U9660 (N_9660,N_8790,N_8694);
nor U9661 (N_9661,N_8330,N_8329);
or U9662 (N_9662,N_8396,N_8715);
or U9663 (N_9663,N_8546,N_8060);
xnor U9664 (N_9664,N_8618,N_8498);
nor U9665 (N_9665,N_8461,N_8536);
or U9666 (N_9666,N_8520,N_8204);
or U9667 (N_9667,N_8047,N_8157);
nor U9668 (N_9668,N_8020,N_8359);
nor U9669 (N_9669,N_8326,N_8939);
xor U9670 (N_9670,N_8542,N_8868);
and U9671 (N_9671,N_8823,N_8524);
nor U9672 (N_9672,N_8605,N_8908);
and U9673 (N_9673,N_8405,N_8595);
or U9674 (N_9674,N_8185,N_8195);
nor U9675 (N_9675,N_8799,N_8070);
nor U9676 (N_9676,N_8058,N_8806);
nand U9677 (N_9677,N_8586,N_8987);
nor U9678 (N_9678,N_8644,N_8135);
nor U9679 (N_9679,N_8554,N_8927);
nand U9680 (N_9680,N_8532,N_8490);
or U9681 (N_9681,N_8739,N_8714);
and U9682 (N_9682,N_8991,N_8214);
xnor U9683 (N_9683,N_8027,N_8546);
nand U9684 (N_9684,N_8355,N_8613);
and U9685 (N_9685,N_8796,N_8042);
and U9686 (N_9686,N_8145,N_8350);
nor U9687 (N_9687,N_8903,N_8426);
or U9688 (N_9688,N_8679,N_8970);
nor U9689 (N_9689,N_8167,N_8535);
or U9690 (N_9690,N_8914,N_8539);
or U9691 (N_9691,N_8728,N_8529);
nor U9692 (N_9692,N_8782,N_8906);
and U9693 (N_9693,N_8431,N_8182);
xor U9694 (N_9694,N_8468,N_8128);
nand U9695 (N_9695,N_8701,N_8048);
and U9696 (N_9696,N_8938,N_8628);
nor U9697 (N_9697,N_8713,N_8221);
and U9698 (N_9698,N_8244,N_8156);
nand U9699 (N_9699,N_8464,N_8866);
xnor U9700 (N_9700,N_8989,N_8847);
nand U9701 (N_9701,N_8283,N_8617);
xnor U9702 (N_9702,N_8409,N_8701);
and U9703 (N_9703,N_8284,N_8151);
or U9704 (N_9704,N_8613,N_8021);
nand U9705 (N_9705,N_8319,N_8917);
and U9706 (N_9706,N_8787,N_8873);
nand U9707 (N_9707,N_8952,N_8460);
nand U9708 (N_9708,N_8674,N_8146);
and U9709 (N_9709,N_8380,N_8891);
nor U9710 (N_9710,N_8753,N_8866);
nor U9711 (N_9711,N_8757,N_8154);
or U9712 (N_9712,N_8744,N_8536);
or U9713 (N_9713,N_8939,N_8094);
or U9714 (N_9714,N_8492,N_8773);
nor U9715 (N_9715,N_8243,N_8934);
and U9716 (N_9716,N_8986,N_8205);
and U9717 (N_9717,N_8576,N_8154);
nor U9718 (N_9718,N_8703,N_8809);
nor U9719 (N_9719,N_8651,N_8639);
xor U9720 (N_9720,N_8866,N_8166);
or U9721 (N_9721,N_8122,N_8793);
xor U9722 (N_9722,N_8641,N_8157);
nor U9723 (N_9723,N_8987,N_8857);
nand U9724 (N_9724,N_8317,N_8305);
or U9725 (N_9725,N_8650,N_8977);
nor U9726 (N_9726,N_8389,N_8515);
and U9727 (N_9727,N_8222,N_8174);
and U9728 (N_9728,N_8476,N_8122);
xnor U9729 (N_9729,N_8029,N_8813);
and U9730 (N_9730,N_8685,N_8038);
or U9731 (N_9731,N_8681,N_8243);
and U9732 (N_9732,N_8263,N_8285);
or U9733 (N_9733,N_8270,N_8678);
and U9734 (N_9734,N_8188,N_8988);
nor U9735 (N_9735,N_8744,N_8117);
nor U9736 (N_9736,N_8634,N_8032);
nand U9737 (N_9737,N_8872,N_8493);
and U9738 (N_9738,N_8742,N_8182);
nand U9739 (N_9739,N_8045,N_8714);
or U9740 (N_9740,N_8783,N_8893);
and U9741 (N_9741,N_8228,N_8372);
or U9742 (N_9742,N_8079,N_8309);
nand U9743 (N_9743,N_8789,N_8713);
nor U9744 (N_9744,N_8794,N_8366);
nand U9745 (N_9745,N_8362,N_8591);
and U9746 (N_9746,N_8909,N_8310);
and U9747 (N_9747,N_8847,N_8767);
and U9748 (N_9748,N_8122,N_8286);
and U9749 (N_9749,N_8340,N_8149);
and U9750 (N_9750,N_8984,N_8060);
and U9751 (N_9751,N_8042,N_8447);
nor U9752 (N_9752,N_8170,N_8573);
xor U9753 (N_9753,N_8089,N_8444);
xnor U9754 (N_9754,N_8340,N_8823);
nand U9755 (N_9755,N_8195,N_8854);
or U9756 (N_9756,N_8005,N_8907);
and U9757 (N_9757,N_8859,N_8687);
or U9758 (N_9758,N_8191,N_8513);
and U9759 (N_9759,N_8731,N_8143);
or U9760 (N_9760,N_8934,N_8737);
nand U9761 (N_9761,N_8909,N_8719);
xnor U9762 (N_9762,N_8925,N_8818);
xnor U9763 (N_9763,N_8822,N_8889);
and U9764 (N_9764,N_8630,N_8590);
nor U9765 (N_9765,N_8106,N_8430);
and U9766 (N_9766,N_8114,N_8620);
or U9767 (N_9767,N_8601,N_8125);
nor U9768 (N_9768,N_8921,N_8952);
nor U9769 (N_9769,N_8158,N_8924);
or U9770 (N_9770,N_8644,N_8641);
nor U9771 (N_9771,N_8592,N_8744);
nand U9772 (N_9772,N_8039,N_8719);
and U9773 (N_9773,N_8189,N_8762);
and U9774 (N_9774,N_8231,N_8665);
and U9775 (N_9775,N_8288,N_8253);
xnor U9776 (N_9776,N_8321,N_8144);
xor U9777 (N_9777,N_8223,N_8792);
and U9778 (N_9778,N_8652,N_8586);
nor U9779 (N_9779,N_8239,N_8454);
or U9780 (N_9780,N_8939,N_8165);
nand U9781 (N_9781,N_8942,N_8132);
nor U9782 (N_9782,N_8721,N_8461);
xnor U9783 (N_9783,N_8565,N_8807);
nor U9784 (N_9784,N_8023,N_8429);
or U9785 (N_9785,N_8074,N_8805);
and U9786 (N_9786,N_8593,N_8200);
or U9787 (N_9787,N_8541,N_8719);
or U9788 (N_9788,N_8065,N_8316);
nor U9789 (N_9789,N_8417,N_8267);
nand U9790 (N_9790,N_8217,N_8326);
nand U9791 (N_9791,N_8905,N_8137);
or U9792 (N_9792,N_8736,N_8000);
and U9793 (N_9793,N_8190,N_8113);
or U9794 (N_9794,N_8240,N_8502);
and U9795 (N_9795,N_8402,N_8703);
nor U9796 (N_9796,N_8507,N_8190);
or U9797 (N_9797,N_8659,N_8580);
nand U9798 (N_9798,N_8155,N_8472);
nand U9799 (N_9799,N_8924,N_8527);
nand U9800 (N_9800,N_8624,N_8071);
nor U9801 (N_9801,N_8629,N_8058);
xnor U9802 (N_9802,N_8394,N_8592);
nor U9803 (N_9803,N_8682,N_8425);
nand U9804 (N_9804,N_8388,N_8385);
nand U9805 (N_9805,N_8972,N_8805);
and U9806 (N_9806,N_8927,N_8590);
nor U9807 (N_9807,N_8113,N_8951);
and U9808 (N_9808,N_8379,N_8061);
or U9809 (N_9809,N_8950,N_8496);
and U9810 (N_9810,N_8483,N_8813);
nand U9811 (N_9811,N_8712,N_8789);
nor U9812 (N_9812,N_8570,N_8899);
nand U9813 (N_9813,N_8882,N_8935);
xnor U9814 (N_9814,N_8228,N_8316);
nor U9815 (N_9815,N_8047,N_8391);
nand U9816 (N_9816,N_8191,N_8441);
xor U9817 (N_9817,N_8817,N_8317);
nand U9818 (N_9818,N_8684,N_8087);
nand U9819 (N_9819,N_8946,N_8086);
nor U9820 (N_9820,N_8725,N_8647);
xor U9821 (N_9821,N_8889,N_8182);
nor U9822 (N_9822,N_8631,N_8553);
and U9823 (N_9823,N_8223,N_8817);
nor U9824 (N_9824,N_8387,N_8192);
or U9825 (N_9825,N_8901,N_8987);
xor U9826 (N_9826,N_8295,N_8585);
or U9827 (N_9827,N_8805,N_8732);
or U9828 (N_9828,N_8366,N_8649);
and U9829 (N_9829,N_8905,N_8436);
or U9830 (N_9830,N_8251,N_8576);
and U9831 (N_9831,N_8131,N_8871);
and U9832 (N_9832,N_8541,N_8733);
or U9833 (N_9833,N_8456,N_8976);
nand U9834 (N_9834,N_8477,N_8398);
nor U9835 (N_9835,N_8254,N_8341);
nor U9836 (N_9836,N_8603,N_8454);
nor U9837 (N_9837,N_8655,N_8058);
and U9838 (N_9838,N_8429,N_8899);
xor U9839 (N_9839,N_8266,N_8227);
xnor U9840 (N_9840,N_8323,N_8184);
nand U9841 (N_9841,N_8841,N_8692);
and U9842 (N_9842,N_8954,N_8770);
nor U9843 (N_9843,N_8278,N_8588);
or U9844 (N_9844,N_8605,N_8126);
nor U9845 (N_9845,N_8437,N_8277);
xor U9846 (N_9846,N_8834,N_8926);
nor U9847 (N_9847,N_8171,N_8806);
or U9848 (N_9848,N_8945,N_8936);
nor U9849 (N_9849,N_8024,N_8850);
nor U9850 (N_9850,N_8361,N_8224);
or U9851 (N_9851,N_8646,N_8660);
or U9852 (N_9852,N_8535,N_8861);
nor U9853 (N_9853,N_8462,N_8815);
or U9854 (N_9854,N_8500,N_8822);
nand U9855 (N_9855,N_8428,N_8440);
nand U9856 (N_9856,N_8784,N_8093);
nor U9857 (N_9857,N_8651,N_8120);
xor U9858 (N_9858,N_8648,N_8482);
and U9859 (N_9859,N_8483,N_8728);
or U9860 (N_9860,N_8762,N_8255);
xnor U9861 (N_9861,N_8364,N_8139);
and U9862 (N_9862,N_8519,N_8436);
xnor U9863 (N_9863,N_8688,N_8530);
or U9864 (N_9864,N_8269,N_8197);
nor U9865 (N_9865,N_8610,N_8992);
and U9866 (N_9866,N_8674,N_8073);
and U9867 (N_9867,N_8356,N_8896);
and U9868 (N_9868,N_8298,N_8112);
or U9869 (N_9869,N_8831,N_8381);
nor U9870 (N_9870,N_8335,N_8371);
or U9871 (N_9871,N_8587,N_8255);
nand U9872 (N_9872,N_8640,N_8631);
or U9873 (N_9873,N_8792,N_8420);
nand U9874 (N_9874,N_8157,N_8463);
xnor U9875 (N_9875,N_8728,N_8119);
nand U9876 (N_9876,N_8718,N_8517);
or U9877 (N_9877,N_8197,N_8261);
or U9878 (N_9878,N_8731,N_8383);
or U9879 (N_9879,N_8254,N_8319);
nand U9880 (N_9880,N_8190,N_8128);
nor U9881 (N_9881,N_8513,N_8508);
and U9882 (N_9882,N_8667,N_8823);
or U9883 (N_9883,N_8981,N_8769);
and U9884 (N_9884,N_8870,N_8739);
nor U9885 (N_9885,N_8429,N_8570);
nand U9886 (N_9886,N_8053,N_8365);
nand U9887 (N_9887,N_8194,N_8980);
xnor U9888 (N_9888,N_8384,N_8728);
or U9889 (N_9889,N_8774,N_8495);
nor U9890 (N_9890,N_8668,N_8113);
nand U9891 (N_9891,N_8119,N_8843);
and U9892 (N_9892,N_8311,N_8742);
nand U9893 (N_9893,N_8746,N_8342);
nand U9894 (N_9894,N_8981,N_8742);
or U9895 (N_9895,N_8023,N_8061);
or U9896 (N_9896,N_8869,N_8744);
or U9897 (N_9897,N_8255,N_8862);
or U9898 (N_9898,N_8676,N_8260);
or U9899 (N_9899,N_8578,N_8438);
or U9900 (N_9900,N_8229,N_8549);
or U9901 (N_9901,N_8427,N_8172);
and U9902 (N_9902,N_8083,N_8147);
and U9903 (N_9903,N_8969,N_8553);
and U9904 (N_9904,N_8083,N_8139);
nand U9905 (N_9905,N_8909,N_8374);
nor U9906 (N_9906,N_8704,N_8410);
and U9907 (N_9907,N_8536,N_8305);
nor U9908 (N_9908,N_8265,N_8980);
nand U9909 (N_9909,N_8842,N_8485);
nor U9910 (N_9910,N_8662,N_8423);
and U9911 (N_9911,N_8455,N_8724);
or U9912 (N_9912,N_8043,N_8318);
and U9913 (N_9913,N_8420,N_8065);
nor U9914 (N_9914,N_8788,N_8656);
nor U9915 (N_9915,N_8694,N_8443);
nand U9916 (N_9916,N_8774,N_8303);
nor U9917 (N_9917,N_8089,N_8136);
nor U9918 (N_9918,N_8142,N_8590);
or U9919 (N_9919,N_8293,N_8209);
or U9920 (N_9920,N_8657,N_8469);
nor U9921 (N_9921,N_8271,N_8698);
nor U9922 (N_9922,N_8542,N_8823);
or U9923 (N_9923,N_8979,N_8804);
or U9924 (N_9924,N_8274,N_8248);
nor U9925 (N_9925,N_8882,N_8708);
or U9926 (N_9926,N_8242,N_8874);
xor U9927 (N_9927,N_8980,N_8336);
nand U9928 (N_9928,N_8191,N_8260);
nor U9929 (N_9929,N_8289,N_8570);
nand U9930 (N_9930,N_8302,N_8437);
and U9931 (N_9931,N_8900,N_8367);
and U9932 (N_9932,N_8339,N_8083);
or U9933 (N_9933,N_8951,N_8079);
or U9934 (N_9934,N_8771,N_8920);
or U9935 (N_9935,N_8476,N_8564);
nor U9936 (N_9936,N_8992,N_8243);
nor U9937 (N_9937,N_8148,N_8287);
nand U9938 (N_9938,N_8154,N_8648);
nor U9939 (N_9939,N_8945,N_8141);
nand U9940 (N_9940,N_8352,N_8279);
or U9941 (N_9941,N_8781,N_8404);
xor U9942 (N_9942,N_8322,N_8302);
and U9943 (N_9943,N_8904,N_8819);
and U9944 (N_9944,N_8863,N_8083);
xor U9945 (N_9945,N_8700,N_8880);
nand U9946 (N_9946,N_8751,N_8898);
nand U9947 (N_9947,N_8833,N_8890);
and U9948 (N_9948,N_8130,N_8410);
and U9949 (N_9949,N_8681,N_8164);
and U9950 (N_9950,N_8956,N_8695);
and U9951 (N_9951,N_8653,N_8620);
nor U9952 (N_9952,N_8487,N_8325);
nor U9953 (N_9953,N_8950,N_8585);
and U9954 (N_9954,N_8949,N_8271);
nor U9955 (N_9955,N_8383,N_8329);
nor U9956 (N_9956,N_8677,N_8316);
xor U9957 (N_9957,N_8691,N_8168);
nor U9958 (N_9958,N_8639,N_8080);
and U9959 (N_9959,N_8414,N_8208);
nor U9960 (N_9960,N_8253,N_8530);
nand U9961 (N_9961,N_8949,N_8270);
and U9962 (N_9962,N_8065,N_8651);
and U9963 (N_9963,N_8238,N_8174);
nand U9964 (N_9964,N_8943,N_8282);
nor U9965 (N_9965,N_8644,N_8297);
nor U9966 (N_9966,N_8223,N_8178);
xnor U9967 (N_9967,N_8857,N_8078);
nand U9968 (N_9968,N_8223,N_8488);
nor U9969 (N_9969,N_8571,N_8411);
and U9970 (N_9970,N_8187,N_8176);
nand U9971 (N_9971,N_8654,N_8639);
and U9972 (N_9972,N_8557,N_8442);
xor U9973 (N_9973,N_8810,N_8451);
and U9974 (N_9974,N_8016,N_8124);
and U9975 (N_9975,N_8772,N_8456);
nor U9976 (N_9976,N_8185,N_8582);
xor U9977 (N_9977,N_8229,N_8842);
nor U9978 (N_9978,N_8252,N_8038);
nor U9979 (N_9979,N_8308,N_8662);
or U9980 (N_9980,N_8204,N_8410);
nand U9981 (N_9981,N_8921,N_8377);
nor U9982 (N_9982,N_8988,N_8511);
xor U9983 (N_9983,N_8207,N_8470);
nand U9984 (N_9984,N_8926,N_8720);
nand U9985 (N_9985,N_8313,N_8635);
xnor U9986 (N_9986,N_8063,N_8210);
and U9987 (N_9987,N_8586,N_8140);
and U9988 (N_9988,N_8521,N_8729);
nand U9989 (N_9989,N_8038,N_8173);
and U9990 (N_9990,N_8640,N_8199);
and U9991 (N_9991,N_8942,N_8796);
and U9992 (N_9992,N_8335,N_8560);
nor U9993 (N_9993,N_8813,N_8733);
nand U9994 (N_9994,N_8196,N_8478);
nand U9995 (N_9995,N_8342,N_8109);
and U9996 (N_9996,N_8566,N_8745);
nand U9997 (N_9997,N_8127,N_8891);
or U9998 (N_9998,N_8513,N_8216);
and U9999 (N_9999,N_8317,N_8327);
nor U10000 (N_10000,N_9445,N_9118);
nand U10001 (N_10001,N_9657,N_9642);
nor U10002 (N_10002,N_9492,N_9192);
xor U10003 (N_10003,N_9344,N_9408);
or U10004 (N_10004,N_9833,N_9935);
and U10005 (N_10005,N_9755,N_9858);
nor U10006 (N_10006,N_9865,N_9355);
and U10007 (N_10007,N_9184,N_9191);
or U10008 (N_10008,N_9212,N_9633);
or U10009 (N_10009,N_9526,N_9233);
and U10010 (N_10010,N_9586,N_9473);
nand U10011 (N_10011,N_9495,N_9121);
nor U10012 (N_10012,N_9245,N_9747);
nand U10013 (N_10013,N_9579,N_9977);
or U10014 (N_10014,N_9683,N_9332);
or U10015 (N_10015,N_9005,N_9839);
nor U10016 (N_10016,N_9599,N_9261);
or U10017 (N_10017,N_9360,N_9841);
or U10018 (N_10018,N_9416,N_9109);
nand U10019 (N_10019,N_9565,N_9793);
nand U10020 (N_10020,N_9139,N_9851);
nor U10021 (N_10021,N_9760,N_9933);
and U10022 (N_10022,N_9291,N_9311);
nor U10023 (N_10023,N_9024,N_9187);
or U10024 (N_10024,N_9295,N_9556);
nor U10025 (N_10025,N_9183,N_9217);
nor U10026 (N_10026,N_9924,N_9477);
xnor U10027 (N_10027,N_9074,N_9255);
or U10028 (N_10028,N_9867,N_9919);
nor U10029 (N_10029,N_9265,N_9016);
xor U10030 (N_10030,N_9736,N_9881);
and U10031 (N_10031,N_9649,N_9509);
and U10032 (N_10032,N_9198,N_9860);
and U10033 (N_10033,N_9425,N_9338);
nor U10034 (N_10034,N_9120,N_9010);
and U10035 (N_10035,N_9426,N_9004);
xnor U10036 (N_10036,N_9915,N_9067);
or U10037 (N_10037,N_9136,N_9123);
and U10038 (N_10038,N_9443,N_9751);
or U10039 (N_10039,N_9316,N_9286);
and U10040 (N_10040,N_9968,N_9487);
nand U10041 (N_10041,N_9038,N_9127);
nand U10042 (N_10042,N_9252,N_9454);
nor U10043 (N_10043,N_9373,N_9668);
or U10044 (N_10044,N_9665,N_9825);
or U10045 (N_10045,N_9208,N_9080);
or U10046 (N_10046,N_9838,N_9959);
nor U10047 (N_10047,N_9718,N_9436);
nand U10048 (N_10048,N_9814,N_9196);
and U10049 (N_10049,N_9965,N_9099);
nand U10050 (N_10050,N_9088,N_9435);
nor U10051 (N_10051,N_9894,N_9060);
nor U10052 (N_10052,N_9412,N_9388);
xor U10053 (N_10053,N_9744,N_9557);
nand U10054 (N_10054,N_9802,N_9882);
nand U10055 (N_10055,N_9446,N_9972);
and U10056 (N_10056,N_9626,N_9485);
and U10057 (N_10057,N_9110,N_9571);
and U10058 (N_10058,N_9876,N_9948);
and U10059 (N_10059,N_9672,N_9409);
nor U10060 (N_10060,N_9214,N_9997);
nor U10061 (N_10061,N_9813,N_9122);
xor U10062 (N_10062,N_9149,N_9155);
xnor U10063 (N_10063,N_9264,N_9078);
nand U10064 (N_10064,N_9030,N_9750);
and U10065 (N_10065,N_9752,N_9336);
and U10066 (N_10066,N_9723,N_9367);
nand U10067 (N_10067,N_9569,N_9674);
nor U10068 (N_10068,N_9070,N_9874);
and U10069 (N_10069,N_9358,N_9743);
nor U10070 (N_10070,N_9541,N_9848);
nand U10071 (N_10071,N_9600,N_9021);
nor U10072 (N_10072,N_9902,N_9352);
and U10073 (N_10073,N_9639,N_9385);
and U10074 (N_10074,N_9577,N_9789);
and U10075 (N_10075,N_9998,N_9239);
or U10076 (N_10076,N_9199,N_9654);
or U10077 (N_10077,N_9133,N_9787);
nand U10078 (N_10078,N_9660,N_9119);
and U10079 (N_10079,N_9234,N_9077);
or U10080 (N_10080,N_9927,N_9730);
nor U10081 (N_10081,N_9921,N_9886);
nand U10082 (N_10082,N_9469,N_9319);
and U10083 (N_10083,N_9975,N_9417);
or U10084 (N_10084,N_9065,N_9189);
nor U10085 (N_10085,N_9700,N_9856);
nor U10086 (N_10086,N_9872,N_9363);
nor U10087 (N_10087,N_9103,N_9903);
and U10088 (N_10088,N_9174,N_9505);
nor U10089 (N_10089,N_9173,N_9457);
nand U10090 (N_10090,N_9990,N_9022);
nand U10091 (N_10091,N_9900,N_9580);
or U10092 (N_10092,N_9731,N_9879);
xor U10093 (N_10093,N_9695,N_9595);
nand U10094 (N_10094,N_9896,N_9000);
and U10095 (N_10095,N_9147,N_9606);
nor U10096 (N_10096,N_9464,N_9800);
nand U10097 (N_10097,N_9152,N_9073);
nor U10098 (N_10098,N_9296,N_9346);
nor U10099 (N_10099,N_9284,N_9738);
or U10100 (N_10100,N_9969,N_9034);
and U10101 (N_10101,N_9510,N_9474);
and U10102 (N_10102,N_9986,N_9148);
or U10103 (N_10103,N_9713,N_9891);
nor U10104 (N_10104,N_9535,N_9341);
nor U10105 (N_10105,N_9039,N_9166);
nor U10106 (N_10106,N_9863,N_9244);
nor U10107 (N_10107,N_9223,N_9524);
or U10108 (N_10108,N_9098,N_9321);
nand U10109 (N_10109,N_9826,N_9514);
nor U10110 (N_10110,N_9923,N_9721);
nand U10111 (N_10111,N_9973,N_9156);
nand U10112 (N_10112,N_9203,N_9768);
nor U10113 (N_10113,N_9953,N_9502);
nor U10114 (N_10114,N_9847,N_9684);
nand U10115 (N_10115,N_9943,N_9353);
nor U10116 (N_10116,N_9936,N_9515);
nor U10117 (N_10117,N_9877,N_9076);
and U10118 (N_10118,N_9281,N_9006);
xnor U10119 (N_10119,N_9185,N_9503);
and U10120 (N_10120,N_9047,N_9609);
nand U10121 (N_10121,N_9082,N_9910);
nor U10122 (N_10122,N_9971,N_9624);
nand U10123 (N_10123,N_9611,N_9162);
or U10124 (N_10124,N_9691,N_9270);
or U10125 (N_10125,N_9266,N_9898);
nand U10126 (N_10126,N_9093,N_9799);
nand U10127 (N_10127,N_9737,N_9932);
and U10128 (N_10128,N_9220,N_9638);
nor U10129 (N_10129,N_9568,N_9688);
xor U10130 (N_10130,N_9576,N_9529);
nand U10131 (N_10131,N_9985,N_9947);
or U10132 (N_10132,N_9844,N_9887);
and U10133 (N_10133,N_9419,N_9717);
nor U10134 (N_10134,N_9928,N_9170);
and U10135 (N_10135,N_9071,N_9072);
and U10136 (N_10136,N_9494,N_9250);
and U10137 (N_10137,N_9622,N_9539);
and U10138 (N_10138,N_9958,N_9728);
nor U10139 (N_10139,N_9091,N_9520);
or U10140 (N_10140,N_9020,N_9329);
nand U10141 (N_10141,N_9940,N_9013);
or U10142 (N_10142,N_9612,N_9132);
xor U10143 (N_10143,N_9774,N_9243);
nor U10144 (N_10144,N_9792,N_9201);
nand U10145 (N_10145,N_9868,N_9584);
nor U10146 (N_10146,N_9931,N_9770);
and U10147 (N_10147,N_9242,N_9008);
xnor U10148 (N_10148,N_9478,N_9262);
and U10149 (N_10149,N_9164,N_9298);
nor U10150 (N_10150,N_9756,N_9432);
and U10151 (N_10151,N_9431,N_9791);
nand U10152 (N_10152,N_9112,N_9089);
or U10153 (N_10153,N_9536,N_9277);
and U10154 (N_10154,N_9075,N_9866);
xor U10155 (N_10155,N_9596,N_9617);
and U10156 (N_10156,N_9330,N_9548);
nand U10157 (N_10157,N_9805,N_9911);
nand U10158 (N_10158,N_9371,N_9517);
nand U10159 (N_10159,N_9427,N_9283);
xnor U10160 (N_10160,N_9983,N_9141);
and U10161 (N_10161,N_9776,N_9249);
nor U10162 (N_10162,N_9202,N_9007);
nand U10163 (N_10163,N_9854,N_9429);
and U10164 (N_10164,N_9402,N_9126);
nand U10165 (N_10165,N_9028,N_9258);
xor U10166 (N_10166,N_9689,N_9117);
nor U10167 (N_10167,N_9914,N_9177);
and U10168 (N_10168,N_9094,N_9922);
nand U10169 (N_10169,N_9168,N_9303);
nor U10170 (N_10170,N_9500,N_9871);
nor U10171 (N_10171,N_9285,N_9583);
and U10172 (N_10172,N_9974,N_9530);
or U10173 (N_10173,N_9131,N_9257);
nor U10174 (N_10174,N_9130,N_9690);
or U10175 (N_10175,N_9267,N_9380);
and U10176 (N_10176,N_9661,N_9328);
and U10177 (N_10177,N_9444,N_9128);
nor U10178 (N_10178,N_9383,N_9835);
xor U10179 (N_10179,N_9241,N_9061);
nand U10180 (N_10180,N_9486,N_9716);
and U10181 (N_10181,N_9205,N_9084);
nand U10182 (N_10182,N_9354,N_9307);
or U10183 (N_10183,N_9056,N_9221);
and U10184 (N_10184,N_9890,N_9729);
nor U10185 (N_10185,N_9146,N_9229);
nor U10186 (N_10186,N_9237,N_9063);
nand U10187 (N_10187,N_9323,N_9154);
nand U10188 (N_10188,N_9979,N_9667);
nand U10189 (N_10189,N_9470,N_9224);
xnor U10190 (N_10190,N_9273,N_9389);
or U10191 (N_10191,N_9562,N_9418);
nor U10192 (N_10192,N_9315,N_9238);
or U10193 (N_10193,N_9398,N_9666);
nor U10194 (N_10194,N_9913,N_9885);
or U10195 (N_10195,N_9036,N_9646);
or U10196 (N_10196,N_9995,N_9925);
nand U10197 (N_10197,N_9857,N_9859);
nand U10198 (N_10198,N_9806,N_9878);
nor U10199 (N_10199,N_9533,N_9727);
or U10200 (N_10200,N_9554,N_9163);
and U10201 (N_10201,N_9846,N_9804);
or U10202 (N_10202,N_9675,N_9193);
or U10203 (N_10203,N_9157,N_9853);
and U10204 (N_10204,N_9897,N_9137);
or U10205 (N_10205,N_9655,N_9538);
and U10206 (N_10206,N_9165,N_9767);
and U10207 (N_10207,N_9829,N_9134);
and U10208 (N_10208,N_9899,N_9780);
nor U10209 (N_10209,N_9961,N_9400);
and U10210 (N_10210,N_9917,N_9403);
nor U10211 (N_10211,N_9382,N_9452);
nand U10212 (N_10212,N_9359,N_9694);
and U10213 (N_10213,N_9081,N_9984);
nand U10214 (N_10214,N_9987,N_9545);
or U10215 (N_10215,N_9345,N_9287);
or U10216 (N_10216,N_9339,N_9050);
nand U10217 (N_10217,N_9994,N_9941);
and U10218 (N_10218,N_9171,N_9379);
nor U10219 (N_10219,N_9439,N_9629);
xor U10220 (N_10220,N_9837,N_9488);
xnor U10221 (N_10221,N_9489,N_9294);
and U10222 (N_10222,N_9957,N_9108);
nand U10223 (N_10223,N_9893,N_9410);
and U10224 (N_10224,N_9951,N_9317);
nor U10225 (N_10225,N_9522,N_9699);
or U10226 (N_10226,N_9288,N_9766);
and U10227 (N_10227,N_9322,N_9591);
and U10228 (N_10228,N_9991,N_9889);
nor U10229 (N_10229,N_9875,N_9479);
nor U10230 (N_10230,N_9635,N_9604);
nor U10231 (N_10231,N_9176,N_9278);
and U10232 (N_10232,N_9715,N_9459);
or U10233 (N_10233,N_9786,N_9821);
nand U10234 (N_10234,N_9546,N_9735);
and U10235 (N_10235,N_9504,N_9930);
nand U10236 (N_10236,N_9926,N_9669);
xor U10237 (N_10237,N_9395,N_9671);
nor U10238 (N_10238,N_9151,N_9032);
nor U10239 (N_10239,N_9777,N_9269);
or U10240 (N_10240,N_9605,N_9864);
or U10241 (N_10241,N_9049,N_9450);
or U10242 (N_10242,N_9200,N_9696);
nor U10243 (N_10243,N_9705,N_9460);
nand U10244 (N_10244,N_9348,N_9681);
and U10245 (N_10245,N_9785,N_9543);
nor U10246 (N_10246,N_9892,N_9746);
and U10247 (N_10247,N_9437,N_9456);
nor U10248 (N_10248,N_9368,N_9788);
and U10249 (N_10249,N_9630,N_9906);
or U10250 (N_10250,N_9782,N_9818);
and U10251 (N_10251,N_9017,N_9748);
nor U10252 (N_10252,N_9350,N_9623);
nand U10253 (N_10253,N_9300,N_9033);
or U10254 (N_10254,N_9194,N_9027);
and U10255 (N_10255,N_9415,N_9945);
and U10256 (N_10256,N_9227,N_9645);
or U10257 (N_10257,N_9506,N_9180);
nor U10258 (N_10258,N_9428,N_9167);
or U10259 (N_10259,N_9678,N_9918);
nand U10260 (N_10260,N_9158,N_9706);
xor U10261 (N_10261,N_9702,N_9779);
xnor U10262 (N_10262,N_9764,N_9362);
nor U10263 (N_10263,N_9337,N_9222);
and U10264 (N_10264,N_9585,N_9026);
and U10265 (N_10265,N_9824,N_9920);
nor U10266 (N_10266,N_9433,N_9083);
nor U10267 (N_10267,N_9324,N_9095);
and U10268 (N_10268,N_9527,N_9686);
nor U10269 (N_10269,N_9320,N_9603);
nor U10270 (N_10270,N_9765,N_9213);
xor U10271 (N_10271,N_9331,N_9516);
nand U10272 (N_10272,N_9401,N_9551);
or U10273 (N_10273,N_9652,N_9364);
or U10274 (N_10274,N_9465,N_9542);
nand U10275 (N_10275,N_9447,N_9830);
nand U10276 (N_10276,N_9904,N_9182);
nor U10277 (N_10277,N_9293,N_9326);
xor U10278 (N_10278,N_9009,N_9231);
nor U10279 (N_10279,N_9497,N_9312);
nor U10280 (N_10280,N_9399,N_9276);
nand U10281 (N_10281,N_9905,N_9901);
nor U10282 (N_10282,N_9944,N_9484);
nor U10283 (N_10283,N_9758,N_9757);
and U10284 (N_10284,N_9632,N_9097);
and U10285 (N_10285,N_9340,N_9811);
or U10286 (N_10286,N_9390,N_9989);
or U10287 (N_10287,N_9387,N_9218);
or U10288 (N_10288,N_9619,N_9434);
nand U10289 (N_10289,N_9796,N_9370);
nand U10290 (N_10290,N_9361,N_9292);
nor U10291 (N_10291,N_9710,N_9570);
and U10292 (N_10292,N_9153,N_9960);
or U10293 (N_10293,N_9513,N_9150);
or U10294 (N_10294,N_9396,N_9111);
nand U10295 (N_10295,N_9140,N_9608);
nand U10296 (N_10296,N_9215,N_9376);
nand U10297 (N_10297,N_9880,N_9204);
nor U10298 (N_10298,N_9762,N_9884);
and U10299 (N_10299,N_9680,N_9698);
or U10300 (N_10300,N_9423,N_9697);
and U10301 (N_10301,N_9421,N_9745);
or U10302 (N_10302,N_9976,N_9781);
xnor U10303 (N_10303,N_9572,N_9453);
and U10304 (N_10304,N_9086,N_9302);
or U10305 (N_10305,N_9929,N_9422);
nor U10306 (N_10306,N_9325,N_9314);
or U10307 (N_10307,N_9734,N_9310);
nor U10308 (N_10308,N_9334,N_9031);
nand U10309 (N_10309,N_9240,N_9618);
nor U10310 (N_10310,N_9801,N_9553);
nand U10311 (N_10311,N_9607,N_9996);
nand U10312 (N_10312,N_9988,N_9692);
nor U10313 (N_10313,N_9406,N_9581);
and U10314 (N_10314,N_9753,N_9308);
and U10315 (N_10315,N_9491,N_9209);
nor U10316 (N_10316,N_9544,N_9849);
and U10317 (N_10317,N_9381,N_9125);
nand U10318 (N_10318,N_9018,N_9175);
nor U10319 (N_10319,N_9057,N_9682);
nand U10320 (N_10320,N_9247,N_9643);
or U10321 (N_10321,N_9301,N_9934);
or U10322 (N_10322,N_9615,N_9869);
nand U10323 (N_10323,N_9335,N_9197);
and U10324 (N_10324,N_9145,N_9739);
and U10325 (N_10325,N_9659,N_9613);
and U10326 (N_10326,N_9820,N_9179);
or U10327 (N_10327,N_9420,N_9366);
or U10328 (N_10328,N_9616,N_9587);
nor U10329 (N_10329,N_9950,N_9405);
nand U10330 (N_10330,N_9161,N_9532);
and U10331 (N_10331,N_9481,N_9963);
and U10332 (N_10332,N_9592,N_9575);
or U10333 (N_10333,N_9594,N_9236);
nor U10334 (N_10334,N_9773,N_9663);
nand U10335 (N_10335,N_9413,N_9783);
nand U10336 (N_10336,N_9138,N_9582);
or U10337 (N_10337,N_9507,N_9519);
or U10338 (N_10338,N_9590,N_9377);
nand U10339 (N_10339,N_9102,N_9949);
nand U10340 (N_10340,N_9512,N_9306);
nand U10341 (N_10341,N_9463,N_9304);
nor U10342 (N_10342,N_9707,N_9823);
xor U10343 (N_10343,N_9498,N_9712);
nor U10344 (N_10344,N_9725,N_9620);
and U10345 (N_10345,N_9054,N_9318);
and U10346 (N_10346,N_9101,N_9828);
or U10347 (N_10347,N_9407,N_9115);
or U10348 (N_10348,N_9563,N_9106);
nand U10349 (N_10349,N_9651,N_9521);
nand U10350 (N_10350,N_9939,N_9219);
nand U10351 (N_10351,N_9169,N_9843);
xor U10352 (N_10352,N_9475,N_9836);
xnor U10353 (N_10353,N_9206,N_9862);
or U10354 (N_10354,N_9327,N_9593);
or U10355 (N_10355,N_9499,N_9794);
and U10356 (N_10356,N_9096,N_9573);
nor U10357 (N_10357,N_9042,N_9525);
or U10358 (N_10358,N_9567,N_9916);
or U10359 (N_10359,N_9614,N_9256);
nor U10360 (N_10360,N_9537,N_9597);
nor U10361 (N_10361,N_9834,N_9430);
or U10362 (N_10362,N_9656,N_9803);
and U10363 (N_10363,N_9845,N_9634);
nor U10364 (N_10364,N_9392,N_9181);
nand U10365 (N_10365,N_9662,N_9810);
and U10366 (N_10366,N_9135,N_9955);
nand U10367 (N_10367,N_9769,N_9547);
nand U10368 (N_10368,N_9374,N_9650);
and U10369 (N_10369,N_9482,N_9722);
nor U10370 (N_10370,N_9448,N_9601);
and U10371 (N_10371,N_9822,N_9564);
nand U10372 (N_10372,N_9003,N_9775);
nor U10373 (N_10373,N_9966,N_9888);
nand U10374 (N_10374,N_9832,N_9347);
nor U10375 (N_10375,N_9978,N_9740);
and U10376 (N_10376,N_9211,N_9907);
or U10377 (N_10377,N_9647,N_9462);
or U10378 (N_10378,N_9272,N_9708);
nor U10379 (N_10379,N_9589,N_9260);
nor U10380 (N_10380,N_9226,N_9411);
and U10381 (N_10381,N_9693,N_9942);
and U10382 (N_10382,N_9952,N_9160);
nand U10383 (N_10383,N_9230,N_9068);
nand U10384 (N_10384,N_9391,N_9357);
nand U10385 (N_10385,N_9046,N_9658);
nor U10386 (N_10386,N_9263,N_9274);
nand U10387 (N_10387,N_9369,N_9704);
nor U10388 (N_10388,N_9908,N_9967);
nand U10389 (N_10389,N_9560,N_9351);
and U10390 (N_10390,N_9384,N_9534);
nand U10391 (N_10391,N_9195,N_9946);
and U10392 (N_10392,N_9784,N_9631);
or U10393 (N_10393,N_9540,N_9029);
or U10394 (N_10394,N_9602,N_9644);
and U10395 (N_10395,N_9912,N_9275);
nor U10396 (N_10396,N_9641,N_9937);
nand U10397 (N_10397,N_9610,N_9778);
xnor U10398 (N_10398,N_9999,N_9962);
and U10399 (N_10399,N_9059,N_9552);
or U10400 (N_10400,N_9051,N_9055);
and U10401 (N_10401,N_9414,N_9225);
and U10402 (N_10402,N_9116,N_9025);
nand U10403 (N_10403,N_9850,N_9523);
and U10404 (N_10404,N_9490,N_9687);
nand U10405 (N_10405,N_9290,N_9559);
or U10406 (N_10406,N_9041,N_9964);
or U10407 (N_10407,N_9842,N_9714);
nor U10408 (N_10408,N_9113,N_9636);
or U10409 (N_10409,N_9812,N_9720);
nand U10410 (N_10410,N_9259,N_9528);
nand U10411 (N_10411,N_9044,N_9466);
and U10412 (N_10412,N_9449,N_9909);
and U10413 (N_10413,N_9982,N_9092);
nand U10414 (N_10414,N_9043,N_9216);
or U10415 (N_10415,N_9471,N_9207);
nand U10416 (N_10416,N_9472,N_9142);
nand U10417 (N_10417,N_9754,N_9129);
and U10418 (N_10418,N_9625,N_9069);
nand U10419 (N_10419,N_9733,N_9701);
xor U10420 (N_10420,N_9365,N_9628);
or U10421 (N_10421,N_9759,N_9297);
xnor U10422 (N_10422,N_9468,N_9627);
xor U10423 (N_10423,N_9980,N_9808);
nand U10424 (N_10424,N_9493,N_9861);
or U10425 (N_10425,N_9852,N_9394);
or U10426 (N_10426,N_9040,N_9188);
xor U10427 (N_10427,N_9483,N_9703);
nand U10428 (N_10428,N_9819,N_9461);
nor U10429 (N_10429,N_9002,N_9124);
nand U10430 (N_10430,N_9114,N_9476);
and U10431 (N_10431,N_9001,N_9079);
or U10432 (N_10432,N_9685,N_9578);
xnor U10433 (N_10433,N_9100,N_9664);
xnor U10434 (N_10434,N_9732,N_9561);
and U10435 (N_10435,N_9232,N_9763);
nor U10436 (N_10436,N_9282,N_9741);
or U10437 (N_10437,N_9105,N_9992);
nand U10438 (N_10438,N_9438,N_9555);
and U10439 (N_10439,N_9235,N_9574);
or U10440 (N_10440,N_9378,N_9015);
and U10441 (N_10441,N_9254,N_9558);
xor U10442 (N_10442,N_9809,N_9840);
nand U10443 (N_10443,N_9305,N_9397);
or U10444 (N_10444,N_9090,N_9045);
and U10445 (N_10445,N_9037,N_9795);
or U10446 (N_10446,N_9404,N_9549);
xnor U10447 (N_10447,N_9143,N_9014);
nor U10448 (N_10448,N_9064,N_9676);
and U10449 (N_10449,N_9816,N_9019);
nor U10450 (N_10450,N_9954,N_9653);
or U10451 (N_10451,N_9313,N_9679);
nand U10452 (N_10452,N_9956,N_9372);
or U10453 (N_10453,N_9451,N_9210);
nor U10454 (N_10454,N_9761,N_9981);
nand U10455 (N_10455,N_9333,N_9279);
and U10456 (N_10456,N_9458,N_9343);
nand U10457 (N_10457,N_9742,N_9228);
nand U10458 (N_10458,N_9356,N_9511);
nor U10459 (N_10459,N_9467,N_9870);
and U10460 (N_10460,N_9066,N_9455);
and U10461 (N_10461,N_9253,N_9062);
nor U10462 (N_10462,N_9807,N_9709);
and U10463 (N_10463,N_9011,N_9531);
nor U10464 (N_10464,N_9719,N_9749);
and U10465 (N_10465,N_9442,N_9790);
and U10466 (N_10466,N_9827,N_9883);
xor U10467 (N_10467,N_9831,N_9724);
nand U10468 (N_10468,N_9817,N_9938);
xnor U10469 (N_10469,N_9797,N_9711);
nor U10470 (N_10470,N_9190,N_9566);
nand U10471 (N_10471,N_9012,N_9159);
or U10472 (N_10472,N_9440,N_9771);
or U10473 (N_10473,N_9726,N_9993);
nor U10474 (N_10474,N_9052,N_9309);
or U10475 (N_10475,N_9375,N_9251);
nor U10476 (N_10476,N_9248,N_9508);
nand U10477 (N_10477,N_9299,N_9648);
nor U10478 (N_10478,N_9271,N_9501);
nor U10479 (N_10479,N_9588,N_9280);
and U10480 (N_10480,N_9970,N_9873);
nand U10481 (N_10481,N_9104,N_9855);
or U10482 (N_10482,N_9058,N_9621);
nor U10483 (N_10483,N_9550,N_9677);
or U10484 (N_10484,N_9172,N_9268);
nor U10485 (N_10485,N_9035,N_9107);
nand U10486 (N_10486,N_9087,N_9441);
xnor U10487 (N_10487,N_9342,N_9053);
and U10488 (N_10488,N_9085,N_9386);
and U10489 (N_10489,N_9798,N_9480);
nand U10490 (N_10490,N_9673,N_9246);
nor U10491 (N_10491,N_9393,N_9178);
nor U10492 (N_10492,N_9815,N_9289);
and U10493 (N_10493,N_9349,N_9772);
nor U10494 (N_10494,N_9518,N_9186);
xnor U10495 (N_10495,N_9637,N_9640);
and U10496 (N_10496,N_9670,N_9023);
nand U10497 (N_10497,N_9424,N_9895);
and U10498 (N_10498,N_9144,N_9048);
or U10499 (N_10499,N_9496,N_9598);
nand U10500 (N_10500,N_9996,N_9910);
or U10501 (N_10501,N_9874,N_9509);
or U10502 (N_10502,N_9138,N_9927);
nand U10503 (N_10503,N_9914,N_9271);
nand U10504 (N_10504,N_9333,N_9582);
and U10505 (N_10505,N_9940,N_9706);
or U10506 (N_10506,N_9847,N_9851);
or U10507 (N_10507,N_9610,N_9811);
and U10508 (N_10508,N_9570,N_9157);
nand U10509 (N_10509,N_9178,N_9285);
xor U10510 (N_10510,N_9450,N_9317);
and U10511 (N_10511,N_9175,N_9548);
nor U10512 (N_10512,N_9725,N_9770);
nand U10513 (N_10513,N_9648,N_9601);
and U10514 (N_10514,N_9538,N_9433);
nor U10515 (N_10515,N_9545,N_9491);
or U10516 (N_10516,N_9912,N_9987);
nand U10517 (N_10517,N_9490,N_9496);
xnor U10518 (N_10518,N_9660,N_9644);
or U10519 (N_10519,N_9368,N_9751);
nor U10520 (N_10520,N_9923,N_9397);
xnor U10521 (N_10521,N_9962,N_9585);
nor U10522 (N_10522,N_9554,N_9898);
or U10523 (N_10523,N_9283,N_9162);
and U10524 (N_10524,N_9684,N_9106);
nand U10525 (N_10525,N_9999,N_9996);
nor U10526 (N_10526,N_9556,N_9987);
or U10527 (N_10527,N_9099,N_9011);
nand U10528 (N_10528,N_9152,N_9376);
and U10529 (N_10529,N_9407,N_9265);
xnor U10530 (N_10530,N_9714,N_9855);
and U10531 (N_10531,N_9804,N_9944);
or U10532 (N_10532,N_9016,N_9267);
nand U10533 (N_10533,N_9938,N_9833);
or U10534 (N_10534,N_9201,N_9964);
or U10535 (N_10535,N_9738,N_9458);
or U10536 (N_10536,N_9865,N_9425);
or U10537 (N_10537,N_9405,N_9921);
or U10538 (N_10538,N_9516,N_9185);
nand U10539 (N_10539,N_9301,N_9018);
and U10540 (N_10540,N_9997,N_9186);
nor U10541 (N_10541,N_9558,N_9539);
or U10542 (N_10542,N_9241,N_9585);
and U10543 (N_10543,N_9946,N_9916);
and U10544 (N_10544,N_9107,N_9717);
nand U10545 (N_10545,N_9609,N_9490);
nor U10546 (N_10546,N_9239,N_9199);
or U10547 (N_10547,N_9640,N_9785);
nand U10548 (N_10548,N_9061,N_9769);
xnor U10549 (N_10549,N_9935,N_9899);
nor U10550 (N_10550,N_9962,N_9657);
or U10551 (N_10551,N_9792,N_9806);
or U10552 (N_10552,N_9199,N_9638);
nor U10553 (N_10553,N_9496,N_9482);
nor U10554 (N_10554,N_9156,N_9019);
nand U10555 (N_10555,N_9450,N_9069);
xor U10556 (N_10556,N_9282,N_9562);
xnor U10557 (N_10557,N_9504,N_9310);
or U10558 (N_10558,N_9010,N_9396);
or U10559 (N_10559,N_9074,N_9740);
or U10560 (N_10560,N_9836,N_9561);
nand U10561 (N_10561,N_9959,N_9350);
xor U10562 (N_10562,N_9254,N_9221);
or U10563 (N_10563,N_9626,N_9822);
or U10564 (N_10564,N_9172,N_9371);
nand U10565 (N_10565,N_9044,N_9504);
nand U10566 (N_10566,N_9821,N_9214);
nand U10567 (N_10567,N_9175,N_9977);
nor U10568 (N_10568,N_9029,N_9161);
xor U10569 (N_10569,N_9185,N_9910);
and U10570 (N_10570,N_9457,N_9570);
or U10571 (N_10571,N_9471,N_9672);
or U10572 (N_10572,N_9491,N_9494);
and U10573 (N_10573,N_9951,N_9591);
nor U10574 (N_10574,N_9649,N_9089);
and U10575 (N_10575,N_9810,N_9600);
or U10576 (N_10576,N_9424,N_9130);
nor U10577 (N_10577,N_9740,N_9082);
nand U10578 (N_10578,N_9785,N_9484);
nor U10579 (N_10579,N_9245,N_9968);
and U10580 (N_10580,N_9598,N_9348);
or U10581 (N_10581,N_9008,N_9578);
or U10582 (N_10582,N_9679,N_9971);
nor U10583 (N_10583,N_9426,N_9136);
nand U10584 (N_10584,N_9957,N_9161);
xnor U10585 (N_10585,N_9046,N_9108);
nand U10586 (N_10586,N_9169,N_9898);
or U10587 (N_10587,N_9301,N_9556);
or U10588 (N_10588,N_9652,N_9979);
nand U10589 (N_10589,N_9099,N_9098);
nand U10590 (N_10590,N_9186,N_9956);
and U10591 (N_10591,N_9250,N_9485);
and U10592 (N_10592,N_9038,N_9486);
xnor U10593 (N_10593,N_9924,N_9680);
or U10594 (N_10594,N_9464,N_9558);
nor U10595 (N_10595,N_9755,N_9513);
nor U10596 (N_10596,N_9920,N_9312);
nor U10597 (N_10597,N_9042,N_9643);
xor U10598 (N_10598,N_9269,N_9211);
nor U10599 (N_10599,N_9207,N_9173);
nor U10600 (N_10600,N_9348,N_9467);
and U10601 (N_10601,N_9337,N_9708);
nand U10602 (N_10602,N_9478,N_9215);
xor U10603 (N_10603,N_9931,N_9912);
xor U10604 (N_10604,N_9372,N_9903);
xnor U10605 (N_10605,N_9814,N_9481);
nor U10606 (N_10606,N_9130,N_9505);
nand U10607 (N_10607,N_9205,N_9322);
nand U10608 (N_10608,N_9971,N_9160);
or U10609 (N_10609,N_9243,N_9299);
nand U10610 (N_10610,N_9222,N_9105);
and U10611 (N_10611,N_9956,N_9258);
nand U10612 (N_10612,N_9031,N_9936);
or U10613 (N_10613,N_9177,N_9198);
nor U10614 (N_10614,N_9064,N_9111);
and U10615 (N_10615,N_9696,N_9477);
or U10616 (N_10616,N_9777,N_9575);
or U10617 (N_10617,N_9010,N_9736);
or U10618 (N_10618,N_9401,N_9283);
and U10619 (N_10619,N_9953,N_9565);
and U10620 (N_10620,N_9630,N_9676);
nand U10621 (N_10621,N_9418,N_9326);
nor U10622 (N_10622,N_9319,N_9096);
or U10623 (N_10623,N_9546,N_9007);
or U10624 (N_10624,N_9860,N_9933);
nor U10625 (N_10625,N_9064,N_9950);
nand U10626 (N_10626,N_9572,N_9391);
nand U10627 (N_10627,N_9381,N_9868);
nand U10628 (N_10628,N_9010,N_9288);
or U10629 (N_10629,N_9500,N_9481);
nor U10630 (N_10630,N_9955,N_9891);
nor U10631 (N_10631,N_9027,N_9685);
nand U10632 (N_10632,N_9577,N_9174);
nor U10633 (N_10633,N_9079,N_9787);
or U10634 (N_10634,N_9528,N_9886);
nor U10635 (N_10635,N_9785,N_9869);
nor U10636 (N_10636,N_9654,N_9028);
and U10637 (N_10637,N_9096,N_9675);
nor U10638 (N_10638,N_9576,N_9789);
and U10639 (N_10639,N_9248,N_9540);
nand U10640 (N_10640,N_9336,N_9379);
or U10641 (N_10641,N_9073,N_9454);
nand U10642 (N_10642,N_9932,N_9584);
nand U10643 (N_10643,N_9399,N_9232);
xnor U10644 (N_10644,N_9110,N_9118);
nor U10645 (N_10645,N_9460,N_9926);
nand U10646 (N_10646,N_9758,N_9613);
and U10647 (N_10647,N_9517,N_9809);
and U10648 (N_10648,N_9983,N_9965);
xor U10649 (N_10649,N_9419,N_9305);
and U10650 (N_10650,N_9098,N_9113);
nor U10651 (N_10651,N_9104,N_9924);
and U10652 (N_10652,N_9185,N_9630);
nor U10653 (N_10653,N_9109,N_9352);
xnor U10654 (N_10654,N_9047,N_9920);
or U10655 (N_10655,N_9147,N_9217);
nor U10656 (N_10656,N_9760,N_9924);
xnor U10657 (N_10657,N_9341,N_9920);
or U10658 (N_10658,N_9828,N_9935);
nand U10659 (N_10659,N_9071,N_9927);
nand U10660 (N_10660,N_9003,N_9901);
xor U10661 (N_10661,N_9518,N_9502);
and U10662 (N_10662,N_9660,N_9539);
and U10663 (N_10663,N_9197,N_9726);
or U10664 (N_10664,N_9340,N_9892);
nand U10665 (N_10665,N_9612,N_9320);
and U10666 (N_10666,N_9794,N_9052);
nor U10667 (N_10667,N_9000,N_9171);
nand U10668 (N_10668,N_9624,N_9437);
or U10669 (N_10669,N_9236,N_9910);
and U10670 (N_10670,N_9355,N_9891);
and U10671 (N_10671,N_9017,N_9553);
nor U10672 (N_10672,N_9997,N_9521);
and U10673 (N_10673,N_9225,N_9073);
nand U10674 (N_10674,N_9369,N_9505);
xnor U10675 (N_10675,N_9644,N_9761);
and U10676 (N_10676,N_9361,N_9753);
nand U10677 (N_10677,N_9200,N_9632);
nand U10678 (N_10678,N_9815,N_9814);
nor U10679 (N_10679,N_9767,N_9558);
nand U10680 (N_10680,N_9901,N_9636);
nand U10681 (N_10681,N_9032,N_9146);
nor U10682 (N_10682,N_9707,N_9333);
nor U10683 (N_10683,N_9024,N_9002);
nor U10684 (N_10684,N_9759,N_9144);
or U10685 (N_10685,N_9676,N_9437);
nor U10686 (N_10686,N_9861,N_9321);
or U10687 (N_10687,N_9751,N_9383);
nor U10688 (N_10688,N_9622,N_9493);
nor U10689 (N_10689,N_9795,N_9473);
nor U10690 (N_10690,N_9928,N_9590);
and U10691 (N_10691,N_9197,N_9940);
nand U10692 (N_10692,N_9956,N_9355);
and U10693 (N_10693,N_9023,N_9745);
nand U10694 (N_10694,N_9497,N_9725);
nand U10695 (N_10695,N_9159,N_9848);
or U10696 (N_10696,N_9441,N_9372);
nand U10697 (N_10697,N_9438,N_9902);
nand U10698 (N_10698,N_9239,N_9302);
or U10699 (N_10699,N_9345,N_9145);
and U10700 (N_10700,N_9076,N_9623);
nand U10701 (N_10701,N_9644,N_9193);
nor U10702 (N_10702,N_9526,N_9252);
and U10703 (N_10703,N_9081,N_9278);
or U10704 (N_10704,N_9696,N_9721);
xor U10705 (N_10705,N_9439,N_9490);
nor U10706 (N_10706,N_9623,N_9801);
nand U10707 (N_10707,N_9242,N_9374);
and U10708 (N_10708,N_9247,N_9297);
nor U10709 (N_10709,N_9915,N_9651);
or U10710 (N_10710,N_9577,N_9498);
nor U10711 (N_10711,N_9101,N_9145);
nand U10712 (N_10712,N_9741,N_9075);
nor U10713 (N_10713,N_9691,N_9616);
nor U10714 (N_10714,N_9278,N_9142);
nor U10715 (N_10715,N_9246,N_9041);
nand U10716 (N_10716,N_9398,N_9184);
nor U10717 (N_10717,N_9881,N_9567);
nor U10718 (N_10718,N_9711,N_9160);
nor U10719 (N_10719,N_9941,N_9900);
nor U10720 (N_10720,N_9202,N_9077);
xor U10721 (N_10721,N_9138,N_9886);
or U10722 (N_10722,N_9556,N_9350);
xor U10723 (N_10723,N_9818,N_9763);
nand U10724 (N_10724,N_9217,N_9173);
nand U10725 (N_10725,N_9649,N_9094);
or U10726 (N_10726,N_9974,N_9188);
or U10727 (N_10727,N_9692,N_9939);
nand U10728 (N_10728,N_9330,N_9101);
or U10729 (N_10729,N_9666,N_9721);
nor U10730 (N_10730,N_9027,N_9626);
nor U10731 (N_10731,N_9347,N_9815);
nand U10732 (N_10732,N_9897,N_9896);
and U10733 (N_10733,N_9211,N_9120);
and U10734 (N_10734,N_9396,N_9060);
or U10735 (N_10735,N_9735,N_9079);
xnor U10736 (N_10736,N_9239,N_9093);
nand U10737 (N_10737,N_9398,N_9939);
nor U10738 (N_10738,N_9643,N_9579);
and U10739 (N_10739,N_9509,N_9718);
or U10740 (N_10740,N_9682,N_9862);
nor U10741 (N_10741,N_9278,N_9862);
xor U10742 (N_10742,N_9623,N_9259);
or U10743 (N_10743,N_9957,N_9612);
nand U10744 (N_10744,N_9830,N_9564);
nand U10745 (N_10745,N_9715,N_9337);
nand U10746 (N_10746,N_9309,N_9176);
or U10747 (N_10747,N_9995,N_9504);
nand U10748 (N_10748,N_9385,N_9729);
xor U10749 (N_10749,N_9531,N_9920);
nor U10750 (N_10750,N_9972,N_9753);
nor U10751 (N_10751,N_9642,N_9388);
nor U10752 (N_10752,N_9995,N_9077);
nand U10753 (N_10753,N_9946,N_9258);
or U10754 (N_10754,N_9824,N_9164);
or U10755 (N_10755,N_9024,N_9394);
and U10756 (N_10756,N_9505,N_9295);
and U10757 (N_10757,N_9616,N_9621);
nor U10758 (N_10758,N_9506,N_9624);
xor U10759 (N_10759,N_9524,N_9518);
nor U10760 (N_10760,N_9013,N_9833);
nand U10761 (N_10761,N_9710,N_9851);
or U10762 (N_10762,N_9188,N_9407);
or U10763 (N_10763,N_9364,N_9029);
xnor U10764 (N_10764,N_9002,N_9184);
and U10765 (N_10765,N_9359,N_9115);
nand U10766 (N_10766,N_9273,N_9222);
nand U10767 (N_10767,N_9361,N_9060);
or U10768 (N_10768,N_9568,N_9600);
nand U10769 (N_10769,N_9794,N_9121);
nand U10770 (N_10770,N_9566,N_9191);
xnor U10771 (N_10771,N_9005,N_9277);
nand U10772 (N_10772,N_9254,N_9213);
or U10773 (N_10773,N_9875,N_9122);
and U10774 (N_10774,N_9383,N_9924);
nor U10775 (N_10775,N_9728,N_9456);
and U10776 (N_10776,N_9633,N_9448);
nand U10777 (N_10777,N_9448,N_9690);
nor U10778 (N_10778,N_9799,N_9210);
nand U10779 (N_10779,N_9946,N_9441);
xor U10780 (N_10780,N_9752,N_9726);
nand U10781 (N_10781,N_9588,N_9014);
or U10782 (N_10782,N_9669,N_9005);
or U10783 (N_10783,N_9312,N_9416);
and U10784 (N_10784,N_9256,N_9943);
xor U10785 (N_10785,N_9553,N_9434);
or U10786 (N_10786,N_9946,N_9216);
or U10787 (N_10787,N_9828,N_9033);
nand U10788 (N_10788,N_9183,N_9622);
nor U10789 (N_10789,N_9868,N_9941);
nand U10790 (N_10790,N_9766,N_9529);
nor U10791 (N_10791,N_9140,N_9734);
and U10792 (N_10792,N_9103,N_9152);
nand U10793 (N_10793,N_9096,N_9344);
nand U10794 (N_10794,N_9467,N_9426);
nor U10795 (N_10795,N_9288,N_9700);
or U10796 (N_10796,N_9369,N_9701);
nor U10797 (N_10797,N_9254,N_9072);
nor U10798 (N_10798,N_9890,N_9378);
or U10799 (N_10799,N_9002,N_9435);
xor U10800 (N_10800,N_9945,N_9352);
nor U10801 (N_10801,N_9799,N_9123);
or U10802 (N_10802,N_9466,N_9544);
or U10803 (N_10803,N_9145,N_9428);
or U10804 (N_10804,N_9078,N_9079);
or U10805 (N_10805,N_9886,N_9856);
nor U10806 (N_10806,N_9115,N_9287);
xor U10807 (N_10807,N_9200,N_9612);
or U10808 (N_10808,N_9116,N_9561);
nand U10809 (N_10809,N_9950,N_9870);
or U10810 (N_10810,N_9631,N_9334);
nor U10811 (N_10811,N_9773,N_9218);
nor U10812 (N_10812,N_9185,N_9361);
and U10813 (N_10813,N_9616,N_9240);
and U10814 (N_10814,N_9598,N_9788);
nand U10815 (N_10815,N_9910,N_9266);
nand U10816 (N_10816,N_9401,N_9358);
xor U10817 (N_10817,N_9318,N_9192);
nand U10818 (N_10818,N_9166,N_9773);
nor U10819 (N_10819,N_9361,N_9729);
nor U10820 (N_10820,N_9738,N_9639);
or U10821 (N_10821,N_9783,N_9569);
nand U10822 (N_10822,N_9015,N_9322);
nand U10823 (N_10823,N_9919,N_9599);
nor U10824 (N_10824,N_9548,N_9899);
nand U10825 (N_10825,N_9744,N_9387);
and U10826 (N_10826,N_9216,N_9332);
nor U10827 (N_10827,N_9605,N_9815);
nor U10828 (N_10828,N_9921,N_9311);
or U10829 (N_10829,N_9091,N_9401);
or U10830 (N_10830,N_9057,N_9062);
and U10831 (N_10831,N_9318,N_9457);
nor U10832 (N_10832,N_9457,N_9982);
or U10833 (N_10833,N_9561,N_9259);
nand U10834 (N_10834,N_9214,N_9875);
and U10835 (N_10835,N_9504,N_9013);
xnor U10836 (N_10836,N_9423,N_9076);
and U10837 (N_10837,N_9723,N_9725);
nor U10838 (N_10838,N_9778,N_9940);
and U10839 (N_10839,N_9505,N_9169);
xor U10840 (N_10840,N_9193,N_9702);
nor U10841 (N_10841,N_9102,N_9154);
or U10842 (N_10842,N_9598,N_9181);
or U10843 (N_10843,N_9578,N_9303);
nor U10844 (N_10844,N_9243,N_9224);
nand U10845 (N_10845,N_9252,N_9276);
or U10846 (N_10846,N_9496,N_9737);
or U10847 (N_10847,N_9104,N_9670);
nand U10848 (N_10848,N_9378,N_9082);
or U10849 (N_10849,N_9698,N_9780);
nand U10850 (N_10850,N_9173,N_9050);
nor U10851 (N_10851,N_9409,N_9096);
or U10852 (N_10852,N_9512,N_9835);
nor U10853 (N_10853,N_9899,N_9151);
nor U10854 (N_10854,N_9267,N_9817);
or U10855 (N_10855,N_9470,N_9522);
or U10856 (N_10856,N_9109,N_9718);
and U10857 (N_10857,N_9451,N_9006);
and U10858 (N_10858,N_9141,N_9797);
and U10859 (N_10859,N_9673,N_9215);
nand U10860 (N_10860,N_9873,N_9768);
nand U10861 (N_10861,N_9209,N_9588);
nor U10862 (N_10862,N_9652,N_9944);
xnor U10863 (N_10863,N_9182,N_9077);
nand U10864 (N_10864,N_9109,N_9298);
and U10865 (N_10865,N_9317,N_9738);
xnor U10866 (N_10866,N_9740,N_9474);
nand U10867 (N_10867,N_9797,N_9156);
nand U10868 (N_10868,N_9849,N_9226);
and U10869 (N_10869,N_9724,N_9303);
nand U10870 (N_10870,N_9034,N_9956);
nor U10871 (N_10871,N_9769,N_9328);
and U10872 (N_10872,N_9208,N_9073);
nor U10873 (N_10873,N_9582,N_9665);
nor U10874 (N_10874,N_9778,N_9896);
nor U10875 (N_10875,N_9359,N_9168);
nand U10876 (N_10876,N_9635,N_9466);
or U10877 (N_10877,N_9250,N_9409);
nor U10878 (N_10878,N_9556,N_9057);
nor U10879 (N_10879,N_9435,N_9362);
nor U10880 (N_10880,N_9563,N_9369);
nand U10881 (N_10881,N_9279,N_9754);
or U10882 (N_10882,N_9144,N_9639);
nand U10883 (N_10883,N_9401,N_9862);
nor U10884 (N_10884,N_9564,N_9689);
nand U10885 (N_10885,N_9389,N_9959);
nor U10886 (N_10886,N_9281,N_9665);
nor U10887 (N_10887,N_9223,N_9373);
or U10888 (N_10888,N_9517,N_9400);
nand U10889 (N_10889,N_9702,N_9123);
nand U10890 (N_10890,N_9294,N_9169);
or U10891 (N_10891,N_9459,N_9324);
and U10892 (N_10892,N_9704,N_9573);
nand U10893 (N_10893,N_9446,N_9741);
nand U10894 (N_10894,N_9531,N_9998);
nand U10895 (N_10895,N_9336,N_9056);
nand U10896 (N_10896,N_9256,N_9176);
or U10897 (N_10897,N_9947,N_9918);
or U10898 (N_10898,N_9286,N_9277);
nor U10899 (N_10899,N_9415,N_9961);
nor U10900 (N_10900,N_9230,N_9110);
and U10901 (N_10901,N_9185,N_9625);
nor U10902 (N_10902,N_9781,N_9082);
xor U10903 (N_10903,N_9829,N_9836);
or U10904 (N_10904,N_9561,N_9035);
or U10905 (N_10905,N_9001,N_9625);
nor U10906 (N_10906,N_9119,N_9817);
nand U10907 (N_10907,N_9882,N_9405);
or U10908 (N_10908,N_9745,N_9132);
nor U10909 (N_10909,N_9753,N_9279);
nand U10910 (N_10910,N_9832,N_9755);
or U10911 (N_10911,N_9395,N_9054);
and U10912 (N_10912,N_9075,N_9679);
nand U10913 (N_10913,N_9007,N_9315);
xor U10914 (N_10914,N_9087,N_9585);
nor U10915 (N_10915,N_9078,N_9061);
or U10916 (N_10916,N_9129,N_9031);
nand U10917 (N_10917,N_9587,N_9193);
or U10918 (N_10918,N_9925,N_9228);
or U10919 (N_10919,N_9199,N_9231);
xnor U10920 (N_10920,N_9176,N_9367);
nand U10921 (N_10921,N_9896,N_9101);
nor U10922 (N_10922,N_9085,N_9881);
nand U10923 (N_10923,N_9047,N_9243);
or U10924 (N_10924,N_9042,N_9221);
and U10925 (N_10925,N_9553,N_9147);
and U10926 (N_10926,N_9471,N_9321);
or U10927 (N_10927,N_9193,N_9748);
nor U10928 (N_10928,N_9785,N_9976);
and U10929 (N_10929,N_9829,N_9146);
nor U10930 (N_10930,N_9372,N_9817);
and U10931 (N_10931,N_9987,N_9579);
and U10932 (N_10932,N_9734,N_9135);
and U10933 (N_10933,N_9866,N_9669);
and U10934 (N_10934,N_9406,N_9124);
nor U10935 (N_10935,N_9412,N_9509);
and U10936 (N_10936,N_9430,N_9728);
and U10937 (N_10937,N_9277,N_9981);
nor U10938 (N_10938,N_9959,N_9504);
nand U10939 (N_10939,N_9450,N_9737);
and U10940 (N_10940,N_9320,N_9496);
and U10941 (N_10941,N_9928,N_9187);
nor U10942 (N_10942,N_9143,N_9687);
nor U10943 (N_10943,N_9028,N_9027);
nand U10944 (N_10944,N_9213,N_9175);
or U10945 (N_10945,N_9990,N_9896);
nor U10946 (N_10946,N_9886,N_9255);
and U10947 (N_10947,N_9621,N_9808);
nand U10948 (N_10948,N_9737,N_9700);
or U10949 (N_10949,N_9170,N_9212);
nand U10950 (N_10950,N_9823,N_9715);
nand U10951 (N_10951,N_9182,N_9979);
nand U10952 (N_10952,N_9253,N_9352);
nand U10953 (N_10953,N_9786,N_9062);
nand U10954 (N_10954,N_9404,N_9544);
and U10955 (N_10955,N_9777,N_9731);
nand U10956 (N_10956,N_9948,N_9902);
and U10957 (N_10957,N_9299,N_9466);
nor U10958 (N_10958,N_9117,N_9383);
or U10959 (N_10959,N_9212,N_9235);
nand U10960 (N_10960,N_9767,N_9138);
and U10961 (N_10961,N_9412,N_9218);
xor U10962 (N_10962,N_9188,N_9760);
and U10963 (N_10963,N_9947,N_9562);
and U10964 (N_10964,N_9621,N_9594);
nor U10965 (N_10965,N_9736,N_9785);
nor U10966 (N_10966,N_9055,N_9211);
or U10967 (N_10967,N_9714,N_9059);
and U10968 (N_10968,N_9535,N_9127);
nor U10969 (N_10969,N_9754,N_9959);
xnor U10970 (N_10970,N_9898,N_9788);
nor U10971 (N_10971,N_9375,N_9326);
or U10972 (N_10972,N_9921,N_9039);
nand U10973 (N_10973,N_9687,N_9002);
and U10974 (N_10974,N_9264,N_9675);
or U10975 (N_10975,N_9375,N_9487);
nand U10976 (N_10976,N_9402,N_9347);
and U10977 (N_10977,N_9488,N_9886);
nand U10978 (N_10978,N_9690,N_9106);
nor U10979 (N_10979,N_9987,N_9044);
or U10980 (N_10980,N_9728,N_9450);
xnor U10981 (N_10981,N_9685,N_9477);
nand U10982 (N_10982,N_9113,N_9600);
nor U10983 (N_10983,N_9851,N_9866);
nor U10984 (N_10984,N_9785,N_9255);
or U10985 (N_10985,N_9968,N_9674);
nor U10986 (N_10986,N_9165,N_9761);
nor U10987 (N_10987,N_9794,N_9792);
or U10988 (N_10988,N_9536,N_9483);
nand U10989 (N_10989,N_9999,N_9536);
or U10990 (N_10990,N_9917,N_9654);
and U10991 (N_10991,N_9933,N_9971);
nand U10992 (N_10992,N_9133,N_9136);
nor U10993 (N_10993,N_9284,N_9473);
nor U10994 (N_10994,N_9145,N_9508);
xnor U10995 (N_10995,N_9478,N_9209);
nand U10996 (N_10996,N_9172,N_9605);
or U10997 (N_10997,N_9020,N_9759);
nand U10998 (N_10998,N_9836,N_9843);
or U10999 (N_10999,N_9805,N_9137);
xor U11000 (N_11000,N_10320,N_10304);
or U11001 (N_11001,N_10290,N_10129);
and U11002 (N_11002,N_10429,N_10526);
nand U11003 (N_11003,N_10525,N_10686);
or U11004 (N_11004,N_10330,N_10203);
nor U11005 (N_11005,N_10744,N_10997);
xor U11006 (N_11006,N_10133,N_10113);
xor U11007 (N_11007,N_10472,N_10705);
nand U11008 (N_11008,N_10976,N_10549);
nand U11009 (N_11009,N_10636,N_10794);
nor U11010 (N_11010,N_10460,N_10223);
and U11011 (N_11011,N_10539,N_10079);
nor U11012 (N_11012,N_10088,N_10229);
nor U11013 (N_11013,N_10697,N_10781);
nor U11014 (N_11014,N_10598,N_10842);
or U11015 (N_11015,N_10166,N_10798);
xor U11016 (N_11016,N_10625,N_10639);
nor U11017 (N_11017,N_10482,N_10207);
or U11018 (N_11018,N_10974,N_10851);
nor U11019 (N_11019,N_10544,N_10873);
nor U11020 (N_11020,N_10312,N_10628);
or U11021 (N_11021,N_10154,N_10260);
xnor U11022 (N_11022,N_10713,N_10247);
or U11023 (N_11023,N_10978,N_10144);
nor U11024 (N_11024,N_10097,N_10339);
nor U11025 (N_11025,N_10618,N_10131);
and U11026 (N_11026,N_10022,N_10655);
or U11027 (N_11027,N_10008,N_10871);
and U11028 (N_11028,N_10437,N_10680);
nand U11029 (N_11029,N_10013,N_10522);
nor U11030 (N_11030,N_10666,N_10099);
or U11031 (N_11031,N_10523,N_10483);
and U11032 (N_11032,N_10742,N_10753);
nand U11033 (N_11033,N_10117,N_10867);
nor U11034 (N_11034,N_10956,N_10622);
or U11035 (N_11035,N_10623,N_10121);
and U11036 (N_11036,N_10371,N_10361);
and U11037 (N_11037,N_10733,N_10961);
and U11038 (N_11038,N_10863,N_10775);
nor U11039 (N_11039,N_10137,N_10127);
and U11040 (N_11040,N_10769,N_10704);
and U11041 (N_11041,N_10413,N_10949);
or U11042 (N_11042,N_10856,N_10679);
and U11043 (N_11043,N_10737,N_10998);
nand U11044 (N_11044,N_10224,N_10888);
or U11045 (N_11045,N_10760,N_10476);
and U11046 (N_11046,N_10126,N_10003);
nand U11047 (N_11047,N_10102,N_10311);
xnor U11048 (N_11048,N_10046,N_10351);
or U11049 (N_11049,N_10726,N_10086);
and U11050 (N_11050,N_10272,N_10870);
or U11051 (N_11051,N_10411,N_10477);
xor U11052 (N_11052,N_10327,N_10261);
and U11053 (N_11053,N_10254,N_10595);
or U11054 (N_11054,N_10575,N_10735);
or U11055 (N_11055,N_10635,N_10907);
or U11056 (N_11056,N_10891,N_10903);
and U11057 (N_11057,N_10354,N_10196);
nor U11058 (N_11058,N_10555,N_10514);
or U11059 (N_11059,N_10853,N_10823);
and U11060 (N_11060,N_10346,N_10227);
nand U11061 (N_11061,N_10170,N_10093);
xnor U11062 (N_11062,N_10999,N_10931);
nor U11063 (N_11063,N_10080,N_10119);
or U11064 (N_11064,N_10717,N_10112);
nor U11065 (N_11065,N_10558,N_10064);
or U11066 (N_11066,N_10110,N_10085);
or U11067 (N_11067,N_10634,N_10955);
nor U11068 (N_11068,N_10410,N_10861);
or U11069 (N_11069,N_10389,N_10285);
nor U11070 (N_11070,N_10100,N_10538);
nand U11071 (N_11071,N_10052,N_10958);
nor U11072 (N_11072,N_10583,N_10859);
nand U11073 (N_11073,N_10845,N_10837);
and U11074 (N_11074,N_10439,N_10681);
nor U11075 (N_11075,N_10528,N_10259);
and U11076 (N_11076,N_10458,N_10417);
nand U11077 (N_11077,N_10731,N_10778);
nor U11078 (N_11078,N_10214,N_10569);
or U11079 (N_11079,N_10282,N_10128);
xnor U11080 (N_11080,N_10901,N_10266);
or U11081 (N_11081,N_10248,N_10554);
xnor U11082 (N_11082,N_10606,N_10225);
nand U11083 (N_11083,N_10492,N_10445);
xnor U11084 (N_11084,N_10846,N_10768);
xor U11085 (N_11085,N_10373,N_10649);
xnor U11086 (N_11086,N_10572,N_10299);
nand U11087 (N_11087,N_10637,N_10919);
and U11088 (N_11088,N_10217,N_10834);
nand U11089 (N_11089,N_10688,N_10155);
and U11090 (N_11090,N_10141,N_10825);
and U11091 (N_11091,N_10589,N_10084);
nand U11092 (N_11092,N_10167,N_10762);
nor U11093 (N_11093,N_10576,N_10720);
xor U11094 (N_11094,N_10940,N_10292);
nand U11095 (N_11095,N_10358,N_10750);
or U11096 (N_11096,N_10537,N_10216);
and U11097 (N_11097,N_10935,N_10199);
xor U11098 (N_11098,N_10519,N_10190);
xnor U11099 (N_11099,N_10468,N_10685);
and U11100 (N_11100,N_10215,N_10741);
and U11101 (N_11101,N_10049,N_10255);
nand U11102 (N_11102,N_10467,N_10075);
nor U11103 (N_11103,N_10048,N_10890);
nand U11104 (N_11104,N_10847,N_10063);
or U11105 (N_11105,N_10341,N_10964);
nand U11106 (N_11106,N_10026,N_10153);
nand U11107 (N_11107,N_10811,N_10699);
nor U11108 (N_11108,N_10213,N_10306);
and U11109 (N_11109,N_10944,N_10758);
and U11110 (N_11110,N_10568,N_10719);
xnor U11111 (N_11111,N_10060,N_10721);
or U11112 (N_11112,N_10140,N_10151);
nand U11113 (N_11113,N_10953,N_10201);
nor U11114 (N_11114,N_10548,N_10258);
and U11115 (N_11115,N_10738,N_10420);
and U11116 (N_11116,N_10451,N_10197);
and U11117 (N_11117,N_10596,N_10160);
or U11118 (N_11118,N_10789,N_10473);
and U11119 (N_11119,N_10743,N_10995);
nand U11120 (N_11120,N_10210,N_10072);
or U11121 (N_11121,N_10546,N_10783);
nand U11122 (N_11122,N_10303,N_10186);
nand U11123 (N_11123,N_10673,N_10883);
nand U11124 (N_11124,N_10340,N_10096);
nand U11125 (N_11125,N_10545,N_10319);
xnor U11126 (N_11126,N_10456,N_10307);
or U11127 (N_11127,N_10313,N_10323);
and U11128 (N_11128,N_10943,N_10150);
and U11129 (N_11129,N_10442,N_10403);
xnor U11130 (N_11130,N_10560,N_10984);
nor U11131 (N_11131,N_10565,N_10332);
or U11132 (N_11132,N_10050,N_10130);
and U11133 (N_11133,N_10386,N_10629);
and U11134 (N_11134,N_10378,N_10700);
nand U11135 (N_11135,N_10408,N_10108);
nand U11136 (N_11136,N_10503,N_10138);
nand U11137 (N_11137,N_10593,N_10054);
and U11138 (N_11138,N_10232,N_10550);
and U11139 (N_11139,N_10993,N_10181);
and U11140 (N_11140,N_10136,N_10563);
or U11141 (N_11141,N_10684,N_10109);
and U11142 (N_11142,N_10933,N_10579);
nand U11143 (N_11143,N_10626,N_10763);
nand U11144 (N_11144,N_10582,N_10275);
or U11145 (N_11145,N_10941,N_10019);
and U11146 (N_11146,N_10776,N_10643);
and U11147 (N_11147,N_10391,N_10469);
or U11148 (N_11148,N_10092,N_10271);
nor U11149 (N_11149,N_10376,N_10338);
or U11150 (N_11150,N_10671,N_10114);
nand U11151 (N_11151,N_10496,N_10372);
nor U11152 (N_11152,N_10965,N_10158);
nand U11153 (N_11153,N_10401,N_10954);
and U11154 (N_11154,N_10132,N_10461);
or U11155 (N_11155,N_10250,N_10145);
xnor U11156 (N_11156,N_10914,N_10693);
nand U11157 (N_11157,N_10913,N_10447);
nor U11158 (N_11158,N_10043,N_10218);
nand U11159 (N_11159,N_10270,N_10818);
nand U11160 (N_11160,N_10345,N_10074);
nand U11161 (N_11161,N_10318,N_10297);
or U11162 (N_11162,N_10650,N_10240);
nand U11163 (N_11163,N_10848,N_10055);
nand U11164 (N_11164,N_10288,N_10773);
nand U11165 (N_11165,N_10016,N_10077);
nor U11166 (N_11166,N_10355,N_10424);
nor U11167 (N_11167,N_10360,N_10957);
nor U11168 (N_11168,N_10910,N_10497);
nor U11169 (N_11169,N_10499,N_10594);
xnor U11170 (N_11170,N_10703,N_10148);
nand U11171 (N_11171,N_10716,N_10877);
or U11172 (N_11172,N_10193,N_10101);
nand U11173 (N_11173,N_10381,N_10187);
nor U11174 (N_11174,N_10142,N_10992);
and U11175 (N_11175,N_10784,N_10939);
nor U11176 (N_11176,N_10233,N_10106);
and U11177 (N_11177,N_10159,N_10176);
nand U11178 (N_11178,N_10172,N_10464);
nand U11179 (N_11179,N_10161,N_10070);
xor U11180 (N_11180,N_10895,N_10751);
nand U11181 (N_11181,N_10543,N_10805);
xor U11182 (N_11182,N_10308,N_10926);
nand U11183 (N_11183,N_10342,N_10486);
xnor U11184 (N_11184,N_10745,N_10921);
nor U11185 (N_11185,N_10397,N_10676);
xor U11186 (N_11186,N_10588,N_10804);
or U11187 (N_11187,N_10843,N_10529);
or U11188 (N_11188,N_10951,N_10146);
and U11189 (N_11189,N_10431,N_10103);
or U11190 (N_11190,N_10032,N_10959);
and U11191 (N_11191,N_10475,N_10209);
or U11192 (N_11192,N_10506,N_10868);
nand U11193 (N_11193,N_10395,N_10310);
and U11194 (N_11194,N_10819,N_10239);
nor U11195 (N_11195,N_10337,N_10645);
nand U11196 (N_11196,N_10015,N_10485);
nor U11197 (N_11197,N_10936,N_10017);
or U11198 (N_11198,N_10348,N_10164);
nand U11199 (N_11199,N_10566,N_10143);
and U11200 (N_11200,N_10231,N_10552);
and U11201 (N_11201,N_10149,N_10041);
and U11202 (N_11202,N_10922,N_10257);
and U11203 (N_11203,N_10090,N_10918);
nand U11204 (N_11204,N_10899,N_10898);
and U11205 (N_11205,N_10585,N_10988);
and U11206 (N_11206,N_10644,N_10010);
or U11207 (N_11207,N_10392,N_10840);
and U11208 (N_11208,N_10038,N_10707);
and U11209 (N_11209,N_10387,N_10967);
nand U11210 (N_11210,N_10968,N_10996);
nor U11211 (N_11211,N_10865,N_10706);
and U11212 (N_11212,N_10991,N_10236);
nand U11213 (N_11213,N_10178,N_10157);
nand U11214 (N_11214,N_10527,N_10604);
and U11215 (N_11215,N_10581,N_10449);
nor U11216 (N_11216,N_10897,N_10094);
nor U11217 (N_11217,N_10450,N_10578);
and U11218 (N_11218,N_10284,N_10564);
or U11219 (N_11219,N_10530,N_10653);
nand U11220 (N_11220,N_10709,N_10889);
xnor U11221 (N_11221,N_10324,N_10396);
and U11222 (N_11222,N_10535,N_10540);
nand U11223 (N_11223,N_10872,N_10690);
or U11224 (N_11224,N_10368,N_10524);
xor U11225 (N_11225,N_10321,N_10180);
nand U11226 (N_11226,N_10630,N_10884);
nand U11227 (N_11227,N_10394,N_10416);
nand U11228 (N_11228,N_10816,N_10452);
nor U11229 (N_11229,N_10034,N_10983);
and U11230 (N_11230,N_10711,N_10390);
nand U11231 (N_11231,N_10068,N_10826);
and U11232 (N_11232,N_10646,N_10894);
nand U11233 (N_11233,N_10256,N_10296);
nand U11234 (N_11234,N_10876,N_10274);
nor U11235 (N_11235,N_10230,N_10802);
nand U11236 (N_11236,N_10702,N_10852);
nand U11237 (N_11237,N_10613,N_10577);
or U11238 (N_11238,N_10814,N_10370);
nand U11239 (N_11239,N_10491,N_10438);
nand U11240 (N_11240,N_10832,N_10300);
or U11241 (N_11241,N_10426,N_10208);
and U11242 (N_11242,N_10498,N_10007);
and U11243 (N_11243,N_10466,N_10617);
nor U11244 (N_11244,N_10163,N_10156);
nand U11245 (N_11245,N_10262,N_10675);
xor U11246 (N_11246,N_10356,N_10031);
xnor U11247 (N_11247,N_10878,N_10810);
nor U11248 (N_11248,N_10651,N_10632);
nor U11249 (N_11249,N_10200,N_10624);
nor U11250 (N_11250,N_10631,N_10509);
nand U11251 (N_11251,N_10279,N_10844);
nand U11252 (N_11252,N_10906,N_10045);
nand U11253 (N_11253,N_10985,N_10694);
nor U11254 (N_11254,N_10202,N_10795);
nand U11255 (N_11255,N_10267,N_10542);
or U11256 (N_11256,N_10642,N_10835);
nand U11257 (N_11257,N_10620,N_10018);
nand U11258 (N_11258,N_10375,N_10807);
nand U11259 (N_11259,N_10947,N_10615);
nand U11260 (N_11260,N_10404,N_10611);
nor U11261 (N_11261,N_10994,N_10069);
nand U11262 (N_11262,N_10436,N_10035);
and U11263 (N_11263,N_10571,N_10302);
and U11264 (N_11264,N_10065,N_10756);
nor U11265 (N_11265,N_10665,N_10518);
xnor U11266 (N_11266,N_10195,N_10505);
xor U11267 (N_11267,N_10353,N_10402);
nor U11268 (N_11268,N_10421,N_10977);
nor U11269 (N_11269,N_10425,N_10463);
xor U11270 (N_11270,N_10772,N_10674);
and U11271 (N_11271,N_10603,N_10547);
xnor U11272 (N_11272,N_10656,N_10759);
or U11273 (N_11273,N_10771,N_10030);
nor U11274 (N_11274,N_10559,N_10281);
nand U11275 (N_11275,N_10470,N_10095);
or U11276 (N_11276,N_10882,N_10111);
or U11277 (N_11277,N_10291,N_10335);
nor U11278 (N_11278,N_10029,N_10407);
xnor U11279 (N_11279,N_10553,N_10886);
nor U11280 (N_11280,N_10504,N_10365);
xor U11281 (N_11281,N_10171,N_10067);
or U11282 (N_11282,N_10076,N_10183);
nor U11283 (N_11283,N_10139,N_10607);
or U11284 (N_11284,N_10244,N_10124);
nand U11285 (N_11285,N_10206,N_10599);
nand U11286 (N_11286,N_10715,N_10602);
or U11287 (N_11287,N_10083,N_10732);
and U11288 (N_11288,N_10147,N_10708);
nand U11289 (N_11289,N_10293,N_10587);
nor U11290 (N_11290,N_10057,N_10557);
or U11291 (N_11291,N_10520,N_10409);
or U11292 (N_11292,N_10989,N_10115);
and U11293 (N_11293,N_10765,N_10692);
nor U11294 (N_11294,N_10739,N_10892);
or U11295 (N_11295,N_10945,N_10608);
nor U11296 (N_11296,N_10930,N_10808);
or U11297 (N_11297,N_10226,N_10462);
nand U11298 (N_11298,N_10276,N_10317);
nand U11299 (N_11299,N_10659,N_10830);
xor U11300 (N_11300,N_10382,N_10162);
and U11301 (N_11301,N_10415,N_10836);
nand U11302 (N_11302,N_10986,N_10736);
or U11303 (N_11303,N_10273,N_10289);
nand U11304 (N_11304,N_10383,N_10480);
and U11305 (N_11305,N_10435,N_10934);
or U11306 (N_11306,N_10073,N_10800);
and U11307 (N_11307,N_10803,N_10268);
xor U11308 (N_11308,N_10712,N_10508);
and U11309 (N_11309,N_10513,N_10969);
nand U11310 (N_11310,N_10591,N_10238);
nand U11311 (N_11311,N_10185,N_10047);
nor U11312 (N_11312,N_10219,N_10107);
or U11313 (N_11313,N_10400,N_10328);
and U11314 (N_11314,N_10797,N_10793);
nand U11315 (N_11315,N_10222,N_10748);
and U11316 (N_11316,N_10446,N_10517);
and U11317 (N_11317,N_10089,N_10362);
or U11318 (N_11318,N_10962,N_10740);
xnor U11319 (N_11319,N_10384,N_10600);
and U11320 (N_11320,N_10277,N_10455);
and U11321 (N_11321,N_10044,N_10305);
nor U11322 (N_11322,N_10858,N_10567);
nand U11323 (N_11323,N_10885,N_10001);
nand U11324 (N_11324,N_10761,N_10039);
nand U11325 (N_11325,N_10790,N_10658);
and U11326 (N_11326,N_10388,N_10314);
nand U11327 (N_11327,N_10828,N_10009);
or U11328 (N_11328,N_10824,N_10561);
xnor U11329 (N_11329,N_10799,N_10269);
nor U11330 (N_11330,N_10812,N_10347);
or U11331 (N_11331,N_10125,N_10612);
nor U11332 (N_11332,N_10349,N_10501);
or U11333 (N_11333,N_10942,N_10025);
nor U11334 (N_11334,N_10908,N_10511);
nor U11335 (N_11335,N_10621,N_10746);
or U11336 (N_11336,N_10904,N_10601);
nand U11337 (N_11337,N_10614,N_10718);
nor U11338 (N_11338,N_10874,N_10012);
or U11339 (N_11339,N_10654,N_10813);
nor U11340 (N_11340,N_10662,N_10923);
xor U11341 (N_11341,N_10343,N_10211);
and U11342 (N_11342,N_10573,N_10249);
nor U11343 (N_11343,N_10478,N_10664);
nor U11344 (N_11344,N_10364,N_10489);
and U11345 (N_11345,N_10443,N_10754);
nor U11346 (N_11346,N_10037,N_10605);
nand U11347 (N_11347,N_10459,N_10188);
and U11348 (N_11348,N_10418,N_10963);
nor U11349 (N_11349,N_10900,N_10021);
xor U11350 (N_11350,N_10980,N_10586);
and U11351 (N_11351,N_10875,N_10040);
or U11352 (N_11352,N_10670,N_10329);
and U11353 (N_11353,N_10764,N_10817);
and U11354 (N_11354,N_10309,N_10487);
nand U11355 (N_11355,N_10228,N_10831);
xor U11356 (N_11356,N_10854,N_10058);
nor U11357 (N_11357,N_10787,N_10641);
or U11358 (N_11358,N_10689,N_10087);
and U11359 (N_11359,N_10752,N_10184);
nor U11360 (N_11360,N_10326,N_10253);
xnor U11361 (N_11361,N_10414,N_10280);
nand U11362 (N_11362,N_10952,N_10454);
and U11363 (N_11363,N_10377,N_10647);
nor U11364 (N_11364,N_10234,N_10105);
nor U11365 (N_11365,N_10120,N_10966);
and U11366 (N_11366,N_10152,N_10204);
nor U11367 (N_11367,N_10672,N_10682);
or U11368 (N_11368,N_10465,N_10359);
or U11369 (N_11369,N_10915,N_10194);
nand U11370 (N_11370,N_10880,N_10857);
and U11371 (N_11371,N_10028,N_10433);
or U11372 (N_11372,N_10827,N_10484);
xor U11373 (N_11373,N_10950,N_10011);
and U11374 (N_11374,N_10441,N_10448);
nor U11375 (N_11375,N_10027,N_10325);
xnor U11376 (N_11376,N_10367,N_10168);
nand U11377 (N_11377,N_10352,N_10412);
nand U11378 (N_11378,N_10512,N_10173);
nor U11379 (N_11379,N_10869,N_10474);
or U11380 (N_11380,N_10283,N_10082);
or U11381 (N_11381,N_10165,N_10488);
nor U11382 (N_11382,N_10023,N_10809);
nand U11383 (N_11383,N_10785,N_10766);
or U11384 (N_11384,N_10979,N_10398);
xnor U11385 (N_11385,N_10061,N_10864);
and U11386 (N_11386,N_10722,N_10695);
nor U11387 (N_11387,N_10322,N_10887);
xnor U11388 (N_11388,N_10104,N_10495);
xor U11389 (N_11389,N_10434,N_10987);
and U11390 (N_11390,N_10521,N_10850);
nor U11391 (N_11391,N_10911,N_10432);
and U11392 (N_11392,N_10902,N_10515);
nor U11393 (N_11393,N_10205,N_10344);
and U11394 (N_11394,N_10749,N_10286);
and U11395 (N_11395,N_10000,N_10696);
nand U11396 (N_11396,N_10453,N_10374);
or U11397 (N_11397,N_10242,N_10879);
nor U11398 (N_11398,N_10905,N_10516);
and U11399 (N_11399,N_10042,N_10938);
xor U11400 (N_11400,N_10551,N_10782);
xor U11401 (N_11401,N_10796,N_10972);
or U11402 (N_11402,N_10971,N_10331);
nand U11403 (N_11403,N_10062,N_10369);
nand U11404 (N_11404,N_10334,N_10687);
and U11405 (N_11405,N_10541,N_10929);
nor U11406 (N_11406,N_10246,N_10815);
or U11407 (N_11407,N_10990,N_10235);
nor U11408 (N_11408,N_10059,N_10592);
nor U11409 (N_11409,N_10301,N_10405);
nand U11410 (N_11410,N_10081,N_10801);
nor U11411 (N_11411,N_10767,N_10728);
or U11412 (N_11412,N_10493,N_10385);
and U11413 (N_11413,N_10893,N_10657);
nand U11414 (N_11414,N_10066,N_10263);
and U11415 (N_11415,N_10507,N_10002);
or U11416 (N_11416,N_10574,N_10982);
nor U11417 (N_11417,N_10652,N_10116);
and U11418 (N_11418,N_10924,N_10531);
nand U11419 (N_11419,N_10755,N_10841);
nand U11420 (N_11420,N_10294,N_10118);
nor U11421 (N_11421,N_10806,N_10532);
nor U11422 (N_11422,N_10562,N_10265);
and U11423 (N_11423,N_10036,N_10287);
or U11424 (N_11424,N_10419,N_10777);
nor U11425 (N_11425,N_10315,N_10502);
nand U11426 (N_11426,N_10710,N_10723);
nor U11427 (N_11427,N_10033,N_10440);
nor U11428 (N_11428,N_10406,N_10701);
and U11429 (N_11429,N_10500,N_10298);
or U11430 (N_11430,N_10379,N_10336);
xnor U11431 (N_11431,N_10660,N_10881);
xnor U11432 (N_11432,N_10698,N_10534);
nand U11433 (N_11433,N_10004,N_10734);
or U11434 (N_11434,N_10177,N_10838);
and U11435 (N_11435,N_10134,N_10981);
and U11436 (N_11436,N_10757,N_10243);
or U11437 (N_11437,N_10932,N_10430);
nand U11438 (N_11438,N_10422,N_10822);
nand U11439 (N_11439,N_10916,N_10198);
xor U11440 (N_11440,N_10536,N_10786);
and U11441 (N_11441,N_10423,N_10174);
nor U11442 (N_11442,N_10091,N_10098);
or U11443 (N_11443,N_10730,N_10829);
xnor U11444 (N_11444,N_10678,N_10024);
and U11445 (N_11445,N_10975,N_10774);
nor U11446 (N_11446,N_10399,N_10237);
nor U11447 (N_11447,N_10191,N_10350);
or U11448 (N_11448,N_10669,N_10727);
nand U11449 (N_11449,N_10490,N_10169);
and U11450 (N_11450,N_10780,N_10252);
nand U11451 (N_11451,N_10724,N_10471);
and U11452 (N_11452,N_10820,N_10444);
xor U11453 (N_11453,N_10648,N_10855);
or U11454 (N_11454,N_10363,N_10071);
nand U11455 (N_11455,N_10122,N_10616);
or U11456 (N_11456,N_10479,N_10220);
and U11457 (N_11457,N_10770,N_10380);
or U11458 (N_11458,N_10182,N_10481);
nor U11459 (N_11459,N_10946,N_10691);
and U11460 (N_11460,N_10917,N_10192);
nand U11461 (N_11461,N_10584,N_10912);
nor U11462 (N_11462,N_10960,N_10006);
nor U11463 (N_11463,N_10970,N_10427);
nand U11464 (N_11464,N_10580,N_10245);
or U11465 (N_11465,N_10627,N_10792);
or U11466 (N_11466,N_10927,N_10920);
nor U11467 (N_11467,N_10357,N_10937);
and U11468 (N_11468,N_10189,N_10973);
and U11469 (N_11469,N_10849,N_10619);
and U11470 (N_11470,N_10866,N_10677);
xnor U11471 (N_11471,N_10725,N_10909);
xnor U11472 (N_11472,N_10925,N_10640);
or U11473 (N_11473,N_10494,N_10510);
nand U11474 (N_11474,N_10779,N_10667);
nor U11475 (N_11475,N_10278,N_10316);
or U11476 (N_11476,N_10221,N_10590);
xnor U11477 (N_11477,N_10791,N_10241);
nor U11478 (N_11478,N_10860,N_10747);
nand U11479 (N_11479,N_10175,N_10663);
nand U11480 (N_11480,N_10661,N_10948);
or U11481 (N_11481,N_10729,N_10428);
or U11482 (N_11482,N_10457,N_10928);
nor U11483 (N_11483,N_10333,N_10862);
nand U11484 (N_11484,N_10633,N_10056);
nor U11485 (N_11485,N_10714,N_10556);
and U11486 (N_11486,N_10020,N_10833);
nor U11487 (N_11487,N_10668,N_10366);
nor U11488 (N_11488,N_10896,N_10264);
nor U11489 (N_11489,N_10788,N_10251);
xnor U11490 (N_11490,N_10123,N_10212);
nor U11491 (N_11491,N_10533,N_10393);
xor U11492 (N_11492,N_10839,N_10014);
nand U11493 (N_11493,N_10597,N_10005);
and U11494 (N_11494,N_10610,N_10638);
or U11495 (N_11495,N_10051,N_10179);
nor U11496 (N_11496,N_10683,N_10078);
or U11497 (N_11497,N_10570,N_10053);
and U11498 (N_11498,N_10135,N_10821);
nor U11499 (N_11499,N_10295,N_10609);
nor U11500 (N_11500,N_10012,N_10214);
or U11501 (N_11501,N_10049,N_10940);
and U11502 (N_11502,N_10468,N_10053);
or U11503 (N_11503,N_10369,N_10882);
nand U11504 (N_11504,N_10420,N_10663);
nand U11505 (N_11505,N_10607,N_10589);
nor U11506 (N_11506,N_10807,N_10011);
or U11507 (N_11507,N_10049,N_10039);
and U11508 (N_11508,N_10475,N_10589);
and U11509 (N_11509,N_10780,N_10118);
nor U11510 (N_11510,N_10899,N_10344);
or U11511 (N_11511,N_10842,N_10515);
and U11512 (N_11512,N_10598,N_10447);
or U11513 (N_11513,N_10754,N_10010);
or U11514 (N_11514,N_10507,N_10483);
nand U11515 (N_11515,N_10300,N_10509);
or U11516 (N_11516,N_10461,N_10366);
and U11517 (N_11517,N_10887,N_10285);
nor U11518 (N_11518,N_10662,N_10948);
xor U11519 (N_11519,N_10752,N_10728);
and U11520 (N_11520,N_10973,N_10491);
and U11521 (N_11521,N_10506,N_10188);
nor U11522 (N_11522,N_10069,N_10752);
nand U11523 (N_11523,N_10003,N_10802);
nor U11524 (N_11524,N_10129,N_10447);
nand U11525 (N_11525,N_10758,N_10028);
and U11526 (N_11526,N_10311,N_10049);
or U11527 (N_11527,N_10418,N_10703);
nor U11528 (N_11528,N_10699,N_10365);
or U11529 (N_11529,N_10799,N_10931);
nor U11530 (N_11530,N_10877,N_10131);
or U11531 (N_11531,N_10060,N_10170);
and U11532 (N_11532,N_10343,N_10650);
nor U11533 (N_11533,N_10508,N_10398);
nor U11534 (N_11534,N_10289,N_10826);
or U11535 (N_11535,N_10308,N_10579);
nand U11536 (N_11536,N_10793,N_10316);
xor U11537 (N_11537,N_10353,N_10654);
nor U11538 (N_11538,N_10099,N_10845);
nor U11539 (N_11539,N_10880,N_10782);
and U11540 (N_11540,N_10814,N_10106);
nor U11541 (N_11541,N_10330,N_10272);
nor U11542 (N_11542,N_10297,N_10748);
or U11543 (N_11543,N_10821,N_10726);
or U11544 (N_11544,N_10726,N_10251);
nand U11545 (N_11545,N_10453,N_10733);
or U11546 (N_11546,N_10523,N_10252);
and U11547 (N_11547,N_10931,N_10600);
nand U11548 (N_11548,N_10760,N_10464);
or U11549 (N_11549,N_10409,N_10710);
and U11550 (N_11550,N_10916,N_10088);
nor U11551 (N_11551,N_10417,N_10573);
or U11552 (N_11552,N_10217,N_10015);
or U11553 (N_11553,N_10844,N_10310);
nand U11554 (N_11554,N_10049,N_10634);
nor U11555 (N_11555,N_10677,N_10589);
or U11556 (N_11556,N_10810,N_10655);
nand U11557 (N_11557,N_10282,N_10678);
nor U11558 (N_11558,N_10888,N_10952);
or U11559 (N_11559,N_10044,N_10420);
nand U11560 (N_11560,N_10082,N_10179);
xor U11561 (N_11561,N_10552,N_10717);
nand U11562 (N_11562,N_10308,N_10804);
and U11563 (N_11563,N_10097,N_10260);
and U11564 (N_11564,N_10004,N_10472);
or U11565 (N_11565,N_10606,N_10999);
or U11566 (N_11566,N_10929,N_10047);
nand U11567 (N_11567,N_10340,N_10903);
or U11568 (N_11568,N_10276,N_10257);
nand U11569 (N_11569,N_10166,N_10087);
and U11570 (N_11570,N_10175,N_10476);
nor U11571 (N_11571,N_10153,N_10489);
nor U11572 (N_11572,N_10315,N_10208);
nor U11573 (N_11573,N_10524,N_10495);
and U11574 (N_11574,N_10202,N_10835);
nand U11575 (N_11575,N_10377,N_10992);
and U11576 (N_11576,N_10309,N_10294);
and U11577 (N_11577,N_10593,N_10991);
nand U11578 (N_11578,N_10886,N_10868);
nor U11579 (N_11579,N_10692,N_10367);
and U11580 (N_11580,N_10169,N_10675);
and U11581 (N_11581,N_10655,N_10064);
nand U11582 (N_11582,N_10741,N_10702);
nand U11583 (N_11583,N_10804,N_10081);
and U11584 (N_11584,N_10083,N_10231);
or U11585 (N_11585,N_10974,N_10521);
nand U11586 (N_11586,N_10656,N_10478);
and U11587 (N_11587,N_10839,N_10267);
xor U11588 (N_11588,N_10575,N_10120);
xor U11589 (N_11589,N_10246,N_10477);
and U11590 (N_11590,N_10218,N_10829);
or U11591 (N_11591,N_10282,N_10171);
or U11592 (N_11592,N_10719,N_10545);
nor U11593 (N_11593,N_10840,N_10171);
or U11594 (N_11594,N_10556,N_10027);
nand U11595 (N_11595,N_10784,N_10600);
nand U11596 (N_11596,N_10933,N_10693);
nor U11597 (N_11597,N_10979,N_10578);
or U11598 (N_11598,N_10120,N_10283);
nand U11599 (N_11599,N_10931,N_10409);
nand U11600 (N_11600,N_10249,N_10841);
nor U11601 (N_11601,N_10201,N_10378);
and U11602 (N_11602,N_10398,N_10415);
and U11603 (N_11603,N_10616,N_10386);
nor U11604 (N_11604,N_10493,N_10487);
nor U11605 (N_11605,N_10046,N_10422);
xnor U11606 (N_11606,N_10100,N_10350);
nand U11607 (N_11607,N_10133,N_10211);
nor U11608 (N_11608,N_10307,N_10251);
nand U11609 (N_11609,N_10764,N_10304);
and U11610 (N_11610,N_10887,N_10656);
and U11611 (N_11611,N_10594,N_10964);
xnor U11612 (N_11612,N_10944,N_10647);
or U11613 (N_11613,N_10822,N_10925);
or U11614 (N_11614,N_10863,N_10542);
nor U11615 (N_11615,N_10693,N_10862);
nand U11616 (N_11616,N_10880,N_10124);
or U11617 (N_11617,N_10433,N_10323);
nand U11618 (N_11618,N_10966,N_10944);
or U11619 (N_11619,N_10518,N_10600);
or U11620 (N_11620,N_10095,N_10369);
nor U11621 (N_11621,N_10775,N_10791);
or U11622 (N_11622,N_10557,N_10073);
nor U11623 (N_11623,N_10332,N_10131);
xor U11624 (N_11624,N_10168,N_10320);
or U11625 (N_11625,N_10806,N_10608);
nor U11626 (N_11626,N_10887,N_10988);
nor U11627 (N_11627,N_10629,N_10525);
nand U11628 (N_11628,N_10776,N_10299);
or U11629 (N_11629,N_10328,N_10037);
and U11630 (N_11630,N_10482,N_10313);
nand U11631 (N_11631,N_10652,N_10470);
nor U11632 (N_11632,N_10085,N_10336);
nand U11633 (N_11633,N_10977,N_10818);
or U11634 (N_11634,N_10568,N_10174);
or U11635 (N_11635,N_10396,N_10918);
nor U11636 (N_11636,N_10563,N_10118);
nand U11637 (N_11637,N_10939,N_10374);
and U11638 (N_11638,N_10237,N_10889);
nor U11639 (N_11639,N_10678,N_10173);
nand U11640 (N_11640,N_10348,N_10521);
xor U11641 (N_11641,N_10796,N_10354);
xnor U11642 (N_11642,N_10057,N_10351);
or U11643 (N_11643,N_10666,N_10863);
nor U11644 (N_11644,N_10341,N_10507);
nor U11645 (N_11645,N_10604,N_10010);
or U11646 (N_11646,N_10734,N_10627);
or U11647 (N_11647,N_10476,N_10828);
nor U11648 (N_11648,N_10836,N_10335);
or U11649 (N_11649,N_10778,N_10125);
and U11650 (N_11650,N_10598,N_10168);
or U11651 (N_11651,N_10399,N_10132);
or U11652 (N_11652,N_10628,N_10174);
nand U11653 (N_11653,N_10610,N_10454);
xor U11654 (N_11654,N_10977,N_10569);
nor U11655 (N_11655,N_10533,N_10537);
xnor U11656 (N_11656,N_10266,N_10457);
nor U11657 (N_11657,N_10016,N_10209);
nand U11658 (N_11658,N_10789,N_10103);
or U11659 (N_11659,N_10131,N_10432);
or U11660 (N_11660,N_10277,N_10951);
or U11661 (N_11661,N_10005,N_10567);
and U11662 (N_11662,N_10445,N_10796);
nand U11663 (N_11663,N_10581,N_10691);
nor U11664 (N_11664,N_10814,N_10651);
nor U11665 (N_11665,N_10219,N_10816);
and U11666 (N_11666,N_10043,N_10339);
and U11667 (N_11667,N_10582,N_10635);
or U11668 (N_11668,N_10755,N_10486);
or U11669 (N_11669,N_10941,N_10208);
nand U11670 (N_11670,N_10495,N_10253);
nor U11671 (N_11671,N_10856,N_10121);
nor U11672 (N_11672,N_10192,N_10953);
xnor U11673 (N_11673,N_10375,N_10475);
or U11674 (N_11674,N_10377,N_10964);
or U11675 (N_11675,N_10261,N_10837);
nor U11676 (N_11676,N_10635,N_10941);
nor U11677 (N_11677,N_10878,N_10303);
or U11678 (N_11678,N_10870,N_10740);
or U11679 (N_11679,N_10697,N_10189);
xnor U11680 (N_11680,N_10037,N_10856);
xor U11681 (N_11681,N_10609,N_10869);
or U11682 (N_11682,N_10117,N_10744);
nor U11683 (N_11683,N_10541,N_10290);
xnor U11684 (N_11684,N_10328,N_10100);
or U11685 (N_11685,N_10578,N_10708);
xnor U11686 (N_11686,N_10469,N_10771);
and U11687 (N_11687,N_10308,N_10250);
xor U11688 (N_11688,N_10729,N_10361);
nand U11689 (N_11689,N_10848,N_10127);
nor U11690 (N_11690,N_10661,N_10999);
and U11691 (N_11691,N_10098,N_10821);
nand U11692 (N_11692,N_10074,N_10844);
nand U11693 (N_11693,N_10039,N_10128);
or U11694 (N_11694,N_10639,N_10403);
nand U11695 (N_11695,N_10050,N_10689);
nor U11696 (N_11696,N_10156,N_10665);
xnor U11697 (N_11697,N_10679,N_10002);
and U11698 (N_11698,N_10497,N_10587);
and U11699 (N_11699,N_10947,N_10541);
nand U11700 (N_11700,N_10207,N_10580);
xnor U11701 (N_11701,N_10252,N_10929);
nand U11702 (N_11702,N_10424,N_10404);
nor U11703 (N_11703,N_10379,N_10572);
or U11704 (N_11704,N_10398,N_10089);
nor U11705 (N_11705,N_10813,N_10484);
xor U11706 (N_11706,N_10956,N_10418);
nand U11707 (N_11707,N_10742,N_10161);
or U11708 (N_11708,N_10165,N_10974);
nand U11709 (N_11709,N_10836,N_10357);
and U11710 (N_11710,N_10931,N_10076);
nor U11711 (N_11711,N_10735,N_10910);
xor U11712 (N_11712,N_10923,N_10883);
and U11713 (N_11713,N_10079,N_10059);
nor U11714 (N_11714,N_10530,N_10164);
xor U11715 (N_11715,N_10254,N_10967);
and U11716 (N_11716,N_10452,N_10136);
or U11717 (N_11717,N_10402,N_10845);
nand U11718 (N_11718,N_10797,N_10101);
nand U11719 (N_11719,N_10866,N_10409);
nand U11720 (N_11720,N_10516,N_10174);
nand U11721 (N_11721,N_10736,N_10778);
and U11722 (N_11722,N_10242,N_10606);
or U11723 (N_11723,N_10694,N_10339);
and U11724 (N_11724,N_10119,N_10388);
or U11725 (N_11725,N_10296,N_10113);
or U11726 (N_11726,N_10311,N_10611);
and U11727 (N_11727,N_10304,N_10014);
nand U11728 (N_11728,N_10526,N_10698);
nand U11729 (N_11729,N_10302,N_10860);
and U11730 (N_11730,N_10949,N_10529);
and U11731 (N_11731,N_10158,N_10778);
xnor U11732 (N_11732,N_10500,N_10239);
or U11733 (N_11733,N_10964,N_10568);
or U11734 (N_11734,N_10628,N_10435);
and U11735 (N_11735,N_10095,N_10847);
nor U11736 (N_11736,N_10270,N_10984);
or U11737 (N_11737,N_10922,N_10248);
and U11738 (N_11738,N_10684,N_10166);
nand U11739 (N_11739,N_10992,N_10267);
and U11740 (N_11740,N_10264,N_10074);
or U11741 (N_11741,N_10081,N_10013);
and U11742 (N_11742,N_10426,N_10839);
nor U11743 (N_11743,N_10065,N_10392);
and U11744 (N_11744,N_10807,N_10339);
nor U11745 (N_11745,N_10013,N_10141);
nor U11746 (N_11746,N_10755,N_10345);
nand U11747 (N_11747,N_10099,N_10969);
nor U11748 (N_11748,N_10704,N_10669);
and U11749 (N_11749,N_10917,N_10609);
nand U11750 (N_11750,N_10141,N_10821);
or U11751 (N_11751,N_10526,N_10871);
and U11752 (N_11752,N_10985,N_10197);
and U11753 (N_11753,N_10139,N_10957);
nand U11754 (N_11754,N_10543,N_10415);
or U11755 (N_11755,N_10743,N_10887);
nor U11756 (N_11756,N_10409,N_10570);
or U11757 (N_11757,N_10883,N_10186);
nand U11758 (N_11758,N_10177,N_10171);
nor U11759 (N_11759,N_10458,N_10085);
nand U11760 (N_11760,N_10880,N_10737);
or U11761 (N_11761,N_10291,N_10705);
and U11762 (N_11762,N_10764,N_10416);
nor U11763 (N_11763,N_10961,N_10791);
and U11764 (N_11764,N_10545,N_10751);
nor U11765 (N_11765,N_10200,N_10707);
or U11766 (N_11766,N_10910,N_10091);
or U11767 (N_11767,N_10490,N_10631);
nand U11768 (N_11768,N_10962,N_10671);
nor U11769 (N_11769,N_10991,N_10254);
nor U11770 (N_11770,N_10922,N_10352);
or U11771 (N_11771,N_10082,N_10886);
nand U11772 (N_11772,N_10305,N_10746);
and U11773 (N_11773,N_10516,N_10492);
or U11774 (N_11774,N_10723,N_10870);
nand U11775 (N_11775,N_10958,N_10116);
nand U11776 (N_11776,N_10328,N_10257);
or U11777 (N_11777,N_10909,N_10323);
and U11778 (N_11778,N_10823,N_10431);
or U11779 (N_11779,N_10670,N_10276);
nand U11780 (N_11780,N_10322,N_10411);
nand U11781 (N_11781,N_10900,N_10390);
or U11782 (N_11782,N_10873,N_10927);
and U11783 (N_11783,N_10342,N_10547);
or U11784 (N_11784,N_10269,N_10045);
and U11785 (N_11785,N_10705,N_10623);
xnor U11786 (N_11786,N_10913,N_10977);
and U11787 (N_11787,N_10136,N_10514);
and U11788 (N_11788,N_10581,N_10822);
and U11789 (N_11789,N_10498,N_10460);
xnor U11790 (N_11790,N_10853,N_10537);
xnor U11791 (N_11791,N_10749,N_10077);
or U11792 (N_11792,N_10615,N_10987);
xor U11793 (N_11793,N_10187,N_10224);
and U11794 (N_11794,N_10352,N_10065);
and U11795 (N_11795,N_10475,N_10683);
and U11796 (N_11796,N_10373,N_10523);
or U11797 (N_11797,N_10604,N_10389);
nor U11798 (N_11798,N_10253,N_10621);
nor U11799 (N_11799,N_10804,N_10758);
nor U11800 (N_11800,N_10708,N_10340);
or U11801 (N_11801,N_10973,N_10742);
nand U11802 (N_11802,N_10666,N_10444);
and U11803 (N_11803,N_10956,N_10824);
and U11804 (N_11804,N_10320,N_10936);
nand U11805 (N_11805,N_10194,N_10119);
nor U11806 (N_11806,N_10652,N_10892);
and U11807 (N_11807,N_10525,N_10591);
or U11808 (N_11808,N_10240,N_10243);
nand U11809 (N_11809,N_10838,N_10313);
or U11810 (N_11810,N_10393,N_10899);
and U11811 (N_11811,N_10135,N_10485);
or U11812 (N_11812,N_10206,N_10505);
nand U11813 (N_11813,N_10942,N_10422);
nand U11814 (N_11814,N_10434,N_10802);
and U11815 (N_11815,N_10239,N_10491);
and U11816 (N_11816,N_10225,N_10021);
or U11817 (N_11817,N_10977,N_10406);
and U11818 (N_11818,N_10186,N_10619);
nor U11819 (N_11819,N_10838,N_10481);
nand U11820 (N_11820,N_10142,N_10263);
or U11821 (N_11821,N_10569,N_10235);
xor U11822 (N_11822,N_10156,N_10653);
nand U11823 (N_11823,N_10962,N_10254);
and U11824 (N_11824,N_10485,N_10277);
or U11825 (N_11825,N_10874,N_10812);
nand U11826 (N_11826,N_10175,N_10955);
nor U11827 (N_11827,N_10686,N_10259);
nor U11828 (N_11828,N_10676,N_10218);
nand U11829 (N_11829,N_10341,N_10116);
xnor U11830 (N_11830,N_10566,N_10929);
or U11831 (N_11831,N_10245,N_10944);
or U11832 (N_11832,N_10291,N_10447);
xor U11833 (N_11833,N_10852,N_10595);
or U11834 (N_11834,N_10552,N_10970);
nor U11835 (N_11835,N_10304,N_10947);
nor U11836 (N_11836,N_10653,N_10819);
xor U11837 (N_11837,N_10850,N_10361);
and U11838 (N_11838,N_10178,N_10173);
nand U11839 (N_11839,N_10220,N_10366);
and U11840 (N_11840,N_10036,N_10249);
nor U11841 (N_11841,N_10205,N_10709);
nand U11842 (N_11842,N_10190,N_10012);
nor U11843 (N_11843,N_10716,N_10656);
xnor U11844 (N_11844,N_10974,N_10605);
nand U11845 (N_11845,N_10520,N_10644);
nand U11846 (N_11846,N_10896,N_10735);
and U11847 (N_11847,N_10989,N_10786);
nor U11848 (N_11848,N_10769,N_10447);
nor U11849 (N_11849,N_10833,N_10790);
nand U11850 (N_11850,N_10137,N_10576);
nand U11851 (N_11851,N_10775,N_10991);
and U11852 (N_11852,N_10751,N_10790);
or U11853 (N_11853,N_10904,N_10252);
xnor U11854 (N_11854,N_10684,N_10276);
nand U11855 (N_11855,N_10101,N_10604);
and U11856 (N_11856,N_10865,N_10804);
and U11857 (N_11857,N_10431,N_10736);
nand U11858 (N_11858,N_10166,N_10537);
nand U11859 (N_11859,N_10754,N_10771);
and U11860 (N_11860,N_10310,N_10671);
nor U11861 (N_11861,N_10403,N_10689);
or U11862 (N_11862,N_10540,N_10528);
nor U11863 (N_11863,N_10341,N_10442);
or U11864 (N_11864,N_10729,N_10024);
and U11865 (N_11865,N_10224,N_10543);
nand U11866 (N_11866,N_10827,N_10406);
or U11867 (N_11867,N_10549,N_10142);
xnor U11868 (N_11868,N_10566,N_10438);
nor U11869 (N_11869,N_10725,N_10070);
and U11870 (N_11870,N_10621,N_10853);
nand U11871 (N_11871,N_10265,N_10506);
and U11872 (N_11872,N_10425,N_10325);
nor U11873 (N_11873,N_10212,N_10807);
nand U11874 (N_11874,N_10641,N_10955);
nand U11875 (N_11875,N_10147,N_10766);
nor U11876 (N_11876,N_10213,N_10750);
and U11877 (N_11877,N_10140,N_10012);
or U11878 (N_11878,N_10406,N_10964);
and U11879 (N_11879,N_10458,N_10169);
and U11880 (N_11880,N_10031,N_10701);
and U11881 (N_11881,N_10444,N_10487);
nand U11882 (N_11882,N_10617,N_10845);
nor U11883 (N_11883,N_10651,N_10523);
or U11884 (N_11884,N_10733,N_10279);
nor U11885 (N_11885,N_10886,N_10726);
nor U11886 (N_11886,N_10128,N_10643);
and U11887 (N_11887,N_10009,N_10964);
nand U11888 (N_11888,N_10829,N_10464);
or U11889 (N_11889,N_10606,N_10973);
nor U11890 (N_11890,N_10907,N_10448);
and U11891 (N_11891,N_10948,N_10031);
or U11892 (N_11892,N_10221,N_10595);
nor U11893 (N_11893,N_10449,N_10158);
and U11894 (N_11894,N_10063,N_10231);
or U11895 (N_11895,N_10639,N_10530);
and U11896 (N_11896,N_10108,N_10829);
nor U11897 (N_11897,N_10230,N_10756);
or U11898 (N_11898,N_10001,N_10088);
nor U11899 (N_11899,N_10303,N_10606);
nor U11900 (N_11900,N_10242,N_10875);
xnor U11901 (N_11901,N_10941,N_10337);
nor U11902 (N_11902,N_10154,N_10059);
and U11903 (N_11903,N_10237,N_10575);
or U11904 (N_11904,N_10775,N_10708);
nor U11905 (N_11905,N_10622,N_10082);
or U11906 (N_11906,N_10812,N_10237);
nand U11907 (N_11907,N_10301,N_10627);
nor U11908 (N_11908,N_10153,N_10393);
or U11909 (N_11909,N_10313,N_10810);
nor U11910 (N_11910,N_10379,N_10280);
nand U11911 (N_11911,N_10026,N_10118);
nand U11912 (N_11912,N_10875,N_10415);
nor U11913 (N_11913,N_10637,N_10450);
or U11914 (N_11914,N_10608,N_10486);
nor U11915 (N_11915,N_10447,N_10820);
or U11916 (N_11916,N_10093,N_10342);
nand U11917 (N_11917,N_10749,N_10790);
nand U11918 (N_11918,N_10929,N_10080);
nand U11919 (N_11919,N_10270,N_10216);
or U11920 (N_11920,N_10947,N_10110);
or U11921 (N_11921,N_10398,N_10998);
nor U11922 (N_11922,N_10882,N_10739);
nor U11923 (N_11923,N_10154,N_10798);
and U11924 (N_11924,N_10258,N_10999);
or U11925 (N_11925,N_10845,N_10408);
nor U11926 (N_11926,N_10110,N_10557);
nor U11927 (N_11927,N_10088,N_10980);
or U11928 (N_11928,N_10496,N_10701);
nor U11929 (N_11929,N_10575,N_10434);
nor U11930 (N_11930,N_10861,N_10477);
or U11931 (N_11931,N_10137,N_10186);
xor U11932 (N_11932,N_10475,N_10372);
nor U11933 (N_11933,N_10632,N_10677);
nand U11934 (N_11934,N_10481,N_10353);
and U11935 (N_11935,N_10070,N_10185);
and U11936 (N_11936,N_10563,N_10022);
nor U11937 (N_11937,N_10536,N_10318);
nand U11938 (N_11938,N_10908,N_10619);
nand U11939 (N_11939,N_10875,N_10631);
nor U11940 (N_11940,N_10705,N_10300);
nor U11941 (N_11941,N_10772,N_10431);
nor U11942 (N_11942,N_10912,N_10346);
or U11943 (N_11943,N_10712,N_10213);
and U11944 (N_11944,N_10817,N_10097);
nor U11945 (N_11945,N_10749,N_10877);
nor U11946 (N_11946,N_10851,N_10914);
xor U11947 (N_11947,N_10656,N_10741);
nand U11948 (N_11948,N_10300,N_10840);
nand U11949 (N_11949,N_10401,N_10503);
xnor U11950 (N_11950,N_10416,N_10148);
and U11951 (N_11951,N_10113,N_10809);
nor U11952 (N_11952,N_10244,N_10027);
nor U11953 (N_11953,N_10066,N_10700);
and U11954 (N_11954,N_10945,N_10780);
nand U11955 (N_11955,N_10551,N_10569);
or U11956 (N_11956,N_10345,N_10815);
or U11957 (N_11957,N_10222,N_10553);
or U11958 (N_11958,N_10214,N_10033);
nand U11959 (N_11959,N_10970,N_10389);
nor U11960 (N_11960,N_10748,N_10609);
and U11961 (N_11961,N_10694,N_10371);
nand U11962 (N_11962,N_10057,N_10931);
nor U11963 (N_11963,N_10457,N_10923);
and U11964 (N_11964,N_10560,N_10310);
nor U11965 (N_11965,N_10854,N_10445);
nand U11966 (N_11966,N_10214,N_10792);
or U11967 (N_11967,N_10223,N_10041);
or U11968 (N_11968,N_10679,N_10893);
and U11969 (N_11969,N_10105,N_10992);
xor U11970 (N_11970,N_10546,N_10592);
nor U11971 (N_11971,N_10991,N_10560);
or U11972 (N_11972,N_10297,N_10548);
and U11973 (N_11973,N_10220,N_10393);
xnor U11974 (N_11974,N_10417,N_10576);
nor U11975 (N_11975,N_10957,N_10809);
nor U11976 (N_11976,N_10043,N_10809);
nor U11977 (N_11977,N_10585,N_10120);
or U11978 (N_11978,N_10990,N_10556);
or U11979 (N_11979,N_10759,N_10047);
xor U11980 (N_11980,N_10868,N_10994);
and U11981 (N_11981,N_10388,N_10549);
nand U11982 (N_11982,N_10171,N_10038);
or U11983 (N_11983,N_10397,N_10011);
and U11984 (N_11984,N_10703,N_10402);
and U11985 (N_11985,N_10032,N_10542);
or U11986 (N_11986,N_10491,N_10056);
nor U11987 (N_11987,N_10297,N_10151);
or U11988 (N_11988,N_10702,N_10786);
nand U11989 (N_11989,N_10874,N_10272);
nor U11990 (N_11990,N_10178,N_10081);
nor U11991 (N_11991,N_10811,N_10840);
and U11992 (N_11992,N_10280,N_10815);
or U11993 (N_11993,N_10753,N_10779);
nor U11994 (N_11994,N_10256,N_10580);
nand U11995 (N_11995,N_10793,N_10883);
nor U11996 (N_11996,N_10796,N_10985);
nand U11997 (N_11997,N_10009,N_10694);
nor U11998 (N_11998,N_10553,N_10457);
nand U11999 (N_11999,N_10660,N_10169);
or U12000 (N_12000,N_11177,N_11468);
and U12001 (N_12001,N_11519,N_11332);
nand U12002 (N_12002,N_11983,N_11728);
or U12003 (N_12003,N_11247,N_11084);
nor U12004 (N_12004,N_11736,N_11751);
nand U12005 (N_12005,N_11666,N_11484);
and U12006 (N_12006,N_11859,N_11368);
and U12007 (N_12007,N_11581,N_11241);
nor U12008 (N_12008,N_11524,N_11788);
nand U12009 (N_12009,N_11033,N_11020);
nand U12010 (N_12010,N_11779,N_11361);
and U12011 (N_12011,N_11287,N_11659);
or U12012 (N_12012,N_11086,N_11303);
xnor U12013 (N_12013,N_11937,N_11221);
or U12014 (N_12014,N_11562,N_11698);
or U12015 (N_12015,N_11931,N_11275);
or U12016 (N_12016,N_11929,N_11956);
nor U12017 (N_12017,N_11913,N_11024);
and U12018 (N_12018,N_11656,N_11188);
or U12019 (N_12019,N_11336,N_11180);
nand U12020 (N_12020,N_11535,N_11497);
nor U12021 (N_12021,N_11492,N_11844);
nor U12022 (N_12022,N_11193,N_11057);
nand U12023 (N_12023,N_11328,N_11312);
or U12024 (N_12024,N_11610,N_11002);
nor U12025 (N_12025,N_11867,N_11137);
and U12026 (N_12026,N_11419,N_11218);
and U12027 (N_12027,N_11032,N_11110);
or U12028 (N_12028,N_11650,N_11008);
or U12029 (N_12029,N_11989,N_11754);
xor U12030 (N_12030,N_11070,N_11632);
xor U12031 (N_12031,N_11044,N_11596);
or U12032 (N_12032,N_11371,N_11098);
or U12033 (N_12033,N_11104,N_11615);
xnor U12034 (N_12034,N_11403,N_11628);
and U12035 (N_12035,N_11129,N_11012);
and U12036 (N_12036,N_11962,N_11415);
nor U12037 (N_12037,N_11087,N_11470);
nor U12038 (N_12038,N_11880,N_11749);
nand U12039 (N_12039,N_11317,N_11261);
xnor U12040 (N_12040,N_11267,N_11776);
and U12041 (N_12041,N_11392,N_11223);
or U12042 (N_12042,N_11669,N_11256);
or U12043 (N_12043,N_11250,N_11083);
nor U12044 (N_12044,N_11508,N_11542);
nor U12045 (N_12045,N_11925,N_11340);
nor U12046 (N_12046,N_11485,N_11100);
nor U12047 (N_12047,N_11374,N_11244);
nor U12048 (N_12048,N_11427,N_11118);
nand U12049 (N_12049,N_11406,N_11451);
xor U12050 (N_12050,N_11805,N_11832);
or U12051 (N_12051,N_11428,N_11201);
or U12052 (N_12052,N_11220,N_11851);
or U12053 (N_12053,N_11362,N_11639);
and U12054 (N_12054,N_11270,N_11385);
nand U12055 (N_12055,N_11390,N_11498);
nand U12056 (N_12056,N_11953,N_11882);
and U12057 (N_12057,N_11721,N_11023);
and U12058 (N_12058,N_11539,N_11903);
nand U12059 (N_12059,N_11661,N_11949);
or U12060 (N_12060,N_11954,N_11899);
or U12061 (N_12061,N_11101,N_11151);
nand U12062 (N_12062,N_11471,N_11706);
or U12063 (N_12063,N_11119,N_11993);
or U12064 (N_12064,N_11696,N_11109);
xnor U12065 (N_12065,N_11633,N_11856);
nor U12066 (N_12066,N_11147,N_11263);
nor U12067 (N_12067,N_11552,N_11001);
nor U12068 (N_12068,N_11046,N_11528);
and U12069 (N_12069,N_11257,N_11817);
and U12070 (N_12070,N_11394,N_11773);
nand U12071 (N_12071,N_11347,N_11812);
or U12072 (N_12072,N_11836,N_11125);
xor U12073 (N_12073,N_11324,N_11316);
nor U12074 (N_12074,N_11074,N_11797);
xnor U12075 (N_12075,N_11928,N_11740);
or U12076 (N_12076,N_11240,N_11729);
xor U12077 (N_12077,N_11830,N_11387);
and U12078 (N_12078,N_11759,N_11800);
and U12079 (N_12079,N_11814,N_11770);
nand U12080 (N_12080,N_11479,N_11356);
nor U12081 (N_12081,N_11575,N_11208);
xor U12082 (N_12082,N_11062,N_11231);
xnor U12083 (N_12083,N_11169,N_11093);
nand U12084 (N_12084,N_11136,N_11234);
nand U12085 (N_12085,N_11671,N_11771);
nor U12086 (N_12086,N_11393,N_11548);
or U12087 (N_12087,N_11467,N_11107);
and U12088 (N_12088,N_11541,N_11975);
nand U12089 (N_12089,N_11516,N_11888);
or U12090 (N_12090,N_11653,N_11019);
xor U12091 (N_12091,N_11420,N_11727);
xnor U12092 (N_12092,N_11618,N_11963);
or U12093 (N_12093,N_11298,N_11818);
nor U12094 (N_12094,N_11054,N_11922);
xnor U12095 (N_12095,N_11643,N_11785);
or U12096 (N_12096,N_11733,N_11595);
nor U12097 (N_12097,N_11563,N_11277);
and U12098 (N_12098,N_11782,N_11383);
nor U12099 (N_12099,N_11273,N_11571);
or U12100 (N_12100,N_11538,N_11175);
nor U12101 (N_12101,N_11058,N_11053);
nand U12102 (N_12102,N_11682,N_11737);
xor U12103 (N_12103,N_11441,N_11358);
or U12104 (N_12104,N_11911,N_11703);
and U12105 (N_12105,N_11917,N_11052);
or U12106 (N_12106,N_11710,N_11909);
nand U12107 (N_12107,N_11342,N_11846);
or U12108 (N_12108,N_11158,N_11970);
nand U12109 (N_12109,N_11399,N_11602);
xor U12110 (N_12110,N_11629,N_11613);
nand U12111 (N_12111,N_11013,N_11527);
or U12112 (N_12112,N_11081,N_11212);
and U12113 (N_12113,N_11724,N_11640);
xor U12114 (N_12114,N_11570,N_11819);
and U12115 (N_12115,N_11700,N_11007);
nand U12116 (N_12116,N_11743,N_11999);
nor U12117 (N_12117,N_11339,N_11326);
nand U12118 (N_12118,N_11689,N_11364);
and U12119 (N_12119,N_11676,N_11748);
nand U12120 (N_12120,N_11152,N_11233);
nand U12121 (N_12121,N_11413,N_11604);
and U12122 (N_12122,N_11404,N_11139);
xor U12123 (N_12123,N_11480,N_11506);
or U12124 (N_12124,N_11076,N_11133);
nand U12125 (N_12125,N_11799,N_11744);
and U12126 (N_12126,N_11337,N_11915);
nor U12127 (N_12127,N_11434,N_11646);
and U12128 (N_12128,N_11688,N_11554);
and U12129 (N_12129,N_11121,N_11369);
xnor U12130 (N_12130,N_11319,N_11472);
nand U12131 (N_12131,N_11977,N_11955);
or U12132 (N_12132,N_11536,N_11711);
and U12133 (N_12133,N_11483,N_11335);
or U12134 (N_12134,N_11907,N_11938);
nand U12135 (N_12135,N_11105,N_11841);
nand U12136 (N_12136,N_11707,N_11280);
or U12137 (N_12137,N_11855,N_11190);
nor U12138 (N_12138,N_11908,N_11354);
nand U12139 (N_12139,N_11705,N_11474);
and U12140 (N_12140,N_11274,N_11616);
and U12141 (N_12141,N_11936,N_11300);
and U12142 (N_12142,N_11367,N_11685);
and U12143 (N_12143,N_11246,N_11894);
and U12144 (N_12144,N_11806,N_11069);
nand U12145 (N_12145,N_11864,N_11852);
and U12146 (N_12146,N_11224,N_11510);
or U12147 (N_12147,N_11122,N_11626);
nor U12148 (N_12148,N_11278,N_11195);
nand U12149 (N_12149,N_11893,N_11322);
nand U12150 (N_12150,N_11308,N_11652);
nor U12151 (N_12151,N_11589,N_11126);
nand U12152 (N_12152,N_11810,N_11684);
or U12153 (N_12153,N_11041,N_11421);
and U12154 (N_12154,N_11411,N_11886);
nand U12155 (N_12155,N_11833,N_11828);
nand U12156 (N_12156,N_11329,N_11251);
or U12157 (N_12157,N_11725,N_11625);
nor U12158 (N_12158,N_11416,N_11745);
or U12159 (N_12159,N_11934,N_11601);
nor U12160 (N_12160,N_11741,N_11059);
and U12161 (N_12161,N_11478,N_11892);
nor U12162 (N_12162,N_11884,N_11436);
or U12163 (N_12163,N_11591,N_11198);
xnor U12164 (N_12164,N_11798,N_11330);
xor U12165 (N_12165,N_11866,N_11352);
nand U12166 (N_12166,N_11967,N_11793);
and U12167 (N_12167,N_11488,N_11919);
or U12168 (N_12168,N_11772,N_11588);
or U12169 (N_12169,N_11567,N_11163);
xor U12170 (N_12170,N_11526,N_11445);
and U12171 (N_12171,N_11040,N_11765);
nand U12172 (N_12172,N_11191,N_11932);
or U12173 (N_12173,N_11709,N_11149);
nor U12174 (N_12174,N_11540,N_11714);
nor U12175 (N_12175,N_11140,N_11237);
and U12176 (N_12176,N_11973,N_11473);
or U12177 (N_12177,N_11717,N_11437);
nand U12178 (N_12178,N_11612,N_11847);
nand U12179 (N_12179,N_11811,N_11071);
nand U12180 (N_12180,N_11486,N_11944);
nor U12181 (N_12181,N_11637,N_11114);
nand U12182 (N_12182,N_11378,N_11769);
nand U12183 (N_12183,N_11363,N_11873);
xor U12184 (N_12184,N_11285,N_11874);
nor U12185 (N_12185,N_11726,N_11004);
or U12186 (N_12186,N_11144,N_11172);
or U12187 (N_12187,N_11853,N_11469);
nor U12188 (N_12188,N_11550,N_11758);
or U12189 (N_12189,N_11502,N_11216);
and U12190 (N_12190,N_11295,N_11286);
and U12191 (N_12191,N_11649,N_11900);
xnor U12192 (N_12192,N_11870,N_11202);
nand U12193 (N_12193,N_11631,N_11890);
and U12194 (N_12194,N_11410,N_11957);
nor U12195 (N_12195,N_11382,N_11245);
nand U12196 (N_12196,N_11092,N_11547);
or U12197 (N_12197,N_11569,N_11843);
and U12198 (N_12198,N_11720,N_11395);
or U12199 (N_12199,N_11226,N_11658);
nor U12200 (N_12200,N_11826,N_11222);
xnor U12201 (N_12201,N_11127,N_11397);
or U12202 (N_12202,N_11065,N_11493);
nand U12203 (N_12203,N_11630,N_11842);
nor U12204 (N_12204,N_11608,N_11461);
nand U12205 (N_12205,N_11518,N_11296);
or U12206 (N_12206,N_11102,N_11896);
nand U12207 (N_12207,N_11386,N_11947);
nor U12208 (N_12208,N_11080,N_11006);
and U12209 (N_12209,N_11499,N_11732);
and U12210 (N_12210,N_11822,N_11292);
or U12211 (N_12211,N_11790,N_11346);
nand U12212 (N_12212,N_11009,N_11966);
nand U12213 (N_12213,N_11253,N_11227);
nor U12214 (N_12214,N_11138,N_11375);
nand U12215 (N_12215,N_11553,N_11981);
and U12216 (N_12216,N_11439,N_11960);
xnor U12217 (N_12217,N_11863,N_11412);
or U12218 (N_12218,N_11360,N_11108);
nand U12219 (N_12219,N_11804,N_11454);
xnor U12220 (N_12220,N_11171,N_11763);
nand U12221 (N_12221,N_11746,N_11283);
or U12222 (N_12222,N_11066,N_11760);
or U12223 (N_12223,N_11000,N_11865);
or U12224 (N_12224,N_11945,N_11881);
xnor U12225 (N_12225,N_11134,N_11096);
nor U12226 (N_12226,N_11789,N_11444);
and U12227 (N_12227,N_11681,N_11161);
nand U12228 (N_12228,N_11834,N_11091);
nor U12229 (N_12229,N_11657,N_11848);
nor U12230 (N_12230,N_11564,N_11290);
and U12231 (N_12231,N_11897,N_11641);
nor U12232 (N_12232,N_11787,N_11113);
nor U12233 (N_12233,N_11775,N_11574);
or U12234 (N_12234,N_11872,N_11568);
and U12235 (N_12235,N_11145,N_11597);
nor U12236 (N_12236,N_11036,N_11877);
and U12237 (N_12237,N_11460,N_11675);
nand U12238 (N_12238,N_11513,N_11142);
and U12239 (N_12239,N_11898,N_11320);
and U12240 (N_12240,N_11213,N_11606);
nor U12241 (N_12241,N_11225,N_11085);
nor U12242 (N_12242,N_11477,N_11579);
or U12243 (N_12243,N_11803,N_11901);
nor U12244 (N_12244,N_11935,N_11948);
nor U12245 (N_12245,N_11808,N_11585);
nand U12246 (N_12246,N_11672,N_11715);
nor U12247 (N_12247,N_11294,N_11148);
or U12248 (N_12248,N_11941,N_11991);
nor U12249 (N_12249,N_11584,N_11910);
nand U12250 (N_12250,N_11777,N_11174);
and U12251 (N_12251,N_11723,N_11159);
or U12252 (N_12252,N_11166,N_11160);
or U12253 (N_12253,N_11692,N_11796);
nand U12254 (N_12254,N_11203,N_11704);
or U12255 (N_12255,N_11690,N_11505);
and U12256 (N_12256,N_11599,N_11667);
or U12257 (N_12257,N_11665,N_11755);
and U12258 (N_12258,N_11365,N_11774);
nand U12259 (N_12259,N_11614,N_11534);
xor U12260 (N_12260,N_11572,N_11912);
nand U12261 (N_12261,N_11039,N_11210);
or U12262 (N_12262,N_11854,N_11543);
nor U12263 (N_12263,N_11349,N_11959);
or U12264 (N_12264,N_11022,N_11200);
nor U12265 (N_12265,N_11176,N_11401);
nor U12266 (N_12266,N_11974,N_11099);
nor U12267 (N_12267,N_11103,N_11738);
nor U12268 (N_12268,N_11425,N_11146);
or U12269 (N_12269,N_11940,N_11670);
nand U12270 (N_12270,N_11090,N_11164);
and U12271 (N_12271,N_11314,N_11219);
or U12272 (N_12272,N_11338,N_11742);
xor U12273 (N_12273,N_11942,N_11232);
or U12274 (N_12274,N_11402,N_11952);
or U12275 (N_12275,N_11593,N_11475);
or U12276 (N_12276,N_11334,N_11580);
nand U12277 (N_12277,N_11265,N_11544);
or U12278 (N_12278,N_11357,N_11209);
nand U12279 (N_12279,N_11930,N_11752);
nand U12280 (N_12280,N_11838,N_11824);
nand U12281 (N_12281,N_11924,N_11801);
nor U12282 (N_12282,N_11885,N_11079);
or U12283 (N_12283,N_11398,N_11035);
nor U12284 (N_12284,N_11879,N_11345);
and U12285 (N_12285,N_11611,N_11181);
nor U12286 (N_12286,N_11426,N_11279);
nor U12287 (N_12287,N_11123,N_11077);
nor U12288 (N_12288,N_11998,N_11964);
nand U12289 (N_12289,N_11624,N_11400);
or U12290 (N_12290,N_11687,N_11132);
and U12291 (N_12291,N_11654,N_11305);
and U12292 (N_12292,N_11430,N_11409);
nand U12293 (N_12293,N_11405,N_11115);
nand U12294 (N_12294,N_11868,N_11701);
nor U12295 (N_12295,N_11958,N_11487);
and U12296 (N_12296,N_11313,N_11521);
and U12297 (N_12297,N_11075,N_11592);
nand U12298 (N_12298,N_11691,N_11943);
nor U12299 (N_12299,N_11259,N_11282);
and U12300 (N_12300,N_11695,N_11239);
nand U12301 (N_12301,N_11379,N_11926);
nor U12302 (N_12302,N_11056,N_11600);
and U12303 (N_12303,N_11716,N_11556);
nand U12304 (N_12304,N_11179,N_11323);
or U12305 (N_12305,N_11266,N_11289);
nor U12306 (N_12306,N_11533,N_11594);
and U12307 (N_12307,N_11230,N_11235);
and U12308 (N_12308,N_11141,N_11627);
or U12309 (N_12309,N_11713,N_11450);
xor U12310 (N_12310,N_11262,N_11598);
nor U12311 (N_12311,N_11994,N_11781);
and U12312 (N_12312,N_11355,N_11719);
nor U12313 (N_12313,N_11916,N_11809);
and U12314 (N_12314,N_11990,N_11984);
or U12315 (N_12315,N_11921,N_11311);
nor U12316 (N_12316,N_11010,N_11047);
nor U12317 (N_12317,N_11635,N_11228);
and U12318 (N_12318,N_11545,N_11623);
nor U12319 (N_12319,N_11590,N_11353);
nor U12320 (N_12320,N_11423,N_11197);
and U12321 (N_12321,N_11429,N_11673);
and U12322 (N_12322,N_11918,N_11620);
nand U12323 (N_12323,N_11366,N_11578);
nand U12324 (N_12324,N_11016,N_11186);
nor U12325 (N_12325,N_11531,N_11965);
nand U12326 (N_12326,N_11694,N_11184);
xor U12327 (N_12327,N_11862,N_11587);
or U12328 (N_12328,N_11802,N_11753);
or U12329 (N_12329,N_11117,N_11422);
xor U12330 (N_12330,N_11432,N_11061);
xnor U12331 (N_12331,N_11871,N_11979);
and U12332 (N_12332,N_11242,N_11301);
nor U12333 (N_12333,N_11529,N_11525);
nand U12334 (N_12334,N_11391,N_11827);
nand U12335 (N_12335,N_11154,N_11622);
nor U12336 (N_12336,N_11530,N_11546);
or U12337 (N_12337,N_11786,N_11064);
or U12338 (N_12338,N_11414,N_11651);
nand U12339 (N_12339,N_11206,N_11939);
and U12340 (N_12340,N_11557,N_11968);
nand U12341 (N_12341,N_11088,N_11996);
or U12342 (N_12342,N_11150,N_11082);
and U12343 (N_12343,N_11417,N_11243);
nor U12344 (N_12344,N_11214,N_11333);
nand U12345 (N_12345,N_11807,N_11609);
or U12346 (N_12346,N_11747,N_11045);
nor U12347 (N_12347,N_11784,N_11350);
xor U12348 (N_12348,N_11783,N_11517);
or U12349 (N_12349,N_11331,N_11189);
nand U12350 (N_12350,N_11372,N_11351);
nor U12351 (N_12351,N_11522,N_11304);
and U12352 (N_12352,N_11453,N_11048);
nand U12353 (N_12353,N_11211,N_11566);
nand U12354 (N_12354,N_11951,N_11730);
xor U12355 (N_12355,N_11466,N_11995);
or U12356 (N_12356,N_11820,N_11565);
nor U12357 (N_12357,N_11458,N_11731);
xnor U12358 (N_12358,N_11686,N_11252);
nand U12359 (N_12359,N_11549,N_11792);
or U12360 (N_12360,N_11586,N_11858);
nand U12361 (N_12361,N_11238,N_11850);
or U12362 (N_12362,N_11835,N_11043);
or U12363 (N_12363,N_11825,N_11168);
nor U12364 (N_12364,N_11537,N_11389);
nor U12365 (N_12365,N_11645,N_11143);
and U12366 (N_12366,N_11813,N_11097);
nand U12367 (N_12367,N_11271,N_11971);
nor U12368 (N_12368,N_11976,N_11173);
nand U12369 (N_12369,N_11170,N_11302);
and U12370 (N_12370,N_11560,N_11465);
xor U12371 (N_12371,N_11875,N_11923);
and U12372 (N_12372,N_11555,N_11377);
or U12373 (N_12373,N_11734,N_11512);
nand U12374 (N_12374,N_11603,N_11507);
nor U12375 (N_12375,N_11025,N_11424);
and U12376 (N_12376,N_11987,N_11757);
xor U12377 (N_12377,N_11373,N_11038);
nand U12378 (N_12378,N_11205,N_11217);
or U12379 (N_12379,N_11722,N_11481);
xor U12380 (N_12380,N_11260,N_11491);
or U12381 (N_12381,N_11583,N_11291);
and U12382 (N_12382,N_11318,N_11985);
or U12383 (N_12383,N_11457,N_11307);
nand U12384 (N_12384,N_11343,N_11514);
nand U12385 (N_12385,N_11264,N_11327);
or U12386 (N_12386,N_11523,N_11381);
xor U12387 (N_12387,N_11456,N_11462);
or U12388 (N_12388,N_11162,N_11494);
nand U12389 (N_12389,N_11003,N_11559);
nand U12390 (N_12390,N_11876,N_11490);
and U12391 (N_12391,N_11027,N_11914);
nand U12392 (N_12392,N_11840,N_11055);
or U12393 (N_12393,N_11095,N_11452);
nand U12394 (N_12394,N_11376,N_11718);
xnor U12395 (N_12395,N_11795,N_11028);
nor U12396 (N_12396,N_11664,N_11997);
xor U12397 (N_12397,N_11299,N_11920);
or U12398 (N_12398,N_11185,N_11447);
nor U12399 (N_12399,N_11895,N_11577);
nand U12400 (N_12400,N_11482,N_11648);
xor U12401 (N_12401,N_11204,N_11116);
and U12402 (N_12402,N_11605,N_11449);
and U12403 (N_12403,N_11780,N_11750);
nor U12404 (N_12404,N_11455,N_11933);
and U12405 (N_12405,N_11662,N_11018);
nand U12406 (N_12406,N_11255,N_11380);
nand U12407 (N_12407,N_11464,N_11607);
and U12408 (N_12408,N_11845,N_11551);
xnor U12409 (N_12409,N_11702,N_11031);
nor U12410 (N_12410,N_11504,N_11849);
or U12411 (N_12411,N_11120,N_11005);
and U12412 (N_12412,N_11130,N_11644);
xor U12413 (N_12413,N_11905,N_11268);
or U12414 (N_12414,N_11199,N_11988);
and U12415 (N_12415,N_11015,N_11693);
or U12416 (N_12416,N_11438,N_11683);
nand U12417 (N_12417,N_11094,N_11906);
nand U12418 (N_12418,N_11128,N_11857);
nor U12419 (N_12419,N_11050,N_11156);
or U12420 (N_12420,N_11310,N_11660);
nor U12421 (N_12421,N_11167,N_11215);
nand U12422 (N_12422,N_11756,N_11794);
nand U12423 (N_12423,N_11576,N_11764);
or U12424 (N_12424,N_11463,N_11124);
nand U12425 (N_12425,N_11861,N_11236);
and U12426 (N_12426,N_11011,N_11839);
nand U12427 (N_12427,N_11739,N_11297);
nor U12428 (N_12428,N_11677,N_11321);
nor U12429 (N_12429,N_11254,N_11443);
or U12430 (N_12430,N_11674,N_11837);
and U12431 (N_12431,N_11980,N_11778);
xnor U12432 (N_12432,N_11821,N_11207);
or U12433 (N_12433,N_11511,N_11978);
nor U12434 (N_12434,N_11761,N_11249);
nor U12435 (N_12435,N_11388,N_11021);
xor U12436 (N_12436,N_11192,N_11663);
nand U12437 (N_12437,N_11532,N_11068);
or U12438 (N_12438,N_11276,N_11829);
nand U12439 (N_12439,N_11904,N_11946);
or U12440 (N_12440,N_11902,N_11418);
nand U12441 (N_12441,N_11636,N_11131);
nand U12442 (N_12442,N_11992,N_11678);
nor U12443 (N_12443,N_11878,N_11306);
nor U12444 (N_12444,N_11293,N_11489);
nand U12445 (N_12445,N_11972,N_11153);
or U12446 (N_12446,N_11157,N_11655);
or U12447 (N_12447,N_11459,N_11766);
and U12448 (N_12448,N_11344,N_11448);
xor U12449 (N_12449,N_11638,N_11582);
nor U12450 (N_12450,N_11619,N_11768);
and U12451 (N_12451,N_11961,N_11708);
or U12452 (N_12452,N_11816,N_11073);
or U12453 (N_12453,N_11325,N_11509);
nor U12454 (N_12454,N_11823,N_11229);
xnor U12455 (N_12455,N_11634,N_11183);
nand U12456 (N_12456,N_11341,N_11182);
xor U12457 (N_12457,N_11049,N_11284);
nand U12458 (N_12458,N_11433,N_11680);
nand U12459 (N_12459,N_11735,N_11359);
nand U12460 (N_12460,N_11037,N_11178);
xnor U12461 (N_12461,N_11089,N_11515);
or U12462 (N_12462,N_11869,N_11396);
xnor U12463 (N_12463,N_11067,N_11196);
nor U12464 (N_12464,N_11791,N_11815);
nor U12465 (N_12465,N_11520,N_11927);
nor U12466 (N_12466,N_11969,N_11982);
nand U12467 (N_12467,N_11194,N_11621);
xor U12468 (N_12468,N_11647,N_11135);
and U12469 (N_12469,N_11112,N_11281);
nor U12470 (N_12470,N_11558,N_11496);
or U12471 (N_12471,N_11561,N_11889);
nor U12472 (N_12472,N_11891,N_11034);
and U12473 (N_12473,N_11446,N_11106);
nand U12474 (N_12474,N_11440,N_11155);
nor U12475 (N_12475,N_11017,N_11072);
or U12476 (N_12476,N_11501,N_11617);
nor U12477 (N_12477,N_11883,N_11370);
or U12478 (N_12478,N_11762,N_11030);
xor U12479 (N_12479,N_11315,N_11573);
nand U12480 (N_12480,N_11272,N_11679);
nand U12481 (N_12481,N_11063,N_11697);
and U12482 (N_12482,N_11503,N_11029);
xor U12483 (N_12483,N_11668,N_11288);
or U12484 (N_12484,N_11348,N_11500);
or U12485 (N_12485,N_11431,N_11699);
nand U12486 (N_12486,N_11060,N_11384);
or U12487 (N_12487,N_11165,N_11248);
xor U12488 (N_12488,N_11408,N_11767);
nand U12489 (N_12489,N_11476,N_11887);
nor U12490 (N_12490,N_11950,N_11258);
nand U12491 (N_12491,N_11026,N_11407);
and U12492 (N_12492,N_11051,N_11309);
or U12493 (N_12493,N_11831,N_11860);
or U12494 (N_12494,N_11495,N_11712);
and U12495 (N_12495,N_11014,N_11078);
or U12496 (N_12496,N_11111,N_11986);
xor U12497 (N_12497,N_11442,N_11187);
and U12498 (N_12498,N_11269,N_11435);
nand U12499 (N_12499,N_11642,N_11042);
or U12500 (N_12500,N_11046,N_11871);
nor U12501 (N_12501,N_11157,N_11929);
nand U12502 (N_12502,N_11874,N_11392);
or U12503 (N_12503,N_11453,N_11776);
nand U12504 (N_12504,N_11099,N_11407);
nand U12505 (N_12505,N_11579,N_11200);
or U12506 (N_12506,N_11837,N_11113);
nor U12507 (N_12507,N_11090,N_11817);
nor U12508 (N_12508,N_11427,N_11720);
or U12509 (N_12509,N_11573,N_11723);
or U12510 (N_12510,N_11436,N_11169);
and U12511 (N_12511,N_11015,N_11085);
and U12512 (N_12512,N_11393,N_11701);
nand U12513 (N_12513,N_11668,N_11228);
and U12514 (N_12514,N_11964,N_11396);
nor U12515 (N_12515,N_11363,N_11506);
and U12516 (N_12516,N_11718,N_11816);
nand U12517 (N_12517,N_11691,N_11859);
nand U12518 (N_12518,N_11985,N_11429);
nand U12519 (N_12519,N_11073,N_11972);
xor U12520 (N_12520,N_11642,N_11518);
nand U12521 (N_12521,N_11810,N_11274);
or U12522 (N_12522,N_11609,N_11988);
nor U12523 (N_12523,N_11095,N_11167);
and U12524 (N_12524,N_11824,N_11316);
or U12525 (N_12525,N_11690,N_11954);
nand U12526 (N_12526,N_11914,N_11214);
or U12527 (N_12527,N_11862,N_11970);
or U12528 (N_12528,N_11965,N_11827);
nor U12529 (N_12529,N_11996,N_11951);
nor U12530 (N_12530,N_11886,N_11262);
or U12531 (N_12531,N_11453,N_11399);
or U12532 (N_12532,N_11249,N_11647);
nand U12533 (N_12533,N_11155,N_11820);
or U12534 (N_12534,N_11997,N_11343);
and U12535 (N_12535,N_11481,N_11084);
nand U12536 (N_12536,N_11940,N_11750);
xnor U12537 (N_12537,N_11056,N_11814);
xnor U12538 (N_12538,N_11138,N_11237);
or U12539 (N_12539,N_11876,N_11328);
nand U12540 (N_12540,N_11206,N_11359);
and U12541 (N_12541,N_11879,N_11476);
and U12542 (N_12542,N_11072,N_11078);
or U12543 (N_12543,N_11528,N_11144);
and U12544 (N_12544,N_11465,N_11497);
or U12545 (N_12545,N_11997,N_11282);
nor U12546 (N_12546,N_11741,N_11933);
or U12547 (N_12547,N_11919,N_11446);
and U12548 (N_12548,N_11070,N_11423);
nor U12549 (N_12549,N_11266,N_11829);
and U12550 (N_12550,N_11128,N_11416);
nand U12551 (N_12551,N_11106,N_11803);
nor U12552 (N_12552,N_11001,N_11400);
and U12553 (N_12553,N_11692,N_11538);
nor U12554 (N_12554,N_11010,N_11441);
or U12555 (N_12555,N_11508,N_11376);
xor U12556 (N_12556,N_11865,N_11809);
nand U12557 (N_12557,N_11481,N_11009);
and U12558 (N_12558,N_11970,N_11465);
nand U12559 (N_12559,N_11263,N_11642);
nor U12560 (N_12560,N_11122,N_11604);
or U12561 (N_12561,N_11443,N_11621);
or U12562 (N_12562,N_11157,N_11934);
nand U12563 (N_12563,N_11279,N_11828);
nor U12564 (N_12564,N_11136,N_11684);
nor U12565 (N_12565,N_11575,N_11340);
xor U12566 (N_12566,N_11458,N_11325);
or U12567 (N_12567,N_11989,N_11757);
and U12568 (N_12568,N_11588,N_11031);
nand U12569 (N_12569,N_11759,N_11095);
and U12570 (N_12570,N_11953,N_11266);
and U12571 (N_12571,N_11159,N_11945);
nor U12572 (N_12572,N_11584,N_11701);
xor U12573 (N_12573,N_11078,N_11635);
nor U12574 (N_12574,N_11336,N_11981);
and U12575 (N_12575,N_11010,N_11560);
or U12576 (N_12576,N_11206,N_11985);
nand U12577 (N_12577,N_11877,N_11645);
and U12578 (N_12578,N_11448,N_11807);
or U12579 (N_12579,N_11395,N_11369);
and U12580 (N_12580,N_11134,N_11429);
and U12581 (N_12581,N_11177,N_11640);
or U12582 (N_12582,N_11594,N_11134);
nor U12583 (N_12583,N_11772,N_11136);
or U12584 (N_12584,N_11191,N_11965);
nand U12585 (N_12585,N_11582,N_11378);
or U12586 (N_12586,N_11680,N_11339);
or U12587 (N_12587,N_11428,N_11660);
nor U12588 (N_12588,N_11960,N_11551);
nor U12589 (N_12589,N_11323,N_11970);
or U12590 (N_12590,N_11663,N_11537);
or U12591 (N_12591,N_11990,N_11898);
and U12592 (N_12592,N_11938,N_11510);
nand U12593 (N_12593,N_11033,N_11160);
xor U12594 (N_12594,N_11453,N_11715);
or U12595 (N_12595,N_11512,N_11847);
xor U12596 (N_12596,N_11325,N_11695);
nand U12597 (N_12597,N_11287,N_11724);
and U12598 (N_12598,N_11878,N_11010);
or U12599 (N_12599,N_11189,N_11060);
or U12600 (N_12600,N_11221,N_11049);
nor U12601 (N_12601,N_11655,N_11973);
xnor U12602 (N_12602,N_11888,N_11336);
or U12603 (N_12603,N_11826,N_11392);
nor U12604 (N_12604,N_11393,N_11940);
xnor U12605 (N_12605,N_11418,N_11358);
nand U12606 (N_12606,N_11208,N_11974);
xor U12607 (N_12607,N_11442,N_11154);
or U12608 (N_12608,N_11798,N_11095);
or U12609 (N_12609,N_11517,N_11397);
or U12610 (N_12610,N_11058,N_11567);
nor U12611 (N_12611,N_11194,N_11813);
or U12612 (N_12612,N_11279,N_11906);
xnor U12613 (N_12613,N_11985,N_11516);
nor U12614 (N_12614,N_11976,N_11038);
nand U12615 (N_12615,N_11395,N_11646);
nand U12616 (N_12616,N_11293,N_11093);
xor U12617 (N_12617,N_11143,N_11868);
nand U12618 (N_12618,N_11261,N_11668);
nand U12619 (N_12619,N_11360,N_11803);
or U12620 (N_12620,N_11487,N_11162);
nand U12621 (N_12621,N_11968,N_11910);
nor U12622 (N_12622,N_11846,N_11043);
or U12623 (N_12623,N_11148,N_11624);
nand U12624 (N_12624,N_11212,N_11314);
or U12625 (N_12625,N_11078,N_11695);
or U12626 (N_12626,N_11880,N_11156);
nor U12627 (N_12627,N_11490,N_11765);
or U12628 (N_12628,N_11750,N_11819);
xnor U12629 (N_12629,N_11348,N_11230);
or U12630 (N_12630,N_11098,N_11599);
nand U12631 (N_12631,N_11666,N_11523);
or U12632 (N_12632,N_11217,N_11563);
and U12633 (N_12633,N_11630,N_11824);
nand U12634 (N_12634,N_11659,N_11571);
or U12635 (N_12635,N_11463,N_11015);
and U12636 (N_12636,N_11625,N_11660);
or U12637 (N_12637,N_11208,N_11536);
nor U12638 (N_12638,N_11980,N_11954);
or U12639 (N_12639,N_11203,N_11908);
and U12640 (N_12640,N_11509,N_11561);
nor U12641 (N_12641,N_11587,N_11531);
and U12642 (N_12642,N_11587,N_11590);
and U12643 (N_12643,N_11023,N_11063);
xor U12644 (N_12644,N_11421,N_11247);
nand U12645 (N_12645,N_11787,N_11186);
or U12646 (N_12646,N_11908,N_11524);
or U12647 (N_12647,N_11887,N_11491);
nor U12648 (N_12648,N_11163,N_11712);
nand U12649 (N_12649,N_11104,N_11540);
nor U12650 (N_12650,N_11457,N_11356);
or U12651 (N_12651,N_11095,N_11209);
and U12652 (N_12652,N_11621,N_11247);
or U12653 (N_12653,N_11257,N_11533);
and U12654 (N_12654,N_11020,N_11833);
xnor U12655 (N_12655,N_11347,N_11007);
or U12656 (N_12656,N_11185,N_11934);
xnor U12657 (N_12657,N_11173,N_11973);
or U12658 (N_12658,N_11885,N_11200);
or U12659 (N_12659,N_11633,N_11239);
and U12660 (N_12660,N_11063,N_11354);
or U12661 (N_12661,N_11615,N_11959);
and U12662 (N_12662,N_11873,N_11677);
nor U12663 (N_12663,N_11641,N_11514);
nand U12664 (N_12664,N_11878,N_11122);
or U12665 (N_12665,N_11865,N_11607);
and U12666 (N_12666,N_11807,N_11022);
and U12667 (N_12667,N_11290,N_11929);
nand U12668 (N_12668,N_11100,N_11718);
or U12669 (N_12669,N_11242,N_11633);
or U12670 (N_12670,N_11766,N_11479);
nor U12671 (N_12671,N_11076,N_11245);
xnor U12672 (N_12672,N_11661,N_11617);
xnor U12673 (N_12673,N_11447,N_11813);
or U12674 (N_12674,N_11649,N_11479);
or U12675 (N_12675,N_11068,N_11196);
nor U12676 (N_12676,N_11622,N_11776);
nand U12677 (N_12677,N_11160,N_11584);
nand U12678 (N_12678,N_11400,N_11037);
and U12679 (N_12679,N_11179,N_11063);
nand U12680 (N_12680,N_11939,N_11838);
and U12681 (N_12681,N_11842,N_11386);
or U12682 (N_12682,N_11488,N_11243);
nor U12683 (N_12683,N_11723,N_11941);
nor U12684 (N_12684,N_11369,N_11525);
and U12685 (N_12685,N_11670,N_11009);
nor U12686 (N_12686,N_11903,N_11075);
nand U12687 (N_12687,N_11127,N_11852);
and U12688 (N_12688,N_11370,N_11938);
nor U12689 (N_12689,N_11783,N_11814);
or U12690 (N_12690,N_11488,N_11527);
and U12691 (N_12691,N_11749,N_11689);
nor U12692 (N_12692,N_11117,N_11110);
nand U12693 (N_12693,N_11706,N_11653);
and U12694 (N_12694,N_11645,N_11608);
or U12695 (N_12695,N_11819,N_11084);
nor U12696 (N_12696,N_11188,N_11166);
or U12697 (N_12697,N_11876,N_11914);
nor U12698 (N_12698,N_11699,N_11494);
or U12699 (N_12699,N_11521,N_11178);
and U12700 (N_12700,N_11240,N_11508);
or U12701 (N_12701,N_11267,N_11049);
xnor U12702 (N_12702,N_11462,N_11014);
nor U12703 (N_12703,N_11485,N_11801);
nand U12704 (N_12704,N_11517,N_11321);
or U12705 (N_12705,N_11083,N_11074);
xnor U12706 (N_12706,N_11516,N_11909);
nor U12707 (N_12707,N_11860,N_11907);
and U12708 (N_12708,N_11521,N_11088);
and U12709 (N_12709,N_11721,N_11136);
xnor U12710 (N_12710,N_11101,N_11263);
xnor U12711 (N_12711,N_11439,N_11320);
nor U12712 (N_12712,N_11266,N_11235);
nor U12713 (N_12713,N_11884,N_11252);
and U12714 (N_12714,N_11850,N_11335);
nor U12715 (N_12715,N_11449,N_11663);
nor U12716 (N_12716,N_11892,N_11821);
nor U12717 (N_12717,N_11218,N_11350);
nand U12718 (N_12718,N_11173,N_11482);
nand U12719 (N_12719,N_11169,N_11519);
or U12720 (N_12720,N_11390,N_11519);
and U12721 (N_12721,N_11967,N_11990);
nor U12722 (N_12722,N_11960,N_11441);
and U12723 (N_12723,N_11916,N_11576);
nand U12724 (N_12724,N_11846,N_11453);
xor U12725 (N_12725,N_11826,N_11500);
nor U12726 (N_12726,N_11713,N_11860);
nor U12727 (N_12727,N_11055,N_11384);
and U12728 (N_12728,N_11178,N_11719);
or U12729 (N_12729,N_11770,N_11941);
nor U12730 (N_12730,N_11962,N_11865);
and U12731 (N_12731,N_11886,N_11632);
or U12732 (N_12732,N_11605,N_11967);
or U12733 (N_12733,N_11295,N_11660);
nor U12734 (N_12734,N_11835,N_11338);
and U12735 (N_12735,N_11810,N_11302);
or U12736 (N_12736,N_11405,N_11367);
or U12737 (N_12737,N_11117,N_11193);
nor U12738 (N_12738,N_11455,N_11797);
or U12739 (N_12739,N_11643,N_11146);
nand U12740 (N_12740,N_11225,N_11709);
and U12741 (N_12741,N_11024,N_11271);
xnor U12742 (N_12742,N_11706,N_11811);
and U12743 (N_12743,N_11613,N_11619);
nand U12744 (N_12744,N_11273,N_11845);
nor U12745 (N_12745,N_11312,N_11404);
xor U12746 (N_12746,N_11026,N_11946);
xnor U12747 (N_12747,N_11143,N_11218);
nand U12748 (N_12748,N_11145,N_11101);
nor U12749 (N_12749,N_11236,N_11366);
nand U12750 (N_12750,N_11932,N_11314);
or U12751 (N_12751,N_11798,N_11278);
or U12752 (N_12752,N_11039,N_11282);
xor U12753 (N_12753,N_11916,N_11885);
nand U12754 (N_12754,N_11369,N_11575);
nor U12755 (N_12755,N_11988,N_11216);
xnor U12756 (N_12756,N_11734,N_11055);
nor U12757 (N_12757,N_11506,N_11059);
nand U12758 (N_12758,N_11403,N_11770);
nand U12759 (N_12759,N_11964,N_11204);
nor U12760 (N_12760,N_11574,N_11634);
nand U12761 (N_12761,N_11386,N_11107);
or U12762 (N_12762,N_11018,N_11815);
xnor U12763 (N_12763,N_11775,N_11830);
and U12764 (N_12764,N_11683,N_11877);
nor U12765 (N_12765,N_11829,N_11296);
nor U12766 (N_12766,N_11778,N_11568);
and U12767 (N_12767,N_11843,N_11233);
and U12768 (N_12768,N_11382,N_11657);
nor U12769 (N_12769,N_11420,N_11368);
nand U12770 (N_12770,N_11220,N_11153);
or U12771 (N_12771,N_11058,N_11516);
or U12772 (N_12772,N_11599,N_11427);
or U12773 (N_12773,N_11413,N_11400);
and U12774 (N_12774,N_11926,N_11974);
or U12775 (N_12775,N_11238,N_11197);
nor U12776 (N_12776,N_11485,N_11888);
or U12777 (N_12777,N_11344,N_11891);
nand U12778 (N_12778,N_11687,N_11566);
and U12779 (N_12779,N_11331,N_11609);
nand U12780 (N_12780,N_11880,N_11482);
xor U12781 (N_12781,N_11636,N_11304);
xnor U12782 (N_12782,N_11045,N_11945);
and U12783 (N_12783,N_11584,N_11700);
or U12784 (N_12784,N_11421,N_11360);
or U12785 (N_12785,N_11990,N_11391);
or U12786 (N_12786,N_11152,N_11389);
xor U12787 (N_12787,N_11454,N_11074);
or U12788 (N_12788,N_11150,N_11135);
nor U12789 (N_12789,N_11986,N_11201);
nand U12790 (N_12790,N_11520,N_11501);
nand U12791 (N_12791,N_11989,N_11303);
xor U12792 (N_12792,N_11631,N_11474);
and U12793 (N_12793,N_11698,N_11227);
and U12794 (N_12794,N_11977,N_11984);
and U12795 (N_12795,N_11794,N_11368);
or U12796 (N_12796,N_11400,N_11144);
and U12797 (N_12797,N_11368,N_11567);
or U12798 (N_12798,N_11212,N_11227);
nand U12799 (N_12799,N_11430,N_11393);
or U12800 (N_12800,N_11076,N_11961);
and U12801 (N_12801,N_11869,N_11036);
nand U12802 (N_12802,N_11373,N_11766);
or U12803 (N_12803,N_11402,N_11318);
nor U12804 (N_12804,N_11838,N_11670);
or U12805 (N_12805,N_11844,N_11025);
or U12806 (N_12806,N_11637,N_11523);
and U12807 (N_12807,N_11892,N_11304);
nand U12808 (N_12808,N_11681,N_11492);
nor U12809 (N_12809,N_11700,N_11868);
and U12810 (N_12810,N_11568,N_11642);
nor U12811 (N_12811,N_11002,N_11542);
and U12812 (N_12812,N_11685,N_11329);
and U12813 (N_12813,N_11309,N_11463);
nand U12814 (N_12814,N_11962,N_11391);
xnor U12815 (N_12815,N_11065,N_11336);
xor U12816 (N_12816,N_11267,N_11079);
nor U12817 (N_12817,N_11873,N_11634);
and U12818 (N_12818,N_11157,N_11632);
nor U12819 (N_12819,N_11826,N_11164);
nor U12820 (N_12820,N_11876,N_11165);
and U12821 (N_12821,N_11602,N_11005);
nor U12822 (N_12822,N_11931,N_11503);
or U12823 (N_12823,N_11797,N_11597);
nand U12824 (N_12824,N_11689,N_11932);
nor U12825 (N_12825,N_11287,N_11650);
and U12826 (N_12826,N_11460,N_11198);
nand U12827 (N_12827,N_11070,N_11964);
xor U12828 (N_12828,N_11985,N_11480);
and U12829 (N_12829,N_11205,N_11843);
and U12830 (N_12830,N_11626,N_11056);
nand U12831 (N_12831,N_11891,N_11616);
and U12832 (N_12832,N_11651,N_11563);
nand U12833 (N_12833,N_11589,N_11047);
and U12834 (N_12834,N_11003,N_11252);
nor U12835 (N_12835,N_11343,N_11386);
nand U12836 (N_12836,N_11578,N_11337);
nor U12837 (N_12837,N_11631,N_11965);
or U12838 (N_12838,N_11284,N_11967);
and U12839 (N_12839,N_11713,N_11388);
nand U12840 (N_12840,N_11436,N_11637);
and U12841 (N_12841,N_11339,N_11865);
xnor U12842 (N_12842,N_11507,N_11495);
nand U12843 (N_12843,N_11539,N_11312);
and U12844 (N_12844,N_11833,N_11809);
xor U12845 (N_12845,N_11855,N_11616);
and U12846 (N_12846,N_11851,N_11943);
and U12847 (N_12847,N_11035,N_11341);
nand U12848 (N_12848,N_11036,N_11398);
xnor U12849 (N_12849,N_11031,N_11555);
or U12850 (N_12850,N_11581,N_11662);
or U12851 (N_12851,N_11386,N_11750);
nor U12852 (N_12852,N_11878,N_11559);
nor U12853 (N_12853,N_11543,N_11375);
or U12854 (N_12854,N_11437,N_11798);
nand U12855 (N_12855,N_11662,N_11739);
or U12856 (N_12856,N_11078,N_11934);
and U12857 (N_12857,N_11897,N_11025);
nand U12858 (N_12858,N_11830,N_11786);
and U12859 (N_12859,N_11219,N_11189);
and U12860 (N_12860,N_11149,N_11648);
or U12861 (N_12861,N_11099,N_11844);
nand U12862 (N_12862,N_11795,N_11547);
or U12863 (N_12863,N_11061,N_11154);
nand U12864 (N_12864,N_11831,N_11769);
nand U12865 (N_12865,N_11807,N_11385);
nor U12866 (N_12866,N_11265,N_11852);
nand U12867 (N_12867,N_11407,N_11678);
nand U12868 (N_12868,N_11908,N_11356);
and U12869 (N_12869,N_11084,N_11016);
xnor U12870 (N_12870,N_11520,N_11659);
nor U12871 (N_12871,N_11370,N_11434);
xnor U12872 (N_12872,N_11855,N_11691);
or U12873 (N_12873,N_11155,N_11156);
nor U12874 (N_12874,N_11966,N_11453);
nor U12875 (N_12875,N_11719,N_11683);
and U12876 (N_12876,N_11753,N_11151);
xor U12877 (N_12877,N_11412,N_11977);
and U12878 (N_12878,N_11147,N_11853);
and U12879 (N_12879,N_11489,N_11005);
and U12880 (N_12880,N_11372,N_11255);
or U12881 (N_12881,N_11287,N_11554);
nor U12882 (N_12882,N_11888,N_11087);
nand U12883 (N_12883,N_11221,N_11762);
and U12884 (N_12884,N_11896,N_11066);
or U12885 (N_12885,N_11046,N_11056);
nand U12886 (N_12886,N_11602,N_11051);
and U12887 (N_12887,N_11524,N_11309);
and U12888 (N_12888,N_11620,N_11905);
nand U12889 (N_12889,N_11442,N_11495);
xnor U12890 (N_12890,N_11538,N_11510);
and U12891 (N_12891,N_11370,N_11235);
and U12892 (N_12892,N_11933,N_11846);
or U12893 (N_12893,N_11615,N_11390);
nand U12894 (N_12894,N_11551,N_11582);
and U12895 (N_12895,N_11106,N_11942);
or U12896 (N_12896,N_11556,N_11232);
nor U12897 (N_12897,N_11889,N_11836);
or U12898 (N_12898,N_11726,N_11986);
nor U12899 (N_12899,N_11496,N_11483);
or U12900 (N_12900,N_11425,N_11919);
nand U12901 (N_12901,N_11324,N_11563);
nand U12902 (N_12902,N_11028,N_11706);
nor U12903 (N_12903,N_11613,N_11922);
or U12904 (N_12904,N_11399,N_11633);
or U12905 (N_12905,N_11740,N_11057);
xnor U12906 (N_12906,N_11555,N_11319);
or U12907 (N_12907,N_11509,N_11912);
nor U12908 (N_12908,N_11937,N_11172);
or U12909 (N_12909,N_11775,N_11917);
nor U12910 (N_12910,N_11204,N_11951);
xnor U12911 (N_12911,N_11293,N_11815);
nor U12912 (N_12912,N_11707,N_11788);
or U12913 (N_12913,N_11091,N_11576);
or U12914 (N_12914,N_11836,N_11312);
nor U12915 (N_12915,N_11400,N_11234);
and U12916 (N_12916,N_11619,N_11641);
nand U12917 (N_12917,N_11483,N_11819);
nor U12918 (N_12918,N_11443,N_11617);
or U12919 (N_12919,N_11867,N_11091);
or U12920 (N_12920,N_11332,N_11156);
nand U12921 (N_12921,N_11767,N_11764);
and U12922 (N_12922,N_11303,N_11477);
or U12923 (N_12923,N_11315,N_11719);
nand U12924 (N_12924,N_11434,N_11432);
or U12925 (N_12925,N_11949,N_11921);
and U12926 (N_12926,N_11897,N_11892);
nand U12927 (N_12927,N_11772,N_11358);
or U12928 (N_12928,N_11605,N_11280);
or U12929 (N_12929,N_11803,N_11881);
or U12930 (N_12930,N_11780,N_11617);
or U12931 (N_12931,N_11016,N_11517);
or U12932 (N_12932,N_11741,N_11181);
nor U12933 (N_12933,N_11770,N_11590);
and U12934 (N_12934,N_11598,N_11327);
nor U12935 (N_12935,N_11772,N_11932);
nand U12936 (N_12936,N_11799,N_11128);
or U12937 (N_12937,N_11394,N_11245);
nor U12938 (N_12938,N_11871,N_11156);
or U12939 (N_12939,N_11404,N_11684);
or U12940 (N_12940,N_11120,N_11679);
nor U12941 (N_12941,N_11770,N_11988);
nand U12942 (N_12942,N_11921,N_11035);
nor U12943 (N_12943,N_11833,N_11613);
nor U12944 (N_12944,N_11902,N_11384);
or U12945 (N_12945,N_11717,N_11556);
and U12946 (N_12946,N_11038,N_11718);
nand U12947 (N_12947,N_11417,N_11354);
and U12948 (N_12948,N_11898,N_11015);
nand U12949 (N_12949,N_11619,N_11634);
or U12950 (N_12950,N_11478,N_11560);
and U12951 (N_12951,N_11019,N_11788);
and U12952 (N_12952,N_11099,N_11896);
xor U12953 (N_12953,N_11634,N_11867);
nand U12954 (N_12954,N_11654,N_11811);
or U12955 (N_12955,N_11581,N_11939);
and U12956 (N_12956,N_11998,N_11154);
and U12957 (N_12957,N_11349,N_11344);
or U12958 (N_12958,N_11508,N_11409);
or U12959 (N_12959,N_11589,N_11176);
and U12960 (N_12960,N_11369,N_11806);
and U12961 (N_12961,N_11969,N_11700);
nand U12962 (N_12962,N_11740,N_11945);
nor U12963 (N_12963,N_11171,N_11415);
nor U12964 (N_12964,N_11653,N_11789);
nand U12965 (N_12965,N_11319,N_11937);
nand U12966 (N_12966,N_11265,N_11999);
and U12967 (N_12967,N_11849,N_11353);
nor U12968 (N_12968,N_11147,N_11893);
and U12969 (N_12969,N_11867,N_11120);
nand U12970 (N_12970,N_11161,N_11754);
xor U12971 (N_12971,N_11817,N_11488);
xor U12972 (N_12972,N_11352,N_11778);
or U12973 (N_12973,N_11772,N_11957);
nand U12974 (N_12974,N_11554,N_11272);
nor U12975 (N_12975,N_11298,N_11867);
and U12976 (N_12976,N_11576,N_11614);
nand U12977 (N_12977,N_11465,N_11390);
or U12978 (N_12978,N_11820,N_11229);
nand U12979 (N_12979,N_11184,N_11637);
or U12980 (N_12980,N_11543,N_11596);
and U12981 (N_12981,N_11108,N_11136);
and U12982 (N_12982,N_11090,N_11364);
or U12983 (N_12983,N_11982,N_11005);
nor U12984 (N_12984,N_11982,N_11839);
or U12985 (N_12985,N_11981,N_11506);
and U12986 (N_12986,N_11743,N_11500);
nor U12987 (N_12987,N_11193,N_11923);
xor U12988 (N_12988,N_11131,N_11791);
nor U12989 (N_12989,N_11913,N_11486);
and U12990 (N_12990,N_11827,N_11843);
xnor U12991 (N_12991,N_11886,N_11656);
and U12992 (N_12992,N_11033,N_11646);
nand U12993 (N_12993,N_11225,N_11023);
and U12994 (N_12994,N_11047,N_11092);
nor U12995 (N_12995,N_11310,N_11212);
nand U12996 (N_12996,N_11406,N_11733);
and U12997 (N_12997,N_11435,N_11536);
or U12998 (N_12998,N_11649,N_11609);
and U12999 (N_12999,N_11026,N_11698);
and U13000 (N_13000,N_12433,N_12081);
and U13001 (N_13001,N_12037,N_12427);
or U13002 (N_13002,N_12118,N_12809);
nand U13003 (N_13003,N_12766,N_12194);
xor U13004 (N_13004,N_12016,N_12314);
and U13005 (N_13005,N_12483,N_12830);
or U13006 (N_13006,N_12519,N_12922);
and U13007 (N_13007,N_12499,N_12681);
or U13008 (N_13008,N_12803,N_12846);
nand U13009 (N_13009,N_12182,N_12914);
and U13010 (N_13010,N_12690,N_12890);
nand U13011 (N_13011,N_12812,N_12872);
nor U13012 (N_13012,N_12304,N_12878);
nand U13013 (N_13013,N_12357,N_12250);
nor U13014 (N_13014,N_12783,N_12356);
nor U13015 (N_13015,N_12578,N_12736);
and U13016 (N_13016,N_12436,N_12006);
and U13017 (N_13017,N_12232,N_12237);
or U13018 (N_13018,N_12720,N_12571);
nor U13019 (N_13019,N_12343,N_12033);
or U13020 (N_13020,N_12195,N_12397);
or U13021 (N_13021,N_12149,N_12455);
or U13022 (N_13022,N_12818,N_12177);
and U13023 (N_13023,N_12340,N_12497);
or U13024 (N_13024,N_12539,N_12724);
and U13025 (N_13025,N_12695,N_12341);
xnor U13026 (N_13026,N_12053,N_12932);
nor U13027 (N_13027,N_12869,N_12413);
nand U13028 (N_13028,N_12288,N_12209);
xor U13029 (N_13029,N_12089,N_12036);
nor U13030 (N_13030,N_12208,N_12793);
and U13031 (N_13031,N_12800,N_12073);
nor U13032 (N_13032,N_12320,N_12535);
or U13033 (N_13033,N_12408,N_12333);
and U13034 (N_13034,N_12834,N_12757);
nor U13035 (N_13035,N_12911,N_12502);
nor U13036 (N_13036,N_12190,N_12882);
or U13037 (N_13037,N_12284,N_12755);
or U13038 (N_13038,N_12512,N_12920);
nand U13039 (N_13039,N_12907,N_12184);
nand U13040 (N_13040,N_12490,N_12966);
nand U13041 (N_13041,N_12582,N_12739);
nand U13042 (N_13042,N_12127,N_12046);
and U13043 (N_13043,N_12012,N_12857);
nand U13044 (N_13044,N_12405,N_12646);
nor U13045 (N_13045,N_12521,N_12874);
or U13046 (N_13046,N_12344,N_12167);
nand U13047 (N_13047,N_12370,N_12327);
nand U13048 (N_13048,N_12400,N_12431);
or U13049 (N_13049,N_12558,N_12700);
and U13050 (N_13050,N_12530,N_12509);
and U13051 (N_13051,N_12699,N_12640);
nor U13052 (N_13052,N_12226,N_12396);
and U13053 (N_13053,N_12662,N_12274);
or U13054 (N_13054,N_12139,N_12569);
and U13055 (N_13055,N_12454,N_12929);
and U13056 (N_13056,N_12557,N_12321);
or U13057 (N_13057,N_12366,N_12363);
or U13058 (N_13058,N_12084,N_12547);
nor U13059 (N_13059,N_12712,N_12600);
nand U13060 (N_13060,N_12511,N_12166);
xor U13061 (N_13061,N_12948,N_12076);
nor U13062 (N_13062,N_12031,N_12898);
nor U13063 (N_13063,N_12132,N_12923);
xor U13064 (N_13064,N_12187,N_12605);
and U13065 (N_13065,N_12214,N_12252);
and U13066 (N_13066,N_12691,N_12832);
and U13067 (N_13067,N_12633,N_12204);
nor U13068 (N_13068,N_12376,N_12587);
xor U13069 (N_13069,N_12174,N_12771);
nor U13070 (N_13070,N_12611,N_12245);
xnor U13071 (N_13071,N_12030,N_12723);
nand U13072 (N_13072,N_12022,N_12768);
nand U13073 (N_13073,N_12975,N_12667);
nand U13074 (N_13074,N_12150,N_12589);
or U13075 (N_13075,N_12630,N_12570);
nand U13076 (N_13076,N_12153,N_12399);
xnor U13077 (N_13077,N_12129,N_12641);
nor U13078 (N_13078,N_12824,N_12835);
and U13079 (N_13079,N_12109,N_12625);
nor U13080 (N_13080,N_12991,N_12410);
nand U13081 (N_13081,N_12126,N_12688);
nor U13082 (N_13082,N_12541,N_12648);
and U13083 (N_13083,N_12192,N_12220);
and U13084 (N_13084,N_12685,N_12585);
and U13085 (N_13085,N_12336,N_12961);
nor U13086 (N_13086,N_12718,N_12168);
and U13087 (N_13087,N_12934,N_12442);
or U13088 (N_13088,N_12063,N_12988);
and U13089 (N_13089,N_12735,N_12425);
or U13090 (N_13090,N_12249,N_12488);
and U13091 (N_13091,N_12597,N_12360);
or U13092 (N_13092,N_12540,N_12782);
xnor U13093 (N_13093,N_12849,N_12559);
nor U13094 (N_13094,N_12402,N_12075);
or U13095 (N_13095,N_12562,N_12698);
and U13096 (N_13096,N_12337,N_12889);
or U13097 (N_13097,N_12577,N_12877);
and U13098 (N_13098,N_12114,N_12924);
and U13099 (N_13099,N_12394,N_12576);
and U13100 (N_13100,N_12329,N_12574);
and U13101 (N_13101,N_12420,N_12164);
or U13102 (N_13102,N_12467,N_12623);
nor U13103 (N_13103,N_12430,N_12811);
nor U13104 (N_13104,N_12382,N_12631);
nor U13105 (N_13105,N_12026,N_12950);
and U13106 (N_13106,N_12958,N_12134);
or U13107 (N_13107,N_12271,N_12504);
nor U13108 (N_13108,N_12279,N_12044);
or U13109 (N_13109,N_12444,N_12784);
or U13110 (N_13110,N_12886,N_12138);
or U13111 (N_13111,N_12905,N_12959);
nand U13112 (N_13112,N_12638,N_12916);
and U13113 (N_13113,N_12310,N_12203);
or U13114 (N_13114,N_12115,N_12806);
or U13115 (N_13115,N_12738,N_12759);
nand U13116 (N_13116,N_12668,N_12254);
or U13117 (N_13117,N_12014,N_12353);
nor U13118 (N_13118,N_12939,N_12871);
nor U13119 (N_13119,N_12732,N_12428);
or U13120 (N_13120,N_12302,N_12722);
nand U13121 (N_13121,N_12346,N_12101);
or U13122 (N_13122,N_12848,N_12095);
and U13123 (N_13123,N_12477,N_12915);
xnor U13124 (N_13124,N_12642,N_12584);
nor U13125 (N_13125,N_12435,N_12181);
xnor U13126 (N_13126,N_12072,N_12687);
nand U13127 (N_13127,N_12349,N_12083);
and U13128 (N_13128,N_12813,N_12575);
nand U13129 (N_13129,N_12144,N_12035);
nor U13130 (N_13130,N_12615,N_12224);
or U13131 (N_13131,N_12566,N_12946);
or U13132 (N_13132,N_12248,N_12270);
nor U13133 (N_13133,N_12554,N_12380);
nand U13134 (N_13134,N_12120,N_12219);
and U13135 (N_13135,N_12676,N_12828);
or U13136 (N_13136,N_12749,N_12173);
and U13137 (N_13137,N_12021,N_12761);
nand U13138 (N_13138,N_12839,N_12034);
and U13139 (N_13139,N_12125,N_12008);
nor U13140 (N_13140,N_12263,N_12515);
nor U13141 (N_13141,N_12378,N_12289);
nand U13142 (N_13142,N_12419,N_12309);
or U13143 (N_13143,N_12056,N_12969);
or U13144 (N_13144,N_12826,N_12485);
or U13145 (N_13145,N_12240,N_12403);
and U13146 (N_13146,N_12269,N_12185);
and U13147 (N_13147,N_12422,N_12381);
or U13148 (N_13148,N_12737,N_12170);
and U13149 (N_13149,N_12594,N_12217);
xnor U13150 (N_13150,N_12949,N_12017);
and U13151 (N_13151,N_12358,N_12205);
and U13152 (N_13152,N_12618,N_12437);
xnor U13153 (N_13153,N_12029,N_12465);
xor U13154 (N_13154,N_12155,N_12473);
nand U13155 (N_13155,N_12086,N_12567);
nor U13156 (N_13156,N_12677,N_12598);
nand U13157 (N_13157,N_12710,N_12308);
or U13158 (N_13158,N_12891,N_12156);
nand U13159 (N_13159,N_12316,N_12384);
nand U13160 (N_13160,N_12645,N_12788);
or U13161 (N_13161,N_12550,N_12734);
xor U13162 (N_13162,N_12831,N_12227);
nand U13163 (N_13163,N_12019,N_12798);
nand U13164 (N_13164,N_12262,N_12108);
and U13165 (N_13165,N_12507,N_12319);
or U13166 (N_13166,N_12852,N_12171);
and U13167 (N_13167,N_12816,N_12441);
and U13168 (N_13168,N_12944,N_12315);
nand U13169 (N_13169,N_12627,N_12367);
nand U13170 (N_13170,N_12466,N_12280);
nand U13171 (N_13171,N_12368,N_12267);
nand U13172 (N_13172,N_12434,N_12534);
or U13173 (N_13173,N_12635,N_12912);
nor U13174 (N_13174,N_12626,N_12951);
nor U13175 (N_13175,N_12657,N_12801);
or U13176 (N_13176,N_12649,N_12080);
nand U13177 (N_13177,N_12324,N_12840);
nand U13178 (N_13178,N_12896,N_12746);
nor U13179 (N_13179,N_12440,N_12588);
nand U13180 (N_13180,N_12556,N_12930);
nor U13181 (N_13181,N_12258,N_12836);
and U13182 (N_13182,N_12921,N_12706);
nand U13183 (N_13183,N_12078,N_12514);
nand U13184 (N_13184,N_12365,N_12837);
or U13185 (N_13185,N_12062,N_12471);
nor U13186 (N_13186,N_12364,N_12955);
and U13187 (N_13187,N_12850,N_12157);
xnor U13188 (N_13188,N_12389,N_12751);
or U13189 (N_13189,N_12404,N_12526);
xor U13190 (N_13190,N_12462,N_12350);
nor U13191 (N_13191,N_12945,N_12449);
nand U13192 (N_13192,N_12867,N_12145);
and U13193 (N_13193,N_12985,N_12235);
and U13194 (N_13194,N_12953,N_12387);
and U13195 (N_13195,N_12406,N_12842);
nor U13196 (N_13196,N_12496,N_12439);
nor U13197 (N_13197,N_12716,N_12023);
nand U13198 (N_13198,N_12461,N_12229);
and U13199 (N_13199,N_12742,N_12213);
nand U13200 (N_13200,N_12906,N_12133);
or U13201 (N_13201,N_12369,N_12464);
and U13202 (N_13202,N_12978,N_12954);
or U13203 (N_13203,N_12815,N_12272);
and U13204 (N_13204,N_12814,N_12172);
xor U13205 (N_13205,N_12851,N_12457);
nor U13206 (N_13206,N_12298,N_12620);
and U13207 (N_13207,N_12225,N_12656);
and U13208 (N_13208,N_12342,N_12128);
nor U13209 (N_13209,N_12981,N_12257);
nand U13210 (N_13210,N_12982,N_12234);
nor U13211 (N_13211,N_12317,N_12443);
nand U13212 (N_13212,N_12448,N_12158);
nor U13213 (N_13213,N_12838,N_12244);
and U13214 (N_13214,N_12450,N_12117);
xnor U13215 (N_13215,N_12102,N_12903);
and U13216 (N_13216,N_12762,N_12909);
and U13217 (N_13217,N_12242,N_12595);
nand U13218 (N_13218,N_12847,N_12992);
or U13219 (N_13219,N_12392,N_12061);
nand U13220 (N_13220,N_12841,N_12613);
nor U13221 (N_13221,N_12007,N_12100);
or U13222 (N_13222,N_12077,N_12305);
nand U13223 (N_13223,N_12051,N_12962);
nand U13224 (N_13224,N_12074,N_12282);
and U13225 (N_13225,N_12050,N_12609);
nor U13226 (N_13226,N_12199,N_12459);
and U13227 (N_13227,N_12326,N_12917);
and U13228 (N_13228,N_12565,N_12747);
and U13229 (N_13229,N_12794,N_12860);
nand U13230 (N_13230,N_12493,N_12154);
nand U13231 (N_13231,N_12372,N_12931);
and U13232 (N_13232,N_12658,N_12386);
or U13233 (N_13233,N_12058,N_12479);
nand U13234 (N_13234,N_12744,N_12480);
nand U13235 (N_13235,N_12470,N_12379);
nor U13236 (N_13236,N_12947,N_12418);
nand U13237 (N_13237,N_12347,N_12446);
or U13238 (N_13238,N_12278,N_12622);
nor U13239 (N_13239,N_12474,N_12866);
and U13240 (N_13240,N_12354,N_12426);
and U13241 (N_13241,N_12261,N_12659);
and U13242 (N_13242,N_12068,N_12231);
nand U13243 (N_13243,N_12322,N_12236);
and U13244 (N_13244,N_12990,N_12116);
xor U13245 (N_13245,N_12189,N_12335);
nand U13246 (N_13246,N_12111,N_12495);
nand U13247 (N_13247,N_12313,N_12087);
nor U13248 (N_13248,N_12518,N_12827);
nand U13249 (N_13249,N_12865,N_12482);
and U13250 (N_13250,N_12650,N_12876);
nor U13251 (N_13251,N_12501,N_12728);
nand U13252 (N_13252,N_12215,N_12707);
nor U13253 (N_13253,N_12241,N_12879);
nand U13254 (N_13254,N_12206,N_12296);
nand U13255 (N_13255,N_12573,N_12371);
or U13256 (N_13256,N_12748,N_12792);
and U13257 (N_13257,N_12286,N_12107);
and U13258 (N_13258,N_12750,N_12105);
nand U13259 (N_13259,N_12331,N_12445);
and U13260 (N_13260,N_12475,N_12047);
nand U13261 (N_13261,N_12892,N_12989);
nand U13262 (N_13262,N_12415,N_12655);
nor U13263 (N_13263,N_12974,N_12287);
nand U13264 (N_13264,N_12702,N_12745);
nor U13265 (N_13265,N_12020,N_12276);
or U13266 (N_13266,N_12264,N_12458);
nor U13267 (N_13267,N_12057,N_12028);
xnor U13268 (N_13268,N_12377,N_12819);
and U13269 (N_13269,N_12862,N_12469);
nor U13270 (N_13270,N_12726,N_12741);
nor U13271 (N_13271,N_12999,N_12596);
nor U13272 (N_13272,N_12591,N_12719);
or U13273 (N_13273,N_12001,N_12861);
nand U13274 (N_13274,N_12452,N_12683);
and U13275 (N_13275,N_12561,N_12277);
nand U13276 (N_13276,N_12523,N_12135);
or U13277 (N_13277,N_12979,N_12925);
or U13278 (N_13278,N_12715,N_12935);
nand U13279 (N_13279,N_12881,N_12663);
and U13280 (N_13280,N_12079,N_12936);
nor U13281 (N_13281,N_12928,N_12160);
nor U13282 (N_13282,N_12202,N_12524);
or U13283 (N_13283,N_12854,N_12665);
and U13284 (N_13284,N_12713,N_12634);
nor U13285 (N_13285,N_12612,N_12568);
nor U13286 (N_13286,N_12009,N_12243);
nand U13287 (N_13287,N_12619,N_12176);
nand U13288 (N_13288,N_12416,N_12294);
or U13289 (N_13289,N_12610,N_12251);
or U13290 (N_13290,N_12484,N_12345);
and U13291 (N_13291,N_12775,N_12532);
nand U13292 (N_13292,N_12636,N_12423);
xnor U13293 (N_13293,N_12555,N_12110);
nor U13294 (N_13294,N_12897,N_12082);
nand U13295 (N_13295,N_12478,N_12151);
or U13296 (N_13296,N_12772,N_12805);
and U13297 (N_13297,N_12789,N_12513);
nand U13298 (N_13298,N_12283,N_12822);
or U13299 (N_13299,N_12583,N_12614);
or U13300 (N_13300,N_12670,N_12290);
and U13301 (N_13301,N_12510,N_12752);
and U13302 (N_13302,N_12003,N_12303);
and U13303 (N_13303,N_12285,N_12884);
or U13304 (N_13304,N_12904,N_12863);
xor U13305 (N_13305,N_12338,N_12178);
nor U13306 (N_13306,N_12112,N_12845);
nand U13307 (N_13307,N_12045,N_12987);
xor U13308 (N_13308,N_12104,N_12186);
and U13309 (N_13309,N_12230,N_12143);
nor U13310 (N_13310,N_12301,N_12395);
nand U13311 (N_13311,N_12899,N_12391);
nor U13312 (N_13312,N_12407,N_12281);
or U13313 (N_13313,N_12093,N_12528);
nor U13314 (N_13314,N_12255,N_12980);
and U13315 (N_13315,N_12197,N_12639);
nand U13316 (N_13316,N_12743,N_12829);
nor U13317 (N_13317,N_12137,N_12411);
or U13318 (N_13318,N_12684,N_12875);
nand U13319 (N_13319,N_12956,N_12064);
xnor U13320 (N_13320,N_12498,N_12438);
xor U13321 (N_13321,N_12733,N_12682);
and U13322 (N_13322,N_12159,N_12791);
nand U13323 (N_13323,N_12268,N_12606);
nor U13324 (N_13324,N_12998,N_12069);
or U13325 (N_13325,N_12136,N_12628);
and U13326 (N_13326,N_12207,N_12808);
nor U13327 (N_13327,N_12508,N_12339);
nand U13328 (N_13328,N_12776,N_12894);
or U13329 (N_13329,N_12429,N_12858);
and U13330 (N_13330,N_12375,N_12993);
or U13331 (N_13331,N_12810,N_12537);
or U13332 (N_13332,N_12856,N_12853);
nand U13333 (N_13333,N_12629,N_12481);
xor U13334 (N_13334,N_12506,N_12604);
nand U13335 (N_13335,N_12674,N_12210);
and U13336 (N_13336,N_12373,N_12653);
nand U13337 (N_13337,N_12760,N_12844);
and U13338 (N_13338,N_12119,N_12560);
nand U13339 (N_13339,N_12223,N_12096);
and U13340 (N_13340,N_12088,N_12601);
nor U13341 (N_13341,N_12468,N_12753);
nor U13342 (N_13342,N_12703,N_12786);
or U13343 (N_13343,N_12727,N_12253);
and U13344 (N_13344,N_12533,N_12165);
nor U13345 (N_13345,N_12113,N_12553);
nor U13346 (N_13346,N_12312,N_12130);
or U13347 (N_13347,N_12259,N_12266);
or U13348 (N_13348,N_12586,N_12679);
nor U13349 (N_13349,N_12531,N_12632);
xnor U13350 (N_13350,N_12986,N_12579);
xnor U13351 (N_13351,N_12617,N_12997);
or U13352 (N_13352,N_12754,N_12901);
nor U13353 (N_13353,N_12599,N_12769);
and U13354 (N_13354,N_12147,N_12693);
or U13355 (N_13355,N_12233,N_12859);
and U13356 (N_13356,N_12486,N_12273);
nand U13357 (N_13357,N_12201,N_12005);
nand U13358 (N_13358,N_12306,N_12004);
and U13359 (N_13359,N_12054,N_12552);
xnor U13360 (N_13360,N_12895,N_12293);
nor U13361 (N_13361,N_12804,N_12409);
or U13362 (N_13362,N_12071,N_12692);
and U13363 (N_13363,N_12179,N_12142);
nor U13364 (N_13364,N_12359,N_12390);
or U13365 (N_13365,N_12218,N_12580);
nand U13366 (N_13366,N_12246,N_12581);
or U13367 (N_13367,N_12000,N_12374);
nand U13368 (N_13368,N_12542,N_12960);
or U13369 (N_13369,N_12548,N_12038);
nor U13370 (N_13370,N_12291,N_12977);
and U13371 (N_13371,N_12671,N_12527);
nand U13372 (N_13372,N_12694,N_12015);
nand U13373 (N_13373,N_12121,N_12018);
and U13374 (N_13374,N_12549,N_12183);
xor U13375 (N_13375,N_12770,N_12042);
nor U13376 (N_13376,N_12711,N_12654);
xnor U13377 (N_13377,N_12855,N_12424);
or U13378 (N_13378,N_12902,N_12651);
nand U13379 (N_13379,N_12680,N_12664);
or U13380 (N_13380,N_12807,N_12910);
nor U13381 (N_13381,N_12066,N_12059);
nand U13382 (N_13382,N_12968,N_12432);
or U13383 (N_13383,N_12417,N_12311);
and U13384 (N_13384,N_12708,N_12678);
or U13385 (N_13385,N_12672,N_12967);
and U13386 (N_13386,N_12476,N_12091);
or U13387 (N_13387,N_12334,N_12300);
or U13388 (N_13388,N_12146,N_12238);
or U13389 (N_13389,N_12756,N_12529);
and U13390 (N_13390,N_12228,N_12778);
and U13391 (N_13391,N_12608,N_12725);
xnor U13392 (N_13392,N_12065,N_12701);
nor U13393 (N_13393,N_12787,N_12052);
xor U13394 (N_13394,N_12603,N_12593);
and U13395 (N_13395,N_12996,N_12447);
nand U13396 (N_13396,N_12211,N_12048);
nand U13397 (N_13397,N_12323,N_12487);
or U13398 (N_13398,N_12880,N_12103);
nor U13399 (N_13399,N_12942,N_12351);
and U13400 (N_13400,N_12099,N_12758);
or U13401 (N_13401,N_12796,N_12212);
and U13402 (N_13402,N_12090,N_12297);
nor U13403 (N_13403,N_12729,N_12024);
nand U13404 (N_13404,N_12767,N_12401);
or U13405 (N_13405,N_12328,N_12010);
and U13406 (N_13406,N_12140,N_12607);
nor U13407 (N_13407,N_12572,N_12773);
nand U13408 (N_13408,N_12256,N_12491);
nand U13409 (N_13409,N_12870,N_12162);
nand U13410 (N_13410,N_12543,N_12673);
and U13411 (N_13411,N_12785,N_12325);
and U13412 (N_13412,N_12520,N_12002);
nand U13413 (N_13413,N_12131,N_12141);
and U13414 (N_13414,N_12721,N_12348);
and U13415 (N_13415,N_12175,N_12041);
or U13416 (N_13416,N_12123,N_12652);
nor U13417 (N_13417,N_12970,N_12873);
and U13418 (N_13418,N_12964,N_12952);
nor U13419 (N_13419,N_12221,N_12122);
and U13420 (N_13420,N_12193,N_12564);
nor U13421 (N_13421,N_12332,N_12456);
and U13422 (N_13422,N_12973,N_12709);
nand U13423 (N_13423,N_12544,N_12777);
and U13424 (N_13424,N_12799,N_12385);
nor U13425 (N_13425,N_12669,N_12522);
nand U13426 (N_13426,N_12013,N_12689);
xnor U13427 (N_13427,N_12355,N_12025);
nand U13428 (N_13428,N_12265,N_12503);
and U13429 (N_13429,N_12779,N_12994);
nand U13430 (N_13430,N_12505,N_12516);
nand U13431 (N_13431,N_12820,N_12864);
nand U13432 (N_13432,N_12927,N_12163);
nand U13433 (N_13433,N_12200,N_12152);
and U13434 (N_13434,N_12843,N_12887);
and U13435 (N_13435,N_12963,N_12463);
nand U13436 (N_13436,N_12191,N_12421);
and U13437 (N_13437,N_12098,N_12802);
or U13438 (N_13438,N_12647,N_12551);
xnor U13439 (N_13439,N_12971,N_12106);
and U13440 (N_13440,N_12092,N_12060);
and U13441 (N_13441,N_12027,N_12169);
nand U13442 (N_13442,N_12525,N_12032);
nand U13443 (N_13443,N_12918,N_12494);
nor U13444 (N_13444,N_12908,N_12976);
or U13445 (N_13445,N_12295,N_12885);
and U13446 (N_13446,N_12797,N_12995);
or U13447 (N_13447,N_12124,N_12460);
nor U13448 (N_13448,N_12790,N_12666);
or U13449 (N_13449,N_12740,N_12492);
nor U13450 (N_13450,N_12933,N_12957);
xnor U13451 (N_13451,N_12040,N_12868);
nor U13452 (N_13452,N_12913,N_12307);
and U13453 (N_13453,N_12765,N_12188);
nand U13454 (N_13454,N_12893,N_12602);
nor U13455 (N_13455,N_12055,N_12451);
xor U13456 (N_13456,N_12937,N_12616);
nand U13457 (N_13457,N_12299,N_12983);
and U13458 (N_13458,N_12453,N_12965);
and U13459 (N_13459,N_12067,N_12275);
or U13460 (N_13460,N_12239,N_12085);
or U13461 (N_13461,N_12043,N_12825);
xnor U13462 (N_13462,N_12592,N_12330);
and U13463 (N_13463,N_12414,N_12070);
nor U13464 (N_13464,N_12148,N_12517);
nand U13465 (N_13465,N_12546,N_12717);
nand U13466 (N_13466,N_12260,N_12731);
nand U13467 (N_13467,N_12938,N_12943);
or U13468 (N_13468,N_12196,N_12972);
and U13469 (N_13469,N_12318,N_12393);
nand U13470 (N_13470,N_12292,N_12536);
nor U13471 (N_13471,N_12180,N_12926);
xnor U13472 (N_13472,N_12198,N_12637);
xor U13473 (N_13473,N_12780,N_12590);
and U13474 (N_13474,N_12049,N_12388);
nand U13475 (N_13475,N_12714,N_12247);
nor U13476 (N_13476,N_12696,N_12472);
or U13477 (N_13477,N_12888,N_12624);
and U13478 (N_13478,N_12621,N_12704);
nor U13479 (N_13479,N_12763,N_12817);
nor U13480 (N_13480,N_12398,N_12361);
and U13481 (N_13481,N_12883,N_12489);
nand U13482 (N_13482,N_12222,N_12383);
nand U13483 (N_13483,N_12705,N_12940);
nor U13484 (N_13484,N_12352,N_12563);
nor U13485 (N_13485,N_12412,N_12545);
or U13486 (N_13486,N_12941,N_12161);
nor U13487 (N_13487,N_12362,N_12781);
nand U13488 (N_13488,N_12833,N_12823);
and U13489 (N_13489,N_12011,N_12661);
nand U13490 (N_13490,N_12538,N_12919);
nor U13491 (N_13491,N_12795,N_12900);
nand U13492 (N_13492,N_12643,N_12984);
nor U13493 (N_13493,N_12094,N_12764);
nand U13494 (N_13494,N_12686,N_12774);
nor U13495 (N_13495,N_12675,N_12644);
nor U13496 (N_13496,N_12730,N_12097);
nor U13497 (N_13497,N_12660,N_12500);
and U13498 (N_13498,N_12216,N_12821);
or U13499 (N_13499,N_12697,N_12039);
and U13500 (N_13500,N_12048,N_12335);
or U13501 (N_13501,N_12751,N_12011);
and U13502 (N_13502,N_12517,N_12956);
or U13503 (N_13503,N_12041,N_12523);
or U13504 (N_13504,N_12157,N_12243);
and U13505 (N_13505,N_12205,N_12302);
xor U13506 (N_13506,N_12188,N_12330);
or U13507 (N_13507,N_12039,N_12968);
nand U13508 (N_13508,N_12169,N_12753);
nand U13509 (N_13509,N_12777,N_12206);
nor U13510 (N_13510,N_12567,N_12011);
xnor U13511 (N_13511,N_12952,N_12451);
nand U13512 (N_13512,N_12675,N_12589);
xnor U13513 (N_13513,N_12049,N_12702);
nand U13514 (N_13514,N_12281,N_12115);
nor U13515 (N_13515,N_12750,N_12818);
xnor U13516 (N_13516,N_12730,N_12848);
nand U13517 (N_13517,N_12515,N_12670);
nor U13518 (N_13518,N_12632,N_12497);
nor U13519 (N_13519,N_12599,N_12188);
and U13520 (N_13520,N_12243,N_12423);
nand U13521 (N_13521,N_12972,N_12976);
xnor U13522 (N_13522,N_12415,N_12271);
nand U13523 (N_13523,N_12649,N_12216);
nand U13524 (N_13524,N_12231,N_12152);
and U13525 (N_13525,N_12019,N_12527);
nand U13526 (N_13526,N_12950,N_12832);
nand U13527 (N_13527,N_12927,N_12818);
nand U13528 (N_13528,N_12992,N_12780);
nor U13529 (N_13529,N_12028,N_12514);
and U13530 (N_13530,N_12894,N_12436);
and U13531 (N_13531,N_12639,N_12183);
nand U13532 (N_13532,N_12407,N_12140);
nand U13533 (N_13533,N_12329,N_12366);
nor U13534 (N_13534,N_12313,N_12304);
and U13535 (N_13535,N_12451,N_12205);
and U13536 (N_13536,N_12002,N_12051);
and U13537 (N_13537,N_12539,N_12670);
nor U13538 (N_13538,N_12962,N_12626);
or U13539 (N_13539,N_12375,N_12457);
nor U13540 (N_13540,N_12679,N_12425);
nand U13541 (N_13541,N_12165,N_12172);
and U13542 (N_13542,N_12910,N_12065);
nand U13543 (N_13543,N_12627,N_12370);
nand U13544 (N_13544,N_12324,N_12721);
xnor U13545 (N_13545,N_12794,N_12445);
nand U13546 (N_13546,N_12575,N_12930);
nor U13547 (N_13547,N_12773,N_12051);
nor U13548 (N_13548,N_12136,N_12597);
nand U13549 (N_13549,N_12857,N_12835);
or U13550 (N_13550,N_12315,N_12749);
nand U13551 (N_13551,N_12824,N_12645);
and U13552 (N_13552,N_12965,N_12300);
or U13553 (N_13553,N_12505,N_12713);
nor U13554 (N_13554,N_12498,N_12309);
and U13555 (N_13555,N_12609,N_12962);
and U13556 (N_13556,N_12638,N_12878);
nand U13557 (N_13557,N_12320,N_12640);
xnor U13558 (N_13558,N_12575,N_12879);
and U13559 (N_13559,N_12946,N_12476);
or U13560 (N_13560,N_12286,N_12911);
nand U13561 (N_13561,N_12868,N_12984);
nor U13562 (N_13562,N_12528,N_12466);
or U13563 (N_13563,N_12310,N_12308);
nor U13564 (N_13564,N_12712,N_12126);
and U13565 (N_13565,N_12838,N_12990);
nor U13566 (N_13566,N_12502,N_12684);
or U13567 (N_13567,N_12823,N_12755);
and U13568 (N_13568,N_12137,N_12466);
and U13569 (N_13569,N_12807,N_12867);
xor U13570 (N_13570,N_12342,N_12297);
nand U13571 (N_13571,N_12889,N_12746);
nand U13572 (N_13572,N_12603,N_12693);
and U13573 (N_13573,N_12593,N_12324);
nor U13574 (N_13574,N_12507,N_12989);
or U13575 (N_13575,N_12782,N_12634);
or U13576 (N_13576,N_12756,N_12182);
and U13577 (N_13577,N_12655,N_12010);
nand U13578 (N_13578,N_12395,N_12669);
and U13579 (N_13579,N_12116,N_12027);
or U13580 (N_13580,N_12121,N_12301);
and U13581 (N_13581,N_12731,N_12526);
and U13582 (N_13582,N_12044,N_12989);
nor U13583 (N_13583,N_12920,N_12676);
and U13584 (N_13584,N_12178,N_12001);
or U13585 (N_13585,N_12702,N_12436);
nand U13586 (N_13586,N_12180,N_12792);
and U13587 (N_13587,N_12184,N_12562);
or U13588 (N_13588,N_12451,N_12328);
nand U13589 (N_13589,N_12965,N_12495);
xnor U13590 (N_13590,N_12389,N_12650);
nor U13591 (N_13591,N_12060,N_12533);
nand U13592 (N_13592,N_12383,N_12019);
nor U13593 (N_13593,N_12093,N_12514);
or U13594 (N_13594,N_12562,N_12677);
nor U13595 (N_13595,N_12278,N_12527);
or U13596 (N_13596,N_12720,N_12234);
nor U13597 (N_13597,N_12046,N_12870);
and U13598 (N_13598,N_12454,N_12340);
and U13599 (N_13599,N_12622,N_12968);
and U13600 (N_13600,N_12886,N_12565);
or U13601 (N_13601,N_12166,N_12110);
or U13602 (N_13602,N_12902,N_12276);
or U13603 (N_13603,N_12485,N_12775);
or U13604 (N_13604,N_12564,N_12112);
nor U13605 (N_13605,N_12150,N_12381);
xnor U13606 (N_13606,N_12672,N_12359);
or U13607 (N_13607,N_12296,N_12879);
or U13608 (N_13608,N_12120,N_12932);
and U13609 (N_13609,N_12040,N_12231);
or U13610 (N_13610,N_12822,N_12320);
nor U13611 (N_13611,N_12224,N_12555);
nor U13612 (N_13612,N_12665,N_12939);
nand U13613 (N_13613,N_12334,N_12006);
or U13614 (N_13614,N_12028,N_12044);
and U13615 (N_13615,N_12428,N_12835);
and U13616 (N_13616,N_12999,N_12702);
and U13617 (N_13617,N_12725,N_12713);
or U13618 (N_13618,N_12949,N_12665);
nor U13619 (N_13619,N_12972,N_12155);
nand U13620 (N_13620,N_12230,N_12196);
nand U13621 (N_13621,N_12770,N_12653);
nor U13622 (N_13622,N_12348,N_12504);
nor U13623 (N_13623,N_12387,N_12838);
or U13624 (N_13624,N_12203,N_12770);
nor U13625 (N_13625,N_12043,N_12276);
nand U13626 (N_13626,N_12550,N_12761);
and U13627 (N_13627,N_12737,N_12048);
nand U13628 (N_13628,N_12180,N_12965);
nand U13629 (N_13629,N_12098,N_12789);
xnor U13630 (N_13630,N_12406,N_12788);
nor U13631 (N_13631,N_12713,N_12739);
and U13632 (N_13632,N_12876,N_12246);
nand U13633 (N_13633,N_12758,N_12904);
nand U13634 (N_13634,N_12141,N_12482);
nand U13635 (N_13635,N_12114,N_12063);
nand U13636 (N_13636,N_12108,N_12708);
nand U13637 (N_13637,N_12224,N_12123);
or U13638 (N_13638,N_12930,N_12527);
and U13639 (N_13639,N_12350,N_12867);
nor U13640 (N_13640,N_12110,N_12074);
xor U13641 (N_13641,N_12858,N_12293);
nor U13642 (N_13642,N_12202,N_12139);
or U13643 (N_13643,N_12065,N_12634);
or U13644 (N_13644,N_12476,N_12790);
xor U13645 (N_13645,N_12947,N_12622);
and U13646 (N_13646,N_12689,N_12396);
nor U13647 (N_13647,N_12404,N_12545);
and U13648 (N_13648,N_12487,N_12435);
nor U13649 (N_13649,N_12591,N_12691);
or U13650 (N_13650,N_12887,N_12572);
nand U13651 (N_13651,N_12876,N_12745);
nor U13652 (N_13652,N_12130,N_12480);
nand U13653 (N_13653,N_12385,N_12133);
or U13654 (N_13654,N_12399,N_12261);
nand U13655 (N_13655,N_12188,N_12450);
and U13656 (N_13656,N_12040,N_12122);
or U13657 (N_13657,N_12222,N_12322);
or U13658 (N_13658,N_12923,N_12185);
and U13659 (N_13659,N_12825,N_12897);
nand U13660 (N_13660,N_12006,N_12323);
and U13661 (N_13661,N_12822,N_12181);
and U13662 (N_13662,N_12841,N_12493);
and U13663 (N_13663,N_12834,N_12189);
and U13664 (N_13664,N_12608,N_12409);
and U13665 (N_13665,N_12968,N_12754);
nand U13666 (N_13666,N_12219,N_12060);
nor U13667 (N_13667,N_12469,N_12251);
xor U13668 (N_13668,N_12808,N_12289);
nor U13669 (N_13669,N_12557,N_12525);
nand U13670 (N_13670,N_12459,N_12314);
or U13671 (N_13671,N_12575,N_12993);
and U13672 (N_13672,N_12743,N_12974);
xor U13673 (N_13673,N_12933,N_12462);
nand U13674 (N_13674,N_12746,N_12351);
or U13675 (N_13675,N_12343,N_12236);
nor U13676 (N_13676,N_12538,N_12691);
or U13677 (N_13677,N_12433,N_12635);
nor U13678 (N_13678,N_12003,N_12175);
and U13679 (N_13679,N_12769,N_12695);
or U13680 (N_13680,N_12396,N_12425);
nor U13681 (N_13681,N_12980,N_12718);
nand U13682 (N_13682,N_12954,N_12591);
nand U13683 (N_13683,N_12082,N_12559);
nand U13684 (N_13684,N_12844,N_12797);
and U13685 (N_13685,N_12973,N_12070);
and U13686 (N_13686,N_12135,N_12872);
or U13687 (N_13687,N_12587,N_12931);
or U13688 (N_13688,N_12647,N_12418);
nand U13689 (N_13689,N_12610,N_12430);
nand U13690 (N_13690,N_12144,N_12969);
nor U13691 (N_13691,N_12660,N_12291);
xnor U13692 (N_13692,N_12182,N_12079);
nand U13693 (N_13693,N_12690,N_12017);
nor U13694 (N_13694,N_12078,N_12894);
xor U13695 (N_13695,N_12616,N_12555);
or U13696 (N_13696,N_12023,N_12124);
nor U13697 (N_13697,N_12636,N_12114);
nand U13698 (N_13698,N_12401,N_12568);
nor U13699 (N_13699,N_12279,N_12465);
nor U13700 (N_13700,N_12634,N_12130);
and U13701 (N_13701,N_12463,N_12908);
and U13702 (N_13702,N_12657,N_12693);
nor U13703 (N_13703,N_12564,N_12176);
and U13704 (N_13704,N_12909,N_12343);
and U13705 (N_13705,N_12625,N_12537);
nand U13706 (N_13706,N_12110,N_12719);
and U13707 (N_13707,N_12426,N_12329);
and U13708 (N_13708,N_12625,N_12375);
and U13709 (N_13709,N_12662,N_12636);
nor U13710 (N_13710,N_12793,N_12512);
xnor U13711 (N_13711,N_12182,N_12623);
and U13712 (N_13712,N_12573,N_12328);
xnor U13713 (N_13713,N_12348,N_12085);
or U13714 (N_13714,N_12718,N_12424);
nand U13715 (N_13715,N_12691,N_12814);
or U13716 (N_13716,N_12671,N_12340);
and U13717 (N_13717,N_12311,N_12336);
nand U13718 (N_13718,N_12760,N_12567);
nand U13719 (N_13719,N_12605,N_12851);
nor U13720 (N_13720,N_12672,N_12850);
or U13721 (N_13721,N_12072,N_12703);
nor U13722 (N_13722,N_12852,N_12185);
nand U13723 (N_13723,N_12333,N_12911);
or U13724 (N_13724,N_12318,N_12930);
xor U13725 (N_13725,N_12500,N_12873);
and U13726 (N_13726,N_12512,N_12433);
and U13727 (N_13727,N_12368,N_12529);
and U13728 (N_13728,N_12759,N_12544);
nand U13729 (N_13729,N_12195,N_12946);
and U13730 (N_13730,N_12997,N_12076);
xor U13731 (N_13731,N_12062,N_12409);
and U13732 (N_13732,N_12668,N_12979);
and U13733 (N_13733,N_12690,N_12948);
and U13734 (N_13734,N_12751,N_12233);
or U13735 (N_13735,N_12819,N_12297);
and U13736 (N_13736,N_12433,N_12860);
nand U13737 (N_13737,N_12908,N_12834);
nand U13738 (N_13738,N_12828,N_12825);
and U13739 (N_13739,N_12260,N_12846);
nor U13740 (N_13740,N_12653,N_12041);
or U13741 (N_13741,N_12191,N_12121);
nor U13742 (N_13742,N_12368,N_12146);
and U13743 (N_13743,N_12148,N_12468);
nor U13744 (N_13744,N_12905,N_12586);
xnor U13745 (N_13745,N_12065,N_12721);
nor U13746 (N_13746,N_12385,N_12228);
nand U13747 (N_13747,N_12776,N_12180);
nand U13748 (N_13748,N_12261,N_12876);
nor U13749 (N_13749,N_12395,N_12953);
and U13750 (N_13750,N_12950,N_12132);
and U13751 (N_13751,N_12638,N_12294);
nor U13752 (N_13752,N_12513,N_12294);
or U13753 (N_13753,N_12372,N_12684);
nor U13754 (N_13754,N_12276,N_12903);
nor U13755 (N_13755,N_12703,N_12173);
or U13756 (N_13756,N_12040,N_12272);
nor U13757 (N_13757,N_12010,N_12791);
nor U13758 (N_13758,N_12097,N_12130);
nor U13759 (N_13759,N_12203,N_12345);
nand U13760 (N_13760,N_12851,N_12767);
or U13761 (N_13761,N_12271,N_12534);
or U13762 (N_13762,N_12040,N_12985);
nand U13763 (N_13763,N_12887,N_12745);
nand U13764 (N_13764,N_12020,N_12882);
nor U13765 (N_13765,N_12153,N_12852);
xor U13766 (N_13766,N_12452,N_12699);
or U13767 (N_13767,N_12899,N_12653);
nor U13768 (N_13768,N_12589,N_12529);
xor U13769 (N_13769,N_12126,N_12187);
xor U13770 (N_13770,N_12710,N_12296);
and U13771 (N_13771,N_12257,N_12924);
xor U13772 (N_13772,N_12322,N_12823);
nand U13773 (N_13773,N_12338,N_12909);
nand U13774 (N_13774,N_12196,N_12606);
nand U13775 (N_13775,N_12378,N_12394);
and U13776 (N_13776,N_12427,N_12337);
or U13777 (N_13777,N_12333,N_12087);
and U13778 (N_13778,N_12758,N_12909);
nand U13779 (N_13779,N_12386,N_12893);
or U13780 (N_13780,N_12869,N_12939);
xor U13781 (N_13781,N_12666,N_12192);
or U13782 (N_13782,N_12478,N_12899);
xor U13783 (N_13783,N_12176,N_12081);
nand U13784 (N_13784,N_12052,N_12719);
or U13785 (N_13785,N_12364,N_12129);
and U13786 (N_13786,N_12549,N_12837);
xnor U13787 (N_13787,N_12008,N_12070);
nand U13788 (N_13788,N_12768,N_12574);
and U13789 (N_13789,N_12999,N_12268);
nand U13790 (N_13790,N_12893,N_12651);
nor U13791 (N_13791,N_12364,N_12700);
nand U13792 (N_13792,N_12306,N_12657);
xor U13793 (N_13793,N_12314,N_12387);
or U13794 (N_13794,N_12067,N_12883);
nor U13795 (N_13795,N_12904,N_12957);
nand U13796 (N_13796,N_12361,N_12160);
nand U13797 (N_13797,N_12494,N_12689);
or U13798 (N_13798,N_12385,N_12872);
xnor U13799 (N_13799,N_12466,N_12108);
or U13800 (N_13800,N_12374,N_12390);
and U13801 (N_13801,N_12495,N_12542);
nand U13802 (N_13802,N_12532,N_12355);
nor U13803 (N_13803,N_12324,N_12138);
or U13804 (N_13804,N_12340,N_12712);
nand U13805 (N_13805,N_12251,N_12070);
nor U13806 (N_13806,N_12616,N_12413);
and U13807 (N_13807,N_12489,N_12410);
nor U13808 (N_13808,N_12704,N_12103);
xor U13809 (N_13809,N_12406,N_12807);
nor U13810 (N_13810,N_12346,N_12698);
or U13811 (N_13811,N_12366,N_12297);
or U13812 (N_13812,N_12512,N_12117);
nand U13813 (N_13813,N_12658,N_12130);
or U13814 (N_13814,N_12338,N_12680);
nor U13815 (N_13815,N_12346,N_12956);
nor U13816 (N_13816,N_12035,N_12277);
xor U13817 (N_13817,N_12684,N_12224);
nand U13818 (N_13818,N_12357,N_12034);
and U13819 (N_13819,N_12846,N_12500);
nor U13820 (N_13820,N_12649,N_12879);
xnor U13821 (N_13821,N_12995,N_12166);
and U13822 (N_13822,N_12442,N_12892);
xnor U13823 (N_13823,N_12562,N_12027);
nor U13824 (N_13824,N_12748,N_12924);
nand U13825 (N_13825,N_12440,N_12302);
or U13826 (N_13826,N_12628,N_12861);
or U13827 (N_13827,N_12980,N_12189);
and U13828 (N_13828,N_12096,N_12180);
and U13829 (N_13829,N_12105,N_12277);
and U13830 (N_13830,N_12487,N_12791);
and U13831 (N_13831,N_12919,N_12719);
nor U13832 (N_13832,N_12325,N_12775);
nor U13833 (N_13833,N_12428,N_12133);
and U13834 (N_13834,N_12719,N_12814);
nand U13835 (N_13835,N_12575,N_12311);
nand U13836 (N_13836,N_12403,N_12384);
nor U13837 (N_13837,N_12135,N_12294);
and U13838 (N_13838,N_12674,N_12146);
or U13839 (N_13839,N_12623,N_12956);
or U13840 (N_13840,N_12733,N_12643);
xor U13841 (N_13841,N_12524,N_12783);
xor U13842 (N_13842,N_12818,N_12573);
or U13843 (N_13843,N_12454,N_12994);
and U13844 (N_13844,N_12009,N_12109);
and U13845 (N_13845,N_12944,N_12942);
nand U13846 (N_13846,N_12483,N_12178);
nor U13847 (N_13847,N_12216,N_12193);
nor U13848 (N_13848,N_12244,N_12747);
nand U13849 (N_13849,N_12670,N_12593);
nor U13850 (N_13850,N_12579,N_12374);
nor U13851 (N_13851,N_12419,N_12169);
xnor U13852 (N_13852,N_12148,N_12514);
or U13853 (N_13853,N_12768,N_12975);
or U13854 (N_13854,N_12508,N_12929);
xnor U13855 (N_13855,N_12117,N_12790);
or U13856 (N_13856,N_12369,N_12187);
or U13857 (N_13857,N_12281,N_12616);
xnor U13858 (N_13858,N_12295,N_12476);
nor U13859 (N_13859,N_12410,N_12480);
nand U13860 (N_13860,N_12408,N_12956);
and U13861 (N_13861,N_12855,N_12421);
and U13862 (N_13862,N_12492,N_12953);
nor U13863 (N_13863,N_12600,N_12081);
nand U13864 (N_13864,N_12714,N_12032);
or U13865 (N_13865,N_12341,N_12551);
xor U13866 (N_13866,N_12665,N_12303);
or U13867 (N_13867,N_12794,N_12658);
nand U13868 (N_13868,N_12396,N_12676);
nand U13869 (N_13869,N_12377,N_12431);
and U13870 (N_13870,N_12677,N_12302);
or U13871 (N_13871,N_12507,N_12710);
nand U13872 (N_13872,N_12361,N_12214);
nor U13873 (N_13873,N_12387,N_12798);
nand U13874 (N_13874,N_12245,N_12229);
nor U13875 (N_13875,N_12099,N_12207);
nor U13876 (N_13876,N_12072,N_12352);
or U13877 (N_13877,N_12911,N_12852);
nor U13878 (N_13878,N_12935,N_12454);
nor U13879 (N_13879,N_12146,N_12962);
nor U13880 (N_13880,N_12515,N_12380);
nand U13881 (N_13881,N_12123,N_12739);
nand U13882 (N_13882,N_12613,N_12033);
or U13883 (N_13883,N_12263,N_12400);
nor U13884 (N_13884,N_12694,N_12553);
nor U13885 (N_13885,N_12039,N_12324);
or U13886 (N_13886,N_12802,N_12131);
nor U13887 (N_13887,N_12801,N_12683);
or U13888 (N_13888,N_12221,N_12727);
or U13889 (N_13889,N_12652,N_12615);
nand U13890 (N_13890,N_12143,N_12414);
nor U13891 (N_13891,N_12027,N_12951);
or U13892 (N_13892,N_12075,N_12019);
nor U13893 (N_13893,N_12966,N_12739);
nor U13894 (N_13894,N_12106,N_12908);
nor U13895 (N_13895,N_12176,N_12393);
nand U13896 (N_13896,N_12631,N_12378);
nor U13897 (N_13897,N_12495,N_12124);
xor U13898 (N_13898,N_12101,N_12259);
nand U13899 (N_13899,N_12529,N_12521);
and U13900 (N_13900,N_12284,N_12114);
nand U13901 (N_13901,N_12053,N_12764);
nand U13902 (N_13902,N_12664,N_12300);
nand U13903 (N_13903,N_12585,N_12230);
xor U13904 (N_13904,N_12498,N_12055);
and U13905 (N_13905,N_12457,N_12422);
nor U13906 (N_13906,N_12692,N_12127);
nor U13907 (N_13907,N_12452,N_12572);
xnor U13908 (N_13908,N_12414,N_12970);
nor U13909 (N_13909,N_12258,N_12938);
nand U13910 (N_13910,N_12749,N_12436);
nand U13911 (N_13911,N_12139,N_12713);
nor U13912 (N_13912,N_12688,N_12666);
and U13913 (N_13913,N_12790,N_12011);
and U13914 (N_13914,N_12077,N_12943);
or U13915 (N_13915,N_12240,N_12144);
nor U13916 (N_13916,N_12224,N_12986);
nor U13917 (N_13917,N_12809,N_12065);
nor U13918 (N_13918,N_12639,N_12282);
nor U13919 (N_13919,N_12077,N_12142);
or U13920 (N_13920,N_12502,N_12421);
xnor U13921 (N_13921,N_12402,N_12749);
nor U13922 (N_13922,N_12344,N_12358);
nor U13923 (N_13923,N_12145,N_12305);
nand U13924 (N_13924,N_12102,N_12663);
nor U13925 (N_13925,N_12169,N_12031);
nand U13926 (N_13926,N_12177,N_12089);
nor U13927 (N_13927,N_12785,N_12991);
nor U13928 (N_13928,N_12044,N_12204);
or U13929 (N_13929,N_12399,N_12501);
and U13930 (N_13930,N_12464,N_12682);
nor U13931 (N_13931,N_12409,N_12066);
or U13932 (N_13932,N_12052,N_12290);
xnor U13933 (N_13933,N_12340,N_12369);
and U13934 (N_13934,N_12511,N_12419);
nand U13935 (N_13935,N_12390,N_12503);
xnor U13936 (N_13936,N_12057,N_12200);
and U13937 (N_13937,N_12961,N_12038);
and U13938 (N_13938,N_12710,N_12484);
and U13939 (N_13939,N_12170,N_12929);
or U13940 (N_13940,N_12893,N_12812);
or U13941 (N_13941,N_12644,N_12249);
nand U13942 (N_13942,N_12041,N_12289);
nor U13943 (N_13943,N_12485,N_12425);
nand U13944 (N_13944,N_12946,N_12219);
or U13945 (N_13945,N_12185,N_12718);
nor U13946 (N_13946,N_12616,N_12253);
nor U13947 (N_13947,N_12558,N_12233);
and U13948 (N_13948,N_12775,N_12007);
nand U13949 (N_13949,N_12603,N_12833);
xnor U13950 (N_13950,N_12152,N_12939);
or U13951 (N_13951,N_12257,N_12820);
nor U13952 (N_13952,N_12029,N_12274);
xor U13953 (N_13953,N_12135,N_12030);
or U13954 (N_13954,N_12379,N_12485);
nor U13955 (N_13955,N_12033,N_12887);
nor U13956 (N_13956,N_12426,N_12567);
or U13957 (N_13957,N_12468,N_12549);
xor U13958 (N_13958,N_12517,N_12754);
nor U13959 (N_13959,N_12512,N_12235);
nor U13960 (N_13960,N_12348,N_12272);
nor U13961 (N_13961,N_12257,N_12649);
nor U13962 (N_13962,N_12605,N_12982);
nand U13963 (N_13963,N_12428,N_12176);
nor U13964 (N_13964,N_12817,N_12887);
nor U13965 (N_13965,N_12449,N_12166);
and U13966 (N_13966,N_12330,N_12339);
nor U13967 (N_13967,N_12164,N_12360);
nor U13968 (N_13968,N_12298,N_12348);
xor U13969 (N_13969,N_12576,N_12430);
and U13970 (N_13970,N_12047,N_12407);
xnor U13971 (N_13971,N_12359,N_12997);
and U13972 (N_13972,N_12627,N_12977);
or U13973 (N_13973,N_12902,N_12241);
nand U13974 (N_13974,N_12553,N_12224);
nand U13975 (N_13975,N_12212,N_12483);
or U13976 (N_13976,N_12747,N_12660);
xor U13977 (N_13977,N_12392,N_12913);
nor U13978 (N_13978,N_12033,N_12424);
nand U13979 (N_13979,N_12606,N_12164);
nor U13980 (N_13980,N_12375,N_12272);
nor U13981 (N_13981,N_12553,N_12669);
nand U13982 (N_13982,N_12824,N_12915);
nand U13983 (N_13983,N_12542,N_12799);
or U13984 (N_13984,N_12942,N_12856);
and U13985 (N_13985,N_12117,N_12843);
xnor U13986 (N_13986,N_12052,N_12318);
nand U13987 (N_13987,N_12577,N_12141);
nand U13988 (N_13988,N_12768,N_12684);
nor U13989 (N_13989,N_12056,N_12225);
nor U13990 (N_13990,N_12478,N_12535);
nor U13991 (N_13991,N_12890,N_12706);
nor U13992 (N_13992,N_12283,N_12189);
xnor U13993 (N_13993,N_12645,N_12997);
nand U13994 (N_13994,N_12603,N_12112);
or U13995 (N_13995,N_12686,N_12760);
and U13996 (N_13996,N_12581,N_12266);
xnor U13997 (N_13997,N_12504,N_12050);
or U13998 (N_13998,N_12797,N_12889);
nor U13999 (N_13999,N_12415,N_12956);
nand U14000 (N_14000,N_13531,N_13532);
and U14001 (N_14001,N_13544,N_13733);
or U14002 (N_14002,N_13795,N_13934);
xor U14003 (N_14003,N_13212,N_13200);
xor U14004 (N_14004,N_13654,N_13957);
nand U14005 (N_14005,N_13898,N_13618);
and U14006 (N_14006,N_13490,N_13278);
and U14007 (N_14007,N_13009,N_13002);
xor U14008 (N_14008,N_13605,N_13555);
nor U14009 (N_14009,N_13901,N_13725);
nand U14010 (N_14010,N_13546,N_13098);
nor U14011 (N_14011,N_13420,N_13863);
or U14012 (N_14012,N_13272,N_13767);
nand U14013 (N_14013,N_13864,N_13664);
nor U14014 (N_14014,N_13634,N_13675);
nand U14015 (N_14015,N_13735,N_13802);
nand U14016 (N_14016,N_13261,N_13488);
nor U14017 (N_14017,N_13955,N_13720);
and U14018 (N_14018,N_13855,N_13171);
nand U14019 (N_14019,N_13834,N_13401);
or U14020 (N_14020,N_13086,N_13251);
or U14021 (N_14021,N_13483,N_13335);
nor U14022 (N_14022,N_13011,N_13770);
and U14023 (N_14023,N_13263,N_13260);
nand U14024 (N_14024,N_13637,N_13151);
nand U14025 (N_14025,N_13216,N_13827);
nor U14026 (N_14026,N_13465,N_13785);
or U14027 (N_14027,N_13588,N_13832);
nor U14028 (N_14028,N_13456,N_13110);
xnor U14029 (N_14029,N_13311,N_13611);
nand U14030 (N_14030,N_13027,N_13643);
or U14031 (N_14031,N_13364,N_13942);
nand U14032 (N_14032,N_13852,N_13285);
nand U14033 (N_14033,N_13851,N_13895);
and U14034 (N_14034,N_13803,N_13338);
nor U14035 (N_14035,N_13932,N_13961);
nand U14036 (N_14036,N_13575,N_13615);
or U14037 (N_14037,N_13821,N_13873);
nor U14038 (N_14038,N_13400,N_13585);
nand U14039 (N_14039,N_13826,N_13182);
nor U14040 (N_14040,N_13309,N_13213);
nor U14041 (N_14041,N_13768,N_13199);
nor U14042 (N_14042,N_13917,N_13730);
nor U14043 (N_14043,N_13413,N_13717);
nor U14044 (N_14044,N_13336,N_13220);
and U14045 (N_14045,N_13387,N_13119);
and U14046 (N_14046,N_13244,N_13798);
and U14047 (N_14047,N_13740,N_13576);
nor U14048 (N_14048,N_13810,N_13649);
and U14049 (N_14049,N_13231,N_13485);
nand U14050 (N_14050,N_13640,N_13776);
nor U14051 (N_14051,N_13081,N_13948);
nor U14052 (N_14052,N_13631,N_13983);
and U14053 (N_14053,N_13903,N_13849);
nand U14054 (N_14054,N_13587,N_13202);
and U14055 (N_14055,N_13994,N_13668);
or U14056 (N_14056,N_13923,N_13981);
nand U14057 (N_14057,N_13551,N_13255);
or U14058 (N_14058,N_13842,N_13612);
nand U14059 (N_14059,N_13105,N_13129);
or U14060 (N_14060,N_13678,N_13038);
xor U14061 (N_14061,N_13509,N_13985);
nand U14062 (N_14062,N_13736,N_13931);
nand U14063 (N_14063,N_13807,N_13843);
nor U14064 (N_14064,N_13258,N_13557);
nor U14065 (N_14065,N_13698,N_13040);
nand U14066 (N_14066,N_13629,N_13714);
nand U14067 (N_14067,N_13166,N_13833);
nor U14068 (N_14068,N_13788,N_13159);
or U14069 (N_14069,N_13277,N_13134);
or U14070 (N_14070,N_13327,N_13369);
nor U14071 (N_14071,N_13458,N_13941);
or U14072 (N_14072,N_13750,N_13131);
or U14073 (N_14073,N_13878,N_13390);
and U14074 (N_14074,N_13326,N_13223);
nor U14075 (N_14075,N_13150,N_13621);
or U14076 (N_14076,N_13179,N_13759);
or U14077 (N_14077,N_13092,N_13404);
and U14078 (N_14078,N_13609,N_13321);
nand U14079 (N_14079,N_13626,N_13604);
or U14080 (N_14080,N_13867,N_13731);
xor U14081 (N_14081,N_13204,N_13474);
and U14082 (N_14082,N_13076,N_13121);
nand U14083 (N_14083,N_13882,N_13148);
nand U14084 (N_14084,N_13169,N_13058);
and U14085 (N_14085,N_13891,N_13333);
nor U14086 (N_14086,N_13742,N_13446);
or U14087 (N_14087,N_13727,N_13115);
or U14088 (N_14088,N_13493,N_13633);
or U14089 (N_14089,N_13471,N_13636);
or U14090 (N_14090,N_13806,N_13751);
xor U14091 (N_14091,N_13812,N_13118);
or U14092 (N_14092,N_13971,N_13286);
xnor U14093 (N_14093,N_13794,N_13234);
xor U14094 (N_14094,N_13672,N_13848);
or U14095 (N_14095,N_13581,N_13543);
or U14096 (N_14096,N_13738,N_13703);
or U14097 (N_14097,N_13536,N_13256);
xor U14098 (N_14098,N_13303,N_13419);
nor U14099 (N_14099,N_13693,N_13021);
and U14100 (N_14100,N_13180,N_13093);
nor U14101 (N_14101,N_13088,N_13174);
and U14102 (N_14102,N_13702,N_13195);
nor U14103 (N_14103,N_13032,N_13393);
nor U14104 (N_14104,N_13347,N_13349);
or U14105 (N_14105,N_13356,N_13332);
and U14106 (N_14106,N_13044,N_13872);
nor U14107 (N_14107,N_13573,N_13656);
nand U14108 (N_14108,N_13104,N_13793);
nor U14109 (N_14109,N_13667,N_13964);
nand U14110 (N_14110,N_13894,N_13402);
xor U14111 (N_14111,N_13059,N_13632);
xnor U14112 (N_14112,N_13008,N_13235);
or U14113 (N_14113,N_13215,N_13571);
nor U14114 (N_14114,N_13205,N_13958);
and U14115 (N_14115,N_13624,N_13582);
or U14116 (N_14116,N_13201,N_13425);
nor U14117 (N_14117,N_13377,N_13173);
or U14118 (N_14118,N_13719,N_13756);
or U14119 (N_14119,N_13319,N_13679);
nor U14120 (N_14120,N_13214,N_13014);
and U14121 (N_14121,N_13650,N_13914);
nor U14122 (N_14122,N_13315,N_13904);
and U14123 (N_14123,N_13784,N_13448);
nand U14124 (N_14124,N_13113,N_13363);
and U14125 (N_14125,N_13135,N_13950);
or U14126 (N_14126,N_13574,N_13301);
or U14127 (N_14127,N_13055,N_13491);
or U14128 (N_14128,N_13777,N_13190);
nor U14129 (N_14129,N_13760,N_13519);
nand U14130 (N_14130,N_13185,N_13775);
or U14131 (N_14131,N_13397,N_13921);
nand U14132 (N_14132,N_13973,N_13279);
or U14133 (N_14133,N_13391,N_13791);
and U14134 (N_14134,N_13623,N_13498);
nor U14135 (N_14135,N_13949,N_13550);
nor U14136 (N_14136,N_13619,N_13554);
or U14137 (N_14137,N_13562,N_13470);
nand U14138 (N_14138,N_13647,N_13437);
and U14139 (N_14139,N_13886,N_13883);
nor U14140 (N_14140,N_13183,N_13383);
and U14141 (N_14141,N_13007,N_13579);
nand U14142 (N_14142,N_13868,N_13034);
xnor U14143 (N_14143,N_13570,N_13748);
and U14144 (N_14144,N_13281,N_13999);
xnor U14145 (N_14145,N_13783,N_13359);
nor U14146 (N_14146,N_13096,N_13905);
nand U14147 (N_14147,N_13464,N_13811);
and U14148 (N_14148,N_13937,N_13123);
nor U14149 (N_14149,N_13249,N_13757);
nand U14150 (N_14150,N_13682,N_13769);
or U14151 (N_14151,N_13184,N_13595);
or U14152 (N_14152,N_13252,N_13829);
nor U14153 (N_14153,N_13196,N_13068);
nand U14154 (N_14154,N_13023,N_13300);
nor U14155 (N_14155,N_13427,N_13547);
and U14156 (N_14156,N_13762,N_13599);
nor U14157 (N_14157,N_13701,N_13847);
and U14158 (N_14158,N_13893,N_13210);
nand U14159 (N_14159,N_13658,N_13191);
or U14160 (N_14160,N_13389,N_13240);
xor U14161 (N_14161,N_13339,N_13399);
nand U14162 (N_14162,N_13565,N_13408);
or U14163 (N_14163,N_13450,N_13726);
nand U14164 (N_14164,N_13548,N_13126);
or U14165 (N_14165,N_13237,N_13421);
or U14166 (N_14166,N_13495,N_13165);
nor U14167 (N_14167,N_13592,N_13734);
or U14168 (N_14168,N_13688,N_13500);
and U14169 (N_14169,N_13157,N_13870);
nand U14170 (N_14170,N_13017,N_13177);
nor U14171 (N_14171,N_13149,N_13809);
nor U14172 (N_14172,N_13515,N_13954);
or U14173 (N_14173,N_13861,N_13501);
nor U14174 (N_14174,N_13975,N_13771);
xor U14175 (N_14175,N_13057,N_13317);
and U14176 (N_14176,N_13428,N_13225);
nor U14177 (N_14177,N_13854,N_13823);
nor U14178 (N_14178,N_13642,N_13885);
nand U14179 (N_14179,N_13029,N_13228);
nor U14180 (N_14180,N_13245,N_13559);
nor U14181 (N_14181,N_13520,N_13416);
nor U14182 (N_14182,N_13087,N_13350);
nor U14183 (N_14183,N_13927,N_13875);
nand U14184 (N_14184,N_13395,N_13013);
or U14185 (N_14185,N_13704,N_13375);
nand U14186 (N_14186,N_13262,N_13902);
or U14187 (N_14187,N_13250,N_13951);
nor U14188 (N_14188,N_13746,N_13161);
or U14189 (N_14189,N_13597,N_13602);
and U14190 (N_14190,N_13965,N_13845);
or U14191 (N_14191,N_13304,N_13598);
and U14192 (N_14192,N_13489,N_13354);
nand U14193 (N_14193,N_13487,N_13269);
nand U14194 (N_14194,N_13608,N_13473);
nor U14195 (N_14195,N_13324,N_13158);
nand U14196 (N_14196,N_13928,N_13229);
xnor U14197 (N_14197,N_13197,N_13938);
and U14198 (N_14198,N_13265,N_13030);
nor U14199 (N_14199,N_13671,N_13312);
nand U14200 (N_14200,N_13441,N_13695);
nor U14201 (N_14201,N_13696,N_13765);
or U14202 (N_14202,N_13208,N_13306);
and U14203 (N_14203,N_13538,N_13193);
or U14204 (N_14204,N_13295,N_13345);
xor U14205 (N_14205,N_13486,N_13545);
and U14206 (N_14206,N_13314,N_13107);
nor U14207 (N_14207,N_13522,N_13844);
and U14208 (N_14208,N_13167,N_13063);
xnor U14209 (N_14209,N_13403,N_13706);
and U14210 (N_14210,N_13253,N_13974);
nor U14211 (N_14211,N_13496,N_13313);
nor U14212 (N_14212,N_13075,N_13422);
or U14213 (N_14213,N_13139,N_13722);
nand U14214 (N_14214,N_13100,N_13755);
or U14215 (N_14215,N_13510,N_13995);
nor U14216 (N_14216,N_13374,N_13947);
xor U14217 (N_14217,N_13348,N_13050);
and U14218 (N_14218,N_13101,N_13689);
or U14219 (N_14219,N_13933,N_13398);
and U14220 (N_14220,N_13384,N_13153);
or U14221 (N_14221,N_13627,N_13298);
and U14222 (N_14222,N_13737,N_13911);
nand U14223 (N_14223,N_13410,N_13226);
xor U14224 (N_14224,N_13122,N_13127);
nand U14225 (N_14225,N_13963,N_13028);
xor U14226 (N_14226,N_13972,N_13146);
or U14227 (N_14227,N_13521,N_13323);
nand U14228 (N_14228,N_13128,N_13924);
or U14229 (N_14229,N_13516,N_13020);
or U14230 (N_14230,N_13881,N_13082);
and U14231 (N_14231,N_13772,N_13539);
xor U14232 (N_14232,N_13005,N_13724);
xor U14233 (N_14233,N_13584,N_13417);
nand U14234 (N_14234,N_13346,N_13986);
or U14235 (N_14235,N_13787,N_13039);
nor U14236 (N_14236,N_13247,N_13816);
nor U14237 (N_14237,N_13070,N_13207);
nor U14238 (N_14238,N_13687,N_13876);
or U14239 (N_14239,N_13133,N_13935);
or U14240 (N_14240,N_13836,N_13305);
nor U14241 (N_14241,N_13072,N_13080);
or U14242 (N_14242,N_13945,N_13198);
and U14243 (N_14243,N_13376,N_13978);
nor U14244 (N_14244,N_13529,N_13508);
or U14245 (N_14245,N_13172,N_13857);
nor U14246 (N_14246,N_13690,N_13168);
nand U14247 (N_14247,N_13130,N_13908);
or U14248 (N_14248,N_13800,N_13630);
or U14249 (N_14249,N_13424,N_13558);
nand U14250 (N_14250,N_13713,N_13566);
nor U14251 (N_14251,N_13880,N_13163);
nor U14252 (N_14252,N_13064,N_13537);
nor U14253 (N_14253,N_13897,N_13242);
nor U14254 (N_14254,N_13653,N_13916);
or U14255 (N_14255,N_13342,N_13291);
nor U14256 (N_14256,N_13540,N_13114);
and U14257 (N_14257,N_13060,N_13109);
xor U14258 (N_14258,N_13813,N_13381);
and U14259 (N_14259,N_13361,N_13469);
nand U14260 (N_14260,N_13457,N_13188);
nor U14261 (N_14261,N_13353,N_13970);
or U14262 (N_14262,N_13764,N_13953);
and U14263 (N_14263,N_13239,N_13209);
nor U14264 (N_14264,N_13936,N_13367);
and U14265 (N_14265,N_13061,N_13962);
xor U14266 (N_14266,N_13047,N_13357);
and U14267 (N_14267,N_13680,N_13796);
and U14268 (N_14268,N_13890,N_13284);
xor U14269 (N_14269,N_13049,N_13170);
or U14270 (N_14270,N_13528,N_13869);
nand U14271 (N_14271,N_13120,N_13694);
or U14272 (N_14272,N_13418,N_13230);
and U14273 (N_14273,N_13814,N_13415);
and U14274 (N_14274,N_13856,N_13406);
nor U14275 (N_14275,N_13461,N_13429);
xor U14276 (N_14276,N_13739,N_13988);
and U14277 (N_14277,N_13676,N_13665);
nor U14278 (N_14278,N_13639,N_13503);
nor U14279 (N_14279,N_13589,N_13628);
and U14280 (N_14280,N_13344,N_13553);
nor U14281 (N_14281,N_13066,N_13003);
or U14282 (N_14282,N_13340,N_13111);
and U14283 (N_14283,N_13850,N_13318);
nor U14284 (N_14284,N_13266,N_13912);
xor U14285 (N_14285,N_13670,N_13792);
and U14286 (N_14286,N_13246,N_13297);
nand U14287 (N_14287,N_13477,N_13683);
or U14288 (N_14288,N_13046,N_13287);
nor U14289 (N_14289,N_13162,N_13655);
nand U14290 (N_14290,N_13797,N_13711);
and U14291 (N_14291,N_13661,N_13138);
xor U14292 (N_14292,N_13896,N_13155);
nor U14293 (N_14293,N_13433,N_13232);
nor U14294 (N_14294,N_13859,N_13186);
xor U14295 (N_14295,N_13998,N_13513);
xnor U14296 (N_14296,N_13468,N_13037);
nor U14297 (N_14297,N_13892,N_13926);
or U14298 (N_14298,N_13583,N_13572);
nand U14299 (N_14299,N_13673,N_13663);
or U14300 (N_14300,N_13865,N_13745);
and U14301 (N_14301,N_13411,N_13729);
nand U14302 (N_14302,N_13365,N_13817);
or U14303 (N_14303,N_13053,N_13801);
nor U14304 (N_14304,N_13569,N_13681);
nor U14305 (N_14305,N_13296,N_13325);
or U14306 (N_14306,N_13116,N_13164);
or U14307 (N_14307,N_13394,N_13976);
and U14308 (N_14308,N_13106,N_13140);
and U14309 (N_14309,N_13514,N_13979);
or U14310 (N_14310,N_13789,N_13705);
nor U14311 (N_14311,N_13233,N_13016);
nand U14312 (N_14312,N_13102,N_13459);
xor U14313 (N_14313,N_13211,N_13043);
nor U14314 (N_14314,N_13499,N_13045);
xnor U14315 (N_14315,N_13447,N_13292);
and U14316 (N_14316,N_13918,N_13271);
nand U14317 (N_14317,N_13993,N_13054);
nor U14318 (N_14318,N_13646,N_13526);
and U14319 (N_14319,N_13125,N_13463);
and U14320 (N_14320,N_13600,N_13280);
xnor U14321 (N_14321,N_13178,N_13444);
nand U14322 (N_14322,N_13685,N_13659);
or U14323 (N_14323,N_13723,N_13423);
nand U14324 (N_14324,N_13567,N_13079);
xor U14325 (N_14325,N_13586,N_13943);
or U14326 (N_14326,N_13238,N_13328);
and U14327 (N_14327,N_13378,N_13453);
xor U14328 (N_14328,N_13078,N_13430);
or U14329 (N_14329,N_13268,N_13132);
nor U14330 (N_14330,N_13065,N_13984);
nand U14331 (N_14331,N_13635,N_13227);
nor U14332 (N_14332,N_13660,N_13552);
or U14333 (N_14333,N_13930,N_13031);
nand U14334 (N_14334,N_13780,N_13289);
and U14335 (N_14335,N_13077,N_13097);
or U14336 (N_14336,N_13818,N_13530);
nor U14337 (N_14337,N_13095,N_13966);
nand U14338 (N_14338,N_13684,N_13362);
and U14339 (N_14339,N_13142,N_13270);
and U14340 (N_14340,N_13112,N_13992);
or U14341 (N_14341,N_13607,N_13203);
nor U14342 (N_14342,N_13645,N_13952);
and U14343 (N_14343,N_13846,N_13288);
and U14344 (N_14344,N_13438,N_13454);
or U14345 (N_14345,N_13884,N_13243);
or U14346 (N_14346,N_13478,N_13124);
or U14347 (N_14347,N_13094,N_13614);
and U14348 (N_14348,N_13194,N_13386);
xnor U14349 (N_14349,N_13141,N_13944);
or U14350 (N_14350,N_13396,N_13432);
nor U14351 (N_14351,N_13715,N_13380);
or U14352 (N_14352,N_13334,N_13308);
and U14353 (N_14353,N_13541,N_13603);
and U14354 (N_14354,N_13370,N_13577);
and U14355 (N_14355,N_13480,N_13774);
or U14356 (N_14356,N_13699,N_13915);
nor U14357 (N_14357,N_13652,N_13467);
and U14358 (N_14358,N_13090,N_13484);
xor U14359 (N_14359,N_13502,N_13766);
or U14360 (N_14360,N_13535,N_13638);
nor U14361 (N_14361,N_13449,N_13041);
and U14362 (N_14362,N_13455,N_13004);
xor U14363 (N_14363,N_13388,N_13392);
xnor U14364 (N_14364,N_13071,N_13507);
or U14365 (N_14365,N_13154,N_13860);
nor U14366 (N_14366,N_13877,N_13293);
or U14367 (N_14367,N_13435,N_13907);
and U14368 (N_14368,N_13103,N_13475);
and U14369 (N_14369,N_13913,N_13062);
nor U14370 (N_14370,N_13825,N_13241);
nor U14371 (N_14371,N_13236,N_13666);
or U14372 (N_14372,N_13657,N_13648);
or U14373 (N_14373,N_13409,N_13329);
and U14374 (N_14374,N_13561,N_13761);
and U14375 (N_14375,N_13888,N_13822);
or U14376 (N_14376,N_13412,N_13879);
nand U14377 (N_14377,N_13858,N_13527);
nand U14378 (N_14378,N_13316,N_13594);
or U14379 (N_14379,N_13669,N_13781);
nand U14380 (N_14380,N_13929,N_13492);
xor U14381 (N_14381,N_13752,N_13181);
and U14382 (N_14382,N_13442,N_13052);
nor U14383 (N_14383,N_13743,N_13224);
nand U14384 (N_14384,N_13960,N_13074);
nor U14385 (N_14385,N_13371,N_13707);
and U14386 (N_14386,N_13753,N_13728);
nand U14387 (N_14387,N_13721,N_13264);
xor U14388 (N_14388,N_13741,N_13606);
nor U14389 (N_14389,N_13152,N_13221);
nor U14390 (N_14390,N_13290,N_13732);
xnor U14391 (N_14391,N_13593,N_13482);
nor U14392 (N_14392,N_13542,N_13439);
or U14393 (N_14393,N_13322,N_13692);
or U14394 (N_14394,N_13006,N_13804);
or U14395 (N_14395,N_13620,N_13763);
or U14396 (N_14396,N_13549,N_13839);
and U14397 (N_14397,N_13000,N_13959);
and U14398 (N_14398,N_13956,N_13147);
nand U14399 (N_14399,N_13831,N_13479);
nand U14400 (N_14400,N_13275,N_13355);
and U14401 (N_14401,N_13056,N_13815);
nand U14402 (N_14402,N_13431,N_13137);
nor U14403 (N_14403,N_13414,N_13143);
nand U14404 (N_14404,N_13282,N_13434);
or U14405 (N_14405,N_13036,N_13506);
nand U14406 (N_14406,N_13824,N_13259);
nor U14407 (N_14407,N_13524,N_13294);
nand U14408 (N_14408,N_13187,N_13222);
xor U14409 (N_14409,N_13779,N_13989);
xor U14410 (N_14410,N_13819,N_13866);
nor U14411 (N_14411,N_13218,N_13310);
or U14412 (N_14412,N_13590,N_13700);
and U14413 (N_14413,N_13330,N_13254);
or U14414 (N_14414,N_13436,N_13644);
nand U14415 (N_14415,N_13808,N_13782);
nor U14416 (N_14416,N_13662,N_13697);
or U14417 (N_14417,N_13940,N_13440);
or U14418 (N_14418,N_13069,N_13610);
or U14419 (N_14419,N_13920,N_13580);
and U14420 (N_14420,N_13189,N_13835);
nand U14421 (N_14421,N_13048,N_13677);
nor U14422 (N_14422,N_13505,N_13828);
or U14423 (N_14423,N_13523,N_13405);
nor U14424 (N_14424,N_13136,N_13015);
or U14425 (N_14425,N_13625,N_13906);
and U14426 (N_14426,N_13925,N_13091);
or U14427 (N_14427,N_13341,N_13919);
nand U14428 (N_14428,N_13022,N_13982);
nand U14429 (N_14429,N_13085,N_13710);
nand U14430 (N_14430,N_13466,N_13267);
nand U14431 (N_14431,N_13578,N_13462);
nor U14432 (N_14432,N_13372,N_13564);
nand U14433 (N_14433,N_13525,N_13024);
and U14434 (N_14434,N_13331,N_13591);
or U14435 (N_14435,N_13426,N_13373);
nor U14436 (N_14436,N_13067,N_13874);
nor U14437 (N_14437,N_13805,N_13451);
nand U14438 (N_14438,N_13987,N_13144);
nor U14439 (N_14439,N_13820,N_13967);
xnor U14440 (N_14440,N_13997,N_13051);
or U14441 (N_14441,N_13563,N_13651);
nor U14442 (N_14442,N_13990,N_13533);
or U14443 (N_14443,N_13283,N_13830);
nor U14444 (N_14444,N_13010,N_13219);
or U14445 (N_14445,N_13712,N_13601);
or U14446 (N_14446,N_13909,N_13018);
xor U14447 (N_14447,N_13257,N_13360);
nand U14448 (N_14448,N_13176,N_13887);
or U14449 (N_14449,N_13838,N_13556);
nand U14450 (N_14450,N_13276,N_13622);
nand U14451 (N_14451,N_13320,N_13691);
and U14452 (N_14452,N_13476,N_13517);
xor U14453 (N_14453,N_13862,N_13382);
and U14454 (N_14454,N_13799,N_13337);
nand U14455 (N_14455,N_13099,N_13012);
or U14456 (N_14456,N_13175,N_13156);
or U14457 (N_14457,N_13511,N_13922);
xnor U14458 (N_14458,N_13786,N_13351);
or U14459 (N_14459,N_13089,N_13939);
or U14460 (N_14460,N_13718,N_13494);
nand U14461 (N_14461,N_13616,N_13206);
nand U14462 (N_14462,N_13042,N_13744);
nor U14463 (N_14463,N_13025,N_13248);
nor U14464 (N_14464,N_13108,N_13385);
nand U14465 (N_14465,N_13758,N_13871);
nor U14466 (N_14466,N_13217,N_13841);
or U14467 (N_14467,N_13497,N_13837);
or U14468 (N_14468,N_13299,N_13145);
xnor U14469 (N_14469,N_13853,N_13596);
nor U14470 (N_14470,N_13790,N_13192);
and U14471 (N_14471,N_13534,N_13274);
nand U14472 (N_14472,N_13900,N_13358);
nand U14473 (N_14473,N_13343,N_13991);
or U14474 (N_14474,N_13084,N_13366);
xor U14475 (N_14475,N_13307,N_13445);
and U14476 (N_14476,N_13674,N_13033);
or U14477 (N_14477,N_13035,N_13568);
and U14478 (N_14478,N_13560,N_13379);
nor U14479 (N_14479,N_13019,N_13083);
and U14480 (N_14480,N_13996,N_13352);
xor U14481 (N_14481,N_13641,N_13273);
or U14482 (N_14482,N_13001,N_13889);
and U14483 (N_14483,N_13968,N_13481);
nand U14484 (N_14484,N_13747,N_13617);
or U14485 (N_14485,N_13460,N_13026);
nand U14486 (N_14486,N_13910,N_13708);
nor U14487 (N_14487,N_13518,N_13302);
or U14488 (N_14488,N_13368,N_13899);
and U14489 (N_14489,N_13452,N_13709);
nor U14490 (N_14490,N_13778,N_13613);
nor U14491 (N_14491,N_13160,N_13946);
nand U14492 (N_14492,N_13840,N_13980);
nor U14493 (N_14493,N_13073,N_13773);
nor U14494 (N_14494,N_13754,N_13686);
and U14495 (N_14495,N_13117,N_13407);
nor U14496 (N_14496,N_13504,N_13443);
and U14497 (N_14497,N_13977,N_13749);
and U14498 (N_14498,N_13472,N_13512);
and U14499 (N_14499,N_13969,N_13716);
nand U14500 (N_14500,N_13919,N_13221);
or U14501 (N_14501,N_13040,N_13921);
or U14502 (N_14502,N_13744,N_13560);
or U14503 (N_14503,N_13364,N_13487);
nand U14504 (N_14504,N_13996,N_13791);
and U14505 (N_14505,N_13771,N_13520);
or U14506 (N_14506,N_13352,N_13411);
nand U14507 (N_14507,N_13917,N_13762);
and U14508 (N_14508,N_13769,N_13267);
or U14509 (N_14509,N_13272,N_13473);
and U14510 (N_14510,N_13047,N_13943);
nand U14511 (N_14511,N_13277,N_13100);
nor U14512 (N_14512,N_13726,N_13645);
nor U14513 (N_14513,N_13626,N_13816);
or U14514 (N_14514,N_13532,N_13121);
or U14515 (N_14515,N_13067,N_13103);
xnor U14516 (N_14516,N_13583,N_13928);
or U14517 (N_14517,N_13813,N_13426);
nor U14518 (N_14518,N_13563,N_13156);
xnor U14519 (N_14519,N_13266,N_13202);
nand U14520 (N_14520,N_13236,N_13796);
nand U14521 (N_14521,N_13931,N_13807);
nand U14522 (N_14522,N_13813,N_13321);
nand U14523 (N_14523,N_13270,N_13772);
nand U14524 (N_14524,N_13897,N_13964);
or U14525 (N_14525,N_13792,N_13797);
and U14526 (N_14526,N_13417,N_13603);
nor U14527 (N_14527,N_13885,N_13415);
nor U14528 (N_14528,N_13989,N_13975);
nand U14529 (N_14529,N_13703,N_13631);
and U14530 (N_14530,N_13369,N_13345);
or U14531 (N_14531,N_13880,N_13376);
or U14532 (N_14532,N_13184,N_13920);
and U14533 (N_14533,N_13250,N_13480);
or U14534 (N_14534,N_13302,N_13732);
nand U14535 (N_14535,N_13562,N_13904);
and U14536 (N_14536,N_13712,N_13980);
and U14537 (N_14537,N_13509,N_13504);
nand U14538 (N_14538,N_13130,N_13676);
nand U14539 (N_14539,N_13242,N_13398);
or U14540 (N_14540,N_13279,N_13088);
or U14541 (N_14541,N_13683,N_13335);
nand U14542 (N_14542,N_13725,N_13131);
or U14543 (N_14543,N_13389,N_13275);
or U14544 (N_14544,N_13944,N_13440);
and U14545 (N_14545,N_13320,N_13058);
or U14546 (N_14546,N_13956,N_13712);
or U14547 (N_14547,N_13625,N_13230);
nor U14548 (N_14548,N_13530,N_13228);
or U14549 (N_14549,N_13243,N_13857);
xnor U14550 (N_14550,N_13659,N_13469);
nor U14551 (N_14551,N_13645,N_13761);
nand U14552 (N_14552,N_13502,N_13311);
and U14553 (N_14553,N_13142,N_13852);
nor U14554 (N_14554,N_13982,N_13291);
and U14555 (N_14555,N_13764,N_13128);
or U14556 (N_14556,N_13196,N_13308);
or U14557 (N_14557,N_13089,N_13288);
nand U14558 (N_14558,N_13733,N_13926);
or U14559 (N_14559,N_13996,N_13251);
nor U14560 (N_14560,N_13119,N_13841);
nor U14561 (N_14561,N_13356,N_13278);
nor U14562 (N_14562,N_13521,N_13373);
nor U14563 (N_14563,N_13709,N_13825);
nand U14564 (N_14564,N_13240,N_13585);
or U14565 (N_14565,N_13990,N_13871);
or U14566 (N_14566,N_13580,N_13490);
and U14567 (N_14567,N_13274,N_13346);
and U14568 (N_14568,N_13280,N_13840);
nor U14569 (N_14569,N_13708,N_13320);
and U14570 (N_14570,N_13701,N_13843);
nand U14571 (N_14571,N_13642,N_13346);
or U14572 (N_14572,N_13218,N_13375);
nor U14573 (N_14573,N_13544,N_13022);
nor U14574 (N_14574,N_13768,N_13061);
or U14575 (N_14575,N_13392,N_13421);
nor U14576 (N_14576,N_13486,N_13137);
nor U14577 (N_14577,N_13288,N_13536);
and U14578 (N_14578,N_13383,N_13317);
or U14579 (N_14579,N_13699,N_13045);
nand U14580 (N_14580,N_13795,N_13982);
nand U14581 (N_14581,N_13608,N_13485);
nand U14582 (N_14582,N_13387,N_13774);
or U14583 (N_14583,N_13278,N_13887);
xnor U14584 (N_14584,N_13820,N_13529);
and U14585 (N_14585,N_13737,N_13149);
and U14586 (N_14586,N_13255,N_13775);
nand U14587 (N_14587,N_13185,N_13242);
or U14588 (N_14588,N_13948,N_13142);
nand U14589 (N_14589,N_13629,N_13234);
and U14590 (N_14590,N_13663,N_13328);
or U14591 (N_14591,N_13068,N_13435);
xor U14592 (N_14592,N_13929,N_13430);
and U14593 (N_14593,N_13336,N_13836);
nor U14594 (N_14594,N_13799,N_13366);
nand U14595 (N_14595,N_13534,N_13161);
and U14596 (N_14596,N_13496,N_13260);
or U14597 (N_14597,N_13248,N_13747);
and U14598 (N_14598,N_13290,N_13382);
or U14599 (N_14599,N_13100,N_13737);
or U14600 (N_14600,N_13978,N_13769);
and U14601 (N_14601,N_13360,N_13687);
or U14602 (N_14602,N_13743,N_13759);
nand U14603 (N_14603,N_13970,N_13304);
nor U14604 (N_14604,N_13577,N_13906);
or U14605 (N_14605,N_13731,N_13725);
or U14606 (N_14606,N_13639,N_13289);
or U14607 (N_14607,N_13298,N_13002);
and U14608 (N_14608,N_13318,N_13628);
or U14609 (N_14609,N_13102,N_13890);
xnor U14610 (N_14610,N_13984,N_13740);
nand U14611 (N_14611,N_13507,N_13208);
and U14612 (N_14612,N_13394,N_13445);
or U14613 (N_14613,N_13471,N_13195);
nor U14614 (N_14614,N_13232,N_13956);
or U14615 (N_14615,N_13661,N_13872);
or U14616 (N_14616,N_13105,N_13184);
and U14617 (N_14617,N_13420,N_13442);
nand U14618 (N_14618,N_13417,N_13276);
nand U14619 (N_14619,N_13929,N_13420);
nand U14620 (N_14620,N_13536,N_13388);
or U14621 (N_14621,N_13975,N_13671);
nand U14622 (N_14622,N_13843,N_13904);
xor U14623 (N_14623,N_13510,N_13543);
and U14624 (N_14624,N_13661,N_13044);
or U14625 (N_14625,N_13933,N_13565);
and U14626 (N_14626,N_13849,N_13507);
nand U14627 (N_14627,N_13692,N_13597);
or U14628 (N_14628,N_13351,N_13511);
or U14629 (N_14629,N_13337,N_13123);
nand U14630 (N_14630,N_13010,N_13581);
or U14631 (N_14631,N_13651,N_13482);
or U14632 (N_14632,N_13521,N_13636);
nor U14633 (N_14633,N_13540,N_13622);
nor U14634 (N_14634,N_13704,N_13732);
nand U14635 (N_14635,N_13886,N_13334);
xor U14636 (N_14636,N_13738,N_13099);
or U14637 (N_14637,N_13904,N_13026);
or U14638 (N_14638,N_13618,N_13824);
and U14639 (N_14639,N_13373,N_13034);
nand U14640 (N_14640,N_13054,N_13578);
nor U14641 (N_14641,N_13366,N_13437);
nand U14642 (N_14642,N_13118,N_13925);
and U14643 (N_14643,N_13565,N_13183);
nor U14644 (N_14644,N_13281,N_13830);
nor U14645 (N_14645,N_13042,N_13934);
nor U14646 (N_14646,N_13835,N_13092);
xnor U14647 (N_14647,N_13179,N_13979);
nand U14648 (N_14648,N_13937,N_13349);
nor U14649 (N_14649,N_13701,N_13000);
or U14650 (N_14650,N_13236,N_13988);
nand U14651 (N_14651,N_13965,N_13602);
nand U14652 (N_14652,N_13576,N_13610);
nand U14653 (N_14653,N_13638,N_13842);
nand U14654 (N_14654,N_13412,N_13628);
and U14655 (N_14655,N_13373,N_13608);
nand U14656 (N_14656,N_13277,N_13933);
nor U14657 (N_14657,N_13200,N_13981);
nor U14658 (N_14658,N_13829,N_13874);
and U14659 (N_14659,N_13970,N_13244);
and U14660 (N_14660,N_13448,N_13554);
nor U14661 (N_14661,N_13433,N_13375);
and U14662 (N_14662,N_13612,N_13714);
or U14663 (N_14663,N_13058,N_13770);
nand U14664 (N_14664,N_13370,N_13013);
xnor U14665 (N_14665,N_13942,N_13576);
or U14666 (N_14666,N_13665,N_13603);
or U14667 (N_14667,N_13204,N_13886);
nand U14668 (N_14668,N_13893,N_13042);
nor U14669 (N_14669,N_13332,N_13757);
nand U14670 (N_14670,N_13477,N_13337);
nand U14671 (N_14671,N_13803,N_13225);
or U14672 (N_14672,N_13557,N_13525);
and U14673 (N_14673,N_13850,N_13966);
nor U14674 (N_14674,N_13590,N_13445);
nand U14675 (N_14675,N_13124,N_13200);
nor U14676 (N_14676,N_13084,N_13727);
and U14677 (N_14677,N_13544,N_13536);
nand U14678 (N_14678,N_13033,N_13920);
or U14679 (N_14679,N_13289,N_13061);
xnor U14680 (N_14680,N_13028,N_13776);
or U14681 (N_14681,N_13651,N_13095);
and U14682 (N_14682,N_13104,N_13106);
nor U14683 (N_14683,N_13612,N_13403);
nand U14684 (N_14684,N_13502,N_13132);
or U14685 (N_14685,N_13188,N_13668);
nand U14686 (N_14686,N_13947,N_13901);
nand U14687 (N_14687,N_13813,N_13430);
nand U14688 (N_14688,N_13947,N_13413);
or U14689 (N_14689,N_13910,N_13105);
nor U14690 (N_14690,N_13127,N_13362);
nor U14691 (N_14691,N_13124,N_13139);
and U14692 (N_14692,N_13033,N_13704);
xnor U14693 (N_14693,N_13450,N_13397);
nand U14694 (N_14694,N_13025,N_13087);
or U14695 (N_14695,N_13939,N_13155);
or U14696 (N_14696,N_13912,N_13326);
nand U14697 (N_14697,N_13967,N_13644);
nand U14698 (N_14698,N_13536,N_13652);
nor U14699 (N_14699,N_13717,N_13879);
nor U14700 (N_14700,N_13123,N_13324);
or U14701 (N_14701,N_13701,N_13683);
nor U14702 (N_14702,N_13603,N_13862);
nand U14703 (N_14703,N_13701,N_13862);
nor U14704 (N_14704,N_13342,N_13931);
and U14705 (N_14705,N_13392,N_13412);
nand U14706 (N_14706,N_13268,N_13656);
nor U14707 (N_14707,N_13325,N_13696);
nand U14708 (N_14708,N_13963,N_13856);
or U14709 (N_14709,N_13621,N_13197);
or U14710 (N_14710,N_13495,N_13728);
and U14711 (N_14711,N_13424,N_13922);
nand U14712 (N_14712,N_13041,N_13917);
and U14713 (N_14713,N_13116,N_13347);
or U14714 (N_14714,N_13408,N_13379);
and U14715 (N_14715,N_13822,N_13655);
or U14716 (N_14716,N_13027,N_13707);
nor U14717 (N_14717,N_13496,N_13063);
or U14718 (N_14718,N_13618,N_13227);
nand U14719 (N_14719,N_13508,N_13154);
nand U14720 (N_14720,N_13554,N_13362);
nor U14721 (N_14721,N_13547,N_13568);
or U14722 (N_14722,N_13416,N_13156);
and U14723 (N_14723,N_13525,N_13444);
nor U14724 (N_14724,N_13867,N_13236);
nor U14725 (N_14725,N_13768,N_13606);
xnor U14726 (N_14726,N_13083,N_13302);
or U14727 (N_14727,N_13980,N_13304);
nand U14728 (N_14728,N_13008,N_13368);
or U14729 (N_14729,N_13525,N_13054);
nand U14730 (N_14730,N_13473,N_13031);
xnor U14731 (N_14731,N_13574,N_13420);
or U14732 (N_14732,N_13402,N_13794);
nor U14733 (N_14733,N_13955,N_13236);
and U14734 (N_14734,N_13864,N_13497);
nand U14735 (N_14735,N_13203,N_13361);
xnor U14736 (N_14736,N_13322,N_13151);
nor U14737 (N_14737,N_13444,N_13725);
and U14738 (N_14738,N_13194,N_13770);
or U14739 (N_14739,N_13686,N_13042);
and U14740 (N_14740,N_13218,N_13221);
nor U14741 (N_14741,N_13733,N_13275);
or U14742 (N_14742,N_13842,N_13087);
or U14743 (N_14743,N_13026,N_13922);
or U14744 (N_14744,N_13237,N_13374);
nand U14745 (N_14745,N_13471,N_13394);
and U14746 (N_14746,N_13797,N_13179);
xor U14747 (N_14747,N_13170,N_13461);
nand U14748 (N_14748,N_13903,N_13316);
nor U14749 (N_14749,N_13201,N_13282);
or U14750 (N_14750,N_13876,N_13970);
nor U14751 (N_14751,N_13437,N_13546);
or U14752 (N_14752,N_13442,N_13136);
nand U14753 (N_14753,N_13428,N_13328);
or U14754 (N_14754,N_13044,N_13140);
and U14755 (N_14755,N_13194,N_13969);
or U14756 (N_14756,N_13265,N_13296);
nor U14757 (N_14757,N_13494,N_13235);
nand U14758 (N_14758,N_13060,N_13048);
xor U14759 (N_14759,N_13808,N_13866);
nor U14760 (N_14760,N_13489,N_13256);
nand U14761 (N_14761,N_13729,N_13669);
or U14762 (N_14762,N_13069,N_13875);
or U14763 (N_14763,N_13478,N_13876);
xnor U14764 (N_14764,N_13656,N_13453);
and U14765 (N_14765,N_13769,N_13944);
xnor U14766 (N_14766,N_13096,N_13010);
xnor U14767 (N_14767,N_13261,N_13040);
and U14768 (N_14768,N_13069,N_13906);
xnor U14769 (N_14769,N_13022,N_13123);
xnor U14770 (N_14770,N_13908,N_13880);
nor U14771 (N_14771,N_13070,N_13758);
nand U14772 (N_14772,N_13415,N_13709);
nor U14773 (N_14773,N_13204,N_13806);
and U14774 (N_14774,N_13026,N_13481);
nor U14775 (N_14775,N_13027,N_13343);
nand U14776 (N_14776,N_13361,N_13623);
nand U14777 (N_14777,N_13376,N_13025);
nor U14778 (N_14778,N_13837,N_13030);
and U14779 (N_14779,N_13940,N_13345);
or U14780 (N_14780,N_13981,N_13278);
and U14781 (N_14781,N_13143,N_13707);
xor U14782 (N_14782,N_13214,N_13853);
or U14783 (N_14783,N_13309,N_13782);
nor U14784 (N_14784,N_13043,N_13982);
nand U14785 (N_14785,N_13823,N_13212);
nor U14786 (N_14786,N_13732,N_13359);
or U14787 (N_14787,N_13878,N_13889);
and U14788 (N_14788,N_13224,N_13897);
and U14789 (N_14789,N_13998,N_13135);
and U14790 (N_14790,N_13686,N_13348);
nor U14791 (N_14791,N_13541,N_13476);
nor U14792 (N_14792,N_13999,N_13063);
nor U14793 (N_14793,N_13878,N_13067);
and U14794 (N_14794,N_13129,N_13188);
or U14795 (N_14795,N_13044,N_13350);
or U14796 (N_14796,N_13154,N_13986);
or U14797 (N_14797,N_13906,N_13126);
and U14798 (N_14798,N_13260,N_13108);
nor U14799 (N_14799,N_13392,N_13144);
or U14800 (N_14800,N_13836,N_13952);
or U14801 (N_14801,N_13941,N_13944);
nor U14802 (N_14802,N_13732,N_13294);
and U14803 (N_14803,N_13470,N_13254);
nor U14804 (N_14804,N_13879,N_13601);
nand U14805 (N_14805,N_13141,N_13964);
or U14806 (N_14806,N_13365,N_13647);
or U14807 (N_14807,N_13284,N_13975);
nand U14808 (N_14808,N_13892,N_13037);
or U14809 (N_14809,N_13444,N_13577);
or U14810 (N_14810,N_13282,N_13445);
and U14811 (N_14811,N_13485,N_13049);
or U14812 (N_14812,N_13390,N_13229);
nor U14813 (N_14813,N_13327,N_13608);
nor U14814 (N_14814,N_13830,N_13406);
nor U14815 (N_14815,N_13285,N_13260);
nand U14816 (N_14816,N_13009,N_13930);
and U14817 (N_14817,N_13988,N_13759);
nand U14818 (N_14818,N_13146,N_13982);
nor U14819 (N_14819,N_13430,N_13712);
and U14820 (N_14820,N_13006,N_13863);
and U14821 (N_14821,N_13016,N_13063);
or U14822 (N_14822,N_13403,N_13804);
and U14823 (N_14823,N_13642,N_13749);
or U14824 (N_14824,N_13019,N_13393);
nor U14825 (N_14825,N_13337,N_13092);
nand U14826 (N_14826,N_13881,N_13739);
or U14827 (N_14827,N_13770,N_13661);
and U14828 (N_14828,N_13413,N_13837);
nor U14829 (N_14829,N_13283,N_13983);
nand U14830 (N_14830,N_13710,N_13866);
nand U14831 (N_14831,N_13311,N_13965);
or U14832 (N_14832,N_13386,N_13321);
and U14833 (N_14833,N_13265,N_13207);
or U14834 (N_14834,N_13963,N_13206);
nor U14835 (N_14835,N_13758,N_13207);
and U14836 (N_14836,N_13449,N_13558);
nor U14837 (N_14837,N_13431,N_13427);
nor U14838 (N_14838,N_13456,N_13259);
or U14839 (N_14839,N_13767,N_13976);
nand U14840 (N_14840,N_13944,N_13710);
nor U14841 (N_14841,N_13390,N_13358);
and U14842 (N_14842,N_13295,N_13820);
and U14843 (N_14843,N_13881,N_13906);
nor U14844 (N_14844,N_13709,N_13654);
xor U14845 (N_14845,N_13289,N_13980);
and U14846 (N_14846,N_13829,N_13298);
nand U14847 (N_14847,N_13153,N_13728);
and U14848 (N_14848,N_13506,N_13609);
or U14849 (N_14849,N_13274,N_13843);
and U14850 (N_14850,N_13390,N_13935);
and U14851 (N_14851,N_13816,N_13502);
and U14852 (N_14852,N_13579,N_13818);
or U14853 (N_14853,N_13187,N_13553);
or U14854 (N_14854,N_13277,N_13839);
and U14855 (N_14855,N_13776,N_13073);
and U14856 (N_14856,N_13860,N_13588);
xnor U14857 (N_14857,N_13492,N_13420);
and U14858 (N_14858,N_13563,N_13021);
xor U14859 (N_14859,N_13296,N_13266);
nor U14860 (N_14860,N_13491,N_13270);
and U14861 (N_14861,N_13593,N_13746);
nor U14862 (N_14862,N_13931,N_13895);
and U14863 (N_14863,N_13352,N_13990);
nor U14864 (N_14864,N_13741,N_13374);
or U14865 (N_14865,N_13340,N_13349);
nand U14866 (N_14866,N_13079,N_13891);
and U14867 (N_14867,N_13186,N_13052);
and U14868 (N_14868,N_13288,N_13891);
nand U14869 (N_14869,N_13801,N_13455);
or U14870 (N_14870,N_13915,N_13865);
and U14871 (N_14871,N_13681,N_13385);
or U14872 (N_14872,N_13572,N_13138);
nand U14873 (N_14873,N_13136,N_13232);
nor U14874 (N_14874,N_13635,N_13548);
or U14875 (N_14875,N_13971,N_13007);
or U14876 (N_14876,N_13390,N_13806);
nor U14877 (N_14877,N_13336,N_13745);
nand U14878 (N_14878,N_13905,N_13883);
nor U14879 (N_14879,N_13482,N_13908);
and U14880 (N_14880,N_13063,N_13871);
xnor U14881 (N_14881,N_13435,N_13077);
xor U14882 (N_14882,N_13861,N_13342);
or U14883 (N_14883,N_13073,N_13487);
or U14884 (N_14884,N_13386,N_13693);
nor U14885 (N_14885,N_13280,N_13806);
and U14886 (N_14886,N_13289,N_13741);
or U14887 (N_14887,N_13623,N_13542);
or U14888 (N_14888,N_13967,N_13522);
and U14889 (N_14889,N_13434,N_13475);
nand U14890 (N_14890,N_13141,N_13990);
nor U14891 (N_14891,N_13199,N_13050);
or U14892 (N_14892,N_13842,N_13290);
and U14893 (N_14893,N_13236,N_13139);
or U14894 (N_14894,N_13950,N_13240);
and U14895 (N_14895,N_13991,N_13470);
or U14896 (N_14896,N_13312,N_13591);
nand U14897 (N_14897,N_13134,N_13670);
or U14898 (N_14898,N_13828,N_13671);
and U14899 (N_14899,N_13478,N_13395);
or U14900 (N_14900,N_13374,N_13207);
xnor U14901 (N_14901,N_13279,N_13675);
nand U14902 (N_14902,N_13714,N_13839);
and U14903 (N_14903,N_13738,N_13529);
and U14904 (N_14904,N_13245,N_13434);
xor U14905 (N_14905,N_13478,N_13316);
xnor U14906 (N_14906,N_13972,N_13984);
nor U14907 (N_14907,N_13093,N_13731);
xor U14908 (N_14908,N_13616,N_13330);
nand U14909 (N_14909,N_13384,N_13045);
nor U14910 (N_14910,N_13227,N_13717);
or U14911 (N_14911,N_13023,N_13482);
nand U14912 (N_14912,N_13192,N_13298);
and U14913 (N_14913,N_13489,N_13693);
or U14914 (N_14914,N_13088,N_13190);
xor U14915 (N_14915,N_13430,N_13249);
xnor U14916 (N_14916,N_13609,N_13435);
and U14917 (N_14917,N_13188,N_13286);
nor U14918 (N_14918,N_13004,N_13710);
xnor U14919 (N_14919,N_13332,N_13539);
or U14920 (N_14920,N_13317,N_13291);
nor U14921 (N_14921,N_13002,N_13834);
xnor U14922 (N_14922,N_13146,N_13020);
nand U14923 (N_14923,N_13724,N_13066);
and U14924 (N_14924,N_13315,N_13844);
xnor U14925 (N_14925,N_13744,N_13106);
nand U14926 (N_14926,N_13507,N_13098);
nor U14927 (N_14927,N_13881,N_13121);
nand U14928 (N_14928,N_13222,N_13071);
or U14929 (N_14929,N_13445,N_13274);
and U14930 (N_14930,N_13077,N_13880);
nor U14931 (N_14931,N_13252,N_13643);
nand U14932 (N_14932,N_13661,N_13667);
nor U14933 (N_14933,N_13866,N_13352);
xnor U14934 (N_14934,N_13510,N_13324);
and U14935 (N_14935,N_13519,N_13497);
or U14936 (N_14936,N_13665,N_13374);
nor U14937 (N_14937,N_13779,N_13706);
nand U14938 (N_14938,N_13764,N_13260);
xnor U14939 (N_14939,N_13030,N_13554);
nor U14940 (N_14940,N_13516,N_13375);
xor U14941 (N_14941,N_13966,N_13252);
nand U14942 (N_14942,N_13343,N_13407);
nand U14943 (N_14943,N_13680,N_13433);
nor U14944 (N_14944,N_13404,N_13612);
or U14945 (N_14945,N_13806,N_13992);
or U14946 (N_14946,N_13632,N_13990);
nor U14947 (N_14947,N_13842,N_13939);
or U14948 (N_14948,N_13024,N_13415);
xor U14949 (N_14949,N_13189,N_13479);
nor U14950 (N_14950,N_13641,N_13142);
or U14951 (N_14951,N_13487,N_13027);
nand U14952 (N_14952,N_13373,N_13780);
nor U14953 (N_14953,N_13153,N_13806);
xor U14954 (N_14954,N_13439,N_13374);
nor U14955 (N_14955,N_13748,N_13913);
and U14956 (N_14956,N_13169,N_13487);
or U14957 (N_14957,N_13112,N_13859);
and U14958 (N_14958,N_13240,N_13489);
xor U14959 (N_14959,N_13574,N_13097);
xor U14960 (N_14960,N_13830,N_13270);
nor U14961 (N_14961,N_13984,N_13563);
nand U14962 (N_14962,N_13955,N_13372);
xor U14963 (N_14963,N_13286,N_13088);
nand U14964 (N_14964,N_13052,N_13017);
and U14965 (N_14965,N_13688,N_13604);
nor U14966 (N_14966,N_13727,N_13895);
and U14967 (N_14967,N_13409,N_13331);
or U14968 (N_14968,N_13768,N_13107);
and U14969 (N_14969,N_13023,N_13261);
or U14970 (N_14970,N_13981,N_13415);
or U14971 (N_14971,N_13073,N_13093);
nor U14972 (N_14972,N_13404,N_13616);
nor U14973 (N_14973,N_13516,N_13704);
and U14974 (N_14974,N_13872,N_13861);
and U14975 (N_14975,N_13264,N_13366);
and U14976 (N_14976,N_13585,N_13467);
nand U14977 (N_14977,N_13128,N_13268);
and U14978 (N_14978,N_13343,N_13560);
nand U14979 (N_14979,N_13691,N_13882);
or U14980 (N_14980,N_13832,N_13909);
or U14981 (N_14981,N_13023,N_13227);
and U14982 (N_14982,N_13303,N_13899);
or U14983 (N_14983,N_13285,N_13163);
and U14984 (N_14984,N_13064,N_13570);
or U14985 (N_14985,N_13319,N_13857);
nor U14986 (N_14986,N_13483,N_13500);
or U14987 (N_14987,N_13954,N_13866);
and U14988 (N_14988,N_13330,N_13492);
or U14989 (N_14989,N_13703,N_13014);
nor U14990 (N_14990,N_13880,N_13974);
nor U14991 (N_14991,N_13005,N_13436);
nor U14992 (N_14992,N_13034,N_13320);
and U14993 (N_14993,N_13495,N_13305);
or U14994 (N_14994,N_13586,N_13440);
or U14995 (N_14995,N_13694,N_13588);
nand U14996 (N_14996,N_13556,N_13856);
nor U14997 (N_14997,N_13751,N_13508);
nor U14998 (N_14998,N_13056,N_13800);
and U14999 (N_14999,N_13849,N_13524);
and UO_0 (O_0,N_14767,N_14155);
and UO_1 (O_1,N_14261,N_14070);
nand UO_2 (O_2,N_14896,N_14209);
nand UO_3 (O_3,N_14804,N_14172);
or UO_4 (O_4,N_14302,N_14388);
or UO_5 (O_5,N_14967,N_14222);
or UO_6 (O_6,N_14174,N_14837);
xor UO_7 (O_7,N_14753,N_14688);
nor UO_8 (O_8,N_14941,N_14642);
nor UO_9 (O_9,N_14267,N_14186);
and UO_10 (O_10,N_14255,N_14788);
nand UO_11 (O_11,N_14615,N_14614);
nor UO_12 (O_12,N_14796,N_14276);
nand UO_13 (O_13,N_14204,N_14177);
and UO_14 (O_14,N_14921,N_14441);
and UO_15 (O_15,N_14666,N_14589);
or UO_16 (O_16,N_14021,N_14555);
or UO_17 (O_17,N_14048,N_14569);
nor UO_18 (O_18,N_14041,N_14827);
or UO_19 (O_19,N_14558,N_14727);
or UO_20 (O_20,N_14277,N_14907);
or UO_21 (O_21,N_14023,N_14774);
nand UO_22 (O_22,N_14449,N_14259);
or UO_23 (O_23,N_14624,N_14805);
and UO_24 (O_24,N_14918,N_14932);
or UO_25 (O_25,N_14447,N_14761);
and UO_26 (O_26,N_14817,N_14996);
and UO_27 (O_27,N_14578,N_14143);
nand UO_28 (O_28,N_14892,N_14163);
and UO_29 (O_29,N_14752,N_14110);
or UO_30 (O_30,N_14438,N_14469);
xnor UO_31 (O_31,N_14972,N_14787);
and UO_32 (O_32,N_14819,N_14062);
and UO_33 (O_33,N_14178,N_14218);
nor UO_34 (O_34,N_14146,N_14510);
and UO_35 (O_35,N_14842,N_14610);
and UO_36 (O_36,N_14889,N_14124);
nand UO_37 (O_37,N_14282,N_14310);
and UO_38 (O_38,N_14010,N_14518);
xor UO_39 (O_39,N_14173,N_14563);
and UO_40 (O_40,N_14106,N_14989);
nor UO_41 (O_41,N_14237,N_14185);
and UO_42 (O_42,N_14170,N_14613);
nor UO_43 (O_43,N_14597,N_14776);
or UO_44 (O_44,N_14730,N_14437);
and UO_45 (O_45,N_14911,N_14052);
nor UO_46 (O_46,N_14379,N_14376);
or UO_47 (O_47,N_14865,N_14870);
or UO_48 (O_48,N_14325,N_14479);
nand UO_49 (O_49,N_14579,N_14271);
xor UO_50 (O_50,N_14554,N_14364);
and UO_51 (O_51,N_14129,N_14621);
nand UO_52 (O_52,N_14335,N_14336);
or UO_53 (O_53,N_14036,N_14121);
xor UO_54 (O_54,N_14337,N_14531);
or UO_55 (O_55,N_14693,N_14927);
and UO_56 (O_56,N_14435,N_14821);
and UO_57 (O_57,N_14287,N_14883);
and UO_58 (O_58,N_14414,N_14047);
nand UO_59 (O_59,N_14694,N_14780);
nand UO_60 (O_60,N_14262,N_14368);
or UO_61 (O_61,N_14130,N_14486);
or UO_62 (O_62,N_14220,N_14734);
nand UO_63 (O_63,N_14723,N_14463);
or UO_64 (O_64,N_14851,N_14028);
nand UO_65 (O_65,N_14478,N_14898);
or UO_66 (O_66,N_14093,N_14566);
and UO_67 (O_67,N_14151,N_14369);
or UO_68 (O_68,N_14427,N_14824);
and UO_69 (O_69,N_14971,N_14659);
or UO_70 (O_70,N_14501,N_14200);
and UO_71 (O_71,N_14548,N_14656);
nor UO_72 (O_72,N_14617,N_14456);
nor UO_73 (O_73,N_14552,N_14961);
xor UO_74 (O_74,N_14061,N_14452);
and UO_75 (O_75,N_14446,N_14138);
nand UO_76 (O_76,N_14114,N_14704);
nor UO_77 (O_77,N_14349,N_14654);
or UO_78 (O_78,N_14912,N_14526);
nor UO_79 (O_79,N_14948,N_14091);
and UO_80 (O_80,N_14493,N_14326);
xor UO_81 (O_81,N_14741,N_14288);
nand UO_82 (O_82,N_14489,N_14327);
or UO_83 (O_83,N_14407,N_14886);
or UO_84 (O_84,N_14116,N_14248);
or UO_85 (O_85,N_14457,N_14131);
or UO_86 (O_86,N_14380,N_14616);
and UO_87 (O_87,N_14286,N_14721);
or UO_88 (O_88,N_14649,N_14540);
and UO_89 (O_89,N_14092,N_14958);
or UO_90 (O_90,N_14674,N_14925);
xnor UO_91 (O_91,N_14137,N_14481);
and UO_92 (O_92,N_14986,N_14076);
xor UO_93 (O_93,N_14549,N_14759);
nor UO_94 (O_94,N_14343,N_14784);
nand UO_95 (O_95,N_14133,N_14279);
nor UO_96 (O_96,N_14534,N_14754);
or UO_97 (O_97,N_14394,N_14063);
xor UO_98 (O_98,N_14987,N_14305);
nand UO_99 (O_99,N_14239,N_14082);
xnor UO_100 (O_100,N_14085,N_14645);
and UO_101 (O_101,N_14460,N_14046);
and UO_102 (O_102,N_14201,N_14722);
nor UO_103 (O_103,N_14386,N_14442);
and UO_104 (O_104,N_14525,N_14777);
or UO_105 (O_105,N_14051,N_14301);
and UO_106 (O_106,N_14652,N_14049);
nor UO_107 (O_107,N_14344,N_14322);
nor UO_108 (O_108,N_14104,N_14715);
and UO_109 (O_109,N_14221,N_14260);
nand UO_110 (O_110,N_14057,N_14791);
and UO_111 (O_111,N_14556,N_14998);
nand UO_112 (O_112,N_14852,N_14040);
nor UO_113 (O_113,N_14038,N_14888);
nor UO_114 (O_114,N_14474,N_14553);
and UO_115 (O_115,N_14572,N_14960);
or UO_116 (O_116,N_14350,N_14814);
or UO_117 (O_117,N_14347,N_14080);
nand UO_118 (O_118,N_14772,N_14696);
nor UO_119 (O_119,N_14581,N_14283);
or UO_120 (O_120,N_14874,N_14733);
xor UO_121 (O_121,N_14988,N_14296);
and UO_122 (O_122,N_14223,N_14084);
nor UO_123 (O_123,N_14194,N_14697);
or UO_124 (O_124,N_14145,N_14381);
nor UO_125 (O_125,N_14582,N_14269);
or UO_126 (O_126,N_14071,N_14630);
nand UO_127 (O_127,N_14319,N_14354);
and UO_128 (O_128,N_14862,N_14903);
or UO_129 (O_129,N_14202,N_14854);
and UO_130 (O_130,N_14933,N_14790);
or UO_131 (O_131,N_14845,N_14664);
nand UO_132 (O_132,N_14564,N_14094);
or UO_133 (O_133,N_14692,N_14901);
xnor UO_134 (O_134,N_14208,N_14400);
xnor UO_135 (O_135,N_14743,N_14669);
and UO_136 (O_136,N_14018,N_14088);
or UO_137 (O_137,N_14308,N_14915);
or UO_138 (O_138,N_14598,N_14370);
and UO_139 (O_139,N_14773,N_14686);
nand UO_140 (O_140,N_14820,N_14251);
xnor UO_141 (O_141,N_14978,N_14466);
and UO_142 (O_142,N_14087,N_14627);
xnor UO_143 (O_143,N_14858,N_14166);
or UO_144 (O_144,N_14662,N_14140);
xor UO_145 (O_145,N_14244,N_14182);
and UO_146 (O_146,N_14532,N_14984);
or UO_147 (O_147,N_14785,N_14207);
and UO_148 (O_148,N_14205,N_14801);
and UO_149 (O_149,N_14332,N_14482);
and UO_150 (O_150,N_14635,N_14517);
or UO_151 (O_151,N_14633,N_14813);
nand UO_152 (O_152,N_14789,N_14026);
or UO_153 (O_153,N_14408,N_14618);
xnor UO_154 (O_154,N_14367,N_14426);
and UO_155 (O_155,N_14410,N_14682);
nor UO_156 (O_156,N_14561,N_14003);
nor UO_157 (O_157,N_14849,N_14317);
and UO_158 (O_158,N_14853,N_14396);
and UO_159 (O_159,N_14089,N_14372);
nand UO_160 (O_160,N_14611,N_14398);
nor UO_161 (O_161,N_14968,N_14521);
nand UO_162 (O_162,N_14899,N_14663);
or UO_163 (O_163,N_14965,N_14066);
and UO_164 (O_164,N_14639,N_14011);
and UO_165 (O_165,N_14966,N_14111);
or UO_166 (O_166,N_14770,N_14815);
or UO_167 (O_167,N_14724,N_14891);
or UO_168 (O_168,N_14775,N_14544);
xor UO_169 (O_169,N_14120,N_14833);
nor UO_170 (O_170,N_14810,N_14538);
or UO_171 (O_171,N_14757,N_14751);
nor UO_172 (O_172,N_14195,N_14428);
nor UO_173 (O_173,N_14963,N_14118);
or UO_174 (O_174,N_14632,N_14991);
nand UO_175 (O_175,N_14959,N_14418);
and UO_176 (O_176,N_14389,N_14885);
nand UO_177 (O_177,N_14651,N_14339);
nand UO_178 (O_178,N_14211,N_14044);
nand UO_179 (O_179,N_14904,N_14069);
or UO_180 (O_180,N_14009,N_14878);
nand UO_181 (O_181,N_14962,N_14060);
nor UO_182 (O_182,N_14409,N_14328);
nand UO_183 (O_183,N_14705,N_14976);
nor UO_184 (O_184,N_14718,N_14828);
and UO_185 (O_185,N_14930,N_14866);
or UO_186 (O_186,N_14939,N_14744);
xor UO_187 (O_187,N_14161,N_14462);
nor UO_188 (O_188,N_14232,N_14315);
nor UO_189 (O_189,N_14760,N_14484);
xnor UO_190 (O_190,N_14545,N_14758);
and UO_191 (O_191,N_14924,N_14020);
nor UO_192 (O_192,N_14203,N_14839);
nand UO_193 (O_193,N_14077,N_14947);
nor UO_194 (O_194,N_14687,N_14808);
nand UO_195 (O_195,N_14740,N_14303);
or UO_196 (O_196,N_14516,N_14952);
nor UO_197 (O_197,N_14800,N_14969);
xnor UO_198 (O_198,N_14864,N_14459);
or UO_199 (O_199,N_14491,N_14236);
nor UO_200 (O_200,N_14811,N_14944);
and UO_201 (O_201,N_14226,N_14294);
nand UO_202 (O_202,N_14241,N_14027);
nand UO_203 (O_203,N_14887,N_14217);
or UO_204 (O_204,N_14850,N_14338);
and UO_205 (O_205,N_14951,N_14846);
xor UO_206 (O_206,N_14162,N_14703);
xor UO_207 (O_207,N_14440,N_14345);
nand UO_208 (O_208,N_14378,N_14698);
or UO_209 (O_209,N_14755,N_14494);
nor UO_210 (O_210,N_14298,N_14189);
or UO_211 (O_211,N_14519,N_14713);
or UO_212 (O_212,N_14604,N_14329);
xor UO_213 (O_213,N_14900,N_14197);
and UO_214 (O_214,N_14000,N_14206);
or UO_215 (O_215,N_14647,N_14942);
or UO_216 (O_216,N_14585,N_14530);
nor UO_217 (O_217,N_14181,N_14880);
or UO_218 (O_218,N_14711,N_14297);
or UO_219 (O_219,N_14893,N_14384);
or UO_220 (O_220,N_14096,N_14031);
nand UO_221 (O_221,N_14596,N_14979);
nor UO_222 (O_222,N_14391,N_14316);
or UO_223 (O_223,N_14567,N_14848);
nor UO_224 (O_224,N_14877,N_14745);
or UO_225 (O_225,N_14421,N_14289);
nor UO_226 (O_226,N_14480,N_14955);
and UO_227 (O_227,N_14081,N_14453);
or UO_228 (O_228,N_14629,N_14580);
nand UO_229 (O_229,N_14263,N_14333);
xnor UO_230 (O_230,N_14304,N_14716);
or UO_231 (O_231,N_14242,N_14524);
nor UO_232 (O_232,N_14926,N_14300);
xnor UO_233 (O_233,N_14679,N_14395);
nor UO_234 (O_234,N_14257,N_14461);
nand UO_235 (O_235,N_14506,N_14823);
xnor UO_236 (O_236,N_14245,N_14274);
or UO_237 (O_237,N_14809,N_14425);
nand UO_238 (O_238,N_14356,N_14358);
xor UO_239 (O_239,N_14132,N_14794);
nand UO_240 (O_240,N_14769,N_14374);
nor UO_241 (O_241,N_14861,N_14342);
nand UO_242 (O_242,N_14284,N_14415);
nor UO_243 (O_243,N_14816,N_14868);
nor UO_244 (O_244,N_14646,N_14869);
or UO_245 (O_245,N_14413,N_14065);
nor UO_246 (O_246,N_14728,N_14323);
nor UO_247 (O_247,N_14341,N_14764);
nor UO_248 (O_248,N_14830,N_14588);
nor UO_249 (O_249,N_14637,N_14500);
or UO_250 (O_250,N_14128,N_14075);
xor UO_251 (O_251,N_14024,N_14002);
nor UO_252 (O_252,N_14914,N_14475);
nand UO_253 (O_253,N_14351,N_14511);
nand UO_254 (O_254,N_14340,N_14254);
nand UO_255 (O_255,N_14055,N_14840);
nand UO_256 (O_256,N_14736,N_14292);
and UO_257 (O_257,N_14677,N_14006);
and UO_258 (O_258,N_14037,N_14643);
nand UO_259 (O_259,N_14829,N_14841);
and UO_260 (O_260,N_14247,N_14763);
or UO_261 (O_261,N_14392,N_14606);
nor UO_262 (O_262,N_14980,N_14625);
nor UO_263 (O_263,N_14600,N_14992);
and UO_264 (O_264,N_14739,N_14331);
xnor UO_265 (O_265,N_14660,N_14512);
nor UO_266 (O_266,N_14935,N_14275);
or UO_267 (O_267,N_14681,N_14224);
or UO_268 (O_268,N_14806,N_14433);
nor UO_269 (O_269,N_14265,N_14917);
or UO_270 (O_270,N_14920,N_14192);
nand UO_271 (O_271,N_14109,N_14346);
and UO_272 (O_272,N_14550,N_14235);
nand UO_273 (O_273,N_14184,N_14432);
nor UO_274 (O_274,N_14831,N_14243);
xor UO_275 (O_275,N_14836,N_14270);
nand UO_276 (O_276,N_14699,N_14802);
and UO_277 (O_277,N_14655,N_14576);
nor UO_278 (O_278,N_14875,N_14882);
or UO_279 (O_279,N_14653,N_14957);
and UO_280 (O_280,N_14467,N_14099);
and UO_281 (O_281,N_14436,N_14256);
and UO_282 (O_282,N_14196,N_14742);
and UO_283 (O_283,N_14210,N_14033);
and UO_284 (O_284,N_14190,N_14231);
and UO_285 (O_285,N_14622,N_14975);
or UO_286 (O_286,N_14108,N_14152);
and UO_287 (O_287,N_14249,N_14720);
xnor UO_288 (O_288,N_14465,N_14122);
xor UO_289 (O_289,N_14199,N_14215);
xnor UO_290 (O_290,N_14586,N_14352);
or UO_291 (O_291,N_14464,N_14357);
and UO_292 (O_292,N_14623,N_14607);
nor UO_293 (O_293,N_14826,N_14946);
xor UO_294 (O_294,N_14039,N_14136);
and UO_295 (O_295,N_14547,N_14844);
and UO_296 (O_296,N_14685,N_14495);
nand UO_297 (O_297,N_14863,N_14154);
or UO_298 (O_298,N_14719,N_14086);
nand UO_299 (O_299,N_14648,N_14107);
or UO_300 (O_300,N_14212,N_14079);
and UO_301 (O_301,N_14363,N_14631);
nand UO_302 (O_302,N_14560,N_14043);
and UO_303 (O_303,N_14726,N_14768);
and UO_304 (O_304,N_14406,N_14045);
nor UO_305 (O_305,N_14872,N_14533);
and UO_306 (O_306,N_14536,N_14451);
and UO_307 (O_307,N_14295,N_14689);
xor UO_308 (O_308,N_14090,N_14233);
nor UO_309 (O_309,N_14216,N_14311);
and UO_310 (O_310,N_14473,N_14574);
and UO_311 (O_311,N_14487,N_14291);
or UO_312 (O_312,N_14429,N_14897);
or UO_313 (O_313,N_14312,N_14034);
and UO_314 (O_314,N_14994,N_14273);
nor UO_315 (O_315,N_14568,N_14683);
nand UO_316 (O_316,N_14838,N_14619);
nand UO_317 (O_317,N_14945,N_14515);
or UO_318 (O_318,N_14101,N_14416);
or UO_319 (O_319,N_14620,N_14147);
nor UO_320 (O_320,N_14584,N_14557);
and UO_321 (O_321,N_14855,N_14505);
xor UO_322 (O_322,N_14025,N_14454);
and UO_323 (O_323,N_14470,N_14268);
nor UO_324 (O_324,N_14458,N_14492);
and UO_325 (O_325,N_14188,N_14321);
nand UO_326 (O_326,N_14701,N_14490);
nand UO_327 (O_327,N_14320,N_14970);
or UO_328 (O_328,N_14165,N_14605);
or UO_329 (O_329,N_14150,N_14562);
nand UO_330 (O_330,N_14149,N_14399);
nand UO_331 (O_331,N_14943,N_14934);
nand UO_332 (O_332,N_14671,N_14359);
nand UO_333 (O_333,N_14097,N_14799);
xnor UO_334 (O_334,N_14471,N_14906);
or UO_335 (O_335,N_14573,N_14468);
and UO_336 (O_336,N_14266,N_14765);
nand UO_337 (O_337,N_14142,N_14056);
nor UO_338 (O_338,N_14483,N_14180);
nor UO_339 (O_339,N_14164,N_14565);
nor UO_340 (O_340,N_14225,N_14832);
xor UO_341 (O_341,N_14064,N_14412);
or UO_342 (O_342,N_14382,N_14587);
and UO_343 (O_343,N_14658,N_14691);
xnor UO_344 (O_344,N_14894,N_14450);
nand UO_345 (O_345,N_14700,N_14977);
nor UO_346 (O_346,N_14529,N_14982);
nor UO_347 (O_347,N_14285,N_14419);
nor UO_348 (O_348,N_14008,N_14141);
nor UO_349 (O_349,N_14191,N_14430);
or UO_350 (O_350,N_14179,N_14153);
nor UO_351 (O_351,N_14258,N_14795);
or UO_352 (O_352,N_14923,N_14058);
nand UO_353 (O_353,N_14603,N_14019);
nor UO_354 (O_354,N_14797,N_14762);
nor UO_355 (O_355,N_14860,N_14238);
and UO_356 (O_356,N_14007,N_14158);
xnor UO_357 (O_357,N_14638,N_14135);
or UO_358 (O_358,N_14929,N_14695);
nand UO_359 (O_359,N_14405,N_14183);
nor UO_360 (O_360,N_14890,N_14909);
xnor UO_361 (O_361,N_14953,N_14876);
and UO_362 (O_362,N_14867,N_14280);
xor UO_363 (O_363,N_14667,N_14353);
nand UO_364 (O_364,N_14847,N_14042);
and UO_365 (O_365,N_14117,N_14417);
nand UO_366 (O_366,N_14910,N_14575);
or UO_367 (O_367,N_14022,N_14227);
nand UO_368 (O_368,N_14781,N_14748);
or UO_369 (O_369,N_14675,N_14067);
nand UO_370 (O_370,N_14001,N_14602);
nand UO_371 (O_371,N_14439,N_14187);
or UO_372 (O_372,N_14938,N_14485);
and UO_373 (O_373,N_14919,N_14908);
or UO_374 (O_374,N_14507,N_14176);
and UO_375 (O_375,N_14626,N_14859);
and UO_376 (O_376,N_14361,N_14825);
or UO_377 (O_377,N_14974,N_14102);
and UO_378 (O_378,N_14240,N_14595);
nor UO_379 (O_379,N_14127,N_14126);
nand UO_380 (O_380,N_14214,N_14937);
nand UO_381 (O_381,N_14148,N_14362);
or UO_382 (O_382,N_14577,N_14710);
or UO_383 (O_383,N_14306,N_14523);
or UO_384 (O_384,N_14113,N_14366);
and UO_385 (O_385,N_14431,N_14074);
xnor UO_386 (O_386,N_14676,N_14144);
and UO_387 (O_387,N_14005,N_14445);
or UO_388 (O_388,N_14193,N_14073);
nor UO_389 (O_389,N_14420,N_14375);
nor UO_390 (O_390,N_14059,N_14160);
nor UO_391 (O_391,N_14747,N_14348);
nor UO_392 (O_392,N_14657,N_14502);
nor UO_393 (O_393,N_14159,N_14404);
or UO_394 (O_394,N_14355,N_14029);
and UO_395 (O_395,N_14520,N_14252);
nor UO_396 (O_396,N_14360,N_14542);
nand UO_397 (O_397,N_14973,N_14509);
or UO_398 (O_398,N_14035,N_14168);
or UO_399 (O_399,N_14095,N_14856);
xor UO_400 (O_400,N_14213,N_14871);
nand UO_401 (O_401,N_14068,N_14541);
nor UO_402 (O_402,N_14318,N_14422);
nor UO_403 (O_403,N_14246,N_14725);
nor UO_404 (O_404,N_14735,N_14756);
and UO_405 (O_405,N_14403,N_14738);
nand UO_406 (O_406,N_14766,N_14175);
or UO_407 (O_407,N_14293,N_14964);
and UO_408 (O_408,N_14644,N_14443);
xor UO_409 (O_409,N_14684,N_14707);
nor UO_410 (O_410,N_14640,N_14936);
nor UO_411 (O_411,N_14783,N_14551);
nand UO_412 (O_412,N_14546,N_14902);
and UO_413 (O_413,N_14609,N_14717);
or UO_414 (O_414,N_14004,N_14672);
nand UO_415 (O_415,N_14714,N_14702);
nor UO_416 (O_416,N_14497,N_14737);
or UO_417 (O_417,N_14881,N_14393);
nor UO_418 (O_418,N_14650,N_14535);
or UO_419 (O_419,N_14641,N_14499);
nor UO_420 (O_420,N_14778,N_14309);
nor UO_421 (O_421,N_14083,N_14636);
and UO_422 (O_422,N_14608,N_14746);
and UO_423 (O_423,N_14601,N_14171);
or UO_424 (O_424,N_14385,N_14583);
nor UO_425 (O_425,N_14940,N_14234);
or UO_426 (O_426,N_14570,N_14250);
nand UO_427 (O_427,N_14712,N_14455);
nand UO_428 (O_428,N_14528,N_14423);
nor UO_429 (O_429,N_14013,N_14931);
or UO_430 (O_430,N_14112,N_14954);
nand UO_431 (O_431,N_14812,N_14476);
nand UO_432 (O_432,N_14012,N_14264);
or UO_433 (O_433,N_14612,N_14228);
nand UO_434 (O_434,N_14559,N_14324);
nand UO_435 (O_435,N_14749,N_14661);
and UO_436 (O_436,N_14014,N_14105);
nand UO_437 (O_437,N_14290,N_14017);
or UO_438 (O_438,N_14990,N_14330);
and UO_439 (O_439,N_14950,N_14673);
or UO_440 (O_440,N_14508,N_14299);
or UO_441 (O_441,N_14504,N_14477);
xnor UO_442 (O_442,N_14782,N_14670);
or UO_443 (O_443,N_14371,N_14072);
nand UO_444 (O_444,N_14818,N_14169);
nand UO_445 (O_445,N_14985,N_14157);
nand UO_446 (O_446,N_14402,N_14313);
or UO_447 (O_447,N_14134,N_14843);
nor UO_448 (O_448,N_14424,N_14592);
nand UO_449 (O_449,N_14928,N_14078);
nor UO_450 (O_450,N_14709,N_14680);
and UO_451 (O_451,N_14905,N_14390);
or UO_452 (O_452,N_14729,N_14373);
or UO_453 (O_453,N_14628,N_14678);
or UO_454 (O_454,N_14771,N_14387);
nand UO_455 (O_455,N_14543,N_14750);
nor UO_456 (O_456,N_14731,N_14198);
xor UO_457 (O_457,N_14834,N_14377);
nor UO_458 (O_458,N_14956,N_14103);
and UO_459 (O_459,N_14281,N_14498);
nand UO_460 (O_460,N_14230,N_14448);
nor UO_461 (O_461,N_14593,N_14016);
nand UO_462 (O_462,N_14708,N_14513);
nand UO_463 (O_463,N_14522,N_14125);
or UO_464 (O_464,N_14690,N_14895);
or UO_465 (O_465,N_14949,N_14807);
and UO_466 (O_466,N_14496,N_14822);
and UO_467 (O_467,N_14253,N_14571);
nor UO_468 (O_468,N_14397,N_14732);
nor UO_469 (O_469,N_14995,N_14098);
nand UO_470 (O_470,N_14054,N_14444);
and UO_471 (O_471,N_14314,N_14053);
nor UO_472 (O_472,N_14115,N_14050);
nand UO_473 (O_473,N_14786,N_14993);
or UO_474 (O_474,N_14873,N_14307);
and UO_475 (O_475,N_14139,N_14668);
nand UO_476 (O_476,N_14913,N_14983);
nand UO_477 (O_477,N_14916,N_14594);
nand UO_478 (O_478,N_14272,N_14032);
or UO_479 (O_479,N_14030,N_14365);
xor UO_480 (O_480,N_14879,N_14334);
nor UO_481 (O_481,N_14857,N_14590);
nor UO_482 (O_482,N_14401,N_14119);
and UO_483 (O_483,N_14015,N_14884);
nand UO_484 (O_484,N_14997,N_14514);
and UO_485 (O_485,N_14634,N_14539);
nor UO_486 (O_486,N_14229,N_14434);
nand UO_487 (O_487,N_14999,N_14599);
nand UO_488 (O_488,N_14779,N_14591);
nor UO_489 (O_489,N_14100,N_14167);
nand UO_490 (O_490,N_14798,N_14922);
nand UO_491 (O_491,N_14537,N_14156);
or UO_492 (O_492,N_14123,N_14706);
nand UO_493 (O_493,N_14219,N_14981);
or UO_494 (O_494,N_14278,N_14411);
or UO_495 (O_495,N_14793,N_14472);
xor UO_496 (O_496,N_14792,N_14503);
and UO_497 (O_497,N_14383,N_14665);
nand UO_498 (O_498,N_14835,N_14488);
nor UO_499 (O_499,N_14803,N_14527);
or UO_500 (O_500,N_14851,N_14212);
xor UO_501 (O_501,N_14429,N_14016);
nor UO_502 (O_502,N_14119,N_14186);
or UO_503 (O_503,N_14207,N_14025);
nor UO_504 (O_504,N_14825,N_14814);
nand UO_505 (O_505,N_14382,N_14499);
or UO_506 (O_506,N_14166,N_14796);
xnor UO_507 (O_507,N_14205,N_14646);
and UO_508 (O_508,N_14437,N_14651);
nand UO_509 (O_509,N_14732,N_14014);
nor UO_510 (O_510,N_14282,N_14572);
nor UO_511 (O_511,N_14586,N_14421);
or UO_512 (O_512,N_14243,N_14415);
or UO_513 (O_513,N_14351,N_14851);
nor UO_514 (O_514,N_14701,N_14797);
nand UO_515 (O_515,N_14663,N_14273);
and UO_516 (O_516,N_14924,N_14917);
or UO_517 (O_517,N_14624,N_14069);
or UO_518 (O_518,N_14649,N_14370);
nor UO_519 (O_519,N_14562,N_14892);
nor UO_520 (O_520,N_14755,N_14400);
nand UO_521 (O_521,N_14525,N_14358);
or UO_522 (O_522,N_14330,N_14371);
and UO_523 (O_523,N_14548,N_14981);
and UO_524 (O_524,N_14290,N_14078);
or UO_525 (O_525,N_14285,N_14685);
and UO_526 (O_526,N_14842,N_14667);
xor UO_527 (O_527,N_14895,N_14265);
nor UO_528 (O_528,N_14072,N_14825);
and UO_529 (O_529,N_14428,N_14457);
nand UO_530 (O_530,N_14569,N_14556);
xor UO_531 (O_531,N_14081,N_14839);
and UO_532 (O_532,N_14164,N_14452);
nand UO_533 (O_533,N_14678,N_14459);
nand UO_534 (O_534,N_14203,N_14292);
nor UO_535 (O_535,N_14948,N_14257);
and UO_536 (O_536,N_14793,N_14314);
and UO_537 (O_537,N_14797,N_14014);
nor UO_538 (O_538,N_14935,N_14538);
or UO_539 (O_539,N_14777,N_14469);
nor UO_540 (O_540,N_14830,N_14483);
and UO_541 (O_541,N_14331,N_14932);
or UO_542 (O_542,N_14701,N_14193);
xor UO_543 (O_543,N_14868,N_14481);
or UO_544 (O_544,N_14821,N_14480);
xor UO_545 (O_545,N_14474,N_14750);
xnor UO_546 (O_546,N_14716,N_14250);
nand UO_547 (O_547,N_14304,N_14240);
nor UO_548 (O_548,N_14515,N_14600);
nor UO_549 (O_549,N_14127,N_14369);
or UO_550 (O_550,N_14890,N_14762);
nand UO_551 (O_551,N_14569,N_14916);
nand UO_552 (O_552,N_14912,N_14298);
nand UO_553 (O_553,N_14141,N_14110);
or UO_554 (O_554,N_14209,N_14939);
nor UO_555 (O_555,N_14458,N_14119);
xor UO_556 (O_556,N_14182,N_14597);
and UO_557 (O_557,N_14875,N_14207);
and UO_558 (O_558,N_14669,N_14115);
and UO_559 (O_559,N_14665,N_14299);
nor UO_560 (O_560,N_14831,N_14123);
or UO_561 (O_561,N_14101,N_14016);
or UO_562 (O_562,N_14863,N_14259);
or UO_563 (O_563,N_14031,N_14160);
nor UO_564 (O_564,N_14688,N_14336);
and UO_565 (O_565,N_14840,N_14258);
nor UO_566 (O_566,N_14997,N_14865);
nor UO_567 (O_567,N_14600,N_14296);
and UO_568 (O_568,N_14177,N_14408);
or UO_569 (O_569,N_14831,N_14009);
and UO_570 (O_570,N_14031,N_14235);
nand UO_571 (O_571,N_14014,N_14039);
nand UO_572 (O_572,N_14616,N_14825);
or UO_573 (O_573,N_14114,N_14534);
or UO_574 (O_574,N_14844,N_14849);
nor UO_575 (O_575,N_14706,N_14309);
or UO_576 (O_576,N_14213,N_14521);
nor UO_577 (O_577,N_14140,N_14932);
nand UO_578 (O_578,N_14871,N_14082);
and UO_579 (O_579,N_14838,N_14867);
nor UO_580 (O_580,N_14357,N_14422);
xnor UO_581 (O_581,N_14690,N_14593);
or UO_582 (O_582,N_14597,N_14388);
xor UO_583 (O_583,N_14654,N_14516);
or UO_584 (O_584,N_14446,N_14873);
and UO_585 (O_585,N_14056,N_14705);
or UO_586 (O_586,N_14294,N_14217);
and UO_587 (O_587,N_14809,N_14035);
or UO_588 (O_588,N_14035,N_14470);
nand UO_589 (O_589,N_14812,N_14593);
or UO_590 (O_590,N_14391,N_14635);
nand UO_591 (O_591,N_14482,N_14764);
nor UO_592 (O_592,N_14169,N_14049);
nand UO_593 (O_593,N_14723,N_14819);
or UO_594 (O_594,N_14491,N_14308);
and UO_595 (O_595,N_14113,N_14135);
nor UO_596 (O_596,N_14714,N_14321);
nor UO_597 (O_597,N_14462,N_14951);
xnor UO_598 (O_598,N_14298,N_14342);
and UO_599 (O_599,N_14586,N_14253);
nand UO_600 (O_600,N_14854,N_14103);
and UO_601 (O_601,N_14906,N_14921);
or UO_602 (O_602,N_14262,N_14270);
nand UO_603 (O_603,N_14925,N_14169);
or UO_604 (O_604,N_14771,N_14432);
and UO_605 (O_605,N_14005,N_14888);
or UO_606 (O_606,N_14900,N_14049);
and UO_607 (O_607,N_14399,N_14550);
and UO_608 (O_608,N_14033,N_14776);
xnor UO_609 (O_609,N_14169,N_14080);
or UO_610 (O_610,N_14712,N_14538);
nand UO_611 (O_611,N_14332,N_14096);
nand UO_612 (O_612,N_14652,N_14525);
xor UO_613 (O_613,N_14106,N_14245);
and UO_614 (O_614,N_14853,N_14632);
or UO_615 (O_615,N_14181,N_14571);
or UO_616 (O_616,N_14247,N_14364);
or UO_617 (O_617,N_14592,N_14018);
xor UO_618 (O_618,N_14471,N_14068);
nand UO_619 (O_619,N_14095,N_14050);
xor UO_620 (O_620,N_14313,N_14723);
nor UO_621 (O_621,N_14655,N_14303);
nand UO_622 (O_622,N_14620,N_14435);
xor UO_623 (O_623,N_14669,N_14081);
nor UO_624 (O_624,N_14575,N_14357);
nor UO_625 (O_625,N_14852,N_14711);
nor UO_626 (O_626,N_14278,N_14250);
or UO_627 (O_627,N_14925,N_14464);
nand UO_628 (O_628,N_14249,N_14200);
nor UO_629 (O_629,N_14143,N_14530);
nor UO_630 (O_630,N_14581,N_14349);
and UO_631 (O_631,N_14637,N_14001);
nand UO_632 (O_632,N_14528,N_14777);
nand UO_633 (O_633,N_14075,N_14986);
xnor UO_634 (O_634,N_14593,N_14242);
and UO_635 (O_635,N_14335,N_14247);
nand UO_636 (O_636,N_14064,N_14084);
nand UO_637 (O_637,N_14052,N_14745);
nand UO_638 (O_638,N_14710,N_14449);
and UO_639 (O_639,N_14628,N_14772);
and UO_640 (O_640,N_14356,N_14412);
nor UO_641 (O_641,N_14704,N_14720);
nand UO_642 (O_642,N_14940,N_14106);
xor UO_643 (O_643,N_14330,N_14709);
or UO_644 (O_644,N_14155,N_14873);
or UO_645 (O_645,N_14690,N_14731);
and UO_646 (O_646,N_14113,N_14455);
and UO_647 (O_647,N_14342,N_14449);
nand UO_648 (O_648,N_14990,N_14473);
nand UO_649 (O_649,N_14796,N_14002);
or UO_650 (O_650,N_14824,N_14236);
nor UO_651 (O_651,N_14641,N_14757);
nor UO_652 (O_652,N_14326,N_14434);
and UO_653 (O_653,N_14106,N_14825);
nand UO_654 (O_654,N_14266,N_14292);
and UO_655 (O_655,N_14952,N_14073);
xor UO_656 (O_656,N_14391,N_14096);
nand UO_657 (O_657,N_14285,N_14774);
or UO_658 (O_658,N_14175,N_14832);
nor UO_659 (O_659,N_14878,N_14879);
xor UO_660 (O_660,N_14271,N_14494);
or UO_661 (O_661,N_14681,N_14816);
nand UO_662 (O_662,N_14147,N_14023);
nor UO_663 (O_663,N_14749,N_14275);
nor UO_664 (O_664,N_14129,N_14123);
nor UO_665 (O_665,N_14881,N_14018);
or UO_666 (O_666,N_14673,N_14361);
and UO_667 (O_667,N_14559,N_14546);
nand UO_668 (O_668,N_14705,N_14960);
and UO_669 (O_669,N_14978,N_14416);
xnor UO_670 (O_670,N_14643,N_14827);
nand UO_671 (O_671,N_14518,N_14936);
nand UO_672 (O_672,N_14306,N_14248);
nand UO_673 (O_673,N_14387,N_14116);
or UO_674 (O_674,N_14175,N_14293);
and UO_675 (O_675,N_14499,N_14803);
and UO_676 (O_676,N_14008,N_14048);
and UO_677 (O_677,N_14999,N_14954);
nor UO_678 (O_678,N_14646,N_14852);
and UO_679 (O_679,N_14050,N_14706);
or UO_680 (O_680,N_14871,N_14516);
or UO_681 (O_681,N_14608,N_14851);
nand UO_682 (O_682,N_14736,N_14910);
or UO_683 (O_683,N_14151,N_14045);
or UO_684 (O_684,N_14973,N_14621);
or UO_685 (O_685,N_14011,N_14256);
and UO_686 (O_686,N_14500,N_14744);
xor UO_687 (O_687,N_14397,N_14078);
nand UO_688 (O_688,N_14769,N_14832);
nand UO_689 (O_689,N_14068,N_14246);
nand UO_690 (O_690,N_14139,N_14791);
and UO_691 (O_691,N_14033,N_14914);
and UO_692 (O_692,N_14898,N_14044);
or UO_693 (O_693,N_14678,N_14525);
or UO_694 (O_694,N_14003,N_14674);
nor UO_695 (O_695,N_14575,N_14021);
nor UO_696 (O_696,N_14570,N_14316);
or UO_697 (O_697,N_14479,N_14893);
and UO_698 (O_698,N_14397,N_14512);
nand UO_699 (O_699,N_14674,N_14015);
nand UO_700 (O_700,N_14300,N_14255);
and UO_701 (O_701,N_14929,N_14247);
or UO_702 (O_702,N_14433,N_14639);
nor UO_703 (O_703,N_14902,N_14984);
and UO_704 (O_704,N_14856,N_14818);
or UO_705 (O_705,N_14411,N_14864);
and UO_706 (O_706,N_14864,N_14521);
and UO_707 (O_707,N_14311,N_14491);
nand UO_708 (O_708,N_14793,N_14738);
xnor UO_709 (O_709,N_14599,N_14152);
nor UO_710 (O_710,N_14566,N_14916);
and UO_711 (O_711,N_14115,N_14328);
nand UO_712 (O_712,N_14146,N_14840);
or UO_713 (O_713,N_14874,N_14696);
and UO_714 (O_714,N_14109,N_14115);
and UO_715 (O_715,N_14074,N_14530);
nand UO_716 (O_716,N_14889,N_14102);
nor UO_717 (O_717,N_14443,N_14964);
or UO_718 (O_718,N_14773,N_14662);
nor UO_719 (O_719,N_14803,N_14181);
nor UO_720 (O_720,N_14269,N_14039);
and UO_721 (O_721,N_14865,N_14224);
nand UO_722 (O_722,N_14312,N_14145);
xor UO_723 (O_723,N_14715,N_14622);
nor UO_724 (O_724,N_14026,N_14639);
nor UO_725 (O_725,N_14586,N_14279);
nand UO_726 (O_726,N_14744,N_14807);
or UO_727 (O_727,N_14281,N_14218);
xor UO_728 (O_728,N_14498,N_14850);
or UO_729 (O_729,N_14268,N_14089);
nor UO_730 (O_730,N_14742,N_14625);
nor UO_731 (O_731,N_14001,N_14862);
and UO_732 (O_732,N_14000,N_14485);
and UO_733 (O_733,N_14428,N_14759);
or UO_734 (O_734,N_14888,N_14588);
nor UO_735 (O_735,N_14316,N_14746);
or UO_736 (O_736,N_14110,N_14241);
nand UO_737 (O_737,N_14595,N_14858);
nor UO_738 (O_738,N_14479,N_14092);
nor UO_739 (O_739,N_14440,N_14949);
xor UO_740 (O_740,N_14233,N_14414);
nor UO_741 (O_741,N_14205,N_14203);
or UO_742 (O_742,N_14240,N_14759);
or UO_743 (O_743,N_14828,N_14383);
xnor UO_744 (O_744,N_14736,N_14022);
or UO_745 (O_745,N_14933,N_14842);
nor UO_746 (O_746,N_14798,N_14904);
xnor UO_747 (O_747,N_14340,N_14490);
or UO_748 (O_748,N_14488,N_14257);
and UO_749 (O_749,N_14307,N_14141);
nor UO_750 (O_750,N_14669,N_14755);
and UO_751 (O_751,N_14691,N_14360);
nand UO_752 (O_752,N_14292,N_14624);
and UO_753 (O_753,N_14180,N_14005);
nand UO_754 (O_754,N_14436,N_14875);
nor UO_755 (O_755,N_14897,N_14262);
and UO_756 (O_756,N_14754,N_14896);
nand UO_757 (O_757,N_14216,N_14463);
nor UO_758 (O_758,N_14527,N_14487);
xnor UO_759 (O_759,N_14296,N_14602);
xnor UO_760 (O_760,N_14579,N_14807);
nor UO_761 (O_761,N_14706,N_14766);
or UO_762 (O_762,N_14204,N_14099);
nor UO_763 (O_763,N_14177,N_14071);
and UO_764 (O_764,N_14427,N_14484);
nand UO_765 (O_765,N_14345,N_14027);
or UO_766 (O_766,N_14444,N_14498);
nand UO_767 (O_767,N_14416,N_14493);
xnor UO_768 (O_768,N_14496,N_14687);
and UO_769 (O_769,N_14709,N_14825);
or UO_770 (O_770,N_14880,N_14071);
nor UO_771 (O_771,N_14310,N_14101);
nand UO_772 (O_772,N_14174,N_14096);
or UO_773 (O_773,N_14301,N_14472);
or UO_774 (O_774,N_14502,N_14150);
and UO_775 (O_775,N_14633,N_14003);
nand UO_776 (O_776,N_14279,N_14371);
and UO_777 (O_777,N_14463,N_14209);
or UO_778 (O_778,N_14213,N_14614);
nand UO_779 (O_779,N_14522,N_14387);
nand UO_780 (O_780,N_14435,N_14775);
or UO_781 (O_781,N_14630,N_14100);
and UO_782 (O_782,N_14212,N_14261);
xor UO_783 (O_783,N_14121,N_14142);
nor UO_784 (O_784,N_14529,N_14876);
and UO_785 (O_785,N_14672,N_14447);
and UO_786 (O_786,N_14643,N_14295);
nand UO_787 (O_787,N_14437,N_14403);
and UO_788 (O_788,N_14250,N_14176);
or UO_789 (O_789,N_14566,N_14691);
and UO_790 (O_790,N_14499,N_14318);
and UO_791 (O_791,N_14592,N_14587);
xnor UO_792 (O_792,N_14202,N_14213);
nor UO_793 (O_793,N_14504,N_14382);
and UO_794 (O_794,N_14751,N_14293);
nand UO_795 (O_795,N_14688,N_14565);
nor UO_796 (O_796,N_14493,N_14944);
nor UO_797 (O_797,N_14779,N_14241);
nor UO_798 (O_798,N_14241,N_14566);
xor UO_799 (O_799,N_14567,N_14785);
nor UO_800 (O_800,N_14146,N_14320);
or UO_801 (O_801,N_14457,N_14622);
or UO_802 (O_802,N_14974,N_14553);
nand UO_803 (O_803,N_14503,N_14043);
nor UO_804 (O_804,N_14704,N_14234);
and UO_805 (O_805,N_14540,N_14819);
or UO_806 (O_806,N_14935,N_14451);
nand UO_807 (O_807,N_14290,N_14275);
nor UO_808 (O_808,N_14060,N_14652);
or UO_809 (O_809,N_14705,N_14582);
nand UO_810 (O_810,N_14623,N_14402);
nand UO_811 (O_811,N_14369,N_14142);
nand UO_812 (O_812,N_14077,N_14257);
nor UO_813 (O_813,N_14371,N_14116);
nand UO_814 (O_814,N_14820,N_14658);
and UO_815 (O_815,N_14317,N_14596);
or UO_816 (O_816,N_14141,N_14258);
nor UO_817 (O_817,N_14230,N_14108);
nor UO_818 (O_818,N_14061,N_14402);
xnor UO_819 (O_819,N_14103,N_14600);
nor UO_820 (O_820,N_14598,N_14948);
nor UO_821 (O_821,N_14644,N_14175);
nand UO_822 (O_822,N_14325,N_14662);
and UO_823 (O_823,N_14949,N_14329);
or UO_824 (O_824,N_14930,N_14636);
or UO_825 (O_825,N_14333,N_14433);
nor UO_826 (O_826,N_14899,N_14042);
xnor UO_827 (O_827,N_14304,N_14382);
or UO_828 (O_828,N_14953,N_14440);
and UO_829 (O_829,N_14949,N_14303);
and UO_830 (O_830,N_14327,N_14616);
nand UO_831 (O_831,N_14896,N_14238);
nor UO_832 (O_832,N_14329,N_14481);
nand UO_833 (O_833,N_14503,N_14864);
and UO_834 (O_834,N_14432,N_14002);
and UO_835 (O_835,N_14254,N_14145);
xnor UO_836 (O_836,N_14924,N_14353);
nand UO_837 (O_837,N_14369,N_14903);
and UO_838 (O_838,N_14674,N_14449);
nand UO_839 (O_839,N_14393,N_14895);
xnor UO_840 (O_840,N_14285,N_14183);
nor UO_841 (O_841,N_14082,N_14837);
and UO_842 (O_842,N_14334,N_14340);
and UO_843 (O_843,N_14471,N_14143);
nand UO_844 (O_844,N_14019,N_14124);
xnor UO_845 (O_845,N_14303,N_14569);
or UO_846 (O_846,N_14261,N_14995);
or UO_847 (O_847,N_14937,N_14648);
and UO_848 (O_848,N_14825,N_14179);
xor UO_849 (O_849,N_14320,N_14562);
nor UO_850 (O_850,N_14174,N_14908);
and UO_851 (O_851,N_14931,N_14123);
nor UO_852 (O_852,N_14557,N_14658);
nand UO_853 (O_853,N_14743,N_14341);
or UO_854 (O_854,N_14328,N_14136);
or UO_855 (O_855,N_14130,N_14732);
and UO_856 (O_856,N_14064,N_14774);
nor UO_857 (O_857,N_14771,N_14608);
or UO_858 (O_858,N_14575,N_14228);
or UO_859 (O_859,N_14778,N_14382);
xnor UO_860 (O_860,N_14359,N_14537);
or UO_861 (O_861,N_14000,N_14804);
or UO_862 (O_862,N_14430,N_14367);
nor UO_863 (O_863,N_14759,N_14439);
or UO_864 (O_864,N_14714,N_14414);
or UO_865 (O_865,N_14247,N_14367);
and UO_866 (O_866,N_14952,N_14375);
nor UO_867 (O_867,N_14946,N_14573);
or UO_868 (O_868,N_14110,N_14815);
nor UO_869 (O_869,N_14331,N_14268);
or UO_870 (O_870,N_14418,N_14825);
nand UO_871 (O_871,N_14582,N_14156);
nand UO_872 (O_872,N_14003,N_14421);
nor UO_873 (O_873,N_14676,N_14031);
nand UO_874 (O_874,N_14572,N_14234);
nor UO_875 (O_875,N_14243,N_14778);
or UO_876 (O_876,N_14433,N_14724);
nand UO_877 (O_877,N_14064,N_14780);
or UO_878 (O_878,N_14976,N_14979);
and UO_879 (O_879,N_14621,N_14341);
or UO_880 (O_880,N_14638,N_14257);
nand UO_881 (O_881,N_14309,N_14006);
xor UO_882 (O_882,N_14055,N_14109);
nand UO_883 (O_883,N_14930,N_14316);
xnor UO_884 (O_884,N_14816,N_14105);
and UO_885 (O_885,N_14331,N_14505);
nor UO_886 (O_886,N_14543,N_14098);
and UO_887 (O_887,N_14545,N_14581);
and UO_888 (O_888,N_14919,N_14304);
and UO_889 (O_889,N_14168,N_14039);
or UO_890 (O_890,N_14666,N_14991);
or UO_891 (O_891,N_14733,N_14154);
or UO_892 (O_892,N_14126,N_14306);
or UO_893 (O_893,N_14139,N_14926);
nor UO_894 (O_894,N_14847,N_14975);
and UO_895 (O_895,N_14784,N_14637);
and UO_896 (O_896,N_14455,N_14746);
or UO_897 (O_897,N_14514,N_14884);
nor UO_898 (O_898,N_14399,N_14882);
nor UO_899 (O_899,N_14059,N_14558);
nand UO_900 (O_900,N_14825,N_14255);
nor UO_901 (O_901,N_14290,N_14120);
and UO_902 (O_902,N_14504,N_14466);
and UO_903 (O_903,N_14352,N_14291);
nand UO_904 (O_904,N_14257,N_14312);
nand UO_905 (O_905,N_14125,N_14970);
and UO_906 (O_906,N_14548,N_14797);
or UO_907 (O_907,N_14610,N_14762);
xnor UO_908 (O_908,N_14022,N_14806);
xnor UO_909 (O_909,N_14407,N_14765);
and UO_910 (O_910,N_14371,N_14417);
and UO_911 (O_911,N_14277,N_14404);
nor UO_912 (O_912,N_14656,N_14433);
and UO_913 (O_913,N_14097,N_14586);
and UO_914 (O_914,N_14475,N_14265);
or UO_915 (O_915,N_14933,N_14121);
and UO_916 (O_916,N_14189,N_14078);
xnor UO_917 (O_917,N_14576,N_14415);
xnor UO_918 (O_918,N_14608,N_14664);
nand UO_919 (O_919,N_14422,N_14865);
nand UO_920 (O_920,N_14554,N_14378);
nor UO_921 (O_921,N_14111,N_14722);
xor UO_922 (O_922,N_14978,N_14533);
or UO_923 (O_923,N_14438,N_14332);
nand UO_924 (O_924,N_14000,N_14889);
and UO_925 (O_925,N_14443,N_14841);
or UO_926 (O_926,N_14991,N_14086);
nor UO_927 (O_927,N_14063,N_14743);
nor UO_928 (O_928,N_14852,N_14487);
or UO_929 (O_929,N_14483,N_14292);
or UO_930 (O_930,N_14149,N_14594);
and UO_931 (O_931,N_14988,N_14438);
or UO_932 (O_932,N_14299,N_14032);
and UO_933 (O_933,N_14913,N_14008);
or UO_934 (O_934,N_14697,N_14011);
nor UO_935 (O_935,N_14521,N_14072);
nor UO_936 (O_936,N_14158,N_14018);
and UO_937 (O_937,N_14551,N_14556);
nand UO_938 (O_938,N_14836,N_14455);
and UO_939 (O_939,N_14897,N_14190);
nand UO_940 (O_940,N_14272,N_14185);
nor UO_941 (O_941,N_14526,N_14066);
nor UO_942 (O_942,N_14620,N_14774);
or UO_943 (O_943,N_14893,N_14899);
nand UO_944 (O_944,N_14492,N_14693);
nor UO_945 (O_945,N_14188,N_14169);
nor UO_946 (O_946,N_14581,N_14897);
or UO_947 (O_947,N_14010,N_14330);
and UO_948 (O_948,N_14828,N_14899);
and UO_949 (O_949,N_14449,N_14696);
or UO_950 (O_950,N_14935,N_14498);
or UO_951 (O_951,N_14033,N_14496);
nand UO_952 (O_952,N_14615,N_14771);
or UO_953 (O_953,N_14163,N_14596);
nor UO_954 (O_954,N_14971,N_14841);
nand UO_955 (O_955,N_14856,N_14284);
nor UO_956 (O_956,N_14291,N_14208);
nand UO_957 (O_957,N_14005,N_14230);
xnor UO_958 (O_958,N_14119,N_14423);
xor UO_959 (O_959,N_14042,N_14559);
or UO_960 (O_960,N_14156,N_14152);
nand UO_961 (O_961,N_14572,N_14943);
nand UO_962 (O_962,N_14599,N_14391);
and UO_963 (O_963,N_14521,N_14229);
and UO_964 (O_964,N_14364,N_14457);
nand UO_965 (O_965,N_14220,N_14386);
and UO_966 (O_966,N_14106,N_14921);
nand UO_967 (O_967,N_14034,N_14239);
nand UO_968 (O_968,N_14604,N_14738);
xnor UO_969 (O_969,N_14823,N_14471);
or UO_970 (O_970,N_14695,N_14659);
and UO_971 (O_971,N_14473,N_14559);
nand UO_972 (O_972,N_14603,N_14208);
and UO_973 (O_973,N_14289,N_14256);
or UO_974 (O_974,N_14585,N_14784);
nand UO_975 (O_975,N_14927,N_14848);
and UO_976 (O_976,N_14160,N_14731);
or UO_977 (O_977,N_14095,N_14726);
or UO_978 (O_978,N_14068,N_14379);
and UO_979 (O_979,N_14610,N_14172);
and UO_980 (O_980,N_14818,N_14913);
and UO_981 (O_981,N_14772,N_14523);
nand UO_982 (O_982,N_14216,N_14789);
nand UO_983 (O_983,N_14308,N_14457);
nand UO_984 (O_984,N_14963,N_14661);
or UO_985 (O_985,N_14155,N_14397);
nand UO_986 (O_986,N_14818,N_14999);
or UO_987 (O_987,N_14649,N_14679);
xor UO_988 (O_988,N_14347,N_14206);
or UO_989 (O_989,N_14594,N_14476);
or UO_990 (O_990,N_14724,N_14969);
or UO_991 (O_991,N_14552,N_14018);
nand UO_992 (O_992,N_14159,N_14562);
or UO_993 (O_993,N_14023,N_14165);
nand UO_994 (O_994,N_14077,N_14571);
or UO_995 (O_995,N_14646,N_14526);
and UO_996 (O_996,N_14479,N_14014);
nor UO_997 (O_997,N_14800,N_14302);
nor UO_998 (O_998,N_14217,N_14111);
nor UO_999 (O_999,N_14974,N_14453);
nor UO_1000 (O_1000,N_14595,N_14920);
and UO_1001 (O_1001,N_14598,N_14098);
and UO_1002 (O_1002,N_14974,N_14634);
xor UO_1003 (O_1003,N_14283,N_14194);
and UO_1004 (O_1004,N_14295,N_14920);
and UO_1005 (O_1005,N_14414,N_14793);
xor UO_1006 (O_1006,N_14438,N_14349);
nor UO_1007 (O_1007,N_14800,N_14652);
and UO_1008 (O_1008,N_14270,N_14399);
nand UO_1009 (O_1009,N_14766,N_14182);
nand UO_1010 (O_1010,N_14541,N_14534);
and UO_1011 (O_1011,N_14684,N_14101);
nor UO_1012 (O_1012,N_14566,N_14938);
or UO_1013 (O_1013,N_14168,N_14190);
and UO_1014 (O_1014,N_14740,N_14375);
and UO_1015 (O_1015,N_14147,N_14653);
xnor UO_1016 (O_1016,N_14186,N_14284);
or UO_1017 (O_1017,N_14086,N_14587);
and UO_1018 (O_1018,N_14753,N_14006);
or UO_1019 (O_1019,N_14025,N_14950);
nand UO_1020 (O_1020,N_14368,N_14438);
or UO_1021 (O_1021,N_14810,N_14450);
nand UO_1022 (O_1022,N_14107,N_14822);
or UO_1023 (O_1023,N_14722,N_14802);
and UO_1024 (O_1024,N_14061,N_14282);
xor UO_1025 (O_1025,N_14944,N_14590);
xnor UO_1026 (O_1026,N_14457,N_14679);
nor UO_1027 (O_1027,N_14691,N_14480);
and UO_1028 (O_1028,N_14096,N_14535);
nand UO_1029 (O_1029,N_14607,N_14501);
and UO_1030 (O_1030,N_14435,N_14034);
and UO_1031 (O_1031,N_14070,N_14153);
nor UO_1032 (O_1032,N_14912,N_14694);
xor UO_1033 (O_1033,N_14679,N_14830);
and UO_1034 (O_1034,N_14071,N_14186);
nand UO_1035 (O_1035,N_14683,N_14539);
nand UO_1036 (O_1036,N_14435,N_14333);
or UO_1037 (O_1037,N_14727,N_14634);
xor UO_1038 (O_1038,N_14733,N_14302);
nor UO_1039 (O_1039,N_14474,N_14818);
and UO_1040 (O_1040,N_14711,N_14544);
nand UO_1041 (O_1041,N_14341,N_14239);
nand UO_1042 (O_1042,N_14167,N_14867);
or UO_1043 (O_1043,N_14727,N_14719);
nand UO_1044 (O_1044,N_14316,N_14032);
and UO_1045 (O_1045,N_14330,N_14392);
or UO_1046 (O_1046,N_14419,N_14741);
nand UO_1047 (O_1047,N_14585,N_14011);
or UO_1048 (O_1048,N_14398,N_14823);
xnor UO_1049 (O_1049,N_14037,N_14308);
or UO_1050 (O_1050,N_14808,N_14261);
nand UO_1051 (O_1051,N_14769,N_14570);
or UO_1052 (O_1052,N_14538,N_14681);
nand UO_1053 (O_1053,N_14255,N_14701);
nand UO_1054 (O_1054,N_14297,N_14625);
or UO_1055 (O_1055,N_14844,N_14928);
and UO_1056 (O_1056,N_14914,N_14992);
and UO_1057 (O_1057,N_14741,N_14179);
nand UO_1058 (O_1058,N_14822,N_14544);
xor UO_1059 (O_1059,N_14398,N_14929);
and UO_1060 (O_1060,N_14221,N_14843);
nor UO_1061 (O_1061,N_14116,N_14465);
nand UO_1062 (O_1062,N_14455,N_14641);
nor UO_1063 (O_1063,N_14111,N_14949);
and UO_1064 (O_1064,N_14637,N_14264);
and UO_1065 (O_1065,N_14288,N_14208);
nor UO_1066 (O_1066,N_14411,N_14611);
nand UO_1067 (O_1067,N_14025,N_14000);
nor UO_1068 (O_1068,N_14202,N_14100);
nand UO_1069 (O_1069,N_14440,N_14067);
or UO_1070 (O_1070,N_14890,N_14719);
and UO_1071 (O_1071,N_14335,N_14413);
and UO_1072 (O_1072,N_14554,N_14385);
nor UO_1073 (O_1073,N_14009,N_14938);
xnor UO_1074 (O_1074,N_14840,N_14141);
nor UO_1075 (O_1075,N_14719,N_14763);
nand UO_1076 (O_1076,N_14201,N_14950);
nand UO_1077 (O_1077,N_14951,N_14335);
and UO_1078 (O_1078,N_14251,N_14337);
xnor UO_1079 (O_1079,N_14053,N_14640);
and UO_1080 (O_1080,N_14687,N_14471);
and UO_1081 (O_1081,N_14784,N_14130);
nand UO_1082 (O_1082,N_14104,N_14367);
and UO_1083 (O_1083,N_14205,N_14133);
nor UO_1084 (O_1084,N_14665,N_14663);
nor UO_1085 (O_1085,N_14486,N_14822);
xor UO_1086 (O_1086,N_14879,N_14036);
and UO_1087 (O_1087,N_14344,N_14911);
and UO_1088 (O_1088,N_14990,N_14998);
nor UO_1089 (O_1089,N_14860,N_14058);
nand UO_1090 (O_1090,N_14026,N_14371);
and UO_1091 (O_1091,N_14671,N_14341);
and UO_1092 (O_1092,N_14199,N_14736);
and UO_1093 (O_1093,N_14731,N_14997);
nor UO_1094 (O_1094,N_14584,N_14276);
and UO_1095 (O_1095,N_14727,N_14499);
or UO_1096 (O_1096,N_14111,N_14197);
and UO_1097 (O_1097,N_14689,N_14404);
xor UO_1098 (O_1098,N_14110,N_14425);
or UO_1099 (O_1099,N_14734,N_14737);
nand UO_1100 (O_1100,N_14796,N_14885);
or UO_1101 (O_1101,N_14432,N_14780);
or UO_1102 (O_1102,N_14390,N_14349);
nand UO_1103 (O_1103,N_14223,N_14874);
nor UO_1104 (O_1104,N_14438,N_14396);
or UO_1105 (O_1105,N_14097,N_14807);
nor UO_1106 (O_1106,N_14002,N_14008);
xor UO_1107 (O_1107,N_14194,N_14558);
or UO_1108 (O_1108,N_14571,N_14097);
nand UO_1109 (O_1109,N_14064,N_14766);
nand UO_1110 (O_1110,N_14901,N_14564);
or UO_1111 (O_1111,N_14871,N_14927);
and UO_1112 (O_1112,N_14596,N_14256);
nand UO_1113 (O_1113,N_14084,N_14154);
and UO_1114 (O_1114,N_14330,N_14471);
and UO_1115 (O_1115,N_14904,N_14923);
or UO_1116 (O_1116,N_14306,N_14255);
and UO_1117 (O_1117,N_14370,N_14779);
and UO_1118 (O_1118,N_14518,N_14628);
nand UO_1119 (O_1119,N_14615,N_14205);
nor UO_1120 (O_1120,N_14919,N_14650);
xor UO_1121 (O_1121,N_14672,N_14766);
nand UO_1122 (O_1122,N_14078,N_14794);
xnor UO_1123 (O_1123,N_14420,N_14657);
xnor UO_1124 (O_1124,N_14136,N_14729);
nor UO_1125 (O_1125,N_14774,N_14599);
xor UO_1126 (O_1126,N_14803,N_14324);
nand UO_1127 (O_1127,N_14891,N_14845);
and UO_1128 (O_1128,N_14081,N_14675);
nand UO_1129 (O_1129,N_14368,N_14580);
and UO_1130 (O_1130,N_14494,N_14587);
or UO_1131 (O_1131,N_14820,N_14221);
nor UO_1132 (O_1132,N_14425,N_14544);
or UO_1133 (O_1133,N_14479,N_14454);
or UO_1134 (O_1134,N_14342,N_14299);
and UO_1135 (O_1135,N_14513,N_14552);
nor UO_1136 (O_1136,N_14201,N_14755);
and UO_1137 (O_1137,N_14008,N_14004);
or UO_1138 (O_1138,N_14210,N_14613);
or UO_1139 (O_1139,N_14967,N_14466);
xnor UO_1140 (O_1140,N_14250,N_14753);
xor UO_1141 (O_1141,N_14607,N_14049);
xnor UO_1142 (O_1142,N_14461,N_14549);
or UO_1143 (O_1143,N_14874,N_14560);
and UO_1144 (O_1144,N_14277,N_14564);
or UO_1145 (O_1145,N_14313,N_14773);
and UO_1146 (O_1146,N_14988,N_14692);
nor UO_1147 (O_1147,N_14619,N_14024);
nor UO_1148 (O_1148,N_14373,N_14192);
nand UO_1149 (O_1149,N_14467,N_14721);
or UO_1150 (O_1150,N_14811,N_14846);
or UO_1151 (O_1151,N_14458,N_14497);
xor UO_1152 (O_1152,N_14451,N_14448);
or UO_1153 (O_1153,N_14639,N_14079);
nor UO_1154 (O_1154,N_14130,N_14036);
xor UO_1155 (O_1155,N_14932,N_14748);
and UO_1156 (O_1156,N_14219,N_14545);
xnor UO_1157 (O_1157,N_14860,N_14875);
nor UO_1158 (O_1158,N_14957,N_14067);
or UO_1159 (O_1159,N_14910,N_14459);
xnor UO_1160 (O_1160,N_14278,N_14379);
nand UO_1161 (O_1161,N_14749,N_14093);
nor UO_1162 (O_1162,N_14300,N_14129);
xnor UO_1163 (O_1163,N_14907,N_14836);
nor UO_1164 (O_1164,N_14422,N_14125);
nor UO_1165 (O_1165,N_14386,N_14969);
and UO_1166 (O_1166,N_14692,N_14706);
and UO_1167 (O_1167,N_14948,N_14776);
or UO_1168 (O_1168,N_14792,N_14375);
nor UO_1169 (O_1169,N_14979,N_14539);
or UO_1170 (O_1170,N_14251,N_14858);
and UO_1171 (O_1171,N_14503,N_14506);
nand UO_1172 (O_1172,N_14255,N_14847);
nand UO_1173 (O_1173,N_14505,N_14552);
nor UO_1174 (O_1174,N_14759,N_14406);
nand UO_1175 (O_1175,N_14445,N_14508);
nor UO_1176 (O_1176,N_14622,N_14539);
or UO_1177 (O_1177,N_14796,N_14679);
nand UO_1178 (O_1178,N_14498,N_14413);
xor UO_1179 (O_1179,N_14715,N_14289);
or UO_1180 (O_1180,N_14836,N_14846);
and UO_1181 (O_1181,N_14191,N_14527);
nor UO_1182 (O_1182,N_14054,N_14262);
nor UO_1183 (O_1183,N_14015,N_14414);
or UO_1184 (O_1184,N_14063,N_14575);
nor UO_1185 (O_1185,N_14073,N_14407);
or UO_1186 (O_1186,N_14343,N_14881);
and UO_1187 (O_1187,N_14141,N_14439);
nand UO_1188 (O_1188,N_14017,N_14339);
nand UO_1189 (O_1189,N_14680,N_14791);
or UO_1190 (O_1190,N_14882,N_14135);
or UO_1191 (O_1191,N_14345,N_14782);
nand UO_1192 (O_1192,N_14829,N_14528);
and UO_1193 (O_1193,N_14661,N_14739);
or UO_1194 (O_1194,N_14204,N_14065);
nand UO_1195 (O_1195,N_14342,N_14362);
nor UO_1196 (O_1196,N_14673,N_14393);
nand UO_1197 (O_1197,N_14425,N_14984);
nand UO_1198 (O_1198,N_14590,N_14036);
nand UO_1199 (O_1199,N_14486,N_14041);
nand UO_1200 (O_1200,N_14365,N_14419);
and UO_1201 (O_1201,N_14693,N_14235);
xnor UO_1202 (O_1202,N_14592,N_14068);
nor UO_1203 (O_1203,N_14990,N_14364);
or UO_1204 (O_1204,N_14948,N_14241);
and UO_1205 (O_1205,N_14014,N_14332);
nand UO_1206 (O_1206,N_14021,N_14860);
and UO_1207 (O_1207,N_14122,N_14954);
or UO_1208 (O_1208,N_14009,N_14593);
nand UO_1209 (O_1209,N_14071,N_14932);
and UO_1210 (O_1210,N_14650,N_14664);
nor UO_1211 (O_1211,N_14783,N_14424);
xor UO_1212 (O_1212,N_14249,N_14987);
nand UO_1213 (O_1213,N_14446,N_14077);
xor UO_1214 (O_1214,N_14849,N_14806);
xor UO_1215 (O_1215,N_14351,N_14177);
nor UO_1216 (O_1216,N_14572,N_14331);
nor UO_1217 (O_1217,N_14193,N_14384);
nor UO_1218 (O_1218,N_14909,N_14805);
and UO_1219 (O_1219,N_14011,N_14905);
nand UO_1220 (O_1220,N_14284,N_14475);
or UO_1221 (O_1221,N_14046,N_14798);
or UO_1222 (O_1222,N_14747,N_14251);
nor UO_1223 (O_1223,N_14060,N_14611);
and UO_1224 (O_1224,N_14102,N_14861);
and UO_1225 (O_1225,N_14426,N_14293);
nand UO_1226 (O_1226,N_14477,N_14594);
nor UO_1227 (O_1227,N_14225,N_14135);
and UO_1228 (O_1228,N_14372,N_14540);
nand UO_1229 (O_1229,N_14532,N_14514);
nor UO_1230 (O_1230,N_14673,N_14611);
nand UO_1231 (O_1231,N_14235,N_14632);
nor UO_1232 (O_1232,N_14857,N_14589);
or UO_1233 (O_1233,N_14819,N_14752);
nor UO_1234 (O_1234,N_14549,N_14926);
or UO_1235 (O_1235,N_14664,N_14572);
and UO_1236 (O_1236,N_14747,N_14117);
or UO_1237 (O_1237,N_14901,N_14422);
and UO_1238 (O_1238,N_14207,N_14585);
nand UO_1239 (O_1239,N_14089,N_14842);
or UO_1240 (O_1240,N_14941,N_14527);
or UO_1241 (O_1241,N_14240,N_14173);
nand UO_1242 (O_1242,N_14239,N_14575);
nand UO_1243 (O_1243,N_14318,N_14804);
nand UO_1244 (O_1244,N_14020,N_14524);
nand UO_1245 (O_1245,N_14157,N_14712);
or UO_1246 (O_1246,N_14880,N_14653);
and UO_1247 (O_1247,N_14280,N_14848);
and UO_1248 (O_1248,N_14875,N_14364);
nand UO_1249 (O_1249,N_14698,N_14272);
or UO_1250 (O_1250,N_14697,N_14797);
xor UO_1251 (O_1251,N_14922,N_14462);
or UO_1252 (O_1252,N_14690,N_14653);
nand UO_1253 (O_1253,N_14353,N_14073);
nor UO_1254 (O_1254,N_14179,N_14358);
xor UO_1255 (O_1255,N_14209,N_14716);
or UO_1256 (O_1256,N_14276,N_14958);
or UO_1257 (O_1257,N_14554,N_14569);
nand UO_1258 (O_1258,N_14351,N_14977);
xnor UO_1259 (O_1259,N_14158,N_14506);
and UO_1260 (O_1260,N_14739,N_14662);
or UO_1261 (O_1261,N_14515,N_14173);
and UO_1262 (O_1262,N_14555,N_14360);
nor UO_1263 (O_1263,N_14976,N_14057);
xor UO_1264 (O_1264,N_14706,N_14074);
or UO_1265 (O_1265,N_14325,N_14959);
nand UO_1266 (O_1266,N_14800,N_14617);
nand UO_1267 (O_1267,N_14115,N_14066);
nor UO_1268 (O_1268,N_14785,N_14851);
or UO_1269 (O_1269,N_14400,N_14843);
or UO_1270 (O_1270,N_14296,N_14762);
or UO_1271 (O_1271,N_14975,N_14334);
and UO_1272 (O_1272,N_14970,N_14286);
or UO_1273 (O_1273,N_14871,N_14942);
or UO_1274 (O_1274,N_14981,N_14605);
xor UO_1275 (O_1275,N_14128,N_14063);
xor UO_1276 (O_1276,N_14534,N_14027);
or UO_1277 (O_1277,N_14359,N_14016);
nor UO_1278 (O_1278,N_14294,N_14032);
and UO_1279 (O_1279,N_14378,N_14727);
and UO_1280 (O_1280,N_14364,N_14170);
nand UO_1281 (O_1281,N_14743,N_14007);
nor UO_1282 (O_1282,N_14172,N_14949);
or UO_1283 (O_1283,N_14976,N_14041);
and UO_1284 (O_1284,N_14443,N_14829);
and UO_1285 (O_1285,N_14859,N_14999);
nand UO_1286 (O_1286,N_14053,N_14937);
or UO_1287 (O_1287,N_14240,N_14207);
nand UO_1288 (O_1288,N_14695,N_14102);
nand UO_1289 (O_1289,N_14937,N_14906);
and UO_1290 (O_1290,N_14509,N_14227);
and UO_1291 (O_1291,N_14566,N_14688);
nor UO_1292 (O_1292,N_14999,N_14420);
and UO_1293 (O_1293,N_14764,N_14864);
nor UO_1294 (O_1294,N_14681,N_14779);
nand UO_1295 (O_1295,N_14812,N_14338);
nor UO_1296 (O_1296,N_14703,N_14335);
nand UO_1297 (O_1297,N_14353,N_14326);
or UO_1298 (O_1298,N_14408,N_14429);
or UO_1299 (O_1299,N_14485,N_14080);
and UO_1300 (O_1300,N_14993,N_14464);
or UO_1301 (O_1301,N_14026,N_14572);
and UO_1302 (O_1302,N_14816,N_14331);
or UO_1303 (O_1303,N_14336,N_14025);
nand UO_1304 (O_1304,N_14807,N_14103);
xor UO_1305 (O_1305,N_14811,N_14409);
nand UO_1306 (O_1306,N_14717,N_14821);
and UO_1307 (O_1307,N_14255,N_14599);
nor UO_1308 (O_1308,N_14221,N_14856);
nor UO_1309 (O_1309,N_14975,N_14999);
nor UO_1310 (O_1310,N_14628,N_14499);
nand UO_1311 (O_1311,N_14136,N_14597);
nand UO_1312 (O_1312,N_14627,N_14195);
and UO_1313 (O_1313,N_14579,N_14495);
xnor UO_1314 (O_1314,N_14281,N_14811);
nor UO_1315 (O_1315,N_14666,N_14496);
nor UO_1316 (O_1316,N_14504,N_14162);
nor UO_1317 (O_1317,N_14850,N_14226);
nand UO_1318 (O_1318,N_14356,N_14081);
nor UO_1319 (O_1319,N_14572,N_14422);
xor UO_1320 (O_1320,N_14352,N_14626);
and UO_1321 (O_1321,N_14875,N_14376);
nand UO_1322 (O_1322,N_14730,N_14134);
or UO_1323 (O_1323,N_14684,N_14819);
nor UO_1324 (O_1324,N_14107,N_14039);
and UO_1325 (O_1325,N_14079,N_14354);
xnor UO_1326 (O_1326,N_14651,N_14162);
nand UO_1327 (O_1327,N_14028,N_14157);
or UO_1328 (O_1328,N_14668,N_14060);
nor UO_1329 (O_1329,N_14078,N_14150);
or UO_1330 (O_1330,N_14037,N_14182);
nor UO_1331 (O_1331,N_14129,N_14886);
and UO_1332 (O_1332,N_14461,N_14627);
xor UO_1333 (O_1333,N_14688,N_14662);
nor UO_1334 (O_1334,N_14697,N_14999);
nor UO_1335 (O_1335,N_14932,N_14037);
nand UO_1336 (O_1336,N_14413,N_14925);
nor UO_1337 (O_1337,N_14059,N_14527);
nand UO_1338 (O_1338,N_14285,N_14011);
nor UO_1339 (O_1339,N_14713,N_14328);
nand UO_1340 (O_1340,N_14165,N_14784);
and UO_1341 (O_1341,N_14957,N_14902);
or UO_1342 (O_1342,N_14973,N_14182);
and UO_1343 (O_1343,N_14694,N_14106);
nor UO_1344 (O_1344,N_14123,N_14334);
and UO_1345 (O_1345,N_14734,N_14524);
or UO_1346 (O_1346,N_14381,N_14155);
and UO_1347 (O_1347,N_14198,N_14536);
nor UO_1348 (O_1348,N_14112,N_14843);
and UO_1349 (O_1349,N_14900,N_14667);
and UO_1350 (O_1350,N_14802,N_14314);
nor UO_1351 (O_1351,N_14947,N_14649);
nor UO_1352 (O_1352,N_14967,N_14057);
nand UO_1353 (O_1353,N_14087,N_14018);
nand UO_1354 (O_1354,N_14167,N_14686);
and UO_1355 (O_1355,N_14345,N_14791);
nor UO_1356 (O_1356,N_14411,N_14323);
nor UO_1357 (O_1357,N_14963,N_14772);
nand UO_1358 (O_1358,N_14079,N_14328);
nor UO_1359 (O_1359,N_14892,N_14541);
or UO_1360 (O_1360,N_14560,N_14222);
xnor UO_1361 (O_1361,N_14293,N_14474);
or UO_1362 (O_1362,N_14695,N_14580);
nor UO_1363 (O_1363,N_14606,N_14482);
or UO_1364 (O_1364,N_14666,N_14129);
nor UO_1365 (O_1365,N_14510,N_14379);
and UO_1366 (O_1366,N_14122,N_14562);
or UO_1367 (O_1367,N_14123,N_14075);
and UO_1368 (O_1368,N_14770,N_14681);
and UO_1369 (O_1369,N_14736,N_14198);
or UO_1370 (O_1370,N_14086,N_14035);
nand UO_1371 (O_1371,N_14365,N_14106);
or UO_1372 (O_1372,N_14473,N_14478);
xor UO_1373 (O_1373,N_14368,N_14537);
nand UO_1374 (O_1374,N_14106,N_14412);
xor UO_1375 (O_1375,N_14263,N_14633);
or UO_1376 (O_1376,N_14899,N_14711);
and UO_1377 (O_1377,N_14585,N_14612);
nor UO_1378 (O_1378,N_14196,N_14695);
nor UO_1379 (O_1379,N_14964,N_14402);
nand UO_1380 (O_1380,N_14361,N_14233);
and UO_1381 (O_1381,N_14353,N_14685);
nand UO_1382 (O_1382,N_14647,N_14974);
nor UO_1383 (O_1383,N_14338,N_14763);
or UO_1384 (O_1384,N_14815,N_14119);
and UO_1385 (O_1385,N_14666,N_14205);
and UO_1386 (O_1386,N_14587,N_14930);
nand UO_1387 (O_1387,N_14459,N_14589);
or UO_1388 (O_1388,N_14557,N_14538);
nor UO_1389 (O_1389,N_14950,N_14716);
and UO_1390 (O_1390,N_14867,N_14069);
or UO_1391 (O_1391,N_14445,N_14913);
and UO_1392 (O_1392,N_14455,N_14406);
and UO_1393 (O_1393,N_14455,N_14304);
nor UO_1394 (O_1394,N_14768,N_14478);
and UO_1395 (O_1395,N_14758,N_14952);
and UO_1396 (O_1396,N_14762,N_14779);
nor UO_1397 (O_1397,N_14325,N_14400);
nor UO_1398 (O_1398,N_14777,N_14310);
and UO_1399 (O_1399,N_14746,N_14713);
and UO_1400 (O_1400,N_14879,N_14755);
and UO_1401 (O_1401,N_14659,N_14251);
and UO_1402 (O_1402,N_14799,N_14631);
and UO_1403 (O_1403,N_14942,N_14674);
nor UO_1404 (O_1404,N_14667,N_14128);
or UO_1405 (O_1405,N_14561,N_14788);
nor UO_1406 (O_1406,N_14915,N_14447);
nand UO_1407 (O_1407,N_14301,N_14176);
nand UO_1408 (O_1408,N_14626,N_14278);
or UO_1409 (O_1409,N_14226,N_14845);
nor UO_1410 (O_1410,N_14473,N_14678);
nand UO_1411 (O_1411,N_14157,N_14677);
or UO_1412 (O_1412,N_14240,N_14095);
nand UO_1413 (O_1413,N_14405,N_14736);
xnor UO_1414 (O_1414,N_14723,N_14387);
or UO_1415 (O_1415,N_14120,N_14257);
nor UO_1416 (O_1416,N_14638,N_14778);
nor UO_1417 (O_1417,N_14255,N_14170);
nor UO_1418 (O_1418,N_14695,N_14238);
xnor UO_1419 (O_1419,N_14359,N_14227);
or UO_1420 (O_1420,N_14948,N_14924);
nor UO_1421 (O_1421,N_14333,N_14948);
and UO_1422 (O_1422,N_14137,N_14332);
or UO_1423 (O_1423,N_14314,N_14456);
nand UO_1424 (O_1424,N_14617,N_14980);
nand UO_1425 (O_1425,N_14307,N_14027);
or UO_1426 (O_1426,N_14933,N_14467);
and UO_1427 (O_1427,N_14873,N_14305);
and UO_1428 (O_1428,N_14046,N_14788);
and UO_1429 (O_1429,N_14011,N_14475);
xor UO_1430 (O_1430,N_14883,N_14217);
nand UO_1431 (O_1431,N_14940,N_14323);
nand UO_1432 (O_1432,N_14896,N_14909);
and UO_1433 (O_1433,N_14629,N_14217);
and UO_1434 (O_1434,N_14236,N_14585);
nand UO_1435 (O_1435,N_14006,N_14518);
nor UO_1436 (O_1436,N_14891,N_14212);
xor UO_1437 (O_1437,N_14636,N_14660);
nor UO_1438 (O_1438,N_14084,N_14955);
and UO_1439 (O_1439,N_14107,N_14152);
nand UO_1440 (O_1440,N_14534,N_14578);
or UO_1441 (O_1441,N_14389,N_14464);
or UO_1442 (O_1442,N_14418,N_14994);
xor UO_1443 (O_1443,N_14104,N_14714);
or UO_1444 (O_1444,N_14503,N_14736);
xnor UO_1445 (O_1445,N_14055,N_14022);
and UO_1446 (O_1446,N_14830,N_14996);
and UO_1447 (O_1447,N_14796,N_14213);
nor UO_1448 (O_1448,N_14459,N_14999);
nor UO_1449 (O_1449,N_14538,N_14973);
nor UO_1450 (O_1450,N_14972,N_14683);
or UO_1451 (O_1451,N_14718,N_14185);
and UO_1452 (O_1452,N_14718,N_14537);
nor UO_1453 (O_1453,N_14455,N_14127);
nor UO_1454 (O_1454,N_14162,N_14335);
and UO_1455 (O_1455,N_14129,N_14103);
nor UO_1456 (O_1456,N_14832,N_14491);
nor UO_1457 (O_1457,N_14716,N_14889);
xnor UO_1458 (O_1458,N_14964,N_14401);
xnor UO_1459 (O_1459,N_14844,N_14112);
nand UO_1460 (O_1460,N_14019,N_14748);
nand UO_1461 (O_1461,N_14323,N_14646);
nand UO_1462 (O_1462,N_14989,N_14477);
nand UO_1463 (O_1463,N_14323,N_14510);
nand UO_1464 (O_1464,N_14503,N_14185);
or UO_1465 (O_1465,N_14538,N_14248);
nor UO_1466 (O_1466,N_14838,N_14534);
or UO_1467 (O_1467,N_14175,N_14585);
xnor UO_1468 (O_1468,N_14697,N_14484);
or UO_1469 (O_1469,N_14440,N_14445);
and UO_1470 (O_1470,N_14172,N_14962);
nand UO_1471 (O_1471,N_14612,N_14282);
nand UO_1472 (O_1472,N_14075,N_14462);
nand UO_1473 (O_1473,N_14620,N_14889);
nor UO_1474 (O_1474,N_14047,N_14346);
or UO_1475 (O_1475,N_14112,N_14609);
and UO_1476 (O_1476,N_14477,N_14398);
nor UO_1477 (O_1477,N_14862,N_14220);
nor UO_1478 (O_1478,N_14466,N_14054);
or UO_1479 (O_1479,N_14341,N_14363);
and UO_1480 (O_1480,N_14799,N_14133);
and UO_1481 (O_1481,N_14651,N_14212);
nand UO_1482 (O_1482,N_14158,N_14110);
and UO_1483 (O_1483,N_14971,N_14675);
and UO_1484 (O_1484,N_14599,N_14929);
nor UO_1485 (O_1485,N_14647,N_14542);
xor UO_1486 (O_1486,N_14240,N_14355);
and UO_1487 (O_1487,N_14821,N_14549);
nand UO_1488 (O_1488,N_14252,N_14418);
nor UO_1489 (O_1489,N_14465,N_14705);
nor UO_1490 (O_1490,N_14206,N_14705);
nor UO_1491 (O_1491,N_14449,N_14100);
nand UO_1492 (O_1492,N_14982,N_14980);
and UO_1493 (O_1493,N_14490,N_14334);
nor UO_1494 (O_1494,N_14171,N_14320);
xor UO_1495 (O_1495,N_14928,N_14472);
or UO_1496 (O_1496,N_14539,N_14794);
nand UO_1497 (O_1497,N_14087,N_14533);
nand UO_1498 (O_1498,N_14954,N_14684);
and UO_1499 (O_1499,N_14790,N_14687);
or UO_1500 (O_1500,N_14623,N_14006);
and UO_1501 (O_1501,N_14140,N_14349);
xor UO_1502 (O_1502,N_14290,N_14025);
nor UO_1503 (O_1503,N_14383,N_14093);
and UO_1504 (O_1504,N_14358,N_14292);
nor UO_1505 (O_1505,N_14106,N_14348);
nor UO_1506 (O_1506,N_14345,N_14588);
nand UO_1507 (O_1507,N_14871,N_14741);
nor UO_1508 (O_1508,N_14263,N_14907);
or UO_1509 (O_1509,N_14162,N_14900);
or UO_1510 (O_1510,N_14189,N_14159);
and UO_1511 (O_1511,N_14779,N_14089);
and UO_1512 (O_1512,N_14124,N_14831);
and UO_1513 (O_1513,N_14146,N_14830);
nor UO_1514 (O_1514,N_14824,N_14461);
and UO_1515 (O_1515,N_14884,N_14571);
or UO_1516 (O_1516,N_14998,N_14526);
and UO_1517 (O_1517,N_14022,N_14162);
nand UO_1518 (O_1518,N_14378,N_14671);
xnor UO_1519 (O_1519,N_14828,N_14162);
nand UO_1520 (O_1520,N_14259,N_14753);
nor UO_1521 (O_1521,N_14550,N_14318);
or UO_1522 (O_1522,N_14393,N_14563);
nor UO_1523 (O_1523,N_14507,N_14618);
nand UO_1524 (O_1524,N_14351,N_14448);
nor UO_1525 (O_1525,N_14209,N_14296);
nand UO_1526 (O_1526,N_14756,N_14988);
nor UO_1527 (O_1527,N_14479,N_14982);
nand UO_1528 (O_1528,N_14294,N_14198);
nor UO_1529 (O_1529,N_14298,N_14267);
and UO_1530 (O_1530,N_14600,N_14336);
or UO_1531 (O_1531,N_14856,N_14507);
nand UO_1532 (O_1532,N_14653,N_14556);
nand UO_1533 (O_1533,N_14180,N_14580);
nand UO_1534 (O_1534,N_14390,N_14605);
or UO_1535 (O_1535,N_14709,N_14196);
and UO_1536 (O_1536,N_14872,N_14344);
nor UO_1537 (O_1537,N_14253,N_14727);
xnor UO_1538 (O_1538,N_14095,N_14207);
or UO_1539 (O_1539,N_14959,N_14193);
or UO_1540 (O_1540,N_14284,N_14745);
xnor UO_1541 (O_1541,N_14254,N_14191);
nor UO_1542 (O_1542,N_14579,N_14538);
and UO_1543 (O_1543,N_14140,N_14656);
nand UO_1544 (O_1544,N_14269,N_14849);
xnor UO_1545 (O_1545,N_14062,N_14152);
or UO_1546 (O_1546,N_14436,N_14264);
and UO_1547 (O_1547,N_14785,N_14696);
and UO_1548 (O_1548,N_14102,N_14194);
nor UO_1549 (O_1549,N_14810,N_14695);
nand UO_1550 (O_1550,N_14888,N_14705);
xnor UO_1551 (O_1551,N_14343,N_14460);
and UO_1552 (O_1552,N_14492,N_14005);
nand UO_1553 (O_1553,N_14472,N_14445);
xor UO_1554 (O_1554,N_14534,N_14042);
and UO_1555 (O_1555,N_14928,N_14219);
nor UO_1556 (O_1556,N_14175,N_14688);
and UO_1557 (O_1557,N_14244,N_14462);
and UO_1558 (O_1558,N_14319,N_14383);
nand UO_1559 (O_1559,N_14917,N_14650);
or UO_1560 (O_1560,N_14199,N_14752);
or UO_1561 (O_1561,N_14002,N_14429);
nand UO_1562 (O_1562,N_14504,N_14599);
nor UO_1563 (O_1563,N_14869,N_14277);
nand UO_1564 (O_1564,N_14877,N_14716);
nand UO_1565 (O_1565,N_14468,N_14485);
or UO_1566 (O_1566,N_14994,N_14760);
xnor UO_1567 (O_1567,N_14636,N_14772);
nand UO_1568 (O_1568,N_14350,N_14686);
nor UO_1569 (O_1569,N_14697,N_14351);
nand UO_1570 (O_1570,N_14846,N_14462);
nor UO_1571 (O_1571,N_14722,N_14434);
and UO_1572 (O_1572,N_14315,N_14855);
nand UO_1573 (O_1573,N_14550,N_14579);
and UO_1574 (O_1574,N_14549,N_14442);
or UO_1575 (O_1575,N_14982,N_14971);
nor UO_1576 (O_1576,N_14134,N_14813);
and UO_1577 (O_1577,N_14546,N_14698);
nand UO_1578 (O_1578,N_14455,N_14042);
and UO_1579 (O_1579,N_14297,N_14126);
or UO_1580 (O_1580,N_14524,N_14222);
nand UO_1581 (O_1581,N_14084,N_14106);
nand UO_1582 (O_1582,N_14030,N_14649);
or UO_1583 (O_1583,N_14515,N_14740);
and UO_1584 (O_1584,N_14000,N_14547);
nor UO_1585 (O_1585,N_14187,N_14503);
and UO_1586 (O_1586,N_14206,N_14566);
or UO_1587 (O_1587,N_14411,N_14904);
or UO_1588 (O_1588,N_14310,N_14349);
nand UO_1589 (O_1589,N_14250,N_14586);
nand UO_1590 (O_1590,N_14350,N_14413);
nor UO_1591 (O_1591,N_14927,N_14354);
or UO_1592 (O_1592,N_14494,N_14976);
xnor UO_1593 (O_1593,N_14683,N_14276);
xor UO_1594 (O_1594,N_14715,N_14401);
nand UO_1595 (O_1595,N_14697,N_14242);
or UO_1596 (O_1596,N_14513,N_14983);
or UO_1597 (O_1597,N_14361,N_14683);
nor UO_1598 (O_1598,N_14407,N_14085);
xnor UO_1599 (O_1599,N_14711,N_14631);
xor UO_1600 (O_1600,N_14300,N_14053);
or UO_1601 (O_1601,N_14236,N_14435);
nor UO_1602 (O_1602,N_14628,N_14934);
or UO_1603 (O_1603,N_14358,N_14017);
or UO_1604 (O_1604,N_14941,N_14301);
or UO_1605 (O_1605,N_14639,N_14795);
nand UO_1606 (O_1606,N_14628,N_14713);
and UO_1607 (O_1607,N_14430,N_14696);
and UO_1608 (O_1608,N_14035,N_14290);
nor UO_1609 (O_1609,N_14591,N_14230);
and UO_1610 (O_1610,N_14092,N_14061);
xor UO_1611 (O_1611,N_14529,N_14358);
nand UO_1612 (O_1612,N_14857,N_14242);
and UO_1613 (O_1613,N_14338,N_14004);
and UO_1614 (O_1614,N_14620,N_14633);
or UO_1615 (O_1615,N_14667,N_14148);
and UO_1616 (O_1616,N_14762,N_14044);
xor UO_1617 (O_1617,N_14996,N_14527);
nor UO_1618 (O_1618,N_14901,N_14721);
nand UO_1619 (O_1619,N_14396,N_14307);
nor UO_1620 (O_1620,N_14516,N_14535);
and UO_1621 (O_1621,N_14829,N_14860);
or UO_1622 (O_1622,N_14274,N_14838);
nand UO_1623 (O_1623,N_14915,N_14927);
nor UO_1624 (O_1624,N_14734,N_14956);
and UO_1625 (O_1625,N_14461,N_14730);
xnor UO_1626 (O_1626,N_14754,N_14993);
and UO_1627 (O_1627,N_14120,N_14288);
nand UO_1628 (O_1628,N_14623,N_14907);
or UO_1629 (O_1629,N_14146,N_14202);
and UO_1630 (O_1630,N_14276,N_14827);
or UO_1631 (O_1631,N_14822,N_14409);
and UO_1632 (O_1632,N_14536,N_14821);
and UO_1633 (O_1633,N_14266,N_14824);
nor UO_1634 (O_1634,N_14236,N_14036);
nand UO_1635 (O_1635,N_14829,N_14056);
nand UO_1636 (O_1636,N_14473,N_14370);
xnor UO_1637 (O_1637,N_14624,N_14765);
and UO_1638 (O_1638,N_14720,N_14420);
or UO_1639 (O_1639,N_14455,N_14214);
nand UO_1640 (O_1640,N_14937,N_14251);
nand UO_1641 (O_1641,N_14788,N_14263);
xnor UO_1642 (O_1642,N_14174,N_14246);
nand UO_1643 (O_1643,N_14858,N_14378);
and UO_1644 (O_1644,N_14478,N_14849);
nor UO_1645 (O_1645,N_14969,N_14854);
and UO_1646 (O_1646,N_14717,N_14301);
nor UO_1647 (O_1647,N_14141,N_14476);
and UO_1648 (O_1648,N_14085,N_14813);
or UO_1649 (O_1649,N_14827,N_14315);
nor UO_1650 (O_1650,N_14656,N_14530);
and UO_1651 (O_1651,N_14559,N_14021);
or UO_1652 (O_1652,N_14438,N_14512);
nand UO_1653 (O_1653,N_14966,N_14376);
nor UO_1654 (O_1654,N_14552,N_14876);
nand UO_1655 (O_1655,N_14107,N_14697);
or UO_1656 (O_1656,N_14084,N_14222);
xor UO_1657 (O_1657,N_14561,N_14347);
xnor UO_1658 (O_1658,N_14031,N_14402);
or UO_1659 (O_1659,N_14636,N_14001);
xor UO_1660 (O_1660,N_14298,N_14845);
xnor UO_1661 (O_1661,N_14226,N_14940);
nor UO_1662 (O_1662,N_14167,N_14292);
xor UO_1663 (O_1663,N_14544,N_14571);
or UO_1664 (O_1664,N_14226,N_14708);
and UO_1665 (O_1665,N_14756,N_14856);
and UO_1666 (O_1666,N_14491,N_14455);
or UO_1667 (O_1667,N_14580,N_14610);
nor UO_1668 (O_1668,N_14758,N_14216);
or UO_1669 (O_1669,N_14414,N_14196);
nor UO_1670 (O_1670,N_14463,N_14135);
or UO_1671 (O_1671,N_14467,N_14565);
xnor UO_1672 (O_1672,N_14653,N_14944);
nand UO_1673 (O_1673,N_14946,N_14815);
nor UO_1674 (O_1674,N_14237,N_14884);
nor UO_1675 (O_1675,N_14861,N_14126);
and UO_1676 (O_1676,N_14561,N_14200);
or UO_1677 (O_1677,N_14889,N_14208);
nor UO_1678 (O_1678,N_14374,N_14351);
and UO_1679 (O_1679,N_14275,N_14890);
nand UO_1680 (O_1680,N_14139,N_14434);
nor UO_1681 (O_1681,N_14093,N_14085);
and UO_1682 (O_1682,N_14147,N_14790);
and UO_1683 (O_1683,N_14196,N_14741);
or UO_1684 (O_1684,N_14268,N_14910);
or UO_1685 (O_1685,N_14526,N_14451);
or UO_1686 (O_1686,N_14184,N_14232);
nand UO_1687 (O_1687,N_14418,N_14431);
or UO_1688 (O_1688,N_14944,N_14273);
nand UO_1689 (O_1689,N_14478,N_14459);
and UO_1690 (O_1690,N_14126,N_14229);
or UO_1691 (O_1691,N_14867,N_14372);
nand UO_1692 (O_1692,N_14143,N_14750);
nand UO_1693 (O_1693,N_14360,N_14985);
and UO_1694 (O_1694,N_14497,N_14440);
or UO_1695 (O_1695,N_14001,N_14062);
and UO_1696 (O_1696,N_14664,N_14003);
nand UO_1697 (O_1697,N_14112,N_14444);
or UO_1698 (O_1698,N_14518,N_14141);
nor UO_1699 (O_1699,N_14631,N_14457);
or UO_1700 (O_1700,N_14239,N_14522);
nand UO_1701 (O_1701,N_14953,N_14222);
or UO_1702 (O_1702,N_14228,N_14682);
and UO_1703 (O_1703,N_14153,N_14776);
or UO_1704 (O_1704,N_14947,N_14789);
and UO_1705 (O_1705,N_14229,N_14637);
or UO_1706 (O_1706,N_14464,N_14775);
and UO_1707 (O_1707,N_14221,N_14024);
or UO_1708 (O_1708,N_14188,N_14255);
nor UO_1709 (O_1709,N_14789,N_14140);
or UO_1710 (O_1710,N_14909,N_14310);
nand UO_1711 (O_1711,N_14247,N_14099);
nand UO_1712 (O_1712,N_14667,N_14695);
nand UO_1713 (O_1713,N_14053,N_14359);
or UO_1714 (O_1714,N_14312,N_14186);
or UO_1715 (O_1715,N_14093,N_14628);
nor UO_1716 (O_1716,N_14288,N_14306);
and UO_1717 (O_1717,N_14868,N_14668);
and UO_1718 (O_1718,N_14129,N_14981);
nand UO_1719 (O_1719,N_14419,N_14525);
nand UO_1720 (O_1720,N_14560,N_14864);
nand UO_1721 (O_1721,N_14423,N_14546);
and UO_1722 (O_1722,N_14439,N_14117);
nand UO_1723 (O_1723,N_14460,N_14324);
or UO_1724 (O_1724,N_14735,N_14541);
nor UO_1725 (O_1725,N_14832,N_14217);
nor UO_1726 (O_1726,N_14421,N_14563);
or UO_1727 (O_1727,N_14006,N_14685);
nor UO_1728 (O_1728,N_14534,N_14757);
nor UO_1729 (O_1729,N_14521,N_14263);
nor UO_1730 (O_1730,N_14135,N_14323);
nor UO_1731 (O_1731,N_14713,N_14081);
or UO_1732 (O_1732,N_14999,N_14507);
nand UO_1733 (O_1733,N_14129,N_14849);
or UO_1734 (O_1734,N_14452,N_14459);
nand UO_1735 (O_1735,N_14537,N_14612);
or UO_1736 (O_1736,N_14322,N_14642);
and UO_1737 (O_1737,N_14878,N_14288);
nor UO_1738 (O_1738,N_14209,N_14869);
or UO_1739 (O_1739,N_14353,N_14467);
and UO_1740 (O_1740,N_14642,N_14121);
nand UO_1741 (O_1741,N_14652,N_14772);
xnor UO_1742 (O_1742,N_14987,N_14389);
nor UO_1743 (O_1743,N_14449,N_14068);
nor UO_1744 (O_1744,N_14948,N_14071);
nor UO_1745 (O_1745,N_14945,N_14478);
and UO_1746 (O_1746,N_14215,N_14233);
and UO_1747 (O_1747,N_14883,N_14555);
nor UO_1748 (O_1748,N_14436,N_14219);
nor UO_1749 (O_1749,N_14010,N_14654);
or UO_1750 (O_1750,N_14251,N_14368);
nand UO_1751 (O_1751,N_14001,N_14643);
xnor UO_1752 (O_1752,N_14388,N_14778);
and UO_1753 (O_1753,N_14794,N_14258);
nor UO_1754 (O_1754,N_14512,N_14590);
or UO_1755 (O_1755,N_14731,N_14191);
nor UO_1756 (O_1756,N_14524,N_14999);
and UO_1757 (O_1757,N_14488,N_14071);
nor UO_1758 (O_1758,N_14642,N_14830);
and UO_1759 (O_1759,N_14710,N_14886);
or UO_1760 (O_1760,N_14829,N_14055);
nand UO_1761 (O_1761,N_14993,N_14023);
nor UO_1762 (O_1762,N_14701,N_14245);
nand UO_1763 (O_1763,N_14373,N_14057);
nor UO_1764 (O_1764,N_14433,N_14974);
nand UO_1765 (O_1765,N_14559,N_14252);
nand UO_1766 (O_1766,N_14676,N_14461);
or UO_1767 (O_1767,N_14132,N_14620);
nand UO_1768 (O_1768,N_14254,N_14049);
nor UO_1769 (O_1769,N_14540,N_14297);
or UO_1770 (O_1770,N_14982,N_14985);
nor UO_1771 (O_1771,N_14053,N_14429);
or UO_1772 (O_1772,N_14707,N_14642);
or UO_1773 (O_1773,N_14194,N_14733);
nand UO_1774 (O_1774,N_14499,N_14383);
and UO_1775 (O_1775,N_14567,N_14867);
nand UO_1776 (O_1776,N_14026,N_14283);
xnor UO_1777 (O_1777,N_14338,N_14116);
nor UO_1778 (O_1778,N_14567,N_14696);
xor UO_1779 (O_1779,N_14425,N_14725);
nor UO_1780 (O_1780,N_14070,N_14837);
nand UO_1781 (O_1781,N_14935,N_14889);
nand UO_1782 (O_1782,N_14483,N_14017);
or UO_1783 (O_1783,N_14007,N_14394);
or UO_1784 (O_1784,N_14571,N_14358);
nor UO_1785 (O_1785,N_14651,N_14998);
and UO_1786 (O_1786,N_14538,N_14406);
and UO_1787 (O_1787,N_14355,N_14619);
and UO_1788 (O_1788,N_14369,N_14391);
or UO_1789 (O_1789,N_14595,N_14825);
nor UO_1790 (O_1790,N_14838,N_14396);
nor UO_1791 (O_1791,N_14870,N_14099);
and UO_1792 (O_1792,N_14244,N_14986);
and UO_1793 (O_1793,N_14478,N_14603);
nand UO_1794 (O_1794,N_14685,N_14598);
xor UO_1795 (O_1795,N_14132,N_14140);
or UO_1796 (O_1796,N_14270,N_14912);
nor UO_1797 (O_1797,N_14260,N_14095);
xor UO_1798 (O_1798,N_14509,N_14554);
and UO_1799 (O_1799,N_14356,N_14257);
nor UO_1800 (O_1800,N_14389,N_14532);
nor UO_1801 (O_1801,N_14424,N_14068);
nor UO_1802 (O_1802,N_14310,N_14960);
or UO_1803 (O_1803,N_14095,N_14044);
or UO_1804 (O_1804,N_14033,N_14499);
nor UO_1805 (O_1805,N_14602,N_14687);
nor UO_1806 (O_1806,N_14494,N_14785);
xor UO_1807 (O_1807,N_14226,N_14875);
and UO_1808 (O_1808,N_14491,N_14520);
or UO_1809 (O_1809,N_14757,N_14624);
or UO_1810 (O_1810,N_14570,N_14214);
nand UO_1811 (O_1811,N_14796,N_14961);
and UO_1812 (O_1812,N_14711,N_14664);
nand UO_1813 (O_1813,N_14796,N_14382);
nand UO_1814 (O_1814,N_14267,N_14641);
nand UO_1815 (O_1815,N_14444,N_14467);
nand UO_1816 (O_1816,N_14374,N_14527);
nand UO_1817 (O_1817,N_14472,N_14507);
nand UO_1818 (O_1818,N_14910,N_14109);
xor UO_1819 (O_1819,N_14993,N_14578);
xnor UO_1820 (O_1820,N_14643,N_14600);
xnor UO_1821 (O_1821,N_14689,N_14783);
nor UO_1822 (O_1822,N_14569,N_14051);
or UO_1823 (O_1823,N_14204,N_14153);
nor UO_1824 (O_1824,N_14014,N_14455);
or UO_1825 (O_1825,N_14583,N_14777);
nand UO_1826 (O_1826,N_14689,N_14853);
nor UO_1827 (O_1827,N_14607,N_14315);
or UO_1828 (O_1828,N_14118,N_14411);
nand UO_1829 (O_1829,N_14535,N_14645);
or UO_1830 (O_1830,N_14464,N_14986);
nor UO_1831 (O_1831,N_14463,N_14795);
nor UO_1832 (O_1832,N_14983,N_14204);
or UO_1833 (O_1833,N_14572,N_14778);
or UO_1834 (O_1834,N_14454,N_14762);
and UO_1835 (O_1835,N_14768,N_14676);
nand UO_1836 (O_1836,N_14729,N_14620);
or UO_1837 (O_1837,N_14461,N_14488);
nor UO_1838 (O_1838,N_14514,N_14870);
nor UO_1839 (O_1839,N_14613,N_14556);
or UO_1840 (O_1840,N_14164,N_14339);
and UO_1841 (O_1841,N_14915,N_14175);
or UO_1842 (O_1842,N_14128,N_14031);
or UO_1843 (O_1843,N_14142,N_14626);
or UO_1844 (O_1844,N_14104,N_14554);
and UO_1845 (O_1845,N_14044,N_14241);
or UO_1846 (O_1846,N_14497,N_14392);
and UO_1847 (O_1847,N_14527,N_14044);
and UO_1848 (O_1848,N_14477,N_14023);
or UO_1849 (O_1849,N_14761,N_14083);
and UO_1850 (O_1850,N_14444,N_14191);
nor UO_1851 (O_1851,N_14130,N_14398);
nor UO_1852 (O_1852,N_14116,N_14350);
and UO_1853 (O_1853,N_14257,N_14360);
xor UO_1854 (O_1854,N_14568,N_14869);
or UO_1855 (O_1855,N_14399,N_14248);
or UO_1856 (O_1856,N_14834,N_14135);
nand UO_1857 (O_1857,N_14606,N_14058);
or UO_1858 (O_1858,N_14606,N_14315);
and UO_1859 (O_1859,N_14282,N_14041);
nor UO_1860 (O_1860,N_14841,N_14638);
nor UO_1861 (O_1861,N_14609,N_14885);
or UO_1862 (O_1862,N_14764,N_14053);
nand UO_1863 (O_1863,N_14500,N_14274);
or UO_1864 (O_1864,N_14338,N_14101);
and UO_1865 (O_1865,N_14206,N_14755);
and UO_1866 (O_1866,N_14672,N_14693);
nand UO_1867 (O_1867,N_14403,N_14282);
nand UO_1868 (O_1868,N_14884,N_14923);
and UO_1869 (O_1869,N_14782,N_14729);
xnor UO_1870 (O_1870,N_14984,N_14487);
nand UO_1871 (O_1871,N_14979,N_14004);
or UO_1872 (O_1872,N_14155,N_14402);
and UO_1873 (O_1873,N_14699,N_14957);
or UO_1874 (O_1874,N_14174,N_14949);
nand UO_1875 (O_1875,N_14411,N_14499);
or UO_1876 (O_1876,N_14064,N_14471);
or UO_1877 (O_1877,N_14283,N_14310);
or UO_1878 (O_1878,N_14698,N_14497);
nor UO_1879 (O_1879,N_14955,N_14479);
nand UO_1880 (O_1880,N_14704,N_14468);
and UO_1881 (O_1881,N_14122,N_14301);
nand UO_1882 (O_1882,N_14885,N_14817);
nand UO_1883 (O_1883,N_14021,N_14884);
and UO_1884 (O_1884,N_14076,N_14643);
nor UO_1885 (O_1885,N_14972,N_14419);
or UO_1886 (O_1886,N_14009,N_14199);
or UO_1887 (O_1887,N_14239,N_14494);
xor UO_1888 (O_1888,N_14468,N_14143);
nor UO_1889 (O_1889,N_14174,N_14854);
nor UO_1890 (O_1890,N_14707,N_14109);
or UO_1891 (O_1891,N_14749,N_14283);
or UO_1892 (O_1892,N_14090,N_14800);
or UO_1893 (O_1893,N_14782,N_14450);
or UO_1894 (O_1894,N_14271,N_14663);
nand UO_1895 (O_1895,N_14793,N_14928);
nor UO_1896 (O_1896,N_14904,N_14037);
and UO_1897 (O_1897,N_14338,N_14973);
nand UO_1898 (O_1898,N_14059,N_14317);
and UO_1899 (O_1899,N_14308,N_14356);
nand UO_1900 (O_1900,N_14895,N_14452);
nand UO_1901 (O_1901,N_14477,N_14188);
and UO_1902 (O_1902,N_14333,N_14321);
nand UO_1903 (O_1903,N_14633,N_14338);
nor UO_1904 (O_1904,N_14680,N_14758);
and UO_1905 (O_1905,N_14557,N_14849);
and UO_1906 (O_1906,N_14411,N_14653);
nor UO_1907 (O_1907,N_14912,N_14917);
and UO_1908 (O_1908,N_14061,N_14174);
or UO_1909 (O_1909,N_14980,N_14565);
nand UO_1910 (O_1910,N_14515,N_14366);
and UO_1911 (O_1911,N_14262,N_14349);
nand UO_1912 (O_1912,N_14842,N_14377);
xnor UO_1913 (O_1913,N_14416,N_14119);
and UO_1914 (O_1914,N_14423,N_14067);
nand UO_1915 (O_1915,N_14700,N_14401);
or UO_1916 (O_1916,N_14381,N_14978);
nor UO_1917 (O_1917,N_14192,N_14258);
nand UO_1918 (O_1918,N_14159,N_14776);
nand UO_1919 (O_1919,N_14903,N_14111);
or UO_1920 (O_1920,N_14947,N_14211);
and UO_1921 (O_1921,N_14714,N_14830);
nor UO_1922 (O_1922,N_14690,N_14724);
nor UO_1923 (O_1923,N_14012,N_14475);
nand UO_1924 (O_1924,N_14044,N_14301);
nor UO_1925 (O_1925,N_14878,N_14444);
nor UO_1926 (O_1926,N_14305,N_14655);
and UO_1927 (O_1927,N_14611,N_14463);
or UO_1928 (O_1928,N_14629,N_14845);
nor UO_1929 (O_1929,N_14812,N_14958);
nor UO_1930 (O_1930,N_14773,N_14316);
nand UO_1931 (O_1931,N_14730,N_14937);
or UO_1932 (O_1932,N_14706,N_14336);
and UO_1933 (O_1933,N_14069,N_14380);
xnor UO_1934 (O_1934,N_14337,N_14827);
or UO_1935 (O_1935,N_14354,N_14323);
or UO_1936 (O_1936,N_14172,N_14049);
nor UO_1937 (O_1937,N_14358,N_14235);
and UO_1938 (O_1938,N_14273,N_14854);
xnor UO_1939 (O_1939,N_14203,N_14199);
nand UO_1940 (O_1940,N_14644,N_14844);
and UO_1941 (O_1941,N_14222,N_14746);
nand UO_1942 (O_1942,N_14077,N_14374);
nand UO_1943 (O_1943,N_14299,N_14912);
or UO_1944 (O_1944,N_14524,N_14898);
or UO_1945 (O_1945,N_14687,N_14351);
nand UO_1946 (O_1946,N_14528,N_14629);
or UO_1947 (O_1947,N_14967,N_14384);
nor UO_1948 (O_1948,N_14127,N_14524);
nand UO_1949 (O_1949,N_14141,N_14939);
and UO_1950 (O_1950,N_14110,N_14620);
nand UO_1951 (O_1951,N_14424,N_14924);
nand UO_1952 (O_1952,N_14176,N_14001);
or UO_1953 (O_1953,N_14144,N_14178);
and UO_1954 (O_1954,N_14087,N_14023);
nor UO_1955 (O_1955,N_14580,N_14318);
or UO_1956 (O_1956,N_14033,N_14897);
nor UO_1957 (O_1957,N_14811,N_14494);
nand UO_1958 (O_1958,N_14169,N_14949);
nor UO_1959 (O_1959,N_14506,N_14975);
and UO_1960 (O_1960,N_14022,N_14643);
or UO_1961 (O_1961,N_14107,N_14493);
nor UO_1962 (O_1962,N_14151,N_14833);
nand UO_1963 (O_1963,N_14854,N_14834);
nand UO_1964 (O_1964,N_14425,N_14450);
and UO_1965 (O_1965,N_14706,N_14610);
nor UO_1966 (O_1966,N_14862,N_14972);
nor UO_1967 (O_1967,N_14703,N_14479);
nor UO_1968 (O_1968,N_14432,N_14159);
or UO_1969 (O_1969,N_14936,N_14358);
xnor UO_1970 (O_1970,N_14620,N_14744);
nand UO_1971 (O_1971,N_14774,N_14917);
nand UO_1972 (O_1972,N_14517,N_14279);
and UO_1973 (O_1973,N_14128,N_14740);
xor UO_1974 (O_1974,N_14221,N_14770);
nand UO_1975 (O_1975,N_14272,N_14355);
nor UO_1976 (O_1976,N_14964,N_14010);
and UO_1977 (O_1977,N_14065,N_14421);
and UO_1978 (O_1978,N_14682,N_14194);
nand UO_1979 (O_1979,N_14325,N_14028);
xnor UO_1980 (O_1980,N_14063,N_14078);
nor UO_1981 (O_1981,N_14588,N_14255);
nor UO_1982 (O_1982,N_14248,N_14820);
or UO_1983 (O_1983,N_14804,N_14138);
and UO_1984 (O_1984,N_14364,N_14866);
xnor UO_1985 (O_1985,N_14307,N_14458);
xor UO_1986 (O_1986,N_14866,N_14970);
xor UO_1987 (O_1987,N_14437,N_14615);
or UO_1988 (O_1988,N_14182,N_14020);
nand UO_1989 (O_1989,N_14065,N_14167);
nand UO_1990 (O_1990,N_14515,N_14633);
nand UO_1991 (O_1991,N_14734,N_14413);
and UO_1992 (O_1992,N_14230,N_14018);
nor UO_1993 (O_1993,N_14342,N_14661);
nor UO_1994 (O_1994,N_14385,N_14991);
or UO_1995 (O_1995,N_14421,N_14049);
and UO_1996 (O_1996,N_14116,N_14490);
and UO_1997 (O_1997,N_14403,N_14555);
and UO_1998 (O_1998,N_14524,N_14612);
or UO_1999 (O_1999,N_14919,N_14565);
endmodule