module basic_2500_25000_3000_4_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18861,N_18862,N_18863,N_18864,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19035,N_19036,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19053,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19082,N_19083,N_19084,N_19085,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19255,N_19256,N_19257,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19293,N_19294,N_19295,N_19296,N_19297,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19411,N_19412,N_19413,N_19414,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19456,N_19457,N_19458,N_19459,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19659,N_19660,N_19661,N_19662,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20232,N_20233,N_20234,N_20235,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20394,N_20395,N_20396,N_20397,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20803,N_20804,N_20805,N_20806,N_20807,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21171,N_21172,N_21174,N_21175,N_21176,N_21177,N_21178,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21200,N_21201,N_21202,N_21203,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21336,N_21337,N_21338,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21614,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21853,N_21854,N_21855,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21869,N_21870,N_21871,N_21872,N_21873,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21901,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21996,N_21997,N_21998,N_21999,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22066,N_22068,N_22069,N_22070,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22453,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22476,N_22477,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22606,N_22607,N_22608,N_22609,N_22610,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22772,N_22773,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22787,N_22788,N_22789,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23100,N_23101,N_23102,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23651,N_23652,N_23653,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24039,N_24040,N_24041,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24573,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24609,N_24610,N_24611,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24635,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24869,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_1538,In_1418);
nand U1 (N_1,In_1372,In_967);
and U2 (N_2,In_413,In_1749);
and U3 (N_3,In_2111,In_2480);
xor U4 (N_4,In_2246,In_501);
xor U5 (N_5,In_498,In_745);
nor U6 (N_6,In_797,In_2410);
nand U7 (N_7,In_1820,In_258);
and U8 (N_8,In_1825,In_712);
and U9 (N_9,In_199,In_1872);
or U10 (N_10,In_755,In_2249);
nor U11 (N_11,In_1821,In_2148);
and U12 (N_12,In_1889,In_1900);
nor U13 (N_13,In_2348,In_2220);
xnor U14 (N_14,In_1589,In_2451);
nor U15 (N_15,In_1163,In_2183);
nor U16 (N_16,In_610,In_1436);
xnor U17 (N_17,In_2232,In_185);
and U18 (N_18,In_399,In_17);
nand U19 (N_19,In_1153,In_1009);
or U20 (N_20,In_2474,In_791);
xnor U21 (N_21,In_1050,In_828);
xor U22 (N_22,In_1575,In_565);
xor U23 (N_23,In_2096,In_2021);
xnor U24 (N_24,In_1426,In_603);
and U25 (N_25,In_694,In_1063);
and U26 (N_26,In_1364,In_1099);
and U27 (N_27,In_1524,In_1242);
or U28 (N_28,In_597,In_2364);
nand U29 (N_29,In_1791,In_1542);
nor U30 (N_30,In_1065,In_841);
xor U31 (N_31,In_2282,In_950);
xnor U32 (N_32,In_25,In_545);
or U33 (N_33,In_2456,In_669);
xnor U34 (N_34,In_2238,In_1654);
and U35 (N_35,In_1873,In_162);
nand U36 (N_36,In_1990,In_1579);
xor U37 (N_37,In_261,In_1472);
or U38 (N_38,In_2036,In_1265);
nor U39 (N_39,In_2375,In_2254);
or U40 (N_40,In_2491,In_123);
xnor U41 (N_41,In_1493,In_2022);
or U42 (N_42,In_1862,In_2065);
nor U43 (N_43,In_1371,In_2446);
and U44 (N_44,In_856,In_2035);
and U45 (N_45,In_850,In_590);
nand U46 (N_46,In_2083,In_2122);
or U47 (N_47,In_728,In_1813);
nor U48 (N_48,In_553,In_1156);
nor U49 (N_49,In_2050,In_1963);
and U50 (N_50,In_549,In_2109);
nand U51 (N_51,In_1856,In_1478);
and U52 (N_52,In_1832,In_1802);
xor U53 (N_53,In_666,In_1222);
or U54 (N_54,In_8,In_508);
nand U55 (N_55,In_382,In_426);
nand U56 (N_56,In_1420,In_1836);
nor U57 (N_57,In_1313,In_319);
xor U58 (N_58,In_1494,In_527);
or U59 (N_59,In_686,In_2316);
or U60 (N_60,In_1609,In_352);
and U61 (N_61,In_1535,In_1582);
nand U62 (N_62,In_1578,In_264);
xor U63 (N_63,In_1572,In_2221);
nand U64 (N_64,In_251,In_139);
and U65 (N_65,In_917,In_443);
and U66 (N_66,In_1347,In_108);
nand U67 (N_67,In_2310,In_2098);
nor U68 (N_68,In_751,In_223);
nor U69 (N_69,In_1017,In_302);
xnor U70 (N_70,In_847,In_1714);
nand U71 (N_71,In_1552,In_1845);
or U72 (N_72,In_1505,In_102);
nor U73 (N_73,In_490,In_286);
nor U74 (N_74,In_1893,In_1079);
nor U75 (N_75,In_2139,In_2132);
or U76 (N_76,In_100,In_1783);
nor U77 (N_77,In_132,In_140);
xor U78 (N_78,In_457,In_349);
xor U79 (N_79,In_744,In_485);
or U80 (N_80,In_359,In_853);
or U81 (N_81,In_418,In_2289);
nor U82 (N_82,In_2234,In_2177);
nor U83 (N_83,In_768,In_699);
nand U84 (N_84,In_1119,In_1058);
nor U85 (N_85,In_305,In_188);
nor U86 (N_86,In_294,In_40);
nor U87 (N_87,In_1546,In_354);
and U88 (N_88,In_2453,In_697);
or U89 (N_89,In_406,In_27);
nand U90 (N_90,In_723,In_2360);
or U91 (N_91,In_506,In_400);
and U92 (N_92,In_2058,In_390);
or U93 (N_93,In_1811,In_1988);
nor U94 (N_94,In_1620,In_1249);
or U95 (N_95,In_1155,In_130);
nand U96 (N_96,In_2199,In_2012);
nor U97 (N_97,In_1788,In_980);
nor U98 (N_98,In_1670,In_1742);
nor U99 (N_99,In_1210,In_14);
or U100 (N_100,In_1462,In_907);
and U101 (N_101,In_2019,In_1111);
or U102 (N_102,In_1209,In_1735);
nor U103 (N_103,In_1322,In_1957);
nand U104 (N_104,In_1699,In_2013);
nand U105 (N_105,In_2297,In_480);
xnor U106 (N_106,In_1011,In_1165);
nor U107 (N_107,In_2286,In_156);
or U108 (N_108,In_126,In_2075);
nor U109 (N_109,In_1149,In_1154);
nand U110 (N_110,In_2349,In_2433);
or U111 (N_111,In_557,In_863);
xor U112 (N_112,In_74,In_604);
or U113 (N_113,In_1396,In_205);
and U114 (N_114,In_756,In_781);
nor U115 (N_115,In_2495,In_763);
or U116 (N_116,In_88,In_1930);
nor U117 (N_117,In_635,In_137);
nor U118 (N_118,In_345,In_795);
or U119 (N_119,In_739,In_2396);
nand U120 (N_120,In_2178,In_2329);
nand U121 (N_121,In_1866,In_952);
nor U122 (N_122,In_670,In_2219);
xnor U123 (N_123,In_2413,In_1554);
and U124 (N_124,In_22,In_2452);
nand U125 (N_125,In_1214,In_1675);
and U126 (N_126,In_974,In_81);
or U127 (N_127,In_1199,In_2266);
and U128 (N_128,In_1787,In_1328);
xnor U129 (N_129,In_1905,In_1270);
nor U130 (N_130,In_1230,In_1726);
or U131 (N_131,In_63,In_1687);
xor U132 (N_132,In_1857,In_1281);
and U133 (N_133,In_178,In_1176);
and U134 (N_134,In_1037,In_454);
nand U135 (N_135,In_1122,In_1168);
and U136 (N_136,In_877,In_417);
nor U137 (N_137,In_988,In_2273);
xnor U138 (N_138,In_1728,In_5);
or U139 (N_139,In_957,In_1236);
and U140 (N_140,In_1458,In_1838);
and U141 (N_141,In_634,In_150);
nand U142 (N_142,In_2293,In_379);
nand U143 (N_143,In_1262,In_1036);
xnor U144 (N_144,In_2357,In_978);
and U145 (N_145,In_1485,In_1432);
nor U146 (N_146,In_762,In_2398);
nand U147 (N_147,In_427,In_1019);
xor U148 (N_148,In_1690,In_584);
and U149 (N_149,In_279,In_2130);
nor U150 (N_150,In_249,In_1439);
xnor U151 (N_151,In_281,In_1522);
nor U152 (N_152,In_1745,In_195);
nor U153 (N_153,In_1400,In_98);
nor U154 (N_154,In_2296,In_190);
xnor U155 (N_155,In_1688,In_1875);
xor U156 (N_156,In_1577,In_122);
and U157 (N_157,In_805,In_227);
nor U158 (N_158,In_391,In_1683);
and U159 (N_159,In_1319,In_1401);
and U160 (N_160,In_1084,In_678);
or U161 (N_161,In_82,In_1502);
xor U162 (N_162,In_2113,In_606);
nand U163 (N_163,In_912,In_882);
or U164 (N_164,In_821,In_394);
and U165 (N_165,In_2205,In_840);
xnor U166 (N_166,In_1549,In_1488);
nand U167 (N_167,In_410,In_753);
or U168 (N_168,In_1006,In_520);
xor U169 (N_169,In_87,In_1641);
or U170 (N_170,In_1539,In_552);
nand U171 (N_171,In_1561,In_1061);
and U172 (N_172,In_1588,In_1809);
nor U173 (N_173,In_1012,In_2313);
or U174 (N_174,In_922,In_2270);
nor U175 (N_175,In_541,In_1141);
nor U176 (N_176,In_1747,In_381);
xor U177 (N_177,In_213,In_968);
xnor U178 (N_178,In_2034,In_1890);
xor U179 (N_179,In_1217,In_1151);
nor U180 (N_180,In_2274,In_1438);
nor U181 (N_181,In_1943,In_2179);
and U182 (N_182,In_2124,In_2346);
or U183 (N_183,In_1049,In_892);
xnor U184 (N_184,In_1088,In_1479);
or U185 (N_185,In_422,In_1672);
nor U186 (N_186,In_533,In_2041);
nor U187 (N_187,In_471,In_1105);
and U188 (N_188,In_1080,In_1302);
and U189 (N_189,In_144,In_374);
nor U190 (N_190,In_1174,In_2324);
xor U191 (N_191,In_2020,In_326);
nand U192 (N_192,In_121,In_1570);
nor U193 (N_193,In_519,In_1877);
and U194 (N_194,In_1858,In_511);
and U195 (N_195,In_53,In_1374);
nand U196 (N_196,In_865,In_857);
nand U197 (N_197,In_529,In_1020);
nand U198 (N_198,In_2425,In_1638);
xnor U199 (N_199,In_2067,In_99);
xnor U200 (N_200,In_702,In_2315);
and U201 (N_201,In_11,In_438);
nor U202 (N_202,In_1108,In_2029);
xnor U203 (N_203,In_528,In_2243);
and U204 (N_204,In_2319,In_34);
or U205 (N_205,In_1022,In_1972);
nor U206 (N_206,In_748,In_307);
or U207 (N_207,In_1780,In_367);
and U208 (N_208,In_433,In_2088);
or U209 (N_209,In_2033,In_1334);
or U210 (N_210,In_2217,In_1441);
and U211 (N_211,In_1923,In_2107);
nor U212 (N_212,In_774,In_435);
xnor U213 (N_213,In_1606,In_740);
nand U214 (N_214,In_1311,In_2371);
xnor U215 (N_215,In_2429,In_547);
nand U216 (N_216,In_1078,In_2361);
and U217 (N_217,In_1658,In_1650);
nand U218 (N_218,In_871,In_1786);
and U219 (N_219,In_1186,In_158);
nand U220 (N_220,In_1381,In_1417);
nor U221 (N_221,In_256,In_924);
xnor U222 (N_222,In_1619,In_2247);
or U223 (N_223,In_1451,In_2472);
nor U224 (N_224,In_908,In_66);
or U225 (N_225,In_331,In_535);
nand U226 (N_226,In_1237,In_929);
xnor U227 (N_227,In_802,In_487);
nand U228 (N_228,In_278,In_1275);
xnor U229 (N_229,In_2197,In_210);
or U230 (N_230,In_1693,In_887);
nor U231 (N_231,In_1805,In_784);
nand U232 (N_232,In_465,In_2027);
and U233 (N_233,In_308,In_78);
or U234 (N_234,In_1949,In_591);
nor U235 (N_235,In_2117,In_870);
or U236 (N_236,In_1402,In_742);
and U237 (N_237,In_2216,In_1365);
and U238 (N_238,In_1481,In_69);
or U239 (N_239,In_1770,In_179);
xnor U240 (N_240,In_690,In_1941);
nand U241 (N_241,In_45,In_288);
nor U242 (N_242,In_676,In_2135);
and U243 (N_243,In_4,In_1697);
xor U244 (N_244,In_1536,In_530);
nor U245 (N_245,In_2407,In_2253);
and U246 (N_246,In_1795,In_1766);
nor U247 (N_247,In_1917,In_1031);
and U248 (N_248,In_614,In_726);
and U249 (N_249,In_2261,In_2223);
nor U250 (N_250,In_543,In_103);
xnor U251 (N_251,In_660,In_1405);
and U252 (N_252,In_1898,In_1700);
nor U253 (N_253,In_682,In_1389);
nand U254 (N_254,In_298,In_263);
xor U255 (N_255,In_706,In_270);
and U256 (N_256,In_1404,In_783);
nand U257 (N_257,In_1602,In_2461);
nor U258 (N_258,In_1733,In_478);
and U259 (N_259,In_464,In_155);
nor U260 (N_260,In_641,In_1568);
nor U261 (N_261,In_1789,In_200);
nand U262 (N_262,In_1342,In_1173);
xor U263 (N_263,In_854,In_1777);
nor U264 (N_264,In_194,In_55);
xor U265 (N_265,In_1376,In_564);
nor U266 (N_266,In_383,In_2030);
and U267 (N_267,In_561,In_1066);
nor U268 (N_268,In_1185,In_656);
xor U269 (N_269,In_949,In_348);
nor U270 (N_270,In_2131,In_644);
xor U271 (N_271,In_442,In_2073);
nor U272 (N_272,In_975,In_1920);
nand U273 (N_273,In_1500,In_1495);
nor U274 (N_274,In_215,In_601);
or U275 (N_275,In_1534,In_2342);
or U276 (N_276,In_786,In_482);
xor U277 (N_277,In_536,In_260);
nor U278 (N_278,In_860,In_2385);
and U279 (N_279,In_79,In_1403);
and U280 (N_280,In_1509,In_142);
xor U281 (N_281,In_2275,In_693);
or U282 (N_282,In_1955,In_1999);
nand U283 (N_283,In_1296,In_581);
nand U284 (N_284,In_268,In_698);
xnor U285 (N_285,In_542,In_1617);
or U286 (N_286,In_41,In_1895);
or U287 (N_287,In_611,In_2031);
nor U288 (N_288,In_695,In_2494);
xnor U289 (N_289,In_759,In_1718);
xnor U290 (N_290,In_1909,In_677);
nor U291 (N_291,In_2248,In_562);
and U292 (N_292,In_996,In_1892);
nor U293 (N_293,In_1759,In_350);
nor U294 (N_294,In_28,In_869);
nor U295 (N_295,In_765,In_167);
nor U296 (N_296,In_1684,In_112);
and U297 (N_297,In_159,In_115);
and U298 (N_298,In_979,In_2432);
and U299 (N_299,In_2448,In_1416);
or U300 (N_300,In_1016,In_369);
nand U301 (N_301,In_1419,In_2160);
nor U302 (N_302,In_173,In_626);
or U303 (N_303,In_816,In_1279);
xor U304 (N_304,In_1375,In_954);
nand U305 (N_305,In_789,In_1130);
nand U306 (N_306,In_448,In_2242);
or U307 (N_307,In_211,In_1722);
nor U308 (N_308,In_1682,In_1064);
and U309 (N_309,In_880,In_415);
and U310 (N_310,In_2295,In_1707);
xnor U311 (N_311,In_741,In_1355);
xnor U312 (N_312,In_377,In_1126);
nor U313 (N_313,In_1188,In_1255);
nand U314 (N_314,In_1005,In_1986);
nor U315 (N_315,In_1540,In_2158);
nor U316 (N_316,In_1271,In_475);
nor U317 (N_317,In_1278,In_1286);
xnor U318 (N_318,In_546,In_1197);
nor U319 (N_319,In_1812,In_1600);
xnor U320 (N_320,In_193,In_2490);
xnor U321 (N_321,In_2365,In_2268);
nand U322 (N_322,In_842,In_738);
or U323 (N_323,In_1339,In_505);
and U324 (N_324,In_1213,In_717);
nor U325 (N_325,In_1003,In_537);
nand U326 (N_326,In_1387,In_1719);
or U327 (N_327,In_2047,In_101);
nand U328 (N_328,In_220,In_1706);
nor U329 (N_329,In_2406,In_1198);
nor U330 (N_330,In_884,In_360);
or U331 (N_331,In_244,In_1558);
nand U332 (N_332,In_772,In_868);
nor U333 (N_333,In_2269,In_1627);
nand U334 (N_334,In_515,In_1407);
or U335 (N_335,In_1574,In_2322);
and U336 (N_336,In_1916,In_1659);
xnor U337 (N_337,In_469,In_1263);
nand U338 (N_338,In_2350,In_300);
and U339 (N_339,In_2392,In_813);
nor U340 (N_340,In_1204,In_1459);
nand U341 (N_341,In_970,In_339);
and U342 (N_342,In_1424,In_1656);
xor U343 (N_343,In_1876,In_2231);
xnor U344 (N_344,In_1622,In_2264);
or U345 (N_345,In_1363,In_1959);
nand U346 (N_346,In_1450,In_995);
nand U347 (N_347,In_1482,In_262);
or U348 (N_348,In_107,In_2175);
nand U349 (N_349,In_787,In_1804);
xor U350 (N_350,In_711,In_1545);
xnor U351 (N_351,In_493,In_2184);
or U352 (N_352,In_309,In_60);
nor U353 (N_353,In_114,In_1624);
nand U354 (N_354,In_1447,In_673);
xnor U355 (N_355,In_990,In_737);
nand U356 (N_356,In_1254,In_1140);
or U357 (N_357,In_2009,In_2189);
nand U358 (N_358,In_92,In_1694);
or U359 (N_359,In_1984,In_1598);
or U360 (N_360,In_794,In_2064);
or U361 (N_361,In_2068,In_387);
nand U362 (N_362,In_1928,In_2087);
or U363 (N_363,In_2108,In_1044);
or U364 (N_364,In_449,In_727);
and U365 (N_365,In_1497,In_1052);
xnor U366 (N_366,In_2482,In_1239);
or U367 (N_367,In_72,In_1764);
or U368 (N_368,In_1644,In_187);
xor U369 (N_369,In_2086,In_652);
xnor U370 (N_370,In_109,In_1962);
or U371 (N_371,In_1625,In_2389);
or U372 (N_372,In_648,In_732);
xor U373 (N_373,In_378,In_2468);
and U374 (N_374,In_1531,In_1234);
xnor U375 (N_375,In_643,In_70);
nor U376 (N_376,In_600,In_1685);
or U377 (N_377,In_1580,In_642);
and U378 (N_378,In_1671,In_1038);
nand U379 (N_379,In_1429,In_2478);
xnor U380 (N_380,In_583,In_342);
and U381 (N_381,In_1354,In_152);
and U382 (N_382,In_609,In_290);
nor U383 (N_383,In_1935,In_332);
nand U384 (N_384,In_110,In_1142);
xor U385 (N_385,In_253,In_1618);
or U386 (N_386,In_250,In_687);
or U387 (N_387,In_2442,In_1260);
or U388 (N_388,In_2081,In_1067);
or U389 (N_389,In_1915,In_1705);
and U390 (N_390,In_1740,In_1807);
and U391 (N_391,In_218,In_602);
and U392 (N_392,In_2048,In_916);
xor U393 (N_393,In_2162,In_793);
xor U394 (N_394,In_1712,In_2481);
nor U395 (N_395,In_234,In_1307);
xnor U396 (N_396,In_764,In_754);
or U397 (N_397,In_2118,In_208);
nand U398 (N_398,In_1824,In_1288);
or U399 (N_399,In_274,In_1193);
and U400 (N_400,In_900,In_835);
or U401 (N_401,In_1292,In_1732);
xor U402 (N_402,In_36,In_1258);
xor U403 (N_403,In_472,In_1362);
nand U404 (N_404,In_2203,In_1483);
and U405 (N_405,In_380,In_1903);
nand U406 (N_406,In_1397,In_859);
nand U407 (N_407,In_1072,In_586);
and U408 (N_408,In_2479,In_2103);
nor U409 (N_409,In_1103,In_1135);
or U410 (N_410,In_2016,In_1267);
nor U411 (N_411,In_1390,In_640);
or U412 (N_412,In_1259,In_225);
nor U413 (N_413,In_1569,In_26);
or U414 (N_414,In_799,In_2460);
nor U415 (N_415,In_650,In_133);
xor U416 (N_416,In_2070,In_423);
nand U417 (N_417,In_289,In_999);
nand U418 (N_418,In_2386,In_6);
xnor U419 (N_419,In_1982,In_2260);
nand U420 (N_420,In_1175,In_1094);
nand U421 (N_421,In_269,In_1901);
and U422 (N_422,In_1716,In_920);
and U423 (N_423,In_1781,In_1810);
nor U424 (N_424,In_1116,In_408);
nand U425 (N_425,In_595,In_1253);
nand U426 (N_426,In_1002,In_1703);
nor U427 (N_427,In_2049,In_811);
nand U428 (N_428,In_58,In_843);
xor U429 (N_429,In_1615,In_1218);
nor U430 (N_430,In_1326,In_807);
nor U431 (N_431,In_1384,In_1132);
and U432 (N_432,In_2416,In_2218);
or U433 (N_433,In_452,In_1434);
nand U434 (N_434,In_2492,In_312);
and U435 (N_435,In_2191,In_665);
and U436 (N_436,In_2280,In_684);
nand U437 (N_437,In_2,In_2236);
nor U438 (N_438,In_855,In_1287);
or U439 (N_439,In_940,In_1603);
nand U440 (N_440,In_1018,In_1792);
nand U441 (N_441,In_1849,In_2449);
or U442 (N_442,In_2439,In_10);
and U443 (N_443,In_1106,In_2172);
nand U444 (N_444,In_2422,In_2142);
or U445 (N_445,In_1881,In_1980);
and U446 (N_446,In_1601,In_296);
and U447 (N_447,In_311,In_403);
nand U448 (N_448,In_1991,In_1144);
or U449 (N_449,In_2403,In_2347);
or U450 (N_450,In_800,In_1059);
and U451 (N_451,In_2161,In_555);
xnor U452 (N_452,In_1664,In_68);
nand U453 (N_453,In_146,In_2100);
nor U454 (N_454,In_2330,In_623);
xor U455 (N_455,In_1630,In_153);
nand U456 (N_456,In_1782,In_2204);
or U457 (N_457,In_236,In_334);
or U458 (N_458,In_812,In_177);
or U459 (N_459,In_267,In_50);
nand U460 (N_460,In_143,In_983);
nand U461 (N_461,In_579,In_2190);
or U462 (N_462,In_1632,In_2121);
nor U463 (N_463,In_1743,In_180);
xor U464 (N_464,In_2428,In_1123);
and U465 (N_465,In_2017,In_1921);
or U466 (N_466,In_282,In_1851);
xnor U467 (N_467,In_358,In_982);
and U468 (N_468,In_956,In_538);
nand U469 (N_469,In_1252,In_1551);
and U470 (N_470,In_254,In_513);
nand U471 (N_471,In_560,In_104);
or U472 (N_472,In_1282,In_1771);
and U473 (N_473,In_658,In_631);
nor U474 (N_474,In_2388,In_1169);
nand U475 (N_475,In_1118,In_172);
xor U476 (N_476,In_1994,In_558);
or U477 (N_477,In_761,In_1075);
or U478 (N_478,In_2213,In_1338);
nor U479 (N_479,In_1817,In_531);
nor U480 (N_480,In_2458,In_1280);
nand U481 (N_481,In_284,In_2192);
xnor U482 (N_482,In_1121,In_948);
xnor U483 (N_483,In_2391,In_2344);
nor U484 (N_484,In_1246,In_1518);
nor U485 (N_485,In_1349,In_35);
nor U486 (N_486,In_1027,In_373);
or U487 (N_487,In_421,In_1880);
nor U488 (N_488,In_2046,In_818);
nand U489 (N_489,In_327,In_2136);
or U490 (N_490,In_1415,In_930);
or U491 (N_491,In_509,In_2470);
nor U492 (N_492,In_1492,In_2151);
nand U493 (N_493,In_1350,In_1803);
or U494 (N_494,In_1138,In_1592);
or U495 (N_495,In_1014,In_1793);
nand U496 (N_496,In_1663,In_257);
nand U497 (N_497,In_13,In_1556);
and U498 (N_498,In_1701,In_375);
xnor U499 (N_499,In_874,In_733);
or U500 (N_500,In_1939,In_1445);
and U501 (N_501,In_1547,In_1227);
nor U502 (N_502,In_483,In_1768);
nand U503 (N_503,In_984,In_456);
and U504 (N_504,In_1353,In_2401);
and U505 (N_505,In_1336,In_2423);
nor U506 (N_506,In_2239,In_1076);
and U507 (N_507,In_1467,In_453);
xnor U508 (N_508,In_1651,In_1647);
or U509 (N_509,In_2104,In_237);
nand U510 (N_510,In_649,In_719);
xnor U511 (N_511,In_2339,In_313);
nor U512 (N_512,In_2447,In_1166);
or U513 (N_513,In_1844,In_224);
xor U514 (N_514,In_2302,In_324);
xor U515 (N_515,In_645,In_1104);
nand U516 (N_516,In_838,In_1368);
and U517 (N_517,In_627,In_1143);
nor U518 (N_518,In_2277,In_2164);
or U519 (N_519,In_659,In_2200);
xor U520 (N_520,In_1170,In_2202);
or U521 (N_521,In_436,In_2288);
xnor U522 (N_522,In_890,In_1653);
nand U523 (N_523,In_2182,In_328);
xnor U524 (N_524,In_1047,In_474);
xnor U525 (N_525,In_1680,In_2462);
and U526 (N_526,In_2227,In_1514);
xor U527 (N_527,In_2198,In_1965);
xor U528 (N_528,In_2443,In_801);
or U529 (N_529,In_1136,In_2032);
xnor U530 (N_530,In_1927,In_2489);
xnor U531 (N_531,In_2351,In_1369);
or U532 (N_532,In_1251,In_196);
nand U533 (N_533,In_1593,In_2300);
nand U534 (N_534,In_1504,In_2498);
nor U535 (N_535,In_976,In_1553);
xnor U536 (N_536,In_861,In_1159);
or U537 (N_537,In_434,In_1738);
nor U538 (N_538,In_2186,In_580);
nand U539 (N_539,In_2233,In_1640);
or U540 (N_540,In_1045,In_989);
nand U541 (N_541,In_798,In_1748);
or U542 (N_542,In_1846,In_2362);
nand U543 (N_543,In_12,In_1679);
or U544 (N_544,In_1833,In_629);
nor U545 (N_545,In_2209,In_639);
or U546 (N_546,In_1233,In_1013);
xnor U547 (N_547,In_1392,In_729);
nand U548 (N_548,In_111,In_94);
xor U549 (N_549,In_1989,In_489);
nor U550 (N_550,In_1244,In_276);
nor U551 (N_551,In_1775,In_2466);
xnor U552 (N_552,In_2134,In_612);
nor U553 (N_553,In_2188,In_2263);
nand U554 (N_554,In_1274,In_526);
and U555 (N_555,In_2358,In_496);
nor U556 (N_556,In_986,In_1785);
or U557 (N_557,In_315,In_2467);
and U558 (N_558,In_241,In_2099);
nor U559 (N_559,In_2062,In_1435);
or U560 (N_560,In_1773,In_2379);
nand U561 (N_561,In_2370,In_1674);
xnor U562 (N_562,In_2138,In_1137);
xor U563 (N_563,In_1240,In_1261);
and U564 (N_564,In_637,In_2079);
nand U565 (N_565,In_524,In_317);
and U566 (N_566,In_1189,In_301);
xor U567 (N_567,In_2149,In_1669);
nor U568 (N_568,In_721,In_1790);
and U569 (N_569,In_62,In_1268);
and U570 (N_570,In_1946,In_2037);
nand U571 (N_571,In_2076,In_362);
nor U572 (N_572,In_619,In_47);
xnor U573 (N_573,In_1695,In_2157);
and U574 (N_574,In_1029,In_752);
nand U575 (N_575,In_632,In_181);
xnor U576 (N_576,In_2354,In_2077);
nor U577 (N_577,In_1077,In_2080);
nand U578 (N_578,In_1486,In_824);
nand U579 (N_579,In_1667,In_630);
nand U580 (N_580,In_599,In_933);
nand U581 (N_581,In_2010,In_125);
nor U582 (N_582,In_769,In_1202);
and U583 (N_583,In_2259,In_1883);
nand U584 (N_584,In_1211,In_770);
nand U585 (N_585,In_624,In_1940);
xor U586 (N_586,In_1520,In_405);
xor U587 (N_587,In_2420,In_1041);
or U588 (N_588,In_951,In_2181);
and U589 (N_589,In_335,In_1098);
and U590 (N_590,In_1291,In_1919);
nand U591 (N_591,In_775,In_16);
xnor U592 (N_592,In_700,In_1300);
nor U593 (N_593,In_1333,In_1095);
xnor U594 (N_594,In_2043,In_1506);
xnor U595 (N_595,In_2469,In_522);
nor U596 (N_596,In_1635,In_2267);
nand U597 (N_597,In_1191,In_437);
or U598 (N_598,In_2475,In_1412);
and U599 (N_599,In_903,In_746);
and U600 (N_600,In_295,In_347);
nand U601 (N_601,In_1512,In_731);
nand U602 (N_602,In_2110,In_1131);
and U603 (N_603,In_2169,In_2063);
and U604 (N_604,In_428,In_834);
nor U605 (N_605,In_145,In_1741);
xnor U606 (N_606,In_201,In_576);
nand U607 (N_607,In_285,In_1829);
xor U608 (N_608,In_1888,In_1398);
or U609 (N_609,In_906,In_202);
and U610 (N_610,In_291,In_119);
or U611 (N_611,In_914,In_735);
or U612 (N_612,In_191,In_447);
xnor U613 (N_613,In_2380,In_1293);
nor U614 (N_614,In_671,In_2095);
and U615 (N_615,In_1042,In_1308);
nand U616 (N_616,In_398,In_376);
nand U617 (N_617,In_1661,In_2473);
nor U618 (N_618,In_973,In_1147);
nor U619 (N_619,In_2321,In_1563);
or U620 (N_620,In_1842,In_275);
and U621 (N_621,In_1444,In_1087);
nand U622 (N_622,In_2424,In_306);
nor U623 (N_623,In_1272,In_1345);
nor U624 (N_624,In_2228,In_2214);
xnor U625 (N_625,In_1200,In_239);
and U626 (N_626,In_51,In_1356);
or U627 (N_627,In_2312,In_876);
nor U628 (N_628,In_459,In_2445);
and U629 (N_629,In_2368,In_2171);
and U630 (N_630,In_2044,In_2152);
or U631 (N_631,In_1243,In_1864);
nor U632 (N_632,In_1068,In_1133);
xor U633 (N_633,In_1937,In_1933);
or U634 (N_634,In_803,In_240);
or U635 (N_635,In_2226,In_2165);
or U636 (N_636,In_1508,In_441);
xor U637 (N_637,In_2026,In_1408);
and U638 (N_638,In_1489,In_2206);
nor U639 (N_639,In_2025,In_1784);
nand U640 (N_640,In_2327,In_960);
nor U641 (N_641,In_1951,In_1565);
nor U642 (N_642,In_680,In_1966);
or U643 (N_643,In_310,In_1340);
and U644 (N_644,In_945,In_1961);
nor U645 (N_645,In_1393,In_1830);
and U646 (N_646,In_1865,In_504);
or U647 (N_647,In_1367,In_192);
xor U648 (N_648,In_370,In_1752);
or U649 (N_649,In_862,In_1377);
nor U650 (N_650,In_2015,In_931);
xnor U651 (N_651,In_1823,In_2090);
xor U652 (N_652,In_1457,In_1208);
xnor U653 (N_653,In_1779,In_1885);
nor U654 (N_654,In_724,In_147);
or U655 (N_655,In_1000,In_767);
and U656 (N_656,In_420,In_875);
or U657 (N_657,In_2497,In_24);
nor U658 (N_658,In_1776,In_451);
nand U659 (N_659,In_1399,In_127);
and U660 (N_660,In_1053,In_1526);
or U661 (N_661,In_2251,In_479);
xnor U662 (N_662,In_1320,In_1071);
xor U663 (N_663,In_1530,In_372);
and U664 (N_664,In_889,In_461);
or U665 (N_665,In_2257,In_1932);
or U666 (N_666,In_1225,In_1501);
nand U667 (N_667,In_1613,In_1998);
and U668 (N_668,In_2258,In_316);
nor U669 (N_669,In_2317,In_1060);
and U670 (N_670,In_654,In_363);
and U671 (N_671,In_638,In_1030);
nor U672 (N_672,In_991,In_675);
and U673 (N_673,In_705,In_1573);
xor U674 (N_674,In_2336,In_48);
nor U675 (N_675,In_668,In_2335);
and U676 (N_676,In_2120,In_971);
nor U677 (N_677,In_825,In_57);
and U678 (N_678,In_776,In_314);
or U679 (N_679,In_568,In_833);
xor U680 (N_680,In_337,In_238);
or U681 (N_681,In_1942,In_939);
nand U682 (N_682,In_2262,In_1007);
nand U683 (N_683,In_2408,In_212);
xor U684 (N_684,In_1304,In_1177);
or U685 (N_685,In_1922,In_1767);
nand U686 (N_686,In_2355,In_1351);
nor U687 (N_687,In_1594,In_965);
nand U688 (N_688,In_89,In_2128);
nand U689 (N_689,In_1571,In_2476);
nor U690 (N_690,In_412,In_1870);
nor U691 (N_691,In_2112,In_1182);
xnor U692 (N_692,In_2299,In_2144);
and U693 (N_693,In_997,In_2325);
nand U694 (N_694,In_539,In_1751);
nor U695 (N_695,In_271,In_2212);
and U696 (N_696,In_1179,In_20);
nand U697 (N_697,In_1207,In_872);
xor U698 (N_698,In_2091,In_1455);
xor U699 (N_699,In_1934,In_1090);
nand U700 (N_700,In_1992,In_2272);
or U701 (N_701,In_2040,In_1026);
and U702 (N_702,In_90,In_589);
or U703 (N_703,In_1612,In_2174);
nor U704 (N_704,In_1597,In_1150);
or U705 (N_705,In_228,In_463);
nor U706 (N_706,In_1801,In_2116);
nand U707 (N_707,In_946,In_287);
and U708 (N_708,In_1491,In_926);
and U709 (N_709,In_466,In_607);
and U710 (N_710,In_1128,In_886);
nor U711 (N_711,In_1040,In_1555);
nor U712 (N_712,In_1626,In_2024);
or U713 (N_713,In_280,In_554);
xor U714 (N_714,In_1914,In_852);
xor U715 (N_715,In_484,In_488);
nor U716 (N_716,In_1798,In_304);
or U717 (N_717,In_1034,In_1427);
nor U718 (N_718,In_1477,In_1470);
or U719 (N_719,In_1673,In_622);
nor U720 (N_720,In_2373,In_2180);
nor U721 (N_721,In_1715,In_216);
nor U722 (N_722,In_1083,In_1100);
xnor U723 (N_723,In_2281,In_1523);
nand U724 (N_724,In_1473,In_1190);
and U725 (N_725,In_61,In_2308);
nand U726 (N_726,In_329,In_1378);
or U727 (N_727,In_30,In_964);
xor U728 (N_728,In_1510,In_2028);
nand U729 (N_729,In_551,In_2320);
or U730 (N_730,In_346,In_468);
xnor U731 (N_731,In_2394,In_2241);
nand U732 (N_732,In_1815,In_1314);
nor U733 (N_733,In_2187,In_1655);
and U734 (N_734,In_1448,In_1475);
or U735 (N_735,In_492,In_1769);
nand U736 (N_736,In_371,In_2294);
xor U737 (N_737,In_1139,In_2061);
nand U738 (N_738,In_1382,In_1428);
xor U739 (N_739,In_934,In_708);
and U740 (N_740,In_2417,In_919);
xnor U741 (N_741,In_1484,In_1827);
xnor U742 (N_742,In_1228,In_935);
xnor U743 (N_743,In_184,In_2008);
and U744 (N_744,In_1660,In_2493);
xnor U745 (N_745,In_2436,In_2060);
nor U746 (N_746,In_272,In_1599);
nand U747 (N_747,In_2143,In_1564);
nor U748 (N_748,In_2133,In_76);
xor U749 (N_749,In_936,In_1);
nand U750 (N_750,In_1590,In_2484);
or U751 (N_751,In_1380,In_2066);
nor U752 (N_752,In_1623,In_550);
nand U753 (N_753,In_2283,In_1727);
or U754 (N_754,In_1607,In_500);
nand U755 (N_755,In_667,In_1953);
nor U756 (N_756,In_1936,In_1848);
xnor U757 (N_757,In_1086,In_1195);
or U758 (N_758,In_1360,In_1778);
xnor U759 (N_759,In_1297,In_330);
xor U760 (N_760,In_1414,In_411);
and U761 (N_761,In_1028,In_445);
or U762 (N_762,In_219,In_1290);
nand U763 (N_763,In_1346,In_1051);
or U764 (N_764,In_502,In_796);
xor U765 (N_765,In_2405,In_1960);
nand U766 (N_766,In_32,In_683);
xnor U767 (N_767,In_943,In_1430);
xor U768 (N_768,In_396,In_844);
or U769 (N_769,In_1887,In_356);
xnor U770 (N_770,In_1325,In_2078);
or U771 (N_771,In_2069,In_1996);
or U772 (N_772,In_1985,In_1461);
nand U773 (N_773,In_963,In_1341);
nand U774 (N_774,In_897,In_2156);
nand U775 (N_775,In_918,In_777);
or U776 (N_776,In_1120,In_402);
nor U777 (N_777,In_136,In_618);
or U778 (N_778,In_1276,In_587);
or U779 (N_779,In_749,In_2399);
nand U780 (N_780,In_578,In_1391);
xor U781 (N_781,In_663,In_532);
xnor U782 (N_782,In_1816,In_2363);
nand U783 (N_783,In_820,In_961);
xnor U784 (N_784,In_1808,In_1604);
xnor U785 (N_785,In_894,In_1908);
and U786 (N_786,In_1298,In_1797);
xnor U787 (N_787,In_888,In_303);
or U788 (N_788,In_134,In_151);
xor U789 (N_789,In_2145,In_1273);
or U790 (N_790,In_149,In_2123);
and U791 (N_791,In_1215,In_1091);
nor U792 (N_792,In_743,In_2326);
nand U793 (N_793,In_1152,In_815);
or U794 (N_794,In_1373,In_2240);
or U795 (N_795,In_2072,In_883);
or U796 (N_796,In_1974,In_2285);
nor U797 (N_797,In_18,In_1731);
or U798 (N_798,In_1910,In_52);
or U799 (N_799,In_895,In_141);
nand U800 (N_800,In_1178,In_2369);
and U801 (N_801,In_514,In_848);
and U802 (N_802,In_1911,In_621);
xor U803 (N_803,In_1756,In_2279);
nand U804 (N_804,In_1519,In_2318);
and U805 (N_805,In_1181,In_2252);
nand U806 (N_806,In_230,In_507);
or U807 (N_807,In_2244,In_2042);
and U808 (N_808,In_1721,In_1852);
nand U809 (N_809,In_1528,In_2045);
or U810 (N_810,In_1713,In_1585);
or U811 (N_811,In_221,In_124);
and U812 (N_812,In_1591,In_1361);
nor U813 (N_813,In_1794,In_266);
nor U814 (N_814,In_1025,In_1765);
or U815 (N_815,In_1567,In_2440);
or U816 (N_816,In_161,In_2097);
and U817 (N_817,In_1238,In_2352);
and U818 (N_818,In_2333,In_2002);
or U819 (N_819,In_458,In_681);
or U820 (N_820,In_1662,In_2390);
or U821 (N_821,In_1303,In_885);
nand U822 (N_822,In_1460,In_1248);
and U823 (N_823,In_620,In_1968);
xor U824 (N_824,In_1586,In_1737);
xnor U825 (N_825,In_1843,In_2404);
xor U826 (N_826,In_37,In_2056);
or U827 (N_827,In_1359,In_431);
or U828 (N_828,In_1511,In_2463);
xnor U829 (N_829,In_2059,In_839);
nand U830 (N_830,In_2222,In_2455);
xnor U831 (N_831,In_1410,In_2125);
xor U832 (N_832,In_336,In_867);
nor U833 (N_833,In_2003,In_65);
nand U834 (N_834,In_1950,In_1878);
nand U835 (N_835,In_106,In_2378);
xnor U836 (N_836,In_571,In_2381);
and U837 (N_837,In_1557,In_2341);
xor U838 (N_838,In_836,In_2323);
and U839 (N_839,In_1431,In_1529);
xor U840 (N_840,In_2155,In_2400);
xnor U841 (N_841,In_544,In_168);
nand U842 (N_842,In_277,In_1686);
nand U843 (N_843,In_1394,In_1146);
or U844 (N_844,In_1082,In_259);
nor U845 (N_845,In_1124,In_2094);
or U846 (N_846,In_2211,In_1033);
nand U847 (N_847,In_1956,In_1666);
and U848 (N_848,In_1978,In_548);
nand U849 (N_849,In_84,In_207);
or U850 (N_850,In_679,In_340);
nor U851 (N_851,In_651,In_806);
nand U852 (N_852,In_1463,In_1212);
nand U853 (N_853,In_1521,In_615);
nor U854 (N_854,In_2225,In_1468);
xnor U855 (N_855,In_1648,In_333);
xnor U856 (N_856,In_899,In_1452);
nand U857 (N_857,In_1069,In_2105);
xor U858 (N_858,In_846,In_1583);
xor U859 (N_859,In_736,In_1725);
and U860 (N_860,In_1366,In_2195);
nand U861 (N_861,In_1476,In_56);
nor U862 (N_862,In_1406,In_42);
and U863 (N_863,In_782,In_525);
or U864 (N_864,In_233,In_209);
and U865 (N_865,In_392,In_203);
or U866 (N_866,In_1114,In_704);
or U867 (N_867,In_1107,In_692);
or U868 (N_868,In_1421,In_2014);
nand U869 (N_869,In_1918,In_955);
nand U870 (N_870,In_1498,In_785);
nand U871 (N_871,In_1689,In_1897);
nand U872 (N_872,In_395,In_2102);
and U873 (N_873,In_59,In_2393);
nor U874 (N_874,In_116,In_1621);
nor U875 (N_875,In_2459,In_323);
xor U876 (N_876,In_534,In_1631);
nand U877 (N_877,In_80,In_953);
nand U878 (N_878,In_1206,In_2353);
or U879 (N_879,In_592,In_1250);
nor U880 (N_880,In_636,In_521);
nor U881 (N_881,In_1834,In_657);
or U882 (N_882,In_2071,In_2185);
or U883 (N_883,In_1628,In_998);
xor U884 (N_884,In_760,In_1471);
nor U885 (N_885,In_318,In_2193);
and U886 (N_886,In_2332,In_1912);
xor U887 (N_887,In_958,In_2051);
or U888 (N_888,In_1205,In_2093);
nor U889 (N_889,In_197,In_2431);
nor U890 (N_890,In_1437,In_1001);
or U891 (N_891,In_2305,In_941);
nand U892 (N_892,In_1541,In_425);
nor U893 (N_893,In_129,In_2488);
nand U894 (N_894,In_368,In_1772);
or U895 (N_895,In_858,In_43);
xor U896 (N_896,In_849,In_2115);
nand U897 (N_897,In_2284,In_1958);
or U898 (N_898,In_985,In_1548);
or U899 (N_899,In_2421,In_1456);
nand U900 (N_900,In_491,In_283);
and U901 (N_901,In_416,In_613);
xor U902 (N_902,In_1056,In_64);
nand U903 (N_903,In_384,In_1723);
and U904 (N_904,In_243,In_1969);
nand U905 (N_905,In_2306,In_1422);
and U906 (N_906,In_97,In_817);
xnor U907 (N_907,In_2101,In_2215);
nor U908 (N_908,In_2359,In_1442);
or U909 (N_909,In_1440,In_189);
or U910 (N_910,In_902,In_1183);
nand U911 (N_911,In_1774,In_2054);
nor U912 (N_912,In_429,In_1964);
and U913 (N_913,In_563,In_1868);
nor U914 (N_914,In_1983,In_171);
xnor U915 (N_915,In_231,In_901);
xnor U916 (N_916,In_2201,In_15);
nor U917 (N_917,In_217,In_1973);
nor U918 (N_918,In_851,In_866);
or U919 (N_919,In_718,In_567);
xnor U920 (N_920,In_388,In_2292);
xnor U921 (N_921,In_2150,In_771);
nand U922 (N_922,In_1711,In_175);
and U923 (N_923,In_1466,In_570);
nand U924 (N_924,In_1947,In_2194);
or U925 (N_925,In_2085,In_2230);
xnor U926 (N_926,In_790,In_1677);
nor U927 (N_927,In_987,In_430);
nor U928 (N_928,In_1754,In_947);
xnor U929 (N_929,In_788,In_1926);
or U930 (N_930,In_1649,In_829);
nor U931 (N_931,In_95,In_1317);
nor U932 (N_932,In_1760,In_1102);
or U933 (N_933,In_1004,In_1633);
xor U934 (N_934,In_407,In_2441);
nor U935 (N_935,In_1289,In_1294);
xnor U936 (N_936,In_878,In_497);
and U937 (N_937,In_1464,In_574);
or U938 (N_938,In_1970,In_1231);
or U939 (N_939,In_959,In_1219);
or U940 (N_940,In_1283,In_1344);
or U941 (N_941,In_909,In_1048);
nand U942 (N_942,In_1335,In_734);
nand U943 (N_943,In_1799,In_1423);
or U944 (N_944,In_1235,In_720);
and U945 (N_945,In_1977,In_1092);
nor U946 (N_946,In_166,In_1595);
nand U947 (N_947,In_1474,In_588);
xor U948 (N_948,In_1096,In_826);
nor U949 (N_949,In_344,In_351);
nand U950 (N_950,In_93,In_1015);
or U951 (N_951,In_512,In_204);
nand U952 (N_952,In_2176,In_1074);
and U953 (N_953,In_898,In_881);
or U954 (N_954,In_499,In_248);
xor U955 (N_955,In_750,In_2304);
and U956 (N_956,In_1576,In_2412);
nor U957 (N_957,In_691,In_2345);
nand U958 (N_958,In_2167,In_1709);
nor U959 (N_959,In_1681,In_1196);
and U960 (N_960,In_1201,In_404);
and U961 (N_961,In_1054,In_2356);
xor U962 (N_962,In_1891,In_214);
or U963 (N_963,In_608,In_2052);
and U964 (N_964,In_2454,In_1584);
and U965 (N_965,In_674,In_120);
or U966 (N_966,In_927,In_2168);
xor U967 (N_967,In_1629,In_2337);
nor U968 (N_968,In_2126,In_444);
or U969 (N_969,In_2307,In_1899);
xor U970 (N_970,In_2154,In_1194);
nor U971 (N_971,In_1610,In_2005);
nor U972 (N_972,In_1698,In_1229);
and U973 (N_973,In_1841,In_1763);
nand U974 (N_974,In_1330,In_714);
nand U975 (N_975,In_247,In_2053);
nand U976 (N_976,In_2278,In_2082);
and U977 (N_977,In_896,In_1157);
and U978 (N_978,In_1134,In_1952);
and U979 (N_979,In_1324,In_67);
nor U980 (N_980,In_2224,In_2006);
nor U981 (N_981,In_1062,In_1449);
nand U982 (N_982,In_516,In_2483);
nand U983 (N_983,In_293,In_2255);
xnor U984 (N_984,In_831,In_86);
nor U985 (N_985,In_503,In_364);
and U986 (N_986,In_1869,In_1882);
or U987 (N_987,In_1224,In_341);
nor U988 (N_988,In_1886,In_937);
xnor U989 (N_989,In_1097,In_1544);
nand U990 (N_990,In_1499,In_355);
nand U991 (N_991,In_628,In_44);
or U992 (N_992,In_2084,In_1309);
nand U993 (N_993,In_2415,In_1269);
or U994 (N_994,In_1636,In_1859);
nand U995 (N_995,In_2395,In_1513);
nor U996 (N_996,In_357,In_1645);
xnor U997 (N_997,In_1321,In_2434);
and U998 (N_998,In_1411,In_1967);
nand U999 (N_999,In_9,In_255);
or U1000 (N_1000,In_1357,In_2196);
xnor U1001 (N_1001,In_1753,In_2409);
and U1002 (N_1002,In_1383,In_1223);
nor U1003 (N_1003,In_823,In_969);
and U1004 (N_1004,In_904,In_1750);
nand U1005 (N_1005,In_1085,In_2311);
xnor U1006 (N_1006,In_1944,In_292);
and U1007 (N_1007,In_1516,In_1559);
nand U1008 (N_1008,In_1532,In_1469);
and U1009 (N_1009,In_401,In_462);
nand U1010 (N_1010,In_1316,In_1755);
xor U1011 (N_1011,In_1332,In_703);
and U1012 (N_1012,In_1203,In_1867);
nand U1013 (N_1013,In_414,In_1840);
nor U1014 (N_1014,In_1884,In_1158);
nand U1015 (N_1015,In_1055,In_1527);
and U1016 (N_1016,In_810,In_2438);
nand U1017 (N_1017,In_1691,In_730);
or U1018 (N_1018,In_1277,In_696);
and U1019 (N_1019,In_701,In_229);
or U1020 (N_1020,In_992,In_2287);
nor U1021 (N_1021,In_2114,In_2457);
xnor U1022 (N_1022,In_792,In_2376);
xor U1023 (N_1023,In_647,In_2250);
nor U1024 (N_1024,In_981,In_2437);
or U1025 (N_1025,In_1125,In_655);
nor U1026 (N_1026,In_556,In_455);
xor U1027 (N_1027,In_510,In_170);
xnor U1028 (N_1028,In_75,In_778);
nor U1029 (N_1029,In_440,In_1306);
nor U1030 (N_1030,In_1729,In_893);
xor U1031 (N_1031,In_1863,In_176);
or U1032 (N_1032,In_2159,In_325);
nor U1033 (N_1033,In_1814,In_1835);
or U1034 (N_1034,In_1284,In_2207);
or U1035 (N_1035,In_1854,In_361);
xnor U1036 (N_1036,In_49,In_1370);
nor U1037 (N_1037,In_707,In_389);
nand U1038 (N_1038,In_572,In_1446);
nand U1039 (N_1039,In_1021,In_169);
xnor U1040 (N_1040,In_2499,In_518);
nor U1041 (N_1041,In_1871,In_1596);
or U1042 (N_1042,In_105,In_1358);
and U1043 (N_1043,In_1611,In_495);
nor U1044 (N_1044,In_685,In_809);
xnor U1045 (N_1045,In_662,In_625);
nor U1046 (N_1046,In_1343,In_1035);
and U1047 (N_1047,In_1855,In_206);
and U1048 (N_1048,In_1008,In_1696);
and U1049 (N_1049,In_1537,In_569);
xor U1050 (N_1050,In_2450,In_1757);
xor U1051 (N_1051,In_1285,In_598);
nand U1052 (N_1052,In_1315,In_1692);
or U1053 (N_1053,In_2485,In_1976);
xor U1054 (N_1054,In_1161,In_1192);
xnor U1055 (N_1055,In_226,In_174);
or U1056 (N_1056,In_232,In_2256);
xor U1057 (N_1057,In_1907,In_972);
and U1058 (N_1058,In_1032,In_1507);
nand U1059 (N_1059,In_1874,In_299);
and U1060 (N_1060,In_117,In_1646);
and U1061 (N_1061,In_2140,In_273);
xor U1062 (N_1062,In_944,In_1616);
xnor U1063 (N_1063,In_923,In_446);
nor U1064 (N_1064,In_1702,In_1352);
nor U1065 (N_1065,In_925,In_460);
or U1066 (N_1066,In_477,In_2173);
or U1067 (N_1067,In_1543,In_2074);
and U1068 (N_1068,In_476,In_2245);
xor U1069 (N_1069,In_2419,In_2366);
xnor U1070 (N_1070,In_1503,In_1443);
nor U1071 (N_1071,In_154,In_1160);
or U1072 (N_1072,In_2486,In_2384);
nor U1073 (N_1073,In_1301,In_1226);
nor U1074 (N_1074,In_715,In_1295);
or U1075 (N_1075,In_1800,In_2147);
nor U1076 (N_1076,In_1730,In_2106);
nor U1077 (N_1077,In_928,In_1533);
or U1078 (N_1078,In_1894,In_186);
nand U1079 (N_1079,In_1329,In_1904);
and U1080 (N_1080,In_1453,In_1184);
or U1081 (N_1081,In_1657,In_29);
or U1082 (N_1082,In_2387,In_1101);
and U1083 (N_1083,In_932,In_85);
and U1084 (N_1084,In_1581,In_242);
nor U1085 (N_1085,In_46,In_523);
nand U1086 (N_1086,In_2418,In_2210);
and U1087 (N_1087,In_2229,In_911);
and U1088 (N_1088,In_1433,In_1948);
and U1089 (N_1089,In_1187,In_1480);
or U1090 (N_1090,In_1386,In_2435);
or U1091 (N_1091,In_1465,In_1744);
xor U1092 (N_1092,In_54,In_1318);
and U1093 (N_1093,In_135,In_977);
or U1094 (N_1094,In_1164,In_779);
xnor U1095 (N_1095,In_1117,In_2001);
or U1096 (N_1096,In_1913,In_2011);
nor U1097 (N_1097,In_1180,In_2427);
or U1098 (N_1098,In_1245,In_1853);
nand U1099 (N_1099,In_1093,In_1587);
and U1100 (N_1100,In_2119,In_1637);
or U1101 (N_1101,In_39,In_942);
nor U1102 (N_1102,In_1310,In_830);
and U1103 (N_1103,In_845,In_2271);
or U1104 (N_1104,In_1221,In_905);
nand U1105 (N_1105,In_814,In_1720);
nand U1106 (N_1106,In_1172,In_1818);
nor U1107 (N_1107,In_2170,In_1409);
and U1108 (N_1108,In_2411,In_1642);
and U1109 (N_1109,In_1746,In_2163);
nor U1110 (N_1110,In_397,In_73);
nor U1111 (N_1111,In_1739,In_2334);
and U1112 (N_1112,In_2127,In_1525);
nand U1113 (N_1113,In_1896,In_338);
or U1114 (N_1114,In_1323,In_96);
and U1115 (N_1115,In_2141,In_118);
nor U1116 (N_1116,In_593,In_1327);
nand U1117 (N_1117,In_38,In_1822);
and U1118 (N_1118,In_1232,In_1938);
xnor U1119 (N_1119,In_1736,In_1517);
nand U1120 (N_1120,In_2039,In_2276);
or U1121 (N_1121,In_1676,In_689);
or U1122 (N_1122,In_91,In_31);
nand U1123 (N_1123,In_2477,In_1945);
nor U1124 (N_1124,In_1337,In_716);
or U1125 (N_1125,In_71,In_252);
nand U1126 (N_1126,In_246,In_2338);
nor U1127 (N_1127,In_1388,In_2426);
nor U1128 (N_1128,In_575,In_710);
and U1129 (N_1129,In_808,In_113);
nand U1130 (N_1130,In_832,In_1023);
nand U1131 (N_1131,In_1652,In_1839);
nand U1132 (N_1132,In_1043,In_235);
nor U1133 (N_1133,In_1831,In_1734);
and U1134 (N_1134,In_962,In_915);
nand U1135 (N_1135,In_1758,In_1312);
nand U1136 (N_1136,In_2237,In_2166);
and U1137 (N_1137,In_1073,In_2496);
xor U1138 (N_1138,In_596,In_1024);
nand U1139 (N_1139,In_1039,In_1995);
and U1140 (N_1140,In_1837,In_633);
nand U1141 (N_1141,In_822,In_1264);
or U1142 (N_1142,In_1305,In_321);
or U1143 (N_1143,In_1665,In_688);
nand U1144 (N_1144,In_1331,In_1241);
and U1145 (N_1145,In_2153,In_766);
and U1146 (N_1146,In_725,In_1299);
or U1147 (N_1147,In_2291,In_1256);
or U1148 (N_1148,In_2372,In_1724);
nand U1149 (N_1149,In_473,In_486);
xnor U1150 (N_1150,In_1550,In_713);
xnor U1151 (N_1151,In_594,In_1010);
or U1152 (N_1152,In_163,In_21);
nand U1153 (N_1153,In_77,In_2382);
or U1154 (N_1154,In_470,In_2208);
nand U1155 (N_1155,In_1924,In_1906);
nand U1156 (N_1156,In_424,In_2444);
or U1157 (N_1157,In_891,In_1257);
nor U1158 (N_1158,In_393,In_2004);
xnor U1159 (N_1159,In_131,In_1148);
nand U1160 (N_1160,In_2328,In_165);
xnor U1161 (N_1161,In_2265,In_2018);
and U1162 (N_1162,In_1762,In_966);
xor U1163 (N_1163,In_366,In_1145);
or U1164 (N_1164,In_1997,In_128);
xnor U1165 (N_1165,In_1902,In_1070);
and U1166 (N_1166,In_1515,In_182);
nand U1167 (N_1167,In_1979,In_2397);
xor U1168 (N_1168,In_2414,In_160);
and U1169 (N_1169,In_2374,In_2038);
xnor U1170 (N_1170,In_804,In_1454);
nor U1171 (N_1171,In_1379,In_320);
or U1172 (N_1172,In_559,In_245);
and U1173 (N_1173,In_450,In_577);
or U1174 (N_1174,In_1639,In_2129);
or U1175 (N_1175,In_661,In_481);
nor U1176 (N_1176,In_1109,In_1981);
nor U1177 (N_1177,In_198,In_617);
nand U1178 (N_1178,In_157,In_1861);
or U1179 (N_1179,In_1796,In_2367);
xor U1180 (N_1180,In_1247,In_2089);
xor U1181 (N_1181,In_2402,In_2331);
nor U1182 (N_1182,In_297,In_1266);
xnor U1183 (N_1183,In_1860,In_664);
nand U1184 (N_1184,In_585,In_517);
nor U1185 (N_1185,In_864,In_1113);
nand U1186 (N_1186,In_1925,In_2309);
and U1187 (N_1187,In_1931,In_773);
nand U1188 (N_1188,In_1129,In_1668);
xor U1189 (N_1189,In_1566,In_913);
nor U1190 (N_1190,In_1490,In_2314);
nor U1191 (N_1191,In_646,In_2092);
or U1192 (N_1192,In_1425,In_1112);
nor U1193 (N_1193,In_419,In_873);
xnor U1194 (N_1194,In_1089,In_2303);
nor U1195 (N_1195,In_616,In_1879);
nand U1196 (N_1196,In_1993,In_1704);
and U1197 (N_1197,In_2471,In_879);
nor U1198 (N_1198,In_1046,In_1710);
or U1199 (N_1199,In_2235,In_1608);
nand U1200 (N_1200,In_2057,In_1115);
and U1201 (N_1201,In_1167,In_1987);
nand U1202 (N_1202,In_1819,In_467);
xnor U1203 (N_1203,In_747,In_1708);
nor U1204 (N_1204,In_1971,In_2290);
nor U1205 (N_1205,In_709,In_1127);
nor U1206 (N_1206,In_2301,In_540);
and U1207 (N_1207,In_1717,In_1057);
nand U1208 (N_1208,In_1110,In_386);
and U1209 (N_1209,In_439,In_1678);
nor U1210 (N_1210,In_573,In_2487);
xnor U1211 (N_1211,In_758,In_1413);
and U1212 (N_1212,In_827,In_2055);
or U1213 (N_1213,In_494,In_2298);
and U1214 (N_1214,In_994,In_183);
and U1215 (N_1215,In_1081,In_1975);
nand U1216 (N_1216,In_164,In_1385);
nor U1217 (N_1217,In_148,In_2377);
or U1218 (N_1218,In_138,In_2383);
xor U1219 (N_1219,In_1826,In_1828);
nand U1220 (N_1220,In_322,In_837);
xor U1221 (N_1221,In_365,In_1605);
or U1222 (N_1222,In_23,In_722);
xor U1223 (N_1223,In_2464,In_1850);
nand U1224 (N_1224,In_605,In_1847);
xor U1225 (N_1225,In_1216,In_1348);
or U1226 (N_1226,In_353,In_1560);
xor U1227 (N_1227,In_910,In_1487);
xor U1228 (N_1228,In_672,In_1634);
nor U1229 (N_1229,In_2007,In_1171);
and U1230 (N_1230,In_653,In_1220);
and U1231 (N_1231,In_409,In_1562);
or U1232 (N_1232,In_582,In_1761);
nor U1233 (N_1233,In_3,In_1929);
nor U1234 (N_1234,In_432,In_222);
xor U1235 (N_1235,In_7,In_19);
xor U1236 (N_1236,In_819,In_566);
or U1237 (N_1237,In_2000,In_343);
and U1238 (N_1238,In_2023,In_2465);
nor U1239 (N_1239,In_1162,In_1954);
nor U1240 (N_1240,In_1496,In_1395);
xnor U1241 (N_1241,In_385,In_2146);
or U1242 (N_1242,In_0,In_2137);
xor U1243 (N_1243,In_993,In_2430);
and U1244 (N_1244,In_921,In_1643);
and U1245 (N_1245,In_1806,In_33);
nand U1246 (N_1246,In_2340,In_265);
nand U1247 (N_1247,In_1614,In_757);
nor U1248 (N_1248,In_83,In_938);
xor U1249 (N_1249,In_2343,In_780);
xnor U1250 (N_1250,In_2477,In_2437);
and U1251 (N_1251,In_466,In_122);
or U1252 (N_1252,In_392,In_1008);
and U1253 (N_1253,In_623,In_876);
and U1254 (N_1254,In_246,In_1153);
xor U1255 (N_1255,In_1029,In_782);
and U1256 (N_1256,In_1898,In_2113);
or U1257 (N_1257,In_1982,In_231);
xor U1258 (N_1258,In_2395,In_805);
nor U1259 (N_1259,In_2482,In_5);
xnor U1260 (N_1260,In_1194,In_1952);
nor U1261 (N_1261,In_864,In_2454);
xor U1262 (N_1262,In_950,In_1348);
and U1263 (N_1263,In_1366,In_1807);
xnor U1264 (N_1264,In_1510,In_996);
and U1265 (N_1265,In_1310,In_1474);
or U1266 (N_1266,In_25,In_1295);
and U1267 (N_1267,In_515,In_194);
nand U1268 (N_1268,In_1562,In_939);
xor U1269 (N_1269,In_1086,In_1705);
or U1270 (N_1270,In_938,In_1113);
nand U1271 (N_1271,In_1482,In_407);
xnor U1272 (N_1272,In_49,In_1702);
xor U1273 (N_1273,In_1035,In_2049);
nor U1274 (N_1274,In_1749,In_2495);
nand U1275 (N_1275,In_1387,In_1686);
or U1276 (N_1276,In_952,In_197);
xnor U1277 (N_1277,In_2077,In_2445);
nor U1278 (N_1278,In_1636,In_2160);
xnor U1279 (N_1279,In_1249,In_1603);
and U1280 (N_1280,In_1309,In_367);
and U1281 (N_1281,In_755,In_537);
nand U1282 (N_1282,In_1022,In_1492);
xnor U1283 (N_1283,In_114,In_2404);
and U1284 (N_1284,In_716,In_2055);
nor U1285 (N_1285,In_1046,In_888);
and U1286 (N_1286,In_1073,In_1859);
nor U1287 (N_1287,In_2411,In_1014);
nand U1288 (N_1288,In_2076,In_1990);
or U1289 (N_1289,In_337,In_2279);
nor U1290 (N_1290,In_280,In_2053);
xnor U1291 (N_1291,In_416,In_585);
nor U1292 (N_1292,In_1360,In_983);
nor U1293 (N_1293,In_795,In_313);
or U1294 (N_1294,In_1299,In_2472);
nand U1295 (N_1295,In_2356,In_1031);
or U1296 (N_1296,In_2445,In_1497);
nand U1297 (N_1297,In_1129,In_219);
or U1298 (N_1298,In_521,In_116);
nor U1299 (N_1299,In_1175,In_856);
and U1300 (N_1300,In_930,In_647);
or U1301 (N_1301,In_1636,In_1118);
or U1302 (N_1302,In_1965,In_452);
or U1303 (N_1303,In_2190,In_2032);
nor U1304 (N_1304,In_1207,In_1353);
nor U1305 (N_1305,In_629,In_1388);
nor U1306 (N_1306,In_823,In_464);
nand U1307 (N_1307,In_176,In_1690);
or U1308 (N_1308,In_511,In_2293);
xor U1309 (N_1309,In_991,In_1906);
and U1310 (N_1310,In_823,In_1838);
nand U1311 (N_1311,In_1737,In_1101);
nand U1312 (N_1312,In_1364,In_847);
nand U1313 (N_1313,In_1118,In_2432);
or U1314 (N_1314,In_1456,In_1513);
xnor U1315 (N_1315,In_898,In_2049);
nor U1316 (N_1316,In_785,In_661);
and U1317 (N_1317,In_650,In_157);
or U1318 (N_1318,In_1810,In_1467);
nor U1319 (N_1319,In_1461,In_1554);
and U1320 (N_1320,In_2467,In_828);
xnor U1321 (N_1321,In_918,In_1437);
or U1322 (N_1322,In_1558,In_2339);
nand U1323 (N_1323,In_690,In_609);
nor U1324 (N_1324,In_1409,In_529);
and U1325 (N_1325,In_1864,In_1085);
nand U1326 (N_1326,In_1927,In_880);
xor U1327 (N_1327,In_1004,In_587);
or U1328 (N_1328,In_302,In_1723);
xor U1329 (N_1329,In_459,In_1052);
and U1330 (N_1330,In_120,In_1159);
or U1331 (N_1331,In_2439,In_229);
nand U1332 (N_1332,In_926,In_2479);
and U1333 (N_1333,In_1063,In_863);
nor U1334 (N_1334,In_2288,In_1215);
xor U1335 (N_1335,In_396,In_859);
nor U1336 (N_1336,In_1023,In_2038);
and U1337 (N_1337,In_873,In_2416);
nand U1338 (N_1338,In_2167,In_1475);
or U1339 (N_1339,In_2381,In_1183);
nor U1340 (N_1340,In_2031,In_2436);
nand U1341 (N_1341,In_1220,In_1072);
or U1342 (N_1342,In_1722,In_1187);
nand U1343 (N_1343,In_2029,In_869);
nor U1344 (N_1344,In_1712,In_758);
nand U1345 (N_1345,In_2310,In_1938);
and U1346 (N_1346,In_1730,In_524);
or U1347 (N_1347,In_1314,In_2374);
xnor U1348 (N_1348,In_1340,In_2156);
nand U1349 (N_1349,In_2,In_2099);
and U1350 (N_1350,In_434,In_1612);
or U1351 (N_1351,In_560,In_2221);
nor U1352 (N_1352,In_367,In_1620);
xor U1353 (N_1353,In_653,In_2195);
nor U1354 (N_1354,In_1129,In_176);
nor U1355 (N_1355,In_1362,In_1942);
xnor U1356 (N_1356,In_1704,In_1050);
nand U1357 (N_1357,In_1426,In_1552);
or U1358 (N_1358,In_1723,In_1930);
and U1359 (N_1359,In_883,In_957);
nor U1360 (N_1360,In_511,In_613);
or U1361 (N_1361,In_1047,In_1060);
xor U1362 (N_1362,In_847,In_1367);
nand U1363 (N_1363,In_1900,In_1702);
nand U1364 (N_1364,In_517,In_1495);
xor U1365 (N_1365,In_2103,In_2459);
xor U1366 (N_1366,In_1385,In_1781);
nand U1367 (N_1367,In_2411,In_1514);
or U1368 (N_1368,In_357,In_10);
or U1369 (N_1369,In_957,In_1370);
and U1370 (N_1370,In_760,In_1753);
or U1371 (N_1371,In_2237,In_831);
and U1372 (N_1372,In_2288,In_2253);
nor U1373 (N_1373,In_1092,In_1831);
or U1374 (N_1374,In_236,In_1816);
or U1375 (N_1375,In_480,In_2423);
or U1376 (N_1376,In_101,In_678);
or U1377 (N_1377,In_318,In_1611);
nand U1378 (N_1378,In_1238,In_702);
and U1379 (N_1379,In_888,In_2293);
nand U1380 (N_1380,In_2245,In_1185);
nor U1381 (N_1381,In_2103,In_842);
or U1382 (N_1382,In_1311,In_743);
nor U1383 (N_1383,In_809,In_349);
xnor U1384 (N_1384,In_1821,In_1795);
or U1385 (N_1385,In_1990,In_992);
xnor U1386 (N_1386,In_1277,In_4);
nand U1387 (N_1387,In_37,In_1852);
or U1388 (N_1388,In_1150,In_24);
nor U1389 (N_1389,In_2007,In_2271);
or U1390 (N_1390,In_1283,In_532);
nor U1391 (N_1391,In_1472,In_2039);
nor U1392 (N_1392,In_1937,In_1398);
and U1393 (N_1393,In_834,In_2121);
xnor U1394 (N_1394,In_1770,In_1283);
or U1395 (N_1395,In_936,In_653);
nand U1396 (N_1396,In_692,In_2199);
nand U1397 (N_1397,In_1672,In_1803);
and U1398 (N_1398,In_2472,In_900);
xnor U1399 (N_1399,In_760,In_2308);
and U1400 (N_1400,In_156,In_1904);
nand U1401 (N_1401,In_1618,In_485);
xor U1402 (N_1402,In_1027,In_595);
nand U1403 (N_1403,In_1328,In_1079);
xor U1404 (N_1404,In_635,In_1913);
and U1405 (N_1405,In_1056,In_957);
nand U1406 (N_1406,In_1838,In_1554);
and U1407 (N_1407,In_1808,In_2136);
nand U1408 (N_1408,In_181,In_1139);
and U1409 (N_1409,In_1756,In_93);
xnor U1410 (N_1410,In_1404,In_1691);
xnor U1411 (N_1411,In_1785,In_168);
or U1412 (N_1412,In_2441,In_560);
xor U1413 (N_1413,In_2376,In_1359);
or U1414 (N_1414,In_1774,In_2045);
nand U1415 (N_1415,In_1854,In_1771);
or U1416 (N_1416,In_818,In_1152);
nand U1417 (N_1417,In_2377,In_1286);
xnor U1418 (N_1418,In_1040,In_592);
and U1419 (N_1419,In_404,In_2160);
and U1420 (N_1420,In_1378,In_856);
nor U1421 (N_1421,In_1303,In_1319);
nand U1422 (N_1422,In_2035,In_826);
nor U1423 (N_1423,In_1360,In_1431);
xor U1424 (N_1424,In_941,In_703);
nor U1425 (N_1425,In_1878,In_2336);
xor U1426 (N_1426,In_48,In_1723);
xor U1427 (N_1427,In_98,In_820);
nor U1428 (N_1428,In_2079,In_1048);
and U1429 (N_1429,In_1702,In_2425);
nor U1430 (N_1430,In_1463,In_2065);
or U1431 (N_1431,In_830,In_925);
nor U1432 (N_1432,In_1576,In_1762);
or U1433 (N_1433,In_1649,In_420);
nand U1434 (N_1434,In_874,In_1966);
xor U1435 (N_1435,In_1138,In_1685);
or U1436 (N_1436,In_1795,In_581);
nor U1437 (N_1437,In_763,In_561);
xor U1438 (N_1438,In_1811,In_1009);
or U1439 (N_1439,In_1847,In_2491);
or U1440 (N_1440,In_181,In_1755);
nor U1441 (N_1441,In_1359,In_2021);
xnor U1442 (N_1442,In_835,In_1814);
or U1443 (N_1443,In_831,In_1569);
nand U1444 (N_1444,In_993,In_1427);
xor U1445 (N_1445,In_1523,In_579);
or U1446 (N_1446,In_389,In_1390);
or U1447 (N_1447,In_2381,In_2044);
and U1448 (N_1448,In_566,In_1104);
nand U1449 (N_1449,In_473,In_2024);
and U1450 (N_1450,In_1933,In_1369);
and U1451 (N_1451,In_890,In_208);
or U1452 (N_1452,In_354,In_526);
or U1453 (N_1453,In_635,In_2227);
nor U1454 (N_1454,In_2090,In_1707);
or U1455 (N_1455,In_900,In_2313);
and U1456 (N_1456,In_2108,In_1727);
nand U1457 (N_1457,In_1445,In_2396);
xnor U1458 (N_1458,In_1155,In_396);
and U1459 (N_1459,In_225,In_86);
and U1460 (N_1460,In_1721,In_2149);
nor U1461 (N_1461,In_2282,In_1422);
xor U1462 (N_1462,In_868,In_2049);
nand U1463 (N_1463,In_166,In_1856);
and U1464 (N_1464,In_1770,In_344);
xnor U1465 (N_1465,In_1370,In_1419);
nand U1466 (N_1466,In_2049,In_2290);
or U1467 (N_1467,In_302,In_1400);
nor U1468 (N_1468,In_72,In_276);
xor U1469 (N_1469,In_1097,In_2295);
xor U1470 (N_1470,In_30,In_1186);
nor U1471 (N_1471,In_1173,In_1245);
nand U1472 (N_1472,In_883,In_1006);
nand U1473 (N_1473,In_1367,In_1657);
or U1474 (N_1474,In_1755,In_1916);
nor U1475 (N_1475,In_677,In_2023);
and U1476 (N_1476,In_535,In_382);
and U1477 (N_1477,In_1328,In_2490);
xor U1478 (N_1478,In_1436,In_1649);
nand U1479 (N_1479,In_819,In_70);
xor U1480 (N_1480,In_1096,In_1994);
or U1481 (N_1481,In_1041,In_404);
and U1482 (N_1482,In_1497,In_2437);
nor U1483 (N_1483,In_2074,In_356);
nand U1484 (N_1484,In_174,In_1356);
nand U1485 (N_1485,In_1344,In_1838);
xnor U1486 (N_1486,In_2299,In_1524);
nand U1487 (N_1487,In_1449,In_2219);
nand U1488 (N_1488,In_2441,In_1295);
xnor U1489 (N_1489,In_179,In_1392);
nor U1490 (N_1490,In_366,In_1843);
or U1491 (N_1491,In_733,In_927);
or U1492 (N_1492,In_90,In_1477);
or U1493 (N_1493,In_240,In_535);
and U1494 (N_1494,In_2194,In_1896);
or U1495 (N_1495,In_1880,In_1188);
or U1496 (N_1496,In_2467,In_2249);
nand U1497 (N_1497,In_422,In_2280);
and U1498 (N_1498,In_652,In_465);
xnor U1499 (N_1499,In_956,In_260);
or U1500 (N_1500,In_993,In_2007);
xnor U1501 (N_1501,In_1770,In_545);
and U1502 (N_1502,In_1067,In_609);
nor U1503 (N_1503,In_2001,In_291);
nand U1504 (N_1504,In_2466,In_458);
nand U1505 (N_1505,In_1109,In_371);
nor U1506 (N_1506,In_919,In_236);
xnor U1507 (N_1507,In_2461,In_706);
nand U1508 (N_1508,In_822,In_763);
or U1509 (N_1509,In_381,In_195);
xor U1510 (N_1510,In_1271,In_997);
and U1511 (N_1511,In_255,In_2466);
nor U1512 (N_1512,In_1650,In_2470);
and U1513 (N_1513,In_1827,In_1416);
nand U1514 (N_1514,In_1649,In_1487);
nor U1515 (N_1515,In_1318,In_2185);
nor U1516 (N_1516,In_2498,In_1657);
xnor U1517 (N_1517,In_455,In_1372);
xor U1518 (N_1518,In_1239,In_1548);
xor U1519 (N_1519,In_342,In_2026);
xnor U1520 (N_1520,In_1481,In_2024);
xor U1521 (N_1521,In_202,In_1942);
nor U1522 (N_1522,In_1868,In_1002);
and U1523 (N_1523,In_1316,In_1935);
nor U1524 (N_1524,In_348,In_1080);
and U1525 (N_1525,In_156,In_1125);
or U1526 (N_1526,In_977,In_1709);
or U1527 (N_1527,In_2204,In_925);
nor U1528 (N_1528,In_1185,In_1708);
and U1529 (N_1529,In_1790,In_1430);
nor U1530 (N_1530,In_1681,In_597);
nand U1531 (N_1531,In_501,In_750);
nand U1532 (N_1532,In_992,In_1916);
and U1533 (N_1533,In_2005,In_841);
or U1534 (N_1534,In_2172,In_1222);
nand U1535 (N_1535,In_2116,In_689);
xor U1536 (N_1536,In_243,In_10);
or U1537 (N_1537,In_515,In_1440);
nor U1538 (N_1538,In_82,In_43);
nand U1539 (N_1539,In_401,In_298);
and U1540 (N_1540,In_2021,In_1014);
nand U1541 (N_1541,In_368,In_693);
nor U1542 (N_1542,In_2361,In_2134);
or U1543 (N_1543,In_406,In_2002);
or U1544 (N_1544,In_214,In_417);
nand U1545 (N_1545,In_201,In_2154);
and U1546 (N_1546,In_2392,In_1762);
nor U1547 (N_1547,In_598,In_725);
nor U1548 (N_1548,In_811,In_1061);
xor U1549 (N_1549,In_2109,In_2307);
or U1550 (N_1550,In_1183,In_1422);
or U1551 (N_1551,In_464,In_1814);
xnor U1552 (N_1552,In_166,In_1467);
nand U1553 (N_1553,In_1476,In_2297);
nand U1554 (N_1554,In_379,In_1052);
or U1555 (N_1555,In_204,In_376);
xor U1556 (N_1556,In_1557,In_800);
and U1557 (N_1557,In_2044,In_113);
or U1558 (N_1558,In_263,In_1471);
or U1559 (N_1559,In_586,In_1998);
or U1560 (N_1560,In_1741,In_1011);
or U1561 (N_1561,In_1937,In_665);
nor U1562 (N_1562,In_2360,In_2318);
nand U1563 (N_1563,In_144,In_684);
nor U1564 (N_1564,In_394,In_1907);
nand U1565 (N_1565,In_1402,In_1449);
nor U1566 (N_1566,In_238,In_2433);
nand U1567 (N_1567,In_202,In_2188);
nand U1568 (N_1568,In_1547,In_1241);
xnor U1569 (N_1569,In_1190,In_1628);
nand U1570 (N_1570,In_107,In_799);
nor U1571 (N_1571,In_657,In_1713);
or U1572 (N_1572,In_1346,In_664);
or U1573 (N_1573,In_321,In_940);
and U1574 (N_1574,In_1065,In_847);
or U1575 (N_1575,In_1964,In_415);
and U1576 (N_1576,In_2235,In_1768);
nand U1577 (N_1577,In_696,In_2244);
nor U1578 (N_1578,In_1520,In_1840);
xor U1579 (N_1579,In_1160,In_108);
and U1580 (N_1580,In_1645,In_1954);
nand U1581 (N_1581,In_485,In_1561);
nor U1582 (N_1582,In_1698,In_92);
or U1583 (N_1583,In_2480,In_1980);
xnor U1584 (N_1584,In_1583,In_231);
or U1585 (N_1585,In_2009,In_2284);
nand U1586 (N_1586,In_1108,In_1606);
or U1587 (N_1587,In_394,In_50);
nor U1588 (N_1588,In_567,In_862);
and U1589 (N_1589,In_1532,In_537);
or U1590 (N_1590,In_1344,In_1198);
nor U1591 (N_1591,In_1827,In_1919);
xnor U1592 (N_1592,In_857,In_1437);
nand U1593 (N_1593,In_1924,In_211);
xor U1594 (N_1594,In_672,In_194);
and U1595 (N_1595,In_980,In_904);
nor U1596 (N_1596,In_1786,In_1135);
nor U1597 (N_1597,In_681,In_2080);
or U1598 (N_1598,In_1116,In_1108);
or U1599 (N_1599,In_853,In_1725);
or U1600 (N_1600,In_260,In_856);
xor U1601 (N_1601,In_469,In_2069);
and U1602 (N_1602,In_818,In_2291);
nor U1603 (N_1603,In_1360,In_1351);
nand U1604 (N_1604,In_1725,In_489);
xor U1605 (N_1605,In_753,In_1029);
nand U1606 (N_1606,In_1733,In_1760);
and U1607 (N_1607,In_1501,In_2332);
nor U1608 (N_1608,In_1335,In_706);
nor U1609 (N_1609,In_1610,In_2403);
nor U1610 (N_1610,In_333,In_932);
and U1611 (N_1611,In_402,In_259);
and U1612 (N_1612,In_1502,In_741);
nand U1613 (N_1613,In_343,In_863);
nand U1614 (N_1614,In_261,In_1968);
or U1615 (N_1615,In_2301,In_619);
or U1616 (N_1616,In_776,In_1749);
nand U1617 (N_1617,In_1960,In_662);
nor U1618 (N_1618,In_132,In_2092);
or U1619 (N_1619,In_452,In_461);
and U1620 (N_1620,In_465,In_224);
nand U1621 (N_1621,In_747,In_70);
and U1622 (N_1622,In_725,In_2218);
nor U1623 (N_1623,In_1020,In_1442);
and U1624 (N_1624,In_415,In_2123);
nand U1625 (N_1625,In_218,In_1116);
or U1626 (N_1626,In_1932,In_2124);
nor U1627 (N_1627,In_1682,In_955);
xnor U1628 (N_1628,In_3,In_2161);
and U1629 (N_1629,In_1193,In_1298);
or U1630 (N_1630,In_207,In_419);
xnor U1631 (N_1631,In_1435,In_377);
nor U1632 (N_1632,In_2022,In_1200);
or U1633 (N_1633,In_462,In_829);
nor U1634 (N_1634,In_1805,In_891);
nand U1635 (N_1635,In_1527,In_1877);
nor U1636 (N_1636,In_2317,In_1499);
and U1637 (N_1637,In_1069,In_2187);
nor U1638 (N_1638,In_436,In_1967);
or U1639 (N_1639,In_388,In_1156);
xor U1640 (N_1640,In_2028,In_1081);
xor U1641 (N_1641,In_1402,In_311);
and U1642 (N_1642,In_316,In_1288);
and U1643 (N_1643,In_1133,In_1797);
nand U1644 (N_1644,In_234,In_891);
and U1645 (N_1645,In_136,In_490);
nor U1646 (N_1646,In_725,In_1220);
or U1647 (N_1647,In_1064,In_1186);
nor U1648 (N_1648,In_2010,In_1628);
or U1649 (N_1649,In_1022,In_2112);
or U1650 (N_1650,In_661,In_1134);
nand U1651 (N_1651,In_815,In_1380);
nor U1652 (N_1652,In_702,In_1628);
and U1653 (N_1653,In_512,In_616);
or U1654 (N_1654,In_309,In_1505);
nand U1655 (N_1655,In_1595,In_1889);
or U1656 (N_1656,In_2477,In_229);
or U1657 (N_1657,In_2428,In_432);
or U1658 (N_1658,In_1733,In_1609);
or U1659 (N_1659,In_6,In_267);
nand U1660 (N_1660,In_868,In_2327);
and U1661 (N_1661,In_887,In_1201);
or U1662 (N_1662,In_677,In_820);
nand U1663 (N_1663,In_1529,In_2033);
and U1664 (N_1664,In_2251,In_292);
xnor U1665 (N_1665,In_1095,In_2346);
nand U1666 (N_1666,In_1145,In_129);
and U1667 (N_1667,In_931,In_2182);
or U1668 (N_1668,In_1327,In_300);
nor U1669 (N_1669,In_254,In_1798);
nor U1670 (N_1670,In_757,In_1508);
nand U1671 (N_1671,In_2122,In_672);
xnor U1672 (N_1672,In_1117,In_1134);
nand U1673 (N_1673,In_2161,In_1536);
nand U1674 (N_1674,In_207,In_129);
or U1675 (N_1675,In_2418,In_784);
nand U1676 (N_1676,In_112,In_349);
nor U1677 (N_1677,In_2005,In_1704);
or U1678 (N_1678,In_1008,In_895);
and U1679 (N_1679,In_405,In_1716);
nor U1680 (N_1680,In_1914,In_1292);
or U1681 (N_1681,In_1760,In_1954);
and U1682 (N_1682,In_791,In_1493);
and U1683 (N_1683,In_1870,In_1099);
nor U1684 (N_1684,In_1202,In_1041);
nand U1685 (N_1685,In_1735,In_719);
nand U1686 (N_1686,In_37,In_997);
nor U1687 (N_1687,In_2061,In_1062);
and U1688 (N_1688,In_1921,In_1902);
nor U1689 (N_1689,In_21,In_1922);
nand U1690 (N_1690,In_1150,In_1268);
xor U1691 (N_1691,In_1308,In_536);
nand U1692 (N_1692,In_1129,In_746);
xnor U1693 (N_1693,In_2275,In_1419);
nor U1694 (N_1694,In_1541,In_1501);
nand U1695 (N_1695,In_1086,In_2187);
nand U1696 (N_1696,In_1978,In_1038);
xnor U1697 (N_1697,In_553,In_2248);
or U1698 (N_1698,In_1341,In_2257);
or U1699 (N_1699,In_410,In_1650);
or U1700 (N_1700,In_2048,In_1141);
nor U1701 (N_1701,In_272,In_520);
nand U1702 (N_1702,In_1581,In_1538);
nor U1703 (N_1703,In_1159,In_666);
nand U1704 (N_1704,In_1899,In_687);
nand U1705 (N_1705,In_735,In_2463);
or U1706 (N_1706,In_415,In_328);
nor U1707 (N_1707,In_1114,In_765);
xnor U1708 (N_1708,In_1778,In_965);
nand U1709 (N_1709,In_1236,In_543);
nand U1710 (N_1710,In_1380,In_1892);
and U1711 (N_1711,In_1521,In_223);
or U1712 (N_1712,In_1882,In_2327);
xnor U1713 (N_1713,In_1032,In_1307);
nand U1714 (N_1714,In_1858,In_999);
or U1715 (N_1715,In_1864,In_705);
xnor U1716 (N_1716,In_473,In_522);
and U1717 (N_1717,In_1129,In_210);
and U1718 (N_1718,In_35,In_389);
xor U1719 (N_1719,In_568,In_2156);
or U1720 (N_1720,In_1566,In_2069);
nor U1721 (N_1721,In_539,In_571);
or U1722 (N_1722,In_1380,In_1487);
or U1723 (N_1723,In_1035,In_1020);
nor U1724 (N_1724,In_2066,In_871);
xor U1725 (N_1725,In_2039,In_2214);
nand U1726 (N_1726,In_448,In_677);
or U1727 (N_1727,In_2029,In_1283);
xnor U1728 (N_1728,In_400,In_922);
or U1729 (N_1729,In_1009,In_363);
xnor U1730 (N_1730,In_1499,In_968);
or U1731 (N_1731,In_2160,In_2367);
nand U1732 (N_1732,In_2404,In_1409);
and U1733 (N_1733,In_214,In_2006);
and U1734 (N_1734,In_1649,In_2194);
or U1735 (N_1735,In_2010,In_285);
nand U1736 (N_1736,In_1443,In_1800);
nor U1737 (N_1737,In_1433,In_1867);
nor U1738 (N_1738,In_966,In_2341);
and U1739 (N_1739,In_1629,In_2427);
or U1740 (N_1740,In_126,In_1339);
xor U1741 (N_1741,In_2022,In_717);
xor U1742 (N_1742,In_896,In_465);
and U1743 (N_1743,In_687,In_2318);
nor U1744 (N_1744,In_1860,In_1948);
or U1745 (N_1745,In_447,In_1432);
or U1746 (N_1746,In_1976,In_418);
nor U1747 (N_1747,In_8,In_353);
nor U1748 (N_1748,In_860,In_2283);
and U1749 (N_1749,In_718,In_2314);
xor U1750 (N_1750,In_1515,In_1653);
or U1751 (N_1751,In_2148,In_1948);
nand U1752 (N_1752,In_1541,In_293);
nand U1753 (N_1753,In_1023,In_2429);
nand U1754 (N_1754,In_1021,In_514);
xnor U1755 (N_1755,In_983,In_962);
xor U1756 (N_1756,In_1165,In_2264);
and U1757 (N_1757,In_1233,In_508);
xnor U1758 (N_1758,In_11,In_2193);
or U1759 (N_1759,In_717,In_1208);
and U1760 (N_1760,In_2302,In_1819);
and U1761 (N_1761,In_459,In_2278);
nand U1762 (N_1762,In_434,In_542);
and U1763 (N_1763,In_1586,In_1925);
or U1764 (N_1764,In_939,In_1);
nand U1765 (N_1765,In_130,In_624);
xnor U1766 (N_1766,In_138,In_2153);
xnor U1767 (N_1767,In_333,In_2021);
nand U1768 (N_1768,In_1378,In_1796);
or U1769 (N_1769,In_2292,In_2318);
xor U1770 (N_1770,In_299,In_454);
and U1771 (N_1771,In_2334,In_516);
nand U1772 (N_1772,In_1361,In_2379);
xor U1773 (N_1773,In_615,In_1976);
xor U1774 (N_1774,In_165,In_670);
nand U1775 (N_1775,In_830,In_776);
nand U1776 (N_1776,In_2465,In_665);
or U1777 (N_1777,In_2256,In_2211);
xor U1778 (N_1778,In_1588,In_471);
nand U1779 (N_1779,In_1467,In_1043);
nor U1780 (N_1780,In_1210,In_470);
and U1781 (N_1781,In_455,In_703);
xor U1782 (N_1782,In_2260,In_1114);
or U1783 (N_1783,In_113,In_976);
or U1784 (N_1784,In_844,In_939);
or U1785 (N_1785,In_1312,In_289);
nand U1786 (N_1786,In_2026,In_1161);
xnor U1787 (N_1787,In_734,In_2338);
and U1788 (N_1788,In_2285,In_993);
xnor U1789 (N_1789,In_2031,In_716);
nand U1790 (N_1790,In_1803,In_996);
and U1791 (N_1791,In_54,In_518);
nor U1792 (N_1792,In_2196,In_2077);
xor U1793 (N_1793,In_1743,In_734);
nor U1794 (N_1794,In_923,In_1319);
or U1795 (N_1795,In_859,In_2328);
or U1796 (N_1796,In_376,In_1670);
or U1797 (N_1797,In_1641,In_2036);
nand U1798 (N_1798,In_1287,In_1247);
nor U1799 (N_1799,In_914,In_2223);
nor U1800 (N_1800,In_698,In_1982);
nor U1801 (N_1801,In_1872,In_2281);
and U1802 (N_1802,In_2220,In_397);
or U1803 (N_1803,In_1867,In_1672);
nor U1804 (N_1804,In_939,In_373);
nor U1805 (N_1805,In_317,In_204);
xor U1806 (N_1806,In_348,In_1059);
and U1807 (N_1807,In_141,In_1620);
or U1808 (N_1808,In_1969,In_832);
or U1809 (N_1809,In_894,In_1804);
nand U1810 (N_1810,In_18,In_1088);
nor U1811 (N_1811,In_1968,In_721);
xor U1812 (N_1812,In_2017,In_1407);
or U1813 (N_1813,In_1619,In_883);
nor U1814 (N_1814,In_31,In_316);
nand U1815 (N_1815,In_1689,In_1819);
nor U1816 (N_1816,In_1189,In_808);
nand U1817 (N_1817,In_659,In_2447);
nand U1818 (N_1818,In_684,In_277);
nor U1819 (N_1819,In_2498,In_195);
xor U1820 (N_1820,In_217,In_1640);
and U1821 (N_1821,In_1481,In_2136);
xnor U1822 (N_1822,In_1886,In_344);
and U1823 (N_1823,In_414,In_1184);
or U1824 (N_1824,In_1526,In_1816);
or U1825 (N_1825,In_1485,In_1668);
and U1826 (N_1826,In_1632,In_316);
and U1827 (N_1827,In_959,In_595);
nand U1828 (N_1828,In_414,In_1163);
xnor U1829 (N_1829,In_2182,In_654);
or U1830 (N_1830,In_537,In_285);
nor U1831 (N_1831,In_726,In_1628);
and U1832 (N_1832,In_436,In_240);
and U1833 (N_1833,In_148,In_31);
xor U1834 (N_1834,In_1853,In_1024);
xor U1835 (N_1835,In_990,In_518);
and U1836 (N_1836,In_213,In_1807);
and U1837 (N_1837,In_2211,In_1044);
and U1838 (N_1838,In_768,In_1891);
or U1839 (N_1839,In_2157,In_833);
and U1840 (N_1840,In_2353,In_1919);
or U1841 (N_1841,In_2098,In_2217);
or U1842 (N_1842,In_1,In_686);
and U1843 (N_1843,In_1776,In_609);
nand U1844 (N_1844,In_568,In_2456);
xnor U1845 (N_1845,In_823,In_1130);
and U1846 (N_1846,In_2254,In_2201);
or U1847 (N_1847,In_2227,In_2048);
nor U1848 (N_1848,In_2033,In_273);
nand U1849 (N_1849,In_1354,In_1171);
xor U1850 (N_1850,In_383,In_1081);
nor U1851 (N_1851,In_163,In_1561);
nor U1852 (N_1852,In_1458,In_2067);
and U1853 (N_1853,In_490,In_1625);
nand U1854 (N_1854,In_2075,In_2350);
xnor U1855 (N_1855,In_2362,In_494);
nand U1856 (N_1856,In_2190,In_2042);
xnor U1857 (N_1857,In_27,In_1065);
nor U1858 (N_1858,In_1082,In_799);
nor U1859 (N_1859,In_62,In_856);
xnor U1860 (N_1860,In_910,In_1258);
xnor U1861 (N_1861,In_1101,In_2003);
nand U1862 (N_1862,In_355,In_1958);
nand U1863 (N_1863,In_370,In_1186);
xor U1864 (N_1864,In_1894,In_2044);
xor U1865 (N_1865,In_426,In_2017);
nand U1866 (N_1866,In_1003,In_462);
or U1867 (N_1867,In_1623,In_1089);
xnor U1868 (N_1868,In_2149,In_494);
nand U1869 (N_1869,In_687,In_767);
nor U1870 (N_1870,In_1883,In_2018);
nand U1871 (N_1871,In_103,In_1666);
or U1872 (N_1872,In_971,In_179);
or U1873 (N_1873,In_1964,In_1409);
nand U1874 (N_1874,In_1494,In_2222);
xnor U1875 (N_1875,In_819,In_810);
and U1876 (N_1876,In_2344,In_1580);
and U1877 (N_1877,In_1228,In_980);
nand U1878 (N_1878,In_337,In_1465);
nand U1879 (N_1879,In_876,In_1797);
nand U1880 (N_1880,In_1815,In_1058);
xor U1881 (N_1881,In_129,In_537);
nand U1882 (N_1882,In_1803,In_753);
and U1883 (N_1883,In_712,In_137);
nand U1884 (N_1884,In_1575,In_616);
xor U1885 (N_1885,In_1466,In_1846);
nand U1886 (N_1886,In_2052,In_1731);
nand U1887 (N_1887,In_1567,In_2012);
xnor U1888 (N_1888,In_2347,In_1930);
or U1889 (N_1889,In_792,In_881);
nand U1890 (N_1890,In_1148,In_2473);
or U1891 (N_1891,In_1762,In_1916);
xor U1892 (N_1892,In_333,In_1742);
xnor U1893 (N_1893,In_288,In_342);
nand U1894 (N_1894,In_2423,In_667);
or U1895 (N_1895,In_1871,In_852);
xnor U1896 (N_1896,In_2272,In_1659);
and U1897 (N_1897,In_356,In_298);
nand U1898 (N_1898,In_1857,In_389);
nor U1899 (N_1899,In_557,In_279);
and U1900 (N_1900,In_1359,In_969);
nor U1901 (N_1901,In_1614,In_622);
and U1902 (N_1902,In_2183,In_1811);
nor U1903 (N_1903,In_2044,In_1739);
xnor U1904 (N_1904,In_1856,In_208);
and U1905 (N_1905,In_126,In_404);
and U1906 (N_1906,In_158,In_880);
nor U1907 (N_1907,In_2449,In_1320);
nand U1908 (N_1908,In_1751,In_128);
nor U1909 (N_1909,In_1807,In_17);
nor U1910 (N_1910,In_172,In_1389);
xor U1911 (N_1911,In_965,In_286);
and U1912 (N_1912,In_419,In_92);
nor U1913 (N_1913,In_1875,In_1110);
or U1914 (N_1914,In_1604,In_467);
xor U1915 (N_1915,In_139,In_526);
nand U1916 (N_1916,In_430,In_124);
nor U1917 (N_1917,In_121,In_2167);
or U1918 (N_1918,In_428,In_1625);
and U1919 (N_1919,In_2125,In_2493);
and U1920 (N_1920,In_2410,In_425);
and U1921 (N_1921,In_108,In_2402);
nand U1922 (N_1922,In_878,In_786);
or U1923 (N_1923,In_1467,In_61);
nand U1924 (N_1924,In_955,In_759);
nor U1925 (N_1925,In_541,In_992);
xor U1926 (N_1926,In_300,In_368);
or U1927 (N_1927,In_651,In_2300);
xnor U1928 (N_1928,In_1503,In_1573);
xnor U1929 (N_1929,In_325,In_749);
xnor U1930 (N_1930,In_2037,In_1847);
nand U1931 (N_1931,In_1880,In_32);
nand U1932 (N_1932,In_159,In_1158);
nor U1933 (N_1933,In_527,In_2272);
nor U1934 (N_1934,In_163,In_119);
and U1935 (N_1935,In_1464,In_899);
xor U1936 (N_1936,In_342,In_1344);
or U1937 (N_1937,In_1492,In_1178);
nor U1938 (N_1938,In_746,In_863);
or U1939 (N_1939,In_467,In_1567);
nand U1940 (N_1940,In_1239,In_1319);
xnor U1941 (N_1941,In_2213,In_1471);
or U1942 (N_1942,In_408,In_1515);
nand U1943 (N_1943,In_2128,In_2001);
or U1944 (N_1944,In_921,In_369);
xnor U1945 (N_1945,In_2265,In_558);
and U1946 (N_1946,In_62,In_806);
or U1947 (N_1947,In_1765,In_1915);
and U1948 (N_1948,In_363,In_259);
or U1949 (N_1949,In_234,In_2183);
and U1950 (N_1950,In_25,In_1696);
or U1951 (N_1951,In_2064,In_1850);
nand U1952 (N_1952,In_97,In_421);
and U1953 (N_1953,In_877,In_471);
and U1954 (N_1954,In_6,In_1267);
nor U1955 (N_1955,In_1134,In_2143);
nand U1956 (N_1956,In_27,In_564);
xnor U1957 (N_1957,In_2144,In_1616);
xor U1958 (N_1958,In_2355,In_573);
xor U1959 (N_1959,In_296,In_2181);
and U1960 (N_1960,In_2028,In_1702);
xor U1961 (N_1961,In_1345,In_424);
or U1962 (N_1962,In_1344,In_3);
xnor U1963 (N_1963,In_2336,In_1299);
or U1964 (N_1964,In_1054,In_1535);
nor U1965 (N_1965,In_2388,In_1563);
nor U1966 (N_1966,In_993,In_186);
or U1967 (N_1967,In_2129,In_355);
xor U1968 (N_1968,In_1801,In_87);
nand U1969 (N_1969,In_743,In_959);
nand U1970 (N_1970,In_910,In_76);
xnor U1971 (N_1971,In_1145,In_2413);
and U1972 (N_1972,In_1663,In_350);
xnor U1973 (N_1973,In_1369,In_1868);
and U1974 (N_1974,In_707,In_1382);
or U1975 (N_1975,In_2248,In_1931);
xor U1976 (N_1976,In_977,In_947);
nand U1977 (N_1977,In_529,In_575);
nand U1978 (N_1978,In_2303,In_1986);
and U1979 (N_1979,In_2362,In_1032);
and U1980 (N_1980,In_205,In_2133);
nor U1981 (N_1981,In_829,In_1677);
and U1982 (N_1982,In_838,In_1746);
or U1983 (N_1983,In_1872,In_1250);
and U1984 (N_1984,In_1818,In_8);
xor U1985 (N_1985,In_565,In_1177);
nor U1986 (N_1986,In_1497,In_1961);
nor U1987 (N_1987,In_813,In_2237);
nand U1988 (N_1988,In_2482,In_627);
xor U1989 (N_1989,In_2144,In_1007);
xnor U1990 (N_1990,In_2369,In_284);
xnor U1991 (N_1991,In_701,In_227);
and U1992 (N_1992,In_1022,In_1177);
or U1993 (N_1993,In_2476,In_1832);
xnor U1994 (N_1994,In_1620,In_1580);
nand U1995 (N_1995,In_1865,In_1287);
or U1996 (N_1996,In_1635,In_1334);
or U1997 (N_1997,In_1230,In_1908);
or U1998 (N_1998,In_2436,In_1718);
xor U1999 (N_1999,In_1296,In_1945);
nor U2000 (N_2000,In_1479,In_672);
or U2001 (N_2001,In_132,In_1323);
and U2002 (N_2002,In_1093,In_724);
and U2003 (N_2003,In_2047,In_1396);
and U2004 (N_2004,In_1725,In_644);
nor U2005 (N_2005,In_1055,In_261);
nor U2006 (N_2006,In_1910,In_865);
nor U2007 (N_2007,In_29,In_1909);
xnor U2008 (N_2008,In_443,In_1776);
xnor U2009 (N_2009,In_588,In_2140);
or U2010 (N_2010,In_2323,In_1259);
and U2011 (N_2011,In_660,In_219);
xor U2012 (N_2012,In_552,In_718);
or U2013 (N_2013,In_219,In_1457);
or U2014 (N_2014,In_2285,In_1165);
xnor U2015 (N_2015,In_1928,In_677);
and U2016 (N_2016,In_2262,In_1218);
xor U2017 (N_2017,In_178,In_1669);
nand U2018 (N_2018,In_1598,In_976);
xor U2019 (N_2019,In_230,In_1238);
xnor U2020 (N_2020,In_2106,In_1879);
nand U2021 (N_2021,In_2137,In_1501);
nor U2022 (N_2022,In_1939,In_147);
or U2023 (N_2023,In_320,In_84);
xnor U2024 (N_2024,In_388,In_1120);
or U2025 (N_2025,In_736,In_860);
nand U2026 (N_2026,In_196,In_2427);
nand U2027 (N_2027,In_489,In_1348);
and U2028 (N_2028,In_329,In_1504);
xnor U2029 (N_2029,In_1975,In_812);
xnor U2030 (N_2030,In_1399,In_1820);
or U2031 (N_2031,In_1497,In_1677);
nand U2032 (N_2032,In_2210,In_2380);
or U2033 (N_2033,In_235,In_1470);
and U2034 (N_2034,In_690,In_1820);
and U2035 (N_2035,In_2271,In_639);
nor U2036 (N_2036,In_1943,In_1380);
xor U2037 (N_2037,In_2251,In_725);
nor U2038 (N_2038,In_729,In_1215);
nor U2039 (N_2039,In_288,In_1944);
and U2040 (N_2040,In_1531,In_1910);
or U2041 (N_2041,In_145,In_1376);
nand U2042 (N_2042,In_1858,In_480);
xnor U2043 (N_2043,In_1369,In_772);
nor U2044 (N_2044,In_2213,In_1603);
xnor U2045 (N_2045,In_2150,In_864);
and U2046 (N_2046,In_1244,In_1634);
or U2047 (N_2047,In_1841,In_1715);
and U2048 (N_2048,In_2471,In_742);
nand U2049 (N_2049,In_43,In_2293);
or U2050 (N_2050,In_130,In_288);
or U2051 (N_2051,In_1000,In_1987);
or U2052 (N_2052,In_1062,In_605);
nand U2053 (N_2053,In_922,In_2229);
xor U2054 (N_2054,In_840,In_630);
or U2055 (N_2055,In_2249,In_2496);
xnor U2056 (N_2056,In_1687,In_2316);
nand U2057 (N_2057,In_2139,In_1860);
xor U2058 (N_2058,In_1586,In_568);
nand U2059 (N_2059,In_1848,In_359);
xor U2060 (N_2060,In_2002,In_1053);
or U2061 (N_2061,In_1809,In_2022);
nand U2062 (N_2062,In_161,In_2307);
or U2063 (N_2063,In_634,In_1452);
or U2064 (N_2064,In_2314,In_1892);
and U2065 (N_2065,In_1293,In_654);
nor U2066 (N_2066,In_219,In_953);
nor U2067 (N_2067,In_1903,In_225);
or U2068 (N_2068,In_373,In_1258);
nand U2069 (N_2069,In_1159,In_1612);
and U2070 (N_2070,In_1903,In_742);
xnor U2071 (N_2071,In_95,In_340);
nor U2072 (N_2072,In_1059,In_420);
xnor U2073 (N_2073,In_473,In_596);
nor U2074 (N_2074,In_709,In_164);
nor U2075 (N_2075,In_672,In_417);
and U2076 (N_2076,In_2496,In_246);
xor U2077 (N_2077,In_1812,In_1919);
or U2078 (N_2078,In_364,In_814);
nor U2079 (N_2079,In_2409,In_2041);
nor U2080 (N_2080,In_2280,In_870);
and U2081 (N_2081,In_761,In_1568);
and U2082 (N_2082,In_1321,In_1365);
or U2083 (N_2083,In_1623,In_553);
or U2084 (N_2084,In_1140,In_1566);
or U2085 (N_2085,In_1571,In_11);
nor U2086 (N_2086,In_399,In_263);
and U2087 (N_2087,In_536,In_1951);
nor U2088 (N_2088,In_1708,In_1927);
and U2089 (N_2089,In_1619,In_343);
and U2090 (N_2090,In_682,In_1834);
and U2091 (N_2091,In_1566,In_1220);
or U2092 (N_2092,In_1764,In_507);
xnor U2093 (N_2093,In_908,In_500);
nor U2094 (N_2094,In_1093,In_688);
nor U2095 (N_2095,In_1837,In_1855);
xor U2096 (N_2096,In_1951,In_1182);
nand U2097 (N_2097,In_803,In_1407);
nor U2098 (N_2098,In_449,In_1044);
nor U2099 (N_2099,In_1328,In_1582);
or U2100 (N_2100,In_1609,In_683);
and U2101 (N_2101,In_436,In_2009);
nand U2102 (N_2102,In_1610,In_1385);
nand U2103 (N_2103,In_1702,In_501);
nor U2104 (N_2104,In_997,In_2138);
and U2105 (N_2105,In_216,In_2043);
nand U2106 (N_2106,In_2127,In_1461);
nor U2107 (N_2107,In_1086,In_1988);
or U2108 (N_2108,In_2058,In_226);
and U2109 (N_2109,In_1769,In_1636);
nor U2110 (N_2110,In_2475,In_1242);
xor U2111 (N_2111,In_2372,In_1037);
nand U2112 (N_2112,In_942,In_661);
nand U2113 (N_2113,In_2320,In_2385);
or U2114 (N_2114,In_632,In_1316);
and U2115 (N_2115,In_64,In_1243);
or U2116 (N_2116,In_88,In_535);
nor U2117 (N_2117,In_341,In_977);
nand U2118 (N_2118,In_78,In_1587);
nand U2119 (N_2119,In_908,In_650);
xnor U2120 (N_2120,In_1943,In_793);
or U2121 (N_2121,In_215,In_1289);
or U2122 (N_2122,In_1765,In_1468);
nor U2123 (N_2123,In_1922,In_1470);
or U2124 (N_2124,In_2441,In_274);
xor U2125 (N_2125,In_2156,In_2024);
nor U2126 (N_2126,In_1076,In_417);
xnor U2127 (N_2127,In_2160,In_1852);
nand U2128 (N_2128,In_719,In_216);
xnor U2129 (N_2129,In_207,In_1366);
nand U2130 (N_2130,In_809,In_1779);
and U2131 (N_2131,In_91,In_225);
nor U2132 (N_2132,In_1987,In_1932);
and U2133 (N_2133,In_1911,In_293);
and U2134 (N_2134,In_2022,In_314);
or U2135 (N_2135,In_1046,In_986);
or U2136 (N_2136,In_2173,In_46);
nand U2137 (N_2137,In_2450,In_1199);
or U2138 (N_2138,In_1737,In_581);
nor U2139 (N_2139,In_44,In_929);
nand U2140 (N_2140,In_1002,In_626);
or U2141 (N_2141,In_2198,In_2444);
xor U2142 (N_2142,In_966,In_1567);
nor U2143 (N_2143,In_1279,In_397);
nand U2144 (N_2144,In_683,In_2370);
or U2145 (N_2145,In_797,In_485);
or U2146 (N_2146,In_1854,In_1501);
nand U2147 (N_2147,In_1394,In_2238);
xnor U2148 (N_2148,In_371,In_1449);
and U2149 (N_2149,In_1218,In_204);
xnor U2150 (N_2150,In_606,In_2345);
xnor U2151 (N_2151,In_233,In_715);
xor U2152 (N_2152,In_940,In_735);
nand U2153 (N_2153,In_1507,In_1707);
or U2154 (N_2154,In_1053,In_2352);
nor U2155 (N_2155,In_1597,In_2104);
nand U2156 (N_2156,In_2099,In_414);
and U2157 (N_2157,In_678,In_439);
or U2158 (N_2158,In_1600,In_536);
xor U2159 (N_2159,In_2179,In_465);
and U2160 (N_2160,In_1566,In_609);
nand U2161 (N_2161,In_1941,In_892);
xnor U2162 (N_2162,In_2282,In_1432);
nor U2163 (N_2163,In_1250,In_2197);
nor U2164 (N_2164,In_1082,In_833);
nor U2165 (N_2165,In_535,In_1913);
or U2166 (N_2166,In_963,In_118);
xnor U2167 (N_2167,In_114,In_951);
xnor U2168 (N_2168,In_1454,In_2452);
nor U2169 (N_2169,In_368,In_2126);
xor U2170 (N_2170,In_2186,In_1564);
or U2171 (N_2171,In_478,In_1908);
and U2172 (N_2172,In_1670,In_276);
and U2173 (N_2173,In_1910,In_636);
or U2174 (N_2174,In_2442,In_515);
nand U2175 (N_2175,In_1264,In_1453);
nand U2176 (N_2176,In_1424,In_1257);
nor U2177 (N_2177,In_2447,In_1724);
and U2178 (N_2178,In_943,In_465);
nor U2179 (N_2179,In_474,In_2035);
xnor U2180 (N_2180,In_777,In_2231);
xor U2181 (N_2181,In_855,In_265);
nor U2182 (N_2182,In_2128,In_471);
and U2183 (N_2183,In_152,In_1407);
or U2184 (N_2184,In_743,In_1292);
or U2185 (N_2185,In_2386,In_2363);
and U2186 (N_2186,In_207,In_1003);
nand U2187 (N_2187,In_907,In_210);
nor U2188 (N_2188,In_7,In_1158);
nand U2189 (N_2189,In_1978,In_687);
xor U2190 (N_2190,In_109,In_349);
nor U2191 (N_2191,In_1114,In_1099);
and U2192 (N_2192,In_759,In_2215);
or U2193 (N_2193,In_1062,In_2015);
and U2194 (N_2194,In_1505,In_1470);
or U2195 (N_2195,In_2134,In_1357);
xor U2196 (N_2196,In_607,In_1742);
or U2197 (N_2197,In_1936,In_2113);
xor U2198 (N_2198,In_1684,In_1204);
nor U2199 (N_2199,In_2275,In_1591);
nand U2200 (N_2200,In_161,In_1202);
nor U2201 (N_2201,In_2347,In_1714);
nor U2202 (N_2202,In_1573,In_20);
or U2203 (N_2203,In_638,In_487);
and U2204 (N_2204,In_1052,In_64);
and U2205 (N_2205,In_1489,In_1863);
nor U2206 (N_2206,In_266,In_2441);
nor U2207 (N_2207,In_1482,In_352);
xnor U2208 (N_2208,In_962,In_1552);
or U2209 (N_2209,In_2290,In_594);
nand U2210 (N_2210,In_378,In_2423);
nand U2211 (N_2211,In_1618,In_1122);
xnor U2212 (N_2212,In_62,In_329);
nor U2213 (N_2213,In_1396,In_874);
xor U2214 (N_2214,In_353,In_228);
nand U2215 (N_2215,In_867,In_1442);
and U2216 (N_2216,In_1484,In_1689);
or U2217 (N_2217,In_1152,In_398);
nor U2218 (N_2218,In_981,In_1501);
nor U2219 (N_2219,In_2346,In_1351);
nand U2220 (N_2220,In_711,In_1282);
xnor U2221 (N_2221,In_523,In_879);
xnor U2222 (N_2222,In_2099,In_1811);
and U2223 (N_2223,In_1281,In_1205);
and U2224 (N_2224,In_1333,In_872);
nor U2225 (N_2225,In_1202,In_1730);
xnor U2226 (N_2226,In_2054,In_1730);
xor U2227 (N_2227,In_56,In_116);
xor U2228 (N_2228,In_1983,In_823);
nand U2229 (N_2229,In_1303,In_2189);
xor U2230 (N_2230,In_535,In_98);
and U2231 (N_2231,In_1080,In_545);
nand U2232 (N_2232,In_1629,In_1578);
nor U2233 (N_2233,In_418,In_1997);
or U2234 (N_2234,In_813,In_2285);
xnor U2235 (N_2235,In_2300,In_1488);
and U2236 (N_2236,In_333,In_1163);
and U2237 (N_2237,In_797,In_882);
xor U2238 (N_2238,In_1952,In_2404);
xor U2239 (N_2239,In_647,In_931);
xor U2240 (N_2240,In_1199,In_2053);
nor U2241 (N_2241,In_1886,In_1260);
and U2242 (N_2242,In_1223,In_788);
and U2243 (N_2243,In_212,In_1981);
nor U2244 (N_2244,In_117,In_1756);
nand U2245 (N_2245,In_8,In_750);
nor U2246 (N_2246,In_399,In_1052);
or U2247 (N_2247,In_1227,In_620);
xor U2248 (N_2248,In_375,In_2122);
and U2249 (N_2249,In_1601,In_313);
nand U2250 (N_2250,In_1658,In_109);
xor U2251 (N_2251,In_1336,In_560);
xnor U2252 (N_2252,In_1401,In_1459);
nand U2253 (N_2253,In_1975,In_2405);
nand U2254 (N_2254,In_828,In_2084);
nor U2255 (N_2255,In_2155,In_796);
xnor U2256 (N_2256,In_1177,In_2371);
nor U2257 (N_2257,In_677,In_764);
nor U2258 (N_2258,In_1054,In_1321);
nand U2259 (N_2259,In_1153,In_1356);
xnor U2260 (N_2260,In_960,In_1134);
nand U2261 (N_2261,In_1064,In_971);
xnor U2262 (N_2262,In_900,In_2383);
nand U2263 (N_2263,In_2182,In_464);
and U2264 (N_2264,In_755,In_100);
xor U2265 (N_2265,In_1992,In_260);
and U2266 (N_2266,In_1643,In_1345);
and U2267 (N_2267,In_330,In_2209);
or U2268 (N_2268,In_2270,In_1551);
nand U2269 (N_2269,In_1545,In_656);
or U2270 (N_2270,In_2061,In_2287);
nor U2271 (N_2271,In_2060,In_422);
and U2272 (N_2272,In_1137,In_481);
nor U2273 (N_2273,In_141,In_2382);
nor U2274 (N_2274,In_2398,In_2032);
nor U2275 (N_2275,In_1699,In_1591);
nor U2276 (N_2276,In_2070,In_604);
nor U2277 (N_2277,In_1574,In_1570);
nor U2278 (N_2278,In_255,In_1904);
xor U2279 (N_2279,In_1457,In_704);
or U2280 (N_2280,In_2085,In_1163);
and U2281 (N_2281,In_803,In_666);
nand U2282 (N_2282,In_603,In_1053);
or U2283 (N_2283,In_1904,In_2271);
xnor U2284 (N_2284,In_1265,In_1605);
or U2285 (N_2285,In_1590,In_2437);
and U2286 (N_2286,In_1148,In_324);
and U2287 (N_2287,In_2407,In_236);
xor U2288 (N_2288,In_1840,In_224);
nor U2289 (N_2289,In_536,In_2463);
and U2290 (N_2290,In_1356,In_1662);
and U2291 (N_2291,In_962,In_1329);
or U2292 (N_2292,In_1383,In_1634);
xor U2293 (N_2293,In_1902,In_66);
and U2294 (N_2294,In_2053,In_984);
or U2295 (N_2295,In_1487,In_289);
or U2296 (N_2296,In_1437,In_474);
xor U2297 (N_2297,In_1092,In_1422);
nand U2298 (N_2298,In_987,In_1794);
or U2299 (N_2299,In_2281,In_598);
nor U2300 (N_2300,In_2154,In_568);
nand U2301 (N_2301,In_2203,In_1301);
or U2302 (N_2302,In_496,In_2382);
nand U2303 (N_2303,In_1795,In_1246);
nand U2304 (N_2304,In_1477,In_465);
nand U2305 (N_2305,In_621,In_2155);
xor U2306 (N_2306,In_986,In_731);
or U2307 (N_2307,In_132,In_645);
nor U2308 (N_2308,In_2282,In_1608);
xnor U2309 (N_2309,In_2287,In_1360);
nand U2310 (N_2310,In_1764,In_2326);
or U2311 (N_2311,In_723,In_2187);
and U2312 (N_2312,In_820,In_861);
or U2313 (N_2313,In_1156,In_2345);
xnor U2314 (N_2314,In_341,In_855);
and U2315 (N_2315,In_696,In_321);
or U2316 (N_2316,In_455,In_2204);
nand U2317 (N_2317,In_1286,In_1317);
nor U2318 (N_2318,In_635,In_420);
and U2319 (N_2319,In_1043,In_1094);
nor U2320 (N_2320,In_94,In_2062);
xor U2321 (N_2321,In_1966,In_2340);
nand U2322 (N_2322,In_2190,In_843);
xnor U2323 (N_2323,In_56,In_948);
or U2324 (N_2324,In_1134,In_1091);
nor U2325 (N_2325,In_2298,In_1672);
or U2326 (N_2326,In_1655,In_906);
nor U2327 (N_2327,In_1083,In_1611);
nand U2328 (N_2328,In_1013,In_1393);
or U2329 (N_2329,In_1563,In_2105);
and U2330 (N_2330,In_2470,In_468);
xnor U2331 (N_2331,In_564,In_1449);
nand U2332 (N_2332,In_154,In_366);
and U2333 (N_2333,In_1351,In_1472);
or U2334 (N_2334,In_538,In_925);
nand U2335 (N_2335,In_1016,In_1035);
xor U2336 (N_2336,In_1639,In_839);
and U2337 (N_2337,In_821,In_237);
nand U2338 (N_2338,In_2435,In_824);
nand U2339 (N_2339,In_151,In_148);
and U2340 (N_2340,In_1186,In_1383);
nand U2341 (N_2341,In_2110,In_1096);
nor U2342 (N_2342,In_412,In_2234);
or U2343 (N_2343,In_1590,In_1220);
nor U2344 (N_2344,In_1191,In_1349);
and U2345 (N_2345,In_1152,In_5);
or U2346 (N_2346,In_335,In_297);
and U2347 (N_2347,In_2436,In_1827);
nand U2348 (N_2348,In_1733,In_2398);
and U2349 (N_2349,In_162,In_2281);
or U2350 (N_2350,In_123,In_258);
and U2351 (N_2351,In_765,In_1969);
nand U2352 (N_2352,In_453,In_1736);
nor U2353 (N_2353,In_468,In_491);
or U2354 (N_2354,In_65,In_757);
and U2355 (N_2355,In_957,In_90);
nor U2356 (N_2356,In_825,In_2178);
and U2357 (N_2357,In_2368,In_266);
or U2358 (N_2358,In_2092,In_1008);
and U2359 (N_2359,In_904,In_1590);
nand U2360 (N_2360,In_451,In_543);
xor U2361 (N_2361,In_1773,In_114);
nand U2362 (N_2362,In_1181,In_700);
or U2363 (N_2363,In_1682,In_2203);
nor U2364 (N_2364,In_995,In_2483);
nand U2365 (N_2365,In_69,In_1283);
nor U2366 (N_2366,In_1821,In_63);
nor U2367 (N_2367,In_1605,In_1013);
or U2368 (N_2368,In_251,In_2014);
nor U2369 (N_2369,In_1928,In_998);
nor U2370 (N_2370,In_1379,In_444);
nor U2371 (N_2371,In_127,In_1972);
nand U2372 (N_2372,In_1662,In_1791);
and U2373 (N_2373,In_189,In_596);
or U2374 (N_2374,In_540,In_394);
or U2375 (N_2375,In_557,In_515);
or U2376 (N_2376,In_2307,In_408);
xor U2377 (N_2377,In_2271,In_681);
xnor U2378 (N_2378,In_666,In_1402);
nor U2379 (N_2379,In_431,In_735);
nand U2380 (N_2380,In_550,In_1226);
xor U2381 (N_2381,In_2352,In_1656);
or U2382 (N_2382,In_369,In_34);
nand U2383 (N_2383,In_1343,In_1232);
xnor U2384 (N_2384,In_2211,In_2438);
xor U2385 (N_2385,In_1490,In_972);
xnor U2386 (N_2386,In_2091,In_2322);
or U2387 (N_2387,In_633,In_1569);
xor U2388 (N_2388,In_663,In_1057);
xor U2389 (N_2389,In_586,In_593);
nor U2390 (N_2390,In_1315,In_517);
nor U2391 (N_2391,In_2385,In_237);
nor U2392 (N_2392,In_2467,In_1377);
and U2393 (N_2393,In_884,In_1900);
nand U2394 (N_2394,In_1406,In_838);
and U2395 (N_2395,In_1308,In_327);
xnor U2396 (N_2396,In_294,In_363);
and U2397 (N_2397,In_1716,In_36);
and U2398 (N_2398,In_2292,In_2263);
and U2399 (N_2399,In_868,In_2206);
and U2400 (N_2400,In_1289,In_591);
nand U2401 (N_2401,In_1473,In_2451);
nor U2402 (N_2402,In_1032,In_1129);
and U2403 (N_2403,In_1268,In_723);
and U2404 (N_2404,In_2348,In_1401);
or U2405 (N_2405,In_1327,In_1007);
nand U2406 (N_2406,In_220,In_1414);
nor U2407 (N_2407,In_839,In_1660);
or U2408 (N_2408,In_1268,In_1903);
and U2409 (N_2409,In_692,In_2238);
nor U2410 (N_2410,In_784,In_108);
xor U2411 (N_2411,In_1727,In_438);
xnor U2412 (N_2412,In_1818,In_2407);
nand U2413 (N_2413,In_1163,In_2237);
and U2414 (N_2414,In_1132,In_122);
and U2415 (N_2415,In_1067,In_1686);
or U2416 (N_2416,In_895,In_244);
and U2417 (N_2417,In_1945,In_1483);
and U2418 (N_2418,In_922,In_2485);
nand U2419 (N_2419,In_1152,In_1119);
nor U2420 (N_2420,In_1620,In_2216);
or U2421 (N_2421,In_543,In_1403);
and U2422 (N_2422,In_736,In_2424);
nand U2423 (N_2423,In_1626,In_1328);
xnor U2424 (N_2424,In_2198,In_1071);
nand U2425 (N_2425,In_424,In_1294);
xor U2426 (N_2426,In_1777,In_2247);
or U2427 (N_2427,In_916,In_1863);
or U2428 (N_2428,In_1317,In_531);
and U2429 (N_2429,In_1501,In_637);
xnor U2430 (N_2430,In_1689,In_1300);
nand U2431 (N_2431,In_307,In_1962);
xor U2432 (N_2432,In_1274,In_1691);
and U2433 (N_2433,In_1177,In_1032);
and U2434 (N_2434,In_2070,In_411);
nand U2435 (N_2435,In_1931,In_724);
and U2436 (N_2436,In_2275,In_2064);
nand U2437 (N_2437,In_928,In_51);
and U2438 (N_2438,In_652,In_1380);
and U2439 (N_2439,In_29,In_1059);
xor U2440 (N_2440,In_442,In_1949);
and U2441 (N_2441,In_2282,In_1832);
nor U2442 (N_2442,In_1470,In_1069);
or U2443 (N_2443,In_1072,In_1444);
xnor U2444 (N_2444,In_1457,In_1627);
nand U2445 (N_2445,In_2317,In_1562);
xor U2446 (N_2446,In_892,In_700);
nor U2447 (N_2447,In_104,In_1719);
or U2448 (N_2448,In_269,In_1802);
xnor U2449 (N_2449,In_276,In_1519);
nor U2450 (N_2450,In_1790,In_972);
xnor U2451 (N_2451,In_2144,In_1537);
and U2452 (N_2452,In_1603,In_441);
nand U2453 (N_2453,In_1543,In_869);
nor U2454 (N_2454,In_1833,In_1876);
nand U2455 (N_2455,In_1303,In_2298);
xnor U2456 (N_2456,In_117,In_1874);
and U2457 (N_2457,In_1886,In_112);
nand U2458 (N_2458,In_658,In_1373);
xor U2459 (N_2459,In_1802,In_244);
xnor U2460 (N_2460,In_1660,In_541);
xnor U2461 (N_2461,In_686,In_1035);
nand U2462 (N_2462,In_2334,In_319);
nor U2463 (N_2463,In_2137,In_1295);
or U2464 (N_2464,In_1649,In_2173);
and U2465 (N_2465,In_1936,In_2152);
or U2466 (N_2466,In_1991,In_1898);
nor U2467 (N_2467,In_2340,In_1211);
and U2468 (N_2468,In_2165,In_851);
xnor U2469 (N_2469,In_748,In_984);
and U2470 (N_2470,In_253,In_2486);
and U2471 (N_2471,In_2274,In_1231);
nand U2472 (N_2472,In_2220,In_2199);
or U2473 (N_2473,In_210,In_1721);
and U2474 (N_2474,In_1879,In_1418);
xnor U2475 (N_2475,In_1112,In_2036);
nand U2476 (N_2476,In_1565,In_1882);
xor U2477 (N_2477,In_883,In_858);
or U2478 (N_2478,In_692,In_527);
or U2479 (N_2479,In_1999,In_515);
or U2480 (N_2480,In_604,In_1733);
xnor U2481 (N_2481,In_1707,In_1343);
nand U2482 (N_2482,In_578,In_1395);
or U2483 (N_2483,In_1552,In_887);
xor U2484 (N_2484,In_2232,In_986);
xnor U2485 (N_2485,In_435,In_1597);
nand U2486 (N_2486,In_530,In_1332);
or U2487 (N_2487,In_2212,In_915);
and U2488 (N_2488,In_810,In_865);
nor U2489 (N_2489,In_1230,In_2019);
and U2490 (N_2490,In_1873,In_2080);
nand U2491 (N_2491,In_2196,In_2320);
nor U2492 (N_2492,In_458,In_1827);
and U2493 (N_2493,In_91,In_1340);
and U2494 (N_2494,In_1750,In_1963);
xnor U2495 (N_2495,In_1154,In_616);
and U2496 (N_2496,In_1101,In_1015);
nor U2497 (N_2497,In_2431,In_2420);
xnor U2498 (N_2498,In_1571,In_1478);
nand U2499 (N_2499,In_1682,In_2419);
and U2500 (N_2500,In_675,In_1687);
xor U2501 (N_2501,In_438,In_1146);
and U2502 (N_2502,In_242,In_365);
and U2503 (N_2503,In_206,In_1889);
xnor U2504 (N_2504,In_15,In_987);
or U2505 (N_2505,In_1127,In_1322);
nand U2506 (N_2506,In_1956,In_1238);
or U2507 (N_2507,In_1556,In_1645);
and U2508 (N_2508,In_274,In_1106);
and U2509 (N_2509,In_1592,In_465);
and U2510 (N_2510,In_126,In_2177);
xnor U2511 (N_2511,In_476,In_1146);
nor U2512 (N_2512,In_1255,In_2235);
nor U2513 (N_2513,In_1069,In_1510);
nand U2514 (N_2514,In_1250,In_480);
nand U2515 (N_2515,In_1465,In_1025);
nor U2516 (N_2516,In_188,In_2065);
nand U2517 (N_2517,In_940,In_676);
or U2518 (N_2518,In_1096,In_2334);
xnor U2519 (N_2519,In_1965,In_680);
xor U2520 (N_2520,In_959,In_2401);
or U2521 (N_2521,In_987,In_1729);
nand U2522 (N_2522,In_184,In_2006);
or U2523 (N_2523,In_756,In_388);
xor U2524 (N_2524,In_258,In_1562);
and U2525 (N_2525,In_964,In_2451);
xor U2526 (N_2526,In_500,In_414);
and U2527 (N_2527,In_1265,In_2320);
nand U2528 (N_2528,In_377,In_1639);
nor U2529 (N_2529,In_484,In_1035);
nor U2530 (N_2530,In_209,In_2467);
and U2531 (N_2531,In_111,In_777);
xor U2532 (N_2532,In_779,In_1188);
and U2533 (N_2533,In_1808,In_695);
nand U2534 (N_2534,In_672,In_2193);
xor U2535 (N_2535,In_527,In_2132);
xor U2536 (N_2536,In_1220,In_1290);
xor U2537 (N_2537,In_2334,In_486);
and U2538 (N_2538,In_695,In_1635);
nand U2539 (N_2539,In_193,In_613);
xor U2540 (N_2540,In_908,In_1010);
xor U2541 (N_2541,In_156,In_1648);
and U2542 (N_2542,In_159,In_1967);
nand U2543 (N_2543,In_792,In_1891);
nor U2544 (N_2544,In_1712,In_2132);
and U2545 (N_2545,In_146,In_2226);
xor U2546 (N_2546,In_2160,In_1266);
and U2547 (N_2547,In_1008,In_301);
nand U2548 (N_2548,In_1813,In_2166);
nand U2549 (N_2549,In_1069,In_207);
xnor U2550 (N_2550,In_311,In_1254);
and U2551 (N_2551,In_626,In_1545);
nor U2552 (N_2552,In_1228,In_1931);
nor U2553 (N_2553,In_310,In_137);
or U2554 (N_2554,In_1358,In_2031);
xor U2555 (N_2555,In_124,In_1169);
or U2556 (N_2556,In_401,In_1865);
nand U2557 (N_2557,In_117,In_2466);
nor U2558 (N_2558,In_783,In_2040);
or U2559 (N_2559,In_1400,In_1926);
or U2560 (N_2560,In_1249,In_836);
xnor U2561 (N_2561,In_2436,In_1873);
xor U2562 (N_2562,In_1988,In_1769);
nor U2563 (N_2563,In_20,In_901);
nand U2564 (N_2564,In_1147,In_1165);
or U2565 (N_2565,In_1248,In_2174);
or U2566 (N_2566,In_1714,In_1176);
nand U2567 (N_2567,In_278,In_1858);
xnor U2568 (N_2568,In_1464,In_540);
and U2569 (N_2569,In_566,In_2280);
and U2570 (N_2570,In_1823,In_1449);
xor U2571 (N_2571,In_2061,In_1200);
xnor U2572 (N_2572,In_480,In_1333);
and U2573 (N_2573,In_1286,In_349);
or U2574 (N_2574,In_1703,In_429);
or U2575 (N_2575,In_948,In_1583);
xor U2576 (N_2576,In_1748,In_196);
or U2577 (N_2577,In_15,In_2395);
nand U2578 (N_2578,In_1613,In_1220);
nor U2579 (N_2579,In_118,In_1368);
and U2580 (N_2580,In_1439,In_2000);
or U2581 (N_2581,In_2074,In_106);
and U2582 (N_2582,In_367,In_1341);
nand U2583 (N_2583,In_235,In_919);
or U2584 (N_2584,In_2181,In_1940);
xnor U2585 (N_2585,In_148,In_2287);
xor U2586 (N_2586,In_1378,In_1283);
nand U2587 (N_2587,In_220,In_992);
xor U2588 (N_2588,In_852,In_1494);
nand U2589 (N_2589,In_900,In_2389);
and U2590 (N_2590,In_1474,In_882);
nor U2591 (N_2591,In_155,In_2357);
or U2592 (N_2592,In_401,In_1650);
xor U2593 (N_2593,In_1828,In_317);
nand U2594 (N_2594,In_1281,In_588);
xor U2595 (N_2595,In_615,In_2233);
and U2596 (N_2596,In_535,In_427);
and U2597 (N_2597,In_716,In_1165);
xnor U2598 (N_2598,In_1535,In_2281);
nor U2599 (N_2599,In_1392,In_944);
nand U2600 (N_2600,In_2117,In_1614);
or U2601 (N_2601,In_214,In_1105);
or U2602 (N_2602,In_1483,In_1661);
xnor U2603 (N_2603,In_2173,In_993);
nand U2604 (N_2604,In_747,In_1699);
xor U2605 (N_2605,In_171,In_1071);
nor U2606 (N_2606,In_1413,In_2008);
nand U2607 (N_2607,In_902,In_1818);
xnor U2608 (N_2608,In_2151,In_373);
and U2609 (N_2609,In_54,In_785);
nand U2610 (N_2610,In_562,In_1753);
or U2611 (N_2611,In_1825,In_977);
xnor U2612 (N_2612,In_1585,In_399);
and U2613 (N_2613,In_1982,In_1785);
or U2614 (N_2614,In_904,In_1793);
or U2615 (N_2615,In_758,In_1592);
nand U2616 (N_2616,In_667,In_2278);
nand U2617 (N_2617,In_1599,In_1069);
xnor U2618 (N_2618,In_2067,In_1848);
nor U2619 (N_2619,In_2077,In_671);
nand U2620 (N_2620,In_2175,In_968);
xor U2621 (N_2621,In_2430,In_1315);
xor U2622 (N_2622,In_2017,In_2151);
nand U2623 (N_2623,In_62,In_541);
nand U2624 (N_2624,In_1241,In_2189);
nor U2625 (N_2625,In_1792,In_1689);
nand U2626 (N_2626,In_1226,In_1030);
nor U2627 (N_2627,In_527,In_625);
nor U2628 (N_2628,In_1532,In_2242);
and U2629 (N_2629,In_1964,In_682);
nor U2630 (N_2630,In_465,In_2200);
or U2631 (N_2631,In_2063,In_99);
xor U2632 (N_2632,In_1824,In_2085);
and U2633 (N_2633,In_1695,In_574);
nor U2634 (N_2634,In_1213,In_1666);
xor U2635 (N_2635,In_1278,In_376);
or U2636 (N_2636,In_1796,In_2407);
and U2637 (N_2637,In_2189,In_1245);
nor U2638 (N_2638,In_2267,In_974);
xnor U2639 (N_2639,In_1678,In_505);
nand U2640 (N_2640,In_785,In_1021);
nor U2641 (N_2641,In_904,In_2227);
xnor U2642 (N_2642,In_1372,In_475);
xnor U2643 (N_2643,In_1377,In_1109);
nor U2644 (N_2644,In_719,In_2037);
nor U2645 (N_2645,In_2266,In_846);
xor U2646 (N_2646,In_2014,In_1273);
nand U2647 (N_2647,In_340,In_1735);
nand U2648 (N_2648,In_1482,In_1451);
and U2649 (N_2649,In_2113,In_256);
nor U2650 (N_2650,In_341,In_1963);
or U2651 (N_2651,In_1968,In_633);
xor U2652 (N_2652,In_1729,In_2299);
and U2653 (N_2653,In_234,In_1792);
nor U2654 (N_2654,In_857,In_117);
and U2655 (N_2655,In_1612,In_2467);
nor U2656 (N_2656,In_2174,In_235);
and U2657 (N_2657,In_1084,In_2381);
nand U2658 (N_2658,In_612,In_121);
nor U2659 (N_2659,In_861,In_1272);
and U2660 (N_2660,In_2286,In_1314);
nor U2661 (N_2661,In_1356,In_1515);
and U2662 (N_2662,In_1194,In_555);
xor U2663 (N_2663,In_1800,In_1886);
and U2664 (N_2664,In_1908,In_296);
nand U2665 (N_2665,In_2488,In_461);
or U2666 (N_2666,In_1934,In_1315);
or U2667 (N_2667,In_433,In_2355);
nand U2668 (N_2668,In_1841,In_1017);
and U2669 (N_2669,In_1452,In_704);
nand U2670 (N_2670,In_391,In_477);
or U2671 (N_2671,In_1799,In_662);
xor U2672 (N_2672,In_746,In_94);
nor U2673 (N_2673,In_384,In_2469);
xor U2674 (N_2674,In_1340,In_2442);
or U2675 (N_2675,In_1728,In_1690);
and U2676 (N_2676,In_2036,In_695);
nor U2677 (N_2677,In_2081,In_2023);
nand U2678 (N_2678,In_1950,In_1);
or U2679 (N_2679,In_1275,In_941);
or U2680 (N_2680,In_2010,In_505);
xnor U2681 (N_2681,In_126,In_2135);
or U2682 (N_2682,In_1038,In_1084);
xnor U2683 (N_2683,In_1274,In_533);
xnor U2684 (N_2684,In_78,In_224);
xor U2685 (N_2685,In_1424,In_973);
nor U2686 (N_2686,In_1903,In_2477);
nor U2687 (N_2687,In_2335,In_2253);
or U2688 (N_2688,In_1197,In_2009);
and U2689 (N_2689,In_1330,In_1652);
nand U2690 (N_2690,In_989,In_2481);
xor U2691 (N_2691,In_152,In_319);
xor U2692 (N_2692,In_1968,In_2186);
or U2693 (N_2693,In_341,In_1481);
or U2694 (N_2694,In_1613,In_1886);
and U2695 (N_2695,In_1883,In_928);
or U2696 (N_2696,In_2479,In_101);
or U2697 (N_2697,In_2213,In_1404);
xnor U2698 (N_2698,In_2351,In_1263);
xor U2699 (N_2699,In_1261,In_2229);
or U2700 (N_2700,In_894,In_2053);
xor U2701 (N_2701,In_352,In_2426);
and U2702 (N_2702,In_748,In_2468);
xnor U2703 (N_2703,In_1688,In_1859);
nand U2704 (N_2704,In_1999,In_1501);
nor U2705 (N_2705,In_1429,In_575);
xnor U2706 (N_2706,In_1380,In_1979);
or U2707 (N_2707,In_2287,In_105);
or U2708 (N_2708,In_1715,In_506);
and U2709 (N_2709,In_1518,In_1590);
or U2710 (N_2710,In_2480,In_279);
nor U2711 (N_2711,In_2292,In_882);
and U2712 (N_2712,In_165,In_607);
nor U2713 (N_2713,In_2380,In_2302);
nor U2714 (N_2714,In_2341,In_2064);
nor U2715 (N_2715,In_445,In_1327);
or U2716 (N_2716,In_2377,In_1867);
nand U2717 (N_2717,In_651,In_585);
xnor U2718 (N_2718,In_778,In_1174);
xor U2719 (N_2719,In_1392,In_2013);
nor U2720 (N_2720,In_435,In_1164);
or U2721 (N_2721,In_2151,In_2177);
xnor U2722 (N_2722,In_896,In_2109);
nand U2723 (N_2723,In_468,In_1190);
nor U2724 (N_2724,In_22,In_970);
or U2725 (N_2725,In_2014,In_785);
and U2726 (N_2726,In_627,In_1864);
nand U2727 (N_2727,In_806,In_2228);
or U2728 (N_2728,In_982,In_2026);
or U2729 (N_2729,In_2244,In_1159);
xnor U2730 (N_2730,In_193,In_928);
xor U2731 (N_2731,In_1670,In_104);
or U2732 (N_2732,In_1328,In_1845);
or U2733 (N_2733,In_963,In_429);
xnor U2734 (N_2734,In_1156,In_676);
nand U2735 (N_2735,In_1916,In_1974);
or U2736 (N_2736,In_1089,In_2326);
and U2737 (N_2737,In_43,In_2443);
and U2738 (N_2738,In_402,In_2249);
or U2739 (N_2739,In_456,In_160);
or U2740 (N_2740,In_1555,In_1217);
nor U2741 (N_2741,In_2189,In_1803);
nand U2742 (N_2742,In_1980,In_1676);
or U2743 (N_2743,In_2133,In_754);
nor U2744 (N_2744,In_1376,In_1700);
nor U2745 (N_2745,In_384,In_457);
or U2746 (N_2746,In_260,In_1562);
and U2747 (N_2747,In_585,In_1619);
and U2748 (N_2748,In_570,In_1246);
xor U2749 (N_2749,In_95,In_1339);
nor U2750 (N_2750,In_2069,In_489);
or U2751 (N_2751,In_1313,In_1092);
nand U2752 (N_2752,In_2482,In_1947);
or U2753 (N_2753,In_1567,In_323);
xor U2754 (N_2754,In_726,In_2066);
or U2755 (N_2755,In_2218,In_1951);
nor U2756 (N_2756,In_335,In_1267);
nand U2757 (N_2757,In_2021,In_524);
nor U2758 (N_2758,In_541,In_2498);
xnor U2759 (N_2759,In_992,In_702);
xnor U2760 (N_2760,In_1057,In_2022);
nor U2761 (N_2761,In_1803,In_865);
nand U2762 (N_2762,In_2195,In_2316);
or U2763 (N_2763,In_1375,In_2493);
and U2764 (N_2764,In_311,In_1383);
nor U2765 (N_2765,In_1245,In_2339);
xnor U2766 (N_2766,In_2185,In_1614);
or U2767 (N_2767,In_2165,In_2096);
nor U2768 (N_2768,In_2371,In_1815);
or U2769 (N_2769,In_276,In_1925);
or U2770 (N_2770,In_2343,In_561);
xor U2771 (N_2771,In_927,In_2051);
and U2772 (N_2772,In_1773,In_1250);
nor U2773 (N_2773,In_954,In_700);
or U2774 (N_2774,In_547,In_1109);
nor U2775 (N_2775,In_863,In_252);
or U2776 (N_2776,In_2323,In_1139);
nor U2777 (N_2777,In_440,In_2355);
and U2778 (N_2778,In_699,In_252);
nor U2779 (N_2779,In_1995,In_168);
xor U2780 (N_2780,In_373,In_1004);
xnor U2781 (N_2781,In_2169,In_958);
nor U2782 (N_2782,In_1292,In_1514);
xor U2783 (N_2783,In_1693,In_1181);
nand U2784 (N_2784,In_1477,In_199);
nor U2785 (N_2785,In_2025,In_1225);
xor U2786 (N_2786,In_721,In_72);
nand U2787 (N_2787,In_865,In_2328);
and U2788 (N_2788,In_2353,In_407);
xor U2789 (N_2789,In_1254,In_2032);
or U2790 (N_2790,In_282,In_2087);
xor U2791 (N_2791,In_60,In_2014);
nand U2792 (N_2792,In_524,In_1497);
nor U2793 (N_2793,In_262,In_1542);
nand U2794 (N_2794,In_2094,In_1090);
and U2795 (N_2795,In_541,In_238);
xnor U2796 (N_2796,In_1480,In_732);
xnor U2797 (N_2797,In_1194,In_1360);
xnor U2798 (N_2798,In_827,In_1798);
xor U2799 (N_2799,In_2112,In_2403);
xnor U2800 (N_2800,In_578,In_1521);
nand U2801 (N_2801,In_1228,In_933);
xor U2802 (N_2802,In_1028,In_364);
nand U2803 (N_2803,In_259,In_1861);
or U2804 (N_2804,In_2092,In_550);
xor U2805 (N_2805,In_774,In_1721);
xnor U2806 (N_2806,In_1343,In_1295);
xnor U2807 (N_2807,In_787,In_478);
or U2808 (N_2808,In_1980,In_488);
or U2809 (N_2809,In_158,In_2179);
and U2810 (N_2810,In_1363,In_1636);
nand U2811 (N_2811,In_1323,In_1575);
nand U2812 (N_2812,In_1722,In_25);
nand U2813 (N_2813,In_543,In_475);
nand U2814 (N_2814,In_1665,In_1709);
nor U2815 (N_2815,In_156,In_33);
and U2816 (N_2816,In_254,In_1471);
nor U2817 (N_2817,In_231,In_1410);
and U2818 (N_2818,In_2452,In_1252);
nor U2819 (N_2819,In_1478,In_1647);
or U2820 (N_2820,In_1762,In_1471);
or U2821 (N_2821,In_672,In_1407);
xnor U2822 (N_2822,In_1710,In_1671);
nand U2823 (N_2823,In_1019,In_36);
or U2824 (N_2824,In_1370,In_941);
and U2825 (N_2825,In_2387,In_554);
or U2826 (N_2826,In_744,In_138);
and U2827 (N_2827,In_1173,In_324);
and U2828 (N_2828,In_1963,In_178);
xnor U2829 (N_2829,In_352,In_1646);
nand U2830 (N_2830,In_509,In_503);
nand U2831 (N_2831,In_2001,In_1132);
nand U2832 (N_2832,In_486,In_1473);
and U2833 (N_2833,In_1589,In_105);
nand U2834 (N_2834,In_1529,In_2386);
nand U2835 (N_2835,In_798,In_2072);
nor U2836 (N_2836,In_209,In_910);
nand U2837 (N_2837,In_1466,In_801);
or U2838 (N_2838,In_1453,In_719);
xnor U2839 (N_2839,In_650,In_1);
nand U2840 (N_2840,In_1543,In_488);
nand U2841 (N_2841,In_1484,In_1790);
nand U2842 (N_2842,In_1822,In_217);
and U2843 (N_2843,In_645,In_1925);
xor U2844 (N_2844,In_2084,In_133);
and U2845 (N_2845,In_2128,In_21);
xor U2846 (N_2846,In_1211,In_1473);
nand U2847 (N_2847,In_2401,In_1388);
xnor U2848 (N_2848,In_110,In_2241);
nor U2849 (N_2849,In_2204,In_2005);
or U2850 (N_2850,In_2141,In_2146);
nand U2851 (N_2851,In_804,In_195);
or U2852 (N_2852,In_1108,In_1522);
or U2853 (N_2853,In_1264,In_2390);
or U2854 (N_2854,In_1682,In_1231);
and U2855 (N_2855,In_145,In_324);
nand U2856 (N_2856,In_2382,In_804);
nand U2857 (N_2857,In_2419,In_338);
nor U2858 (N_2858,In_2356,In_1350);
nand U2859 (N_2859,In_1636,In_1299);
nor U2860 (N_2860,In_1770,In_1715);
nand U2861 (N_2861,In_1417,In_1426);
nor U2862 (N_2862,In_2457,In_767);
nand U2863 (N_2863,In_1835,In_2396);
xnor U2864 (N_2864,In_1689,In_175);
xnor U2865 (N_2865,In_465,In_713);
or U2866 (N_2866,In_1649,In_1761);
and U2867 (N_2867,In_2498,In_1861);
xnor U2868 (N_2868,In_1713,In_1570);
nand U2869 (N_2869,In_691,In_160);
or U2870 (N_2870,In_105,In_323);
or U2871 (N_2871,In_902,In_284);
xnor U2872 (N_2872,In_1094,In_669);
or U2873 (N_2873,In_142,In_1441);
nor U2874 (N_2874,In_2280,In_1773);
and U2875 (N_2875,In_1796,In_2287);
and U2876 (N_2876,In_2384,In_2364);
or U2877 (N_2877,In_1739,In_12);
nand U2878 (N_2878,In_1401,In_1562);
or U2879 (N_2879,In_1157,In_72);
nand U2880 (N_2880,In_1126,In_870);
nor U2881 (N_2881,In_1320,In_2072);
and U2882 (N_2882,In_1952,In_363);
nand U2883 (N_2883,In_1214,In_1911);
nand U2884 (N_2884,In_1965,In_1374);
nor U2885 (N_2885,In_1386,In_1536);
and U2886 (N_2886,In_2027,In_1079);
nand U2887 (N_2887,In_636,In_1740);
nand U2888 (N_2888,In_78,In_1334);
nand U2889 (N_2889,In_2038,In_1461);
xor U2890 (N_2890,In_2121,In_360);
or U2891 (N_2891,In_2379,In_1060);
nor U2892 (N_2892,In_728,In_2405);
nand U2893 (N_2893,In_2052,In_649);
xor U2894 (N_2894,In_2413,In_854);
or U2895 (N_2895,In_293,In_750);
and U2896 (N_2896,In_425,In_1900);
and U2897 (N_2897,In_444,In_1207);
xor U2898 (N_2898,In_1352,In_1556);
xnor U2899 (N_2899,In_2058,In_1992);
xnor U2900 (N_2900,In_650,In_1195);
xor U2901 (N_2901,In_403,In_1361);
nor U2902 (N_2902,In_2331,In_305);
or U2903 (N_2903,In_197,In_1700);
nor U2904 (N_2904,In_2131,In_1670);
xnor U2905 (N_2905,In_1570,In_1925);
or U2906 (N_2906,In_2180,In_2183);
or U2907 (N_2907,In_74,In_403);
or U2908 (N_2908,In_1165,In_588);
or U2909 (N_2909,In_1445,In_2112);
and U2910 (N_2910,In_1683,In_1814);
xnor U2911 (N_2911,In_2023,In_1249);
and U2912 (N_2912,In_1437,In_2111);
nand U2913 (N_2913,In_653,In_1486);
xor U2914 (N_2914,In_1323,In_1420);
and U2915 (N_2915,In_2305,In_1006);
nor U2916 (N_2916,In_1462,In_2401);
xnor U2917 (N_2917,In_2468,In_244);
nand U2918 (N_2918,In_501,In_2343);
xnor U2919 (N_2919,In_1308,In_91);
xor U2920 (N_2920,In_848,In_655);
or U2921 (N_2921,In_822,In_1353);
nand U2922 (N_2922,In_1196,In_1096);
or U2923 (N_2923,In_1424,In_2349);
nor U2924 (N_2924,In_2282,In_1008);
or U2925 (N_2925,In_2444,In_249);
or U2926 (N_2926,In_179,In_730);
nand U2927 (N_2927,In_2085,In_1992);
xor U2928 (N_2928,In_1907,In_2313);
or U2929 (N_2929,In_2279,In_2313);
xnor U2930 (N_2930,In_1789,In_923);
nand U2931 (N_2931,In_426,In_1824);
xnor U2932 (N_2932,In_1180,In_475);
or U2933 (N_2933,In_859,In_1996);
nand U2934 (N_2934,In_1695,In_1353);
nor U2935 (N_2935,In_606,In_1067);
or U2936 (N_2936,In_2187,In_1206);
and U2937 (N_2937,In_1422,In_716);
or U2938 (N_2938,In_1421,In_2380);
nor U2939 (N_2939,In_1639,In_1594);
nor U2940 (N_2940,In_486,In_566);
xor U2941 (N_2941,In_1427,In_943);
xor U2942 (N_2942,In_131,In_1040);
and U2943 (N_2943,In_1462,In_796);
and U2944 (N_2944,In_2498,In_1554);
or U2945 (N_2945,In_173,In_1185);
nand U2946 (N_2946,In_2155,In_1354);
nor U2947 (N_2947,In_626,In_1886);
and U2948 (N_2948,In_92,In_1310);
nand U2949 (N_2949,In_714,In_1360);
nor U2950 (N_2950,In_693,In_1706);
nor U2951 (N_2951,In_1733,In_1822);
and U2952 (N_2952,In_542,In_936);
xnor U2953 (N_2953,In_839,In_1215);
nand U2954 (N_2954,In_619,In_674);
nor U2955 (N_2955,In_774,In_1131);
nor U2956 (N_2956,In_2117,In_2144);
nand U2957 (N_2957,In_2084,In_1863);
or U2958 (N_2958,In_2020,In_2164);
or U2959 (N_2959,In_212,In_898);
xor U2960 (N_2960,In_1473,In_1530);
xor U2961 (N_2961,In_283,In_1048);
or U2962 (N_2962,In_1317,In_2107);
xor U2963 (N_2963,In_1514,In_305);
and U2964 (N_2964,In_1732,In_451);
or U2965 (N_2965,In_691,In_2104);
xnor U2966 (N_2966,In_140,In_654);
nand U2967 (N_2967,In_1960,In_620);
and U2968 (N_2968,In_1983,In_2093);
nand U2969 (N_2969,In_9,In_1767);
xor U2970 (N_2970,In_1230,In_1873);
or U2971 (N_2971,In_625,In_792);
nand U2972 (N_2972,In_2481,In_1442);
or U2973 (N_2973,In_1271,In_27);
xor U2974 (N_2974,In_1659,In_1358);
nand U2975 (N_2975,In_2104,In_801);
and U2976 (N_2976,In_342,In_745);
xor U2977 (N_2977,In_39,In_798);
nand U2978 (N_2978,In_132,In_940);
xor U2979 (N_2979,In_869,In_1889);
and U2980 (N_2980,In_1684,In_793);
nand U2981 (N_2981,In_1645,In_752);
nor U2982 (N_2982,In_63,In_432);
nand U2983 (N_2983,In_1998,In_700);
or U2984 (N_2984,In_2322,In_1048);
and U2985 (N_2985,In_679,In_1903);
or U2986 (N_2986,In_868,In_2444);
xnor U2987 (N_2987,In_422,In_2465);
nor U2988 (N_2988,In_942,In_736);
nor U2989 (N_2989,In_2004,In_1303);
xor U2990 (N_2990,In_1881,In_2355);
and U2991 (N_2991,In_1098,In_256);
and U2992 (N_2992,In_2073,In_1761);
nor U2993 (N_2993,In_2163,In_1586);
and U2994 (N_2994,In_2230,In_1486);
or U2995 (N_2995,In_1930,In_546);
xnor U2996 (N_2996,In_300,In_380);
nor U2997 (N_2997,In_1428,In_2045);
nor U2998 (N_2998,In_312,In_983);
or U2999 (N_2999,In_2113,In_190);
or U3000 (N_3000,In_152,In_1385);
xnor U3001 (N_3001,In_410,In_324);
and U3002 (N_3002,In_715,In_1481);
or U3003 (N_3003,In_4,In_1768);
nand U3004 (N_3004,In_1322,In_1498);
nor U3005 (N_3005,In_515,In_419);
and U3006 (N_3006,In_782,In_1406);
nand U3007 (N_3007,In_2372,In_1089);
nor U3008 (N_3008,In_1413,In_1124);
nor U3009 (N_3009,In_971,In_138);
or U3010 (N_3010,In_289,In_2099);
xnor U3011 (N_3011,In_2490,In_1007);
or U3012 (N_3012,In_2428,In_1795);
xnor U3013 (N_3013,In_867,In_399);
and U3014 (N_3014,In_87,In_22);
nor U3015 (N_3015,In_1240,In_500);
and U3016 (N_3016,In_2495,In_286);
or U3017 (N_3017,In_1911,In_79);
or U3018 (N_3018,In_972,In_1268);
nand U3019 (N_3019,In_2434,In_265);
nor U3020 (N_3020,In_1455,In_2036);
nor U3021 (N_3021,In_1709,In_1568);
nand U3022 (N_3022,In_2246,In_2437);
nor U3023 (N_3023,In_286,In_502);
xnor U3024 (N_3024,In_445,In_779);
or U3025 (N_3025,In_2001,In_2009);
nor U3026 (N_3026,In_1939,In_378);
nand U3027 (N_3027,In_385,In_2266);
xor U3028 (N_3028,In_2423,In_1643);
nor U3029 (N_3029,In_1496,In_745);
xor U3030 (N_3030,In_196,In_2435);
nand U3031 (N_3031,In_353,In_918);
xor U3032 (N_3032,In_1271,In_218);
and U3033 (N_3033,In_1740,In_2073);
xor U3034 (N_3034,In_2362,In_1845);
and U3035 (N_3035,In_2142,In_520);
and U3036 (N_3036,In_1622,In_596);
nor U3037 (N_3037,In_897,In_26);
and U3038 (N_3038,In_583,In_2153);
xnor U3039 (N_3039,In_1865,In_671);
and U3040 (N_3040,In_1666,In_2256);
or U3041 (N_3041,In_638,In_2219);
and U3042 (N_3042,In_2135,In_907);
and U3043 (N_3043,In_896,In_902);
xor U3044 (N_3044,In_2218,In_99);
xor U3045 (N_3045,In_1074,In_1821);
and U3046 (N_3046,In_858,In_679);
and U3047 (N_3047,In_2423,In_67);
xnor U3048 (N_3048,In_1584,In_787);
xnor U3049 (N_3049,In_41,In_329);
or U3050 (N_3050,In_572,In_1865);
nor U3051 (N_3051,In_1145,In_726);
nor U3052 (N_3052,In_920,In_682);
nand U3053 (N_3053,In_763,In_563);
or U3054 (N_3054,In_361,In_2099);
nor U3055 (N_3055,In_1088,In_2131);
xnor U3056 (N_3056,In_1299,In_1324);
or U3057 (N_3057,In_858,In_1737);
nand U3058 (N_3058,In_1728,In_319);
xor U3059 (N_3059,In_711,In_1472);
nand U3060 (N_3060,In_1031,In_77);
or U3061 (N_3061,In_2234,In_2473);
and U3062 (N_3062,In_1449,In_637);
nand U3063 (N_3063,In_2055,In_1548);
xor U3064 (N_3064,In_2290,In_1206);
and U3065 (N_3065,In_2494,In_1363);
xor U3066 (N_3066,In_1733,In_1696);
or U3067 (N_3067,In_1700,In_87);
nand U3068 (N_3068,In_683,In_2316);
xor U3069 (N_3069,In_1153,In_1020);
or U3070 (N_3070,In_1506,In_2418);
nor U3071 (N_3071,In_289,In_495);
xor U3072 (N_3072,In_1285,In_94);
nand U3073 (N_3073,In_1068,In_2065);
nor U3074 (N_3074,In_409,In_2034);
and U3075 (N_3075,In_2497,In_2235);
or U3076 (N_3076,In_275,In_1350);
xor U3077 (N_3077,In_1062,In_1251);
nor U3078 (N_3078,In_800,In_1444);
and U3079 (N_3079,In_1996,In_789);
and U3080 (N_3080,In_538,In_2324);
nand U3081 (N_3081,In_931,In_787);
and U3082 (N_3082,In_484,In_1817);
nor U3083 (N_3083,In_2282,In_1367);
nor U3084 (N_3084,In_532,In_1488);
nor U3085 (N_3085,In_47,In_1570);
or U3086 (N_3086,In_1892,In_1923);
or U3087 (N_3087,In_249,In_1463);
or U3088 (N_3088,In_1384,In_2136);
xor U3089 (N_3089,In_2139,In_1223);
nand U3090 (N_3090,In_2211,In_2228);
or U3091 (N_3091,In_527,In_2471);
nand U3092 (N_3092,In_1733,In_1499);
or U3093 (N_3093,In_704,In_821);
nand U3094 (N_3094,In_2312,In_925);
nor U3095 (N_3095,In_678,In_211);
or U3096 (N_3096,In_486,In_1686);
and U3097 (N_3097,In_1655,In_2457);
nand U3098 (N_3098,In_2102,In_2);
xnor U3099 (N_3099,In_480,In_982);
nand U3100 (N_3100,In_734,In_1907);
xnor U3101 (N_3101,In_1555,In_1784);
nand U3102 (N_3102,In_807,In_398);
nand U3103 (N_3103,In_2196,In_463);
nor U3104 (N_3104,In_2149,In_372);
nor U3105 (N_3105,In_1258,In_700);
and U3106 (N_3106,In_1891,In_57);
nor U3107 (N_3107,In_2368,In_1889);
nor U3108 (N_3108,In_535,In_486);
xor U3109 (N_3109,In_2076,In_1200);
nand U3110 (N_3110,In_87,In_1316);
nor U3111 (N_3111,In_656,In_2082);
xnor U3112 (N_3112,In_2128,In_975);
nand U3113 (N_3113,In_1687,In_88);
or U3114 (N_3114,In_1136,In_1104);
and U3115 (N_3115,In_806,In_573);
and U3116 (N_3116,In_2150,In_1683);
nor U3117 (N_3117,In_158,In_2134);
nand U3118 (N_3118,In_2252,In_992);
and U3119 (N_3119,In_500,In_271);
xor U3120 (N_3120,In_1029,In_116);
or U3121 (N_3121,In_682,In_54);
nor U3122 (N_3122,In_1318,In_644);
xnor U3123 (N_3123,In_2339,In_503);
xnor U3124 (N_3124,In_822,In_770);
or U3125 (N_3125,In_1575,In_1497);
nor U3126 (N_3126,In_2268,In_640);
xnor U3127 (N_3127,In_20,In_2046);
xnor U3128 (N_3128,In_1844,In_2217);
or U3129 (N_3129,In_1699,In_2124);
nor U3130 (N_3130,In_1291,In_482);
nand U3131 (N_3131,In_1055,In_1214);
nand U3132 (N_3132,In_348,In_43);
nand U3133 (N_3133,In_1172,In_932);
xnor U3134 (N_3134,In_2441,In_2102);
xor U3135 (N_3135,In_2111,In_1866);
and U3136 (N_3136,In_2168,In_1369);
and U3137 (N_3137,In_1103,In_127);
xnor U3138 (N_3138,In_795,In_1033);
and U3139 (N_3139,In_1839,In_837);
nor U3140 (N_3140,In_258,In_2336);
nor U3141 (N_3141,In_1697,In_2088);
nor U3142 (N_3142,In_315,In_343);
or U3143 (N_3143,In_755,In_1214);
xor U3144 (N_3144,In_1178,In_2324);
xnor U3145 (N_3145,In_1171,In_979);
and U3146 (N_3146,In_563,In_1976);
nand U3147 (N_3147,In_1796,In_1728);
nor U3148 (N_3148,In_28,In_850);
or U3149 (N_3149,In_1716,In_2036);
nor U3150 (N_3150,In_785,In_1526);
xor U3151 (N_3151,In_1487,In_999);
and U3152 (N_3152,In_1850,In_2391);
nand U3153 (N_3153,In_815,In_439);
xnor U3154 (N_3154,In_2006,In_211);
nor U3155 (N_3155,In_769,In_1545);
or U3156 (N_3156,In_1040,In_2417);
nor U3157 (N_3157,In_1360,In_449);
or U3158 (N_3158,In_2410,In_399);
nand U3159 (N_3159,In_836,In_1569);
xor U3160 (N_3160,In_843,In_777);
xor U3161 (N_3161,In_1683,In_1435);
or U3162 (N_3162,In_645,In_339);
or U3163 (N_3163,In_1196,In_1545);
and U3164 (N_3164,In_1203,In_2486);
and U3165 (N_3165,In_1770,In_351);
and U3166 (N_3166,In_913,In_1001);
xnor U3167 (N_3167,In_574,In_1024);
xnor U3168 (N_3168,In_1741,In_393);
or U3169 (N_3169,In_2160,In_2002);
nor U3170 (N_3170,In_1727,In_1033);
and U3171 (N_3171,In_927,In_1342);
nor U3172 (N_3172,In_1487,In_803);
nand U3173 (N_3173,In_1523,In_87);
xnor U3174 (N_3174,In_1935,In_2054);
nor U3175 (N_3175,In_1381,In_1874);
nor U3176 (N_3176,In_1069,In_2120);
or U3177 (N_3177,In_1824,In_2248);
nor U3178 (N_3178,In_543,In_2387);
nor U3179 (N_3179,In_2089,In_466);
and U3180 (N_3180,In_912,In_132);
or U3181 (N_3181,In_1694,In_2074);
nand U3182 (N_3182,In_1591,In_1379);
nand U3183 (N_3183,In_584,In_1026);
and U3184 (N_3184,In_1369,In_707);
or U3185 (N_3185,In_2368,In_422);
or U3186 (N_3186,In_538,In_54);
xnor U3187 (N_3187,In_794,In_117);
nor U3188 (N_3188,In_536,In_761);
nor U3189 (N_3189,In_2378,In_1888);
or U3190 (N_3190,In_248,In_531);
and U3191 (N_3191,In_1702,In_1589);
or U3192 (N_3192,In_1774,In_2163);
or U3193 (N_3193,In_1659,In_1168);
nor U3194 (N_3194,In_440,In_510);
xor U3195 (N_3195,In_2384,In_1447);
nor U3196 (N_3196,In_1769,In_1593);
nor U3197 (N_3197,In_105,In_413);
nor U3198 (N_3198,In_1826,In_586);
xnor U3199 (N_3199,In_994,In_2141);
xnor U3200 (N_3200,In_770,In_1240);
xnor U3201 (N_3201,In_2376,In_1922);
nand U3202 (N_3202,In_227,In_1046);
nor U3203 (N_3203,In_1599,In_1171);
and U3204 (N_3204,In_1487,In_965);
or U3205 (N_3205,In_2129,In_364);
nor U3206 (N_3206,In_773,In_2307);
nand U3207 (N_3207,In_253,In_2117);
nand U3208 (N_3208,In_2239,In_550);
nand U3209 (N_3209,In_2455,In_2095);
xnor U3210 (N_3210,In_1133,In_1577);
nor U3211 (N_3211,In_1327,In_1921);
nor U3212 (N_3212,In_585,In_1579);
nand U3213 (N_3213,In_2193,In_1161);
nand U3214 (N_3214,In_1558,In_1083);
xnor U3215 (N_3215,In_446,In_781);
and U3216 (N_3216,In_123,In_1191);
nand U3217 (N_3217,In_508,In_2241);
and U3218 (N_3218,In_40,In_1630);
nand U3219 (N_3219,In_729,In_2191);
nand U3220 (N_3220,In_2354,In_1584);
xor U3221 (N_3221,In_964,In_571);
or U3222 (N_3222,In_653,In_1456);
xnor U3223 (N_3223,In_908,In_88);
nand U3224 (N_3224,In_566,In_180);
and U3225 (N_3225,In_979,In_164);
nor U3226 (N_3226,In_587,In_2135);
and U3227 (N_3227,In_2095,In_814);
nor U3228 (N_3228,In_2405,In_2433);
and U3229 (N_3229,In_2443,In_693);
nor U3230 (N_3230,In_13,In_28);
nand U3231 (N_3231,In_1968,In_2409);
and U3232 (N_3232,In_971,In_540);
and U3233 (N_3233,In_2310,In_2067);
or U3234 (N_3234,In_658,In_1108);
or U3235 (N_3235,In_1752,In_2198);
or U3236 (N_3236,In_1560,In_380);
nor U3237 (N_3237,In_62,In_955);
nand U3238 (N_3238,In_338,In_195);
nor U3239 (N_3239,In_338,In_1070);
xor U3240 (N_3240,In_611,In_2455);
or U3241 (N_3241,In_170,In_2207);
xnor U3242 (N_3242,In_1622,In_629);
nand U3243 (N_3243,In_1946,In_2120);
nor U3244 (N_3244,In_349,In_1746);
nand U3245 (N_3245,In_146,In_1250);
xor U3246 (N_3246,In_427,In_1096);
and U3247 (N_3247,In_2480,In_1834);
or U3248 (N_3248,In_2453,In_539);
or U3249 (N_3249,In_651,In_969);
nor U3250 (N_3250,In_1047,In_1169);
nor U3251 (N_3251,In_2326,In_102);
and U3252 (N_3252,In_986,In_1142);
nor U3253 (N_3253,In_654,In_398);
xnor U3254 (N_3254,In_2040,In_269);
or U3255 (N_3255,In_392,In_2180);
nand U3256 (N_3256,In_1197,In_103);
and U3257 (N_3257,In_204,In_1340);
nand U3258 (N_3258,In_1784,In_1262);
and U3259 (N_3259,In_983,In_616);
xnor U3260 (N_3260,In_1749,In_1074);
or U3261 (N_3261,In_1461,In_1405);
nand U3262 (N_3262,In_137,In_966);
xor U3263 (N_3263,In_1317,In_1331);
and U3264 (N_3264,In_160,In_1293);
nor U3265 (N_3265,In_1662,In_940);
xnor U3266 (N_3266,In_1381,In_1188);
nor U3267 (N_3267,In_553,In_503);
or U3268 (N_3268,In_1857,In_57);
xor U3269 (N_3269,In_1360,In_2056);
and U3270 (N_3270,In_1376,In_554);
and U3271 (N_3271,In_1230,In_1141);
or U3272 (N_3272,In_826,In_477);
and U3273 (N_3273,In_2135,In_2024);
nor U3274 (N_3274,In_1460,In_749);
nand U3275 (N_3275,In_521,In_183);
and U3276 (N_3276,In_1747,In_1479);
and U3277 (N_3277,In_1798,In_2295);
nand U3278 (N_3278,In_269,In_1127);
nor U3279 (N_3279,In_2118,In_2272);
nor U3280 (N_3280,In_1067,In_795);
and U3281 (N_3281,In_1362,In_1404);
nor U3282 (N_3282,In_1538,In_616);
or U3283 (N_3283,In_251,In_523);
and U3284 (N_3284,In_2471,In_1967);
nor U3285 (N_3285,In_1473,In_980);
or U3286 (N_3286,In_2083,In_1399);
nor U3287 (N_3287,In_17,In_2032);
and U3288 (N_3288,In_2292,In_619);
and U3289 (N_3289,In_974,In_1964);
or U3290 (N_3290,In_2041,In_226);
or U3291 (N_3291,In_2270,In_372);
nand U3292 (N_3292,In_481,In_2269);
nand U3293 (N_3293,In_2301,In_1700);
and U3294 (N_3294,In_2257,In_374);
and U3295 (N_3295,In_2296,In_1199);
nand U3296 (N_3296,In_2178,In_1730);
and U3297 (N_3297,In_2093,In_1489);
nor U3298 (N_3298,In_926,In_1304);
nand U3299 (N_3299,In_91,In_291);
xor U3300 (N_3300,In_862,In_900);
and U3301 (N_3301,In_374,In_39);
and U3302 (N_3302,In_817,In_1756);
or U3303 (N_3303,In_2230,In_1265);
nor U3304 (N_3304,In_1372,In_2465);
or U3305 (N_3305,In_1173,In_442);
nand U3306 (N_3306,In_471,In_293);
and U3307 (N_3307,In_1964,In_1700);
nand U3308 (N_3308,In_775,In_635);
nor U3309 (N_3309,In_869,In_575);
and U3310 (N_3310,In_2258,In_1106);
or U3311 (N_3311,In_1110,In_1155);
and U3312 (N_3312,In_1789,In_101);
nand U3313 (N_3313,In_404,In_1859);
xnor U3314 (N_3314,In_134,In_2406);
nor U3315 (N_3315,In_1996,In_1243);
and U3316 (N_3316,In_1895,In_1678);
xor U3317 (N_3317,In_1418,In_630);
xor U3318 (N_3318,In_533,In_449);
nor U3319 (N_3319,In_1403,In_2466);
or U3320 (N_3320,In_2069,In_2475);
or U3321 (N_3321,In_432,In_1819);
nor U3322 (N_3322,In_1177,In_315);
nand U3323 (N_3323,In_2295,In_1979);
nand U3324 (N_3324,In_923,In_438);
xnor U3325 (N_3325,In_167,In_1115);
or U3326 (N_3326,In_2389,In_958);
or U3327 (N_3327,In_2292,In_547);
xnor U3328 (N_3328,In_1149,In_146);
nand U3329 (N_3329,In_828,In_811);
or U3330 (N_3330,In_2206,In_672);
xnor U3331 (N_3331,In_982,In_1684);
or U3332 (N_3332,In_546,In_2359);
nand U3333 (N_3333,In_179,In_947);
and U3334 (N_3334,In_2316,In_1535);
nor U3335 (N_3335,In_1679,In_2305);
xnor U3336 (N_3336,In_101,In_1888);
nor U3337 (N_3337,In_2036,In_1968);
nand U3338 (N_3338,In_1077,In_631);
nand U3339 (N_3339,In_307,In_900);
nor U3340 (N_3340,In_1954,In_1482);
nor U3341 (N_3341,In_1681,In_2050);
xor U3342 (N_3342,In_867,In_648);
or U3343 (N_3343,In_1868,In_1593);
or U3344 (N_3344,In_1608,In_2303);
xnor U3345 (N_3345,In_896,In_1852);
or U3346 (N_3346,In_1318,In_1043);
nand U3347 (N_3347,In_434,In_1609);
nand U3348 (N_3348,In_767,In_1471);
nor U3349 (N_3349,In_1836,In_661);
or U3350 (N_3350,In_479,In_1875);
or U3351 (N_3351,In_504,In_2052);
nor U3352 (N_3352,In_1545,In_911);
or U3353 (N_3353,In_506,In_782);
nand U3354 (N_3354,In_1135,In_25);
nor U3355 (N_3355,In_1942,In_60);
nand U3356 (N_3356,In_1988,In_1196);
nand U3357 (N_3357,In_2108,In_1080);
and U3358 (N_3358,In_2061,In_1172);
xor U3359 (N_3359,In_152,In_468);
nand U3360 (N_3360,In_48,In_201);
or U3361 (N_3361,In_2486,In_927);
nand U3362 (N_3362,In_1276,In_270);
and U3363 (N_3363,In_297,In_2458);
nand U3364 (N_3364,In_1330,In_1294);
or U3365 (N_3365,In_405,In_2285);
xnor U3366 (N_3366,In_1978,In_1348);
and U3367 (N_3367,In_1649,In_1964);
and U3368 (N_3368,In_525,In_984);
and U3369 (N_3369,In_334,In_1027);
nor U3370 (N_3370,In_2324,In_2119);
nand U3371 (N_3371,In_1076,In_246);
nand U3372 (N_3372,In_270,In_605);
or U3373 (N_3373,In_2042,In_2252);
and U3374 (N_3374,In_2116,In_1039);
nand U3375 (N_3375,In_291,In_2431);
nand U3376 (N_3376,In_571,In_25);
xor U3377 (N_3377,In_412,In_456);
nor U3378 (N_3378,In_2085,In_1175);
nand U3379 (N_3379,In_775,In_356);
nand U3380 (N_3380,In_1073,In_1766);
nor U3381 (N_3381,In_2208,In_2091);
or U3382 (N_3382,In_1252,In_2108);
xor U3383 (N_3383,In_926,In_1779);
nand U3384 (N_3384,In_2264,In_1493);
nand U3385 (N_3385,In_1535,In_2303);
xnor U3386 (N_3386,In_1206,In_1880);
xor U3387 (N_3387,In_1849,In_214);
or U3388 (N_3388,In_1986,In_1394);
nand U3389 (N_3389,In_473,In_2251);
xor U3390 (N_3390,In_510,In_1227);
and U3391 (N_3391,In_1924,In_96);
and U3392 (N_3392,In_1080,In_2416);
and U3393 (N_3393,In_436,In_285);
nand U3394 (N_3394,In_510,In_1096);
nor U3395 (N_3395,In_1818,In_484);
nor U3396 (N_3396,In_2400,In_1115);
nor U3397 (N_3397,In_787,In_1065);
nor U3398 (N_3398,In_1595,In_1233);
or U3399 (N_3399,In_1848,In_50);
nand U3400 (N_3400,In_845,In_274);
and U3401 (N_3401,In_1660,In_1421);
nand U3402 (N_3402,In_2118,In_2353);
and U3403 (N_3403,In_905,In_851);
nor U3404 (N_3404,In_1255,In_2408);
nor U3405 (N_3405,In_1690,In_979);
nand U3406 (N_3406,In_2144,In_1627);
and U3407 (N_3407,In_2429,In_218);
or U3408 (N_3408,In_270,In_1086);
and U3409 (N_3409,In_1025,In_5);
xnor U3410 (N_3410,In_1033,In_1447);
and U3411 (N_3411,In_2183,In_1437);
xor U3412 (N_3412,In_1582,In_2451);
or U3413 (N_3413,In_1349,In_561);
nand U3414 (N_3414,In_1665,In_1162);
or U3415 (N_3415,In_2423,In_655);
and U3416 (N_3416,In_723,In_1069);
nand U3417 (N_3417,In_1666,In_563);
nand U3418 (N_3418,In_374,In_1922);
nand U3419 (N_3419,In_1858,In_1910);
or U3420 (N_3420,In_913,In_1338);
nor U3421 (N_3421,In_1212,In_2228);
and U3422 (N_3422,In_1923,In_1153);
nor U3423 (N_3423,In_557,In_1568);
or U3424 (N_3424,In_469,In_2438);
or U3425 (N_3425,In_597,In_1902);
and U3426 (N_3426,In_50,In_2218);
xor U3427 (N_3427,In_479,In_691);
xor U3428 (N_3428,In_2082,In_819);
and U3429 (N_3429,In_573,In_1477);
nand U3430 (N_3430,In_1618,In_728);
nand U3431 (N_3431,In_1130,In_2147);
nor U3432 (N_3432,In_85,In_1740);
and U3433 (N_3433,In_1673,In_2307);
nor U3434 (N_3434,In_1000,In_81);
nor U3435 (N_3435,In_389,In_435);
and U3436 (N_3436,In_1875,In_1614);
or U3437 (N_3437,In_699,In_308);
or U3438 (N_3438,In_416,In_1533);
nor U3439 (N_3439,In_524,In_950);
xnor U3440 (N_3440,In_1283,In_1325);
xor U3441 (N_3441,In_1598,In_1863);
nor U3442 (N_3442,In_1100,In_1219);
and U3443 (N_3443,In_882,In_1402);
nor U3444 (N_3444,In_1922,In_2352);
nor U3445 (N_3445,In_766,In_1145);
or U3446 (N_3446,In_826,In_1541);
nor U3447 (N_3447,In_598,In_889);
nor U3448 (N_3448,In_765,In_451);
or U3449 (N_3449,In_1342,In_63);
or U3450 (N_3450,In_214,In_2010);
or U3451 (N_3451,In_1873,In_2071);
or U3452 (N_3452,In_689,In_1672);
nor U3453 (N_3453,In_1139,In_1216);
nand U3454 (N_3454,In_1938,In_2020);
nor U3455 (N_3455,In_1783,In_2375);
or U3456 (N_3456,In_1754,In_1122);
nand U3457 (N_3457,In_2195,In_1922);
xor U3458 (N_3458,In_1068,In_981);
xnor U3459 (N_3459,In_708,In_2493);
and U3460 (N_3460,In_1782,In_1454);
and U3461 (N_3461,In_1987,In_682);
and U3462 (N_3462,In_642,In_1808);
nand U3463 (N_3463,In_126,In_2266);
xnor U3464 (N_3464,In_1365,In_164);
nor U3465 (N_3465,In_2168,In_954);
xor U3466 (N_3466,In_1362,In_1014);
nor U3467 (N_3467,In_463,In_1877);
and U3468 (N_3468,In_848,In_109);
and U3469 (N_3469,In_785,In_1835);
nand U3470 (N_3470,In_1942,In_34);
nor U3471 (N_3471,In_91,In_188);
nor U3472 (N_3472,In_2033,In_1620);
nor U3473 (N_3473,In_1666,In_558);
xor U3474 (N_3474,In_842,In_963);
nand U3475 (N_3475,In_861,In_1023);
nor U3476 (N_3476,In_976,In_370);
and U3477 (N_3477,In_315,In_899);
nor U3478 (N_3478,In_238,In_65);
nor U3479 (N_3479,In_1226,In_336);
nor U3480 (N_3480,In_1902,In_332);
xnor U3481 (N_3481,In_65,In_1094);
nor U3482 (N_3482,In_1091,In_1380);
or U3483 (N_3483,In_953,In_388);
nor U3484 (N_3484,In_1527,In_1030);
and U3485 (N_3485,In_1297,In_462);
xor U3486 (N_3486,In_1993,In_366);
nor U3487 (N_3487,In_1059,In_657);
nor U3488 (N_3488,In_349,In_1030);
and U3489 (N_3489,In_1351,In_457);
and U3490 (N_3490,In_1879,In_1398);
nor U3491 (N_3491,In_1673,In_2134);
xor U3492 (N_3492,In_365,In_337);
nor U3493 (N_3493,In_401,In_1342);
xnor U3494 (N_3494,In_556,In_1412);
nand U3495 (N_3495,In_462,In_945);
nor U3496 (N_3496,In_2311,In_1949);
and U3497 (N_3497,In_326,In_2407);
and U3498 (N_3498,In_835,In_1065);
nand U3499 (N_3499,In_1593,In_298);
nor U3500 (N_3500,In_1639,In_1358);
xnor U3501 (N_3501,In_864,In_1492);
nand U3502 (N_3502,In_1170,In_1439);
nor U3503 (N_3503,In_2466,In_1016);
nand U3504 (N_3504,In_541,In_71);
and U3505 (N_3505,In_2468,In_638);
nand U3506 (N_3506,In_1828,In_609);
or U3507 (N_3507,In_402,In_1125);
nor U3508 (N_3508,In_885,In_2447);
or U3509 (N_3509,In_850,In_1357);
xnor U3510 (N_3510,In_2043,In_1291);
and U3511 (N_3511,In_1415,In_2463);
or U3512 (N_3512,In_1347,In_1786);
xor U3513 (N_3513,In_769,In_484);
nand U3514 (N_3514,In_1628,In_2373);
nand U3515 (N_3515,In_1733,In_1019);
and U3516 (N_3516,In_1055,In_815);
xor U3517 (N_3517,In_2447,In_319);
nand U3518 (N_3518,In_299,In_1228);
and U3519 (N_3519,In_1534,In_1061);
xnor U3520 (N_3520,In_1804,In_1960);
nand U3521 (N_3521,In_1750,In_2472);
nand U3522 (N_3522,In_2128,In_814);
xnor U3523 (N_3523,In_915,In_2143);
nor U3524 (N_3524,In_978,In_1057);
nor U3525 (N_3525,In_1249,In_1431);
xor U3526 (N_3526,In_1565,In_1062);
or U3527 (N_3527,In_290,In_37);
xor U3528 (N_3528,In_1672,In_1928);
or U3529 (N_3529,In_826,In_2131);
nor U3530 (N_3530,In_16,In_1036);
nor U3531 (N_3531,In_1570,In_659);
nand U3532 (N_3532,In_701,In_972);
nand U3533 (N_3533,In_1710,In_1879);
nand U3534 (N_3534,In_936,In_371);
or U3535 (N_3535,In_2090,In_2050);
or U3536 (N_3536,In_2330,In_1713);
and U3537 (N_3537,In_1688,In_982);
and U3538 (N_3538,In_276,In_976);
or U3539 (N_3539,In_1788,In_650);
nor U3540 (N_3540,In_1250,In_2017);
nor U3541 (N_3541,In_705,In_103);
and U3542 (N_3542,In_1480,In_395);
or U3543 (N_3543,In_2137,In_418);
nand U3544 (N_3544,In_1118,In_2167);
and U3545 (N_3545,In_1037,In_2348);
or U3546 (N_3546,In_2496,In_1093);
and U3547 (N_3547,In_2496,In_1951);
nor U3548 (N_3548,In_1190,In_1245);
nor U3549 (N_3549,In_412,In_1448);
and U3550 (N_3550,In_173,In_1959);
nand U3551 (N_3551,In_273,In_841);
xor U3552 (N_3552,In_2164,In_2442);
or U3553 (N_3553,In_2011,In_1352);
nor U3554 (N_3554,In_607,In_1653);
xor U3555 (N_3555,In_321,In_1985);
and U3556 (N_3556,In_2317,In_1077);
or U3557 (N_3557,In_2199,In_1393);
or U3558 (N_3558,In_1999,In_466);
or U3559 (N_3559,In_379,In_769);
and U3560 (N_3560,In_1885,In_182);
and U3561 (N_3561,In_1156,In_1567);
xor U3562 (N_3562,In_919,In_243);
xnor U3563 (N_3563,In_1912,In_2128);
nand U3564 (N_3564,In_1424,In_1453);
or U3565 (N_3565,In_1831,In_1869);
or U3566 (N_3566,In_885,In_1466);
nor U3567 (N_3567,In_464,In_1942);
xor U3568 (N_3568,In_296,In_1025);
or U3569 (N_3569,In_789,In_452);
and U3570 (N_3570,In_2454,In_1923);
or U3571 (N_3571,In_1158,In_1885);
nor U3572 (N_3572,In_359,In_1142);
nand U3573 (N_3573,In_1230,In_1353);
or U3574 (N_3574,In_1012,In_191);
nor U3575 (N_3575,In_1703,In_2358);
nor U3576 (N_3576,In_1325,In_2217);
nand U3577 (N_3577,In_876,In_1769);
or U3578 (N_3578,In_675,In_638);
nand U3579 (N_3579,In_1420,In_463);
nor U3580 (N_3580,In_1645,In_918);
nand U3581 (N_3581,In_1797,In_531);
xnor U3582 (N_3582,In_970,In_2495);
nand U3583 (N_3583,In_1444,In_825);
nor U3584 (N_3584,In_1271,In_155);
nor U3585 (N_3585,In_2047,In_1057);
nand U3586 (N_3586,In_1195,In_1271);
nor U3587 (N_3587,In_1956,In_65);
or U3588 (N_3588,In_1849,In_1529);
nand U3589 (N_3589,In_1438,In_1686);
and U3590 (N_3590,In_1018,In_4);
and U3591 (N_3591,In_1490,In_1168);
nand U3592 (N_3592,In_2180,In_59);
and U3593 (N_3593,In_149,In_1256);
and U3594 (N_3594,In_1212,In_1976);
nand U3595 (N_3595,In_1757,In_2288);
or U3596 (N_3596,In_1221,In_1800);
or U3597 (N_3597,In_138,In_1039);
nand U3598 (N_3598,In_764,In_1471);
nor U3599 (N_3599,In_547,In_630);
nor U3600 (N_3600,In_1530,In_477);
nor U3601 (N_3601,In_553,In_1360);
or U3602 (N_3602,In_1151,In_1395);
xnor U3603 (N_3603,In_225,In_2277);
or U3604 (N_3604,In_795,In_2012);
nor U3605 (N_3605,In_1685,In_1865);
nand U3606 (N_3606,In_597,In_2412);
nor U3607 (N_3607,In_62,In_1344);
nand U3608 (N_3608,In_770,In_1378);
and U3609 (N_3609,In_1598,In_1595);
or U3610 (N_3610,In_1416,In_1144);
xor U3611 (N_3611,In_1901,In_2412);
and U3612 (N_3612,In_687,In_61);
nor U3613 (N_3613,In_486,In_1088);
or U3614 (N_3614,In_1210,In_1131);
nor U3615 (N_3615,In_274,In_2197);
or U3616 (N_3616,In_1838,In_973);
and U3617 (N_3617,In_2482,In_2273);
xor U3618 (N_3618,In_2299,In_201);
and U3619 (N_3619,In_2131,In_2206);
nand U3620 (N_3620,In_1188,In_418);
xor U3621 (N_3621,In_2253,In_2452);
nor U3622 (N_3622,In_1116,In_630);
and U3623 (N_3623,In_1303,In_1111);
xor U3624 (N_3624,In_598,In_300);
xnor U3625 (N_3625,In_2239,In_625);
and U3626 (N_3626,In_830,In_1554);
or U3627 (N_3627,In_622,In_276);
xnor U3628 (N_3628,In_1207,In_1275);
nor U3629 (N_3629,In_0,In_1428);
nand U3630 (N_3630,In_603,In_1155);
nand U3631 (N_3631,In_444,In_1355);
xor U3632 (N_3632,In_816,In_2169);
xor U3633 (N_3633,In_312,In_805);
nand U3634 (N_3634,In_1189,In_1441);
nand U3635 (N_3635,In_1280,In_1775);
and U3636 (N_3636,In_434,In_1130);
and U3637 (N_3637,In_203,In_119);
nor U3638 (N_3638,In_95,In_1698);
xnor U3639 (N_3639,In_2043,In_1944);
or U3640 (N_3640,In_349,In_1590);
or U3641 (N_3641,In_1823,In_2214);
xor U3642 (N_3642,In_1,In_2125);
or U3643 (N_3643,In_1529,In_1667);
and U3644 (N_3644,In_773,In_1966);
or U3645 (N_3645,In_1867,In_2005);
xnor U3646 (N_3646,In_1817,In_1553);
and U3647 (N_3647,In_1292,In_529);
nand U3648 (N_3648,In_2361,In_910);
nor U3649 (N_3649,In_2395,In_1989);
nor U3650 (N_3650,In_2097,In_2131);
or U3651 (N_3651,In_1867,In_1482);
or U3652 (N_3652,In_2203,In_1377);
xor U3653 (N_3653,In_1514,In_2427);
and U3654 (N_3654,In_1780,In_99);
and U3655 (N_3655,In_529,In_2105);
nand U3656 (N_3656,In_20,In_1087);
or U3657 (N_3657,In_1361,In_1694);
or U3658 (N_3658,In_787,In_232);
nor U3659 (N_3659,In_152,In_1950);
nor U3660 (N_3660,In_1771,In_729);
nor U3661 (N_3661,In_1731,In_726);
and U3662 (N_3662,In_1527,In_176);
xor U3663 (N_3663,In_1336,In_179);
nand U3664 (N_3664,In_2279,In_68);
nor U3665 (N_3665,In_2082,In_1258);
nand U3666 (N_3666,In_2455,In_485);
nor U3667 (N_3667,In_2493,In_1348);
and U3668 (N_3668,In_331,In_57);
xnor U3669 (N_3669,In_742,In_1246);
and U3670 (N_3670,In_146,In_652);
and U3671 (N_3671,In_2373,In_1033);
nand U3672 (N_3672,In_661,In_2418);
and U3673 (N_3673,In_1950,In_1147);
or U3674 (N_3674,In_1615,In_486);
or U3675 (N_3675,In_2376,In_1352);
nor U3676 (N_3676,In_1818,In_1176);
nand U3677 (N_3677,In_1727,In_2346);
xnor U3678 (N_3678,In_2355,In_1369);
nor U3679 (N_3679,In_500,In_65);
or U3680 (N_3680,In_1787,In_1716);
nor U3681 (N_3681,In_232,In_2489);
nand U3682 (N_3682,In_303,In_1673);
xnor U3683 (N_3683,In_939,In_874);
and U3684 (N_3684,In_1732,In_1872);
xnor U3685 (N_3685,In_111,In_2116);
and U3686 (N_3686,In_2193,In_2159);
xor U3687 (N_3687,In_1987,In_1825);
and U3688 (N_3688,In_1036,In_886);
nor U3689 (N_3689,In_1661,In_2291);
nor U3690 (N_3690,In_109,In_179);
nand U3691 (N_3691,In_1826,In_1218);
nor U3692 (N_3692,In_100,In_1192);
or U3693 (N_3693,In_1495,In_2055);
nor U3694 (N_3694,In_1686,In_1197);
or U3695 (N_3695,In_70,In_607);
or U3696 (N_3696,In_147,In_793);
nor U3697 (N_3697,In_2462,In_814);
xnor U3698 (N_3698,In_1735,In_98);
xnor U3699 (N_3699,In_1954,In_391);
or U3700 (N_3700,In_2127,In_29);
xnor U3701 (N_3701,In_1186,In_617);
nand U3702 (N_3702,In_2312,In_297);
xnor U3703 (N_3703,In_42,In_166);
and U3704 (N_3704,In_923,In_1988);
xnor U3705 (N_3705,In_967,In_680);
nand U3706 (N_3706,In_2336,In_898);
nor U3707 (N_3707,In_749,In_172);
nor U3708 (N_3708,In_543,In_2358);
and U3709 (N_3709,In_167,In_1232);
nand U3710 (N_3710,In_95,In_862);
and U3711 (N_3711,In_1684,In_335);
and U3712 (N_3712,In_434,In_657);
or U3713 (N_3713,In_1307,In_2134);
xnor U3714 (N_3714,In_4,In_1121);
xor U3715 (N_3715,In_917,In_97);
nand U3716 (N_3716,In_437,In_507);
nand U3717 (N_3717,In_2148,In_1774);
and U3718 (N_3718,In_2205,In_1557);
nor U3719 (N_3719,In_399,In_1257);
nor U3720 (N_3720,In_882,In_2294);
xor U3721 (N_3721,In_601,In_1050);
or U3722 (N_3722,In_1561,In_1231);
xor U3723 (N_3723,In_1477,In_1631);
nand U3724 (N_3724,In_1211,In_183);
nor U3725 (N_3725,In_2376,In_1978);
nand U3726 (N_3726,In_1910,In_431);
nand U3727 (N_3727,In_1278,In_1107);
and U3728 (N_3728,In_2124,In_333);
and U3729 (N_3729,In_1561,In_1085);
nor U3730 (N_3730,In_359,In_1624);
nor U3731 (N_3731,In_1624,In_862);
nand U3732 (N_3732,In_1413,In_2466);
and U3733 (N_3733,In_1276,In_293);
xnor U3734 (N_3734,In_2232,In_25);
and U3735 (N_3735,In_1913,In_1029);
and U3736 (N_3736,In_1506,In_1918);
xor U3737 (N_3737,In_249,In_2392);
nor U3738 (N_3738,In_573,In_112);
xor U3739 (N_3739,In_2008,In_416);
or U3740 (N_3740,In_1059,In_2269);
and U3741 (N_3741,In_1511,In_1816);
nand U3742 (N_3742,In_37,In_1137);
and U3743 (N_3743,In_1450,In_16);
xnor U3744 (N_3744,In_1412,In_1197);
nor U3745 (N_3745,In_1488,In_1934);
nor U3746 (N_3746,In_1205,In_1335);
nor U3747 (N_3747,In_1621,In_845);
nand U3748 (N_3748,In_26,In_838);
or U3749 (N_3749,In_1746,In_764);
nor U3750 (N_3750,In_335,In_1423);
xnor U3751 (N_3751,In_1776,In_432);
or U3752 (N_3752,In_1630,In_414);
or U3753 (N_3753,In_1342,In_337);
nor U3754 (N_3754,In_2153,In_509);
and U3755 (N_3755,In_2400,In_2004);
and U3756 (N_3756,In_130,In_1375);
nand U3757 (N_3757,In_1385,In_2381);
xnor U3758 (N_3758,In_1239,In_2418);
and U3759 (N_3759,In_723,In_2299);
or U3760 (N_3760,In_860,In_491);
nand U3761 (N_3761,In_2163,In_407);
nand U3762 (N_3762,In_389,In_233);
nor U3763 (N_3763,In_1577,In_433);
or U3764 (N_3764,In_721,In_959);
or U3765 (N_3765,In_516,In_157);
nor U3766 (N_3766,In_2209,In_1808);
nand U3767 (N_3767,In_764,In_2244);
nor U3768 (N_3768,In_486,In_1494);
nand U3769 (N_3769,In_875,In_2386);
nand U3770 (N_3770,In_718,In_2352);
nand U3771 (N_3771,In_429,In_340);
or U3772 (N_3772,In_515,In_170);
or U3773 (N_3773,In_1447,In_2106);
or U3774 (N_3774,In_2129,In_751);
and U3775 (N_3775,In_21,In_1472);
and U3776 (N_3776,In_198,In_1510);
nor U3777 (N_3777,In_422,In_222);
xor U3778 (N_3778,In_1374,In_1448);
nand U3779 (N_3779,In_1006,In_878);
nor U3780 (N_3780,In_920,In_488);
nand U3781 (N_3781,In_585,In_758);
or U3782 (N_3782,In_945,In_2316);
and U3783 (N_3783,In_136,In_2130);
or U3784 (N_3784,In_1299,In_1875);
xor U3785 (N_3785,In_2370,In_167);
or U3786 (N_3786,In_476,In_336);
nand U3787 (N_3787,In_1728,In_1513);
nor U3788 (N_3788,In_2412,In_1438);
xnor U3789 (N_3789,In_1700,In_2080);
or U3790 (N_3790,In_474,In_2499);
nor U3791 (N_3791,In_1672,In_928);
or U3792 (N_3792,In_1068,In_2173);
xnor U3793 (N_3793,In_1162,In_910);
nor U3794 (N_3794,In_1856,In_1788);
or U3795 (N_3795,In_1932,In_734);
or U3796 (N_3796,In_642,In_407);
xor U3797 (N_3797,In_2179,In_2411);
nand U3798 (N_3798,In_186,In_1997);
or U3799 (N_3799,In_60,In_252);
nand U3800 (N_3800,In_1396,In_1491);
nand U3801 (N_3801,In_1871,In_577);
or U3802 (N_3802,In_2063,In_851);
and U3803 (N_3803,In_1828,In_182);
nand U3804 (N_3804,In_2287,In_2215);
and U3805 (N_3805,In_751,In_529);
and U3806 (N_3806,In_47,In_451);
and U3807 (N_3807,In_2126,In_132);
nand U3808 (N_3808,In_1770,In_2490);
and U3809 (N_3809,In_1061,In_872);
and U3810 (N_3810,In_1428,In_1284);
xnor U3811 (N_3811,In_1245,In_1009);
xor U3812 (N_3812,In_1687,In_1514);
xor U3813 (N_3813,In_522,In_1826);
xor U3814 (N_3814,In_1886,In_2401);
nor U3815 (N_3815,In_891,In_2055);
and U3816 (N_3816,In_330,In_2343);
nand U3817 (N_3817,In_1557,In_105);
nand U3818 (N_3818,In_1199,In_1769);
nor U3819 (N_3819,In_2172,In_1804);
xor U3820 (N_3820,In_890,In_2324);
or U3821 (N_3821,In_1438,In_1221);
xnor U3822 (N_3822,In_1546,In_1594);
nand U3823 (N_3823,In_901,In_1273);
xnor U3824 (N_3824,In_2345,In_425);
xor U3825 (N_3825,In_1438,In_2250);
and U3826 (N_3826,In_698,In_58);
nand U3827 (N_3827,In_143,In_2095);
xor U3828 (N_3828,In_1597,In_253);
or U3829 (N_3829,In_2268,In_1979);
and U3830 (N_3830,In_40,In_1811);
and U3831 (N_3831,In_186,In_211);
and U3832 (N_3832,In_202,In_2027);
nand U3833 (N_3833,In_627,In_702);
or U3834 (N_3834,In_559,In_1949);
nand U3835 (N_3835,In_1721,In_238);
xnor U3836 (N_3836,In_1798,In_1858);
xnor U3837 (N_3837,In_1146,In_870);
nand U3838 (N_3838,In_1090,In_756);
xor U3839 (N_3839,In_1209,In_1188);
or U3840 (N_3840,In_1292,In_1426);
nand U3841 (N_3841,In_1736,In_882);
nor U3842 (N_3842,In_2285,In_923);
or U3843 (N_3843,In_420,In_1948);
nor U3844 (N_3844,In_1897,In_1072);
or U3845 (N_3845,In_684,In_2432);
and U3846 (N_3846,In_281,In_2396);
nor U3847 (N_3847,In_901,In_767);
and U3848 (N_3848,In_1524,In_1276);
nor U3849 (N_3849,In_2334,In_2291);
and U3850 (N_3850,In_1205,In_909);
or U3851 (N_3851,In_1994,In_330);
xnor U3852 (N_3852,In_180,In_2053);
and U3853 (N_3853,In_316,In_671);
or U3854 (N_3854,In_1118,In_186);
and U3855 (N_3855,In_2252,In_638);
and U3856 (N_3856,In_141,In_1943);
nor U3857 (N_3857,In_1278,In_2148);
xnor U3858 (N_3858,In_1970,In_989);
nor U3859 (N_3859,In_2219,In_2286);
and U3860 (N_3860,In_1827,In_934);
or U3861 (N_3861,In_2086,In_1643);
xnor U3862 (N_3862,In_1789,In_1180);
or U3863 (N_3863,In_1919,In_1989);
or U3864 (N_3864,In_1505,In_1391);
nor U3865 (N_3865,In_116,In_1365);
xnor U3866 (N_3866,In_712,In_1296);
nor U3867 (N_3867,In_708,In_781);
or U3868 (N_3868,In_386,In_47);
nor U3869 (N_3869,In_376,In_1478);
and U3870 (N_3870,In_984,In_938);
nor U3871 (N_3871,In_1420,In_1606);
nor U3872 (N_3872,In_209,In_1428);
and U3873 (N_3873,In_1218,In_1703);
or U3874 (N_3874,In_2428,In_1163);
or U3875 (N_3875,In_1229,In_695);
and U3876 (N_3876,In_700,In_1408);
nor U3877 (N_3877,In_2433,In_1128);
or U3878 (N_3878,In_1039,In_2238);
and U3879 (N_3879,In_53,In_78);
nand U3880 (N_3880,In_2445,In_944);
or U3881 (N_3881,In_1657,In_2203);
or U3882 (N_3882,In_1458,In_1352);
xnor U3883 (N_3883,In_1191,In_338);
xor U3884 (N_3884,In_2116,In_2042);
and U3885 (N_3885,In_1840,In_2242);
nand U3886 (N_3886,In_2421,In_1184);
nor U3887 (N_3887,In_962,In_595);
nand U3888 (N_3888,In_1344,In_1280);
nand U3889 (N_3889,In_1970,In_2051);
nand U3890 (N_3890,In_2044,In_1222);
xor U3891 (N_3891,In_1437,In_2162);
nor U3892 (N_3892,In_1326,In_503);
or U3893 (N_3893,In_1488,In_1513);
xor U3894 (N_3894,In_1844,In_105);
nor U3895 (N_3895,In_1992,In_366);
nor U3896 (N_3896,In_1057,In_1139);
nor U3897 (N_3897,In_1528,In_1751);
or U3898 (N_3898,In_1029,In_649);
nor U3899 (N_3899,In_1243,In_1319);
nor U3900 (N_3900,In_848,In_1095);
or U3901 (N_3901,In_2334,In_827);
and U3902 (N_3902,In_1050,In_1531);
or U3903 (N_3903,In_1620,In_890);
and U3904 (N_3904,In_1412,In_1203);
nor U3905 (N_3905,In_2082,In_2262);
nand U3906 (N_3906,In_1851,In_1896);
nand U3907 (N_3907,In_926,In_129);
or U3908 (N_3908,In_1235,In_958);
and U3909 (N_3909,In_2239,In_585);
and U3910 (N_3910,In_129,In_182);
nand U3911 (N_3911,In_481,In_1835);
and U3912 (N_3912,In_293,In_2334);
nor U3913 (N_3913,In_125,In_188);
and U3914 (N_3914,In_886,In_1976);
and U3915 (N_3915,In_563,In_612);
xor U3916 (N_3916,In_2263,In_2223);
nor U3917 (N_3917,In_1298,In_1782);
and U3918 (N_3918,In_491,In_104);
nor U3919 (N_3919,In_2243,In_2495);
xor U3920 (N_3920,In_431,In_217);
xor U3921 (N_3921,In_902,In_1684);
nand U3922 (N_3922,In_2096,In_661);
nand U3923 (N_3923,In_1838,In_1096);
and U3924 (N_3924,In_976,In_1057);
or U3925 (N_3925,In_112,In_1997);
xor U3926 (N_3926,In_625,In_354);
nor U3927 (N_3927,In_181,In_36);
nor U3928 (N_3928,In_178,In_730);
nand U3929 (N_3929,In_1004,In_1058);
xor U3930 (N_3930,In_1880,In_561);
nor U3931 (N_3931,In_2445,In_1538);
nand U3932 (N_3932,In_1697,In_1595);
nand U3933 (N_3933,In_630,In_461);
or U3934 (N_3934,In_1927,In_430);
xnor U3935 (N_3935,In_891,In_391);
and U3936 (N_3936,In_982,In_1128);
and U3937 (N_3937,In_341,In_2113);
and U3938 (N_3938,In_279,In_2364);
nand U3939 (N_3939,In_1034,In_421);
nor U3940 (N_3940,In_2030,In_2295);
nor U3941 (N_3941,In_219,In_1601);
nor U3942 (N_3942,In_1526,In_259);
or U3943 (N_3943,In_573,In_1412);
or U3944 (N_3944,In_1848,In_755);
or U3945 (N_3945,In_1675,In_581);
nor U3946 (N_3946,In_903,In_1237);
nor U3947 (N_3947,In_518,In_1069);
xor U3948 (N_3948,In_2200,In_801);
xnor U3949 (N_3949,In_76,In_1304);
or U3950 (N_3950,In_1152,In_2422);
xnor U3951 (N_3951,In_1515,In_441);
or U3952 (N_3952,In_957,In_1677);
nor U3953 (N_3953,In_641,In_1963);
nand U3954 (N_3954,In_1438,In_404);
or U3955 (N_3955,In_460,In_2470);
or U3956 (N_3956,In_1708,In_465);
and U3957 (N_3957,In_1525,In_723);
nor U3958 (N_3958,In_1954,In_618);
nand U3959 (N_3959,In_1707,In_1239);
or U3960 (N_3960,In_1203,In_2382);
nand U3961 (N_3961,In_2190,In_962);
nor U3962 (N_3962,In_820,In_777);
or U3963 (N_3963,In_989,In_793);
xnor U3964 (N_3964,In_385,In_891);
nor U3965 (N_3965,In_1503,In_549);
nand U3966 (N_3966,In_2166,In_35);
nor U3967 (N_3967,In_2030,In_363);
xnor U3968 (N_3968,In_2375,In_1820);
nand U3969 (N_3969,In_2296,In_459);
nand U3970 (N_3970,In_1166,In_583);
nor U3971 (N_3971,In_619,In_1862);
xnor U3972 (N_3972,In_1536,In_1016);
or U3973 (N_3973,In_928,In_1979);
nand U3974 (N_3974,In_1581,In_214);
nand U3975 (N_3975,In_2286,In_584);
or U3976 (N_3976,In_175,In_883);
and U3977 (N_3977,In_77,In_1819);
or U3978 (N_3978,In_2390,In_60);
and U3979 (N_3979,In_1436,In_2437);
xor U3980 (N_3980,In_981,In_410);
nand U3981 (N_3981,In_1023,In_1648);
nand U3982 (N_3982,In_1607,In_1735);
nor U3983 (N_3983,In_807,In_594);
nand U3984 (N_3984,In_975,In_2137);
and U3985 (N_3985,In_1543,In_1502);
nand U3986 (N_3986,In_64,In_1915);
nor U3987 (N_3987,In_1349,In_1599);
xor U3988 (N_3988,In_1134,In_1396);
or U3989 (N_3989,In_260,In_2433);
nor U3990 (N_3990,In_1846,In_564);
nor U3991 (N_3991,In_910,In_2208);
and U3992 (N_3992,In_2127,In_99);
xnor U3993 (N_3993,In_2419,In_2339);
or U3994 (N_3994,In_2419,In_50);
and U3995 (N_3995,In_861,In_271);
nor U3996 (N_3996,In_1694,In_811);
xor U3997 (N_3997,In_538,In_434);
xor U3998 (N_3998,In_1364,In_1682);
xor U3999 (N_3999,In_1350,In_2322);
and U4000 (N_4000,In_983,In_1741);
nor U4001 (N_4001,In_1843,In_2477);
and U4002 (N_4002,In_1385,In_2089);
or U4003 (N_4003,In_2394,In_1643);
xor U4004 (N_4004,In_2182,In_2006);
and U4005 (N_4005,In_1578,In_2093);
and U4006 (N_4006,In_1714,In_902);
or U4007 (N_4007,In_2127,In_655);
xnor U4008 (N_4008,In_1049,In_1868);
and U4009 (N_4009,In_2387,In_2416);
or U4010 (N_4010,In_1026,In_1006);
xor U4011 (N_4011,In_1067,In_2245);
nand U4012 (N_4012,In_2010,In_327);
or U4013 (N_4013,In_1422,In_1750);
nor U4014 (N_4014,In_1506,In_1545);
or U4015 (N_4015,In_1423,In_915);
or U4016 (N_4016,In_1633,In_1823);
and U4017 (N_4017,In_1246,In_1365);
and U4018 (N_4018,In_510,In_476);
and U4019 (N_4019,In_239,In_1819);
nor U4020 (N_4020,In_1077,In_2493);
and U4021 (N_4021,In_331,In_1252);
and U4022 (N_4022,In_279,In_980);
nor U4023 (N_4023,In_930,In_1923);
xnor U4024 (N_4024,In_1594,In_1217);
or U4025 (N_4025,In_192,In_2008);
nor U4026 (N_4026,In_718,In_1278);
and U4027 (N_4027,In_207,In_2127);
nor U4028 (N_4028,In_669,In_627);
nor U4029 (N_4029,In_695,In_1872);
xnor U4030 (N_4030,In_1263,In_1294);
nand U4031 (N_4031,In_184,In_37);
and U4032 (N_4032,In_2330,In_1129);
and U4033 (N_4033,In_2200,In_1673);
or U4034 (N_4034,In_1365,In_2450);
nor U4035 (N_4035,In_263,In_171);
nand U4036 (N_4036,In_2183,In_2011);
xor U4037 (N_4037,In_1963,In_1841);
and U4038 (N_4038,In_1614,In_238);
and U4039 (N_4039,In_875,In_679);
nand U4040 (N_4040,In_1724,In_2217);
and U4041 (N_4041,In_362,In_1474);
xor U4042 (N_4042,In_2069,In_2313);
or U4043 (N_4043,In_297,In_168);
xor U4044 (N_4044,In_1793,In_784);
xnor U4045 (N_4045,In_1911,In_1528);
or U4046 (N_4046,In_2260,In_2383);
nand U4047 (N_4047,In_546,In_986);
and U4048 (N_4048,In_1935,In_1639);
xor U4049 (N_4049,In_384,In_1225);
nor U4050 (N_4050,In_612,In_2391);
or U4051 (N_4051,In_707,In_2329);
and U4052 (N_4052,In_527,In_118);
or U4053 (N_4053,In_1254,In_695);
and U4054 (N_4054,In_1443,In_162);
xnor U4055 (N_4055,In_962,In_1429);
xnor U4056 (N_4056,In_832,In_1701);
or U4057 (N_4057,In_1713,In_824);
or U4058 (N_4058,In_128,In_1539);
nand U4059 (N_4059,In_734,In_1879);
nor U4060 (N_4060,In_1724,In_1594);
xor U4061 (N_4061,In_2374,In_2253);
or U4062 (N_4062,In_1846,In_1314);
xnor U4063 (N_4063,In_992,In_1385);
nor U4064 (N_4064,In_2495,In_1623);
nor U4065 (N_4065,In_466,In_216);
nand U4066 (N_4066,In_399,In_531);
xnor U4067 (N_4067,In_2204,In_1774);
nand U4068 (N_4068,In_373,In_1772);
xor U4069 (N_4069,In_1608,In_2147);
and U4070 (N_4070,In_99,In_1847);
or U4071 (N_4071,In_823,In_1465);
and U4072 (N_4072,In_2046,In_110);
or U4073 (N_4073,In_1788,In_1776);
nor U4074 (N_4074,In_1766,In_2272);
or U4075 (N_4075,In_1346,In_1423);
or U4076 (N_4076,In_1944,In_957);
nor U4077 (N_4077,In_689,In_538);
xnor U4078 (N_4078,In_1092,In_789);
nand U4079 (N_4079,In_1470,In_1793);
nand U4080 (N_4080,In_2310,In_2185);
xor U4081 (N_4081,In_2397,In_591);
xnor U4082 (N_4082,In_803,In_740);
or U4083 (N_4083,In_866,In_989);
xnor U4084 (N_4084,In_1255,In_1744);
nor U4085 (N_4085,In_1898,In_126);
or U4086 (N_4086,In_1314,In_871);
xnor U4087 (N_4087,In_475,In_1487);
xor U4088 (N_4088,In_1155,In_286);
nor U4089 (N_4089,In_1874,In_1326);
and U4090 (N_4090,In_2257,In_1169);
or U4091 (N_4091,In_990,In_447);
or U4092 (N_4092,In_1765,In_1459);
or U4093 (N_4093,In_1234,In_2333);
and U4094 (N_4094,In_2439,In_1169);
nor U4095 (N_4095,In_634,In_533);
nor U4096 (N_4096,In_362,In_1152);
or U4097 (N_4097,In_1885,In_254);
nand U4098 (N_4098,In_1154,In_737);
or U4099 (N_4099,In_1978,In_157);
xor U4100 (N_4100,In_1397,In_2290);
nand U4101 (N_4101,In_2294,In_1077);
nand U4102 (N_4102,In_485,In_1629);
nand U4103 (N_4103,In_2406,In_281);
nor U4104 (N_4104,In_2387,In_754);
nor U4105 (N_4105,In_740,In_2349);
and U4106 (N_4106,In_560,In_183);
nor U4107 (N_4107,In_731,In_1823);
or U4108 (N_4108,In_1992,In_2481);
or U4109 (N_4109,In_484,In_41);
xnor U4110 (N_4110,In_448,In_2116);
and U4111 (N_4111,In_1366,In_391);
nand U4112 (N_4112,In_2179,In_264);
nand U4113 (N_4113,In_1741,In_284);
nand U4114 (N_4114,In_2109,In_263);
xor U4115 (N_4115,In_285,In_774);
nor U4116 (N_4116,In_1805,In_2425);
nand U4117 (N_4117,In_568,In_97);
and U4118 (N_4118,In_2336,In_875);
or U4119 (N_4119,In_861,In_818);
or U4120 (N_4120,In_1524,In_1003);
and U4121 (N_4121,In_204,In_1998);
nor U4122 (N_4122,In_2305,In_1288);
xnor U4123 (N_4123,In_238,In_1438);
nand U4124 (N_4124,In_1586,In_1591);
xor U4125 (N_4125,In_426,In_1647);
xnor U4126 (N_4126,In_514,In_431);
xor U4127 (N_4127,In_1166,In_813);
nand U4128 (N_4128,In_281,In_510);
and U4129 (N_4129,In_345,In_1106);
nand U4130 (N_4130,In_2257,In_221);
xor U4131 (N_4131,In_456,In_1347);
nand U4132 (N_4132,In_1106,In_300);
nand U4133 (N_4133,In_627,In_1511);
and U4134 (N_4134,In_963,In_684);
nor U4135 (N_4135,In_505,In_1266);
and U4136 (N_4136,In_2238,In_1643);
and U4137 (N_4137,In_451,In_465);
or U4138 (N_4138,In_1389,In_2486);
or U4139 (N_4139,In_1665,In_2200);
or U4140 (N_4140,In_1079,In_1213);
or U4141 (N_4141,In_2202,In_1828);
nand U4142 (N_4142,In_2325,In_295);
and U4143 (N_4143,In_1729,In_322);
xor U4144 (N_4144,In_1259,In_2074);
xnor U4145 (N_4145,In_2420,In_2054);
xnor U4146 (N_4146,In_355,In_2364);
and U4147 (N_4147,In_2,In_2107);
nor U4148 (N_4148,In_2282,In_1068);
or U4149 (N_4149,In_82,In_2245);
xor U4150 (N_4150,In_955,In_34);
or U4151 (N_4151,In_1578,In_558);
or U4152 (N_4152,In_904,In_294);
xor U4153 (N_4153,In_313,In_661);
and U4154 (N_4154,In_1457,In_1663);
xnor U4155 (N_4155,In_19,In_892);
nand U4156 (N_4156,In_640,In_562);
nor U4157 (N_4157,In_1408,In_871);
and U4158 (N_4158,In_2380,In_1785);
xor U4159 (N_4159,In_1403,In_1838);
nor U4160 (N_4160,In_1639,In_2097);
or U4161 (N_4161,In_1260,In_1048);
nor U4162 (N_4162,In_1285,In_917);
nor U4163 (N_4163,In_166,In_1010);
nor U4164 (N_4164,In_897,In_858);
nor U4165 (N_4165,In_339,In_8);
and U4166 (N_4166,In_556,In_1201);
or U4167 (N_4167,In_2469,In_1199);
and U4168 (N_4168,In_1651,In_1414);
nand U4169 (N_4169,In_1609,In_194);
xnor U4170 (N_4170,In_130,In_2276);
nand U4171 (N_4171,In_1588,In_732);
nand U4172 (N_4172,In_1767,In_1040);
xnor U4173 (N_4173,In_2061,In_1232);
nor U4174 (N_4174,In_1700,In_774);
or U4175 (N_4175,In_1911,In_1295);
xnor U4176 (N_4176,In_1989,In_1189);
or U4177 (N_4177,In_465,In_257);
xor U4178 (N_4178,In_1369,In_894);
xor U4179 (N_4179,In_2450,In_1412);
or U4180 (N_4180,In_2109,In_2146);
xnor U4181 (N_4181,In_1272,In_2172);
nand U4182 (N_4182,In_2296,In_1213);
nor U4183 (N_4183,In_979,In_616);
and U4184 (N_4184,In_1099,In_1541);
or U4185 (N_4185,In_1218,In_1951);
nor U4186 (N_4186,In_700,In_235);
nand U4187 (N_4187,In_1462,In_2131);
and U4188 (N_4188,In_946,In_2452);
nand U4189 (N_4189,In_1930,In_2346);
xor U4190 (N_4190,In_420,In_893);
xnor U4191 (N_4191,In_247,In_182);
and U4192 (N_4192,In_1455,In_228);
nor U4193 (N_4193,In_1109,In_882);
and U4194 (N_4194,In_2229,In_1665);
nor U4195 (N_4195,In_75,In_1287);
nor U4196 (N_4196,In_2370,In_885);
nand U4197 (N_4197,In_1105,In_731);
xor U4198 (N_4198,In_805,In_953);
nor U4199 (N_4199,In_854,In_1731);
nor U4200 (N_4200,In_2416,In_1046);
and U4201 (N_4201,In_683,In_825);
nand U4202 (N_4202,In_1351,In_2070);
nand U4203 (N_4203,In_2313,In_2146);
xnor U4204 (N_4204,In_2358,In_1697);
xnor U4205 (N_4205,In_2257,In_837);
nor U4206 (N_4206,In_398,In_1300);
xor U4207 (N_4207,In_1475,In_1345);
or U4208 (N_4208,In_739,In_1041);
or U4209 (N_4209,In_1533,In_1610);
xor U4210 (N_4210,In_133,In_1788);
nand U4211 (N_4211,In_1245,In_278);
xnor U4212 (N_4212,In_2332,In_706);
nand U4213 (N_4213,In_1363,In_2463);
nand U4214 (N_4214,In_377,In_2250);
or U4215 (N_4215,In_1860,In_1271);
xor U4216 (N_4216,In_1061,In_1631);
nor U4217 (N_4217,In_2490,In_1899);
and U4218 (N_4218,In_2422,In_247);
xor U4219 (N_4219,In_1343,In_555);
xnor U4220 (N_4220,In_1,In_1549);
nand U4221 (N_4221,In_442,In_711);
nand U4222 (N_4222,In_1032,In_1645);
and U4223 (N_4223,In_1580,In_21);
nand U4224 (N_4224,In_112,In_720);
xnor U4225 (N_4225,In_2484,In_2330);
xor U4226 (N_4226,In_182,In_1162);
xor U4227 (N_4227,In_1363,In_1102);
and U4228 (N_4228,In_673,In_100);
and U4229 (N_4229,In_440,In_1728);
nor U4230 (N_4230,In_853,In_1101);
nand U4231 (N_4231,In_668,In_81);
xnor U4232 (N_4232,In_154,In_542);
nand U4233 (N_4233,In_784,In_2238);
or U4234 (N_4234,In_551,In_980);
or U4235 (N_4235,In_1074,In_1924);
xor U4236 (N_4236,In_1078,In_1876);
nor U4237 (N_4237,In_695,In_881);
xor U4238 (N_4238,In_377,In_2253);
nor U4239 (N_4239,In_1978,In_1457);
xor U4240 (N_4240,In_1300,In_1581);
and U4241 (N_4241,In_1015,In_1131);
nand U4242 (N_4242,In_801,In_701);
xnor U4243 (N_4243,In_1973,In_1124);
nor U4244 (N_4244,In_1799,In_2143);
or U4245 (N_4245,In_1249,In_1789);
xor U4246 (N_4246,In_2013,In_1354);
nand U4247 (N_4247,In_2484,In_358);
and U4248 (N_4248,In_1769,In_2339);
and U4249 (N_4249,In_975,In_1501);
and U4250 (N_4250,In_834,In_1171);
nor U4251 (N_4251,In_223,In_804);
xnor U4252 (N_4252,In_263,In_113);
or U4253 (N_4253,In_972,In_324);
or U4254 (N_4254,In_396,In_240);
nor U4255 (N_4255,In_1542,In_1075);
nor U4256 (N_4256,In_226,In_538);
or U4257 (N_4257,In_1333,In_786);
nor U4258 (N_4258,In_1854,In_1673);
or U4259 (N_4259,In_717,In_253);
and U4260 (N_4260,In_468,In_1277);
nor U4261 (N_4261,In_1777,In_93);
nor U4262 (N_4262,In_169,In_1033);
and U4263 (N_4263,In_2430,In_2289);
nor U4264 (N_4264,In_2393,In_583);
nor U4265 (N_4265,In_2430,In_907);
and U4266 (N_4266,In_215,In_883);
nand U4267 (N_4267,In_1424,In_743);
and U4268 (N_4268,In_1360,In_2484);
and U4269 (N_4269,In_2066,In_2382);
nor U4270 (N_4270,In_347,In_371);
or U4271 (N_4271,In_2301,In_2229);
nor U4272 (N_4272,In_2428,In_1799);
xor U4273 (N_4273,In_1975,In_373);
nand U4274 (N_4274,In_2352,In_2085);
xor U4275 (N_4275,In_126,In_891);
and U4276 (N_4276,In_1228,In_428);
nand U4277 (N_4277,In_2264,In_2468);
xnor U4278 (N_4278,In_644,In_1396);
and U4279 (N_4279,In_2480,In_490);
or U4280 (N_4280,In_1088,In_2145);
or U4281 (N_4281,In_2389,In_1421);
nor U4282 (N_4282,In_2214,In_2370);
nor U4283 (N_4283,In_904,In_1591);
and U4284 (N_4284,In_1879,In_976);
and U4285 (N_4285,In_656,In_1715);
nor U4286 (N_4286,In_1482,In_898);
xor U4287 (N_4287,In_555,In_1624);
nand U4288 (N_4288,In_2333,In_2168);
nand U4289 (N_4289,In_1315,In_846);
and U4290 (N_4290,In_1903,In_1083);
xnor U4291 (N_4291,In_61,In_1133);
xnor U4292 (N_4292,In_1864,In_1811);
and U4293 (N_4293,In_1877,In_2383);
nand U4294 (N_4294,In_815,In_1235);
nand U4295 (N_4295,In_2438,In_1603);
xnor U4296 (N_4296,In_1903,In_1692);
or U4297 (N_4297,In_123,In_943);
nor U4298 (N_4298,In_142,In_2429);
nor U4299 (N_4299,In_1310,In_795);
and U4300 (N_4300,In_1871,In_1810);
nor U4301 (N_4301,In_2,In_861);
nand U4302 (N_4302,In_184,In_2120);
nor U4303 (N_4303,In_1273,In_346);
nand U4304 (N_4304,In_1894,In_1963);
nand U4305 (N_4305,In_19,In_41);
and U4306 (N_4306,In_144,In_344);
or U4307 (N_4307,In_1948,In_2412);
or U4308 (N_4308,In_608,In_1048);
nor U4309 (N_4309,In_241,In_1532);
nand U4310 (N_4310,In_499,In_970);
and U4311 (N_4311,In_359,In_1999);
nand U4312 (N_4312,In_1483,In_1696);
or U4313 (N_4313,In_575,In_1232);
or U4314 (N_4314,In_1922,In_87);
nand U4315 (N_4315,In_1488,In_1869);
nor U4316 (N_4316,In_1705,In_500);
nand U4317 (N_4317,In_476,In_1721);
and U4318 (N_4318,In_979,In_2409);
and U4319 (N_4319,In_1212,In_1834);
and U4320 (N_4320,In_2493,In_2356);
or U4321 (N_4321,In_1737,In_921);
and U4322 (N_4322,In_964,In_531);
or U4323 (N_4323,In_178,In_573);
nor U4324 (N_4324,In_1225,In_2411);
xnor U4325 (N_4325,In_2367,In_1704);
or U4326 (N_4326,In_2467,In_4);
nor U4327 (N_4327,In_2257,In_2190);
and U4328 (N_4328,In_392,In_1852);
xor U4329 (N_4329,In_386,In_1961);
and U4330 (N_4330,In_297,In_2144);
or U4331 (N_4331,In_1880,In_2015);
or U4332 (N_4332,In_1921,In_755);
nor U4333 (N_4333,In_1712,In_949);
nand U4334 (N_4334,In_56,In_1461);
nand U4335 (N_4335,In_325,In_186);
or U4336 (N_4336,In_14,In_885);
xor U4337 (N_4337,In_1827,In_1040);
or U4338 (N_4338,In_2246,In_1881);
and U4339 (N_4339,In_679,In_1252);
xor U4340 (N_4340,In_2117,In_2291);
xor U4341 (N_4341,In_827,In_1846);
nand U4342 (N_4342,In_845,In_1137);
nand U4343 (N_4343,In_2446,In_708);
or U4344 (N_4344,In_1054,In_146);
xor U4345 (N_4345,In_194,In_128);
nor U4346 (N_4346,In_366,In_2049);
xnor U4347 (N_4347,In_184,In_858);
nand U4348 (N_4348,In_2493,In_741);
and U4349 (N_4349,In_590,In_2468);
xor U4350 (N_4350,In_2136,In_2478);
xor U4351 (N_4351,In_162,In_1993);
nor U4352 (N_4352,In_561,In_1588);
or U4353 (N_4353,In_502,In_2383);
nor U4354 (N_4354,In_949,In_1703);
and U4355 (N_4355,In_1313,In_739);
xor U4356 (N_4356,In_2032,In_1446);
nand U4357 (N_4357,In_1652,In_1649);
nand U4358 (N_4358,In_150,In_1479);
or U4359 (N_4359,In_1944,In_2188);
xnor U4360 (N_4360,In_806,In_1114);
or U4361 (N_4361,In_205,In_1455);
nor U4362 (N_4362,In_2348,In_1765);
xnor U4363 (N_4363,In_803,In_439);
or U4364 (N_4364,In_144,In_109);
or U4365 (N_4365,In_512,In_1406);
nand U4366 (N_4366,In_909,In_470);
nor U4367 (N_4367,In_960,In_1773);
and U4368 (N_4368,In_1796,In_1187);
and U4369 (N_4369,In_648,In_227);
and U4370 (N_4370,In_2308,In_1956);
and U4371 (N_4371,In_1027,In_1558);
xnor U4372 (N_4372,In_125,In_1598);
nor U4373 (N_4373,In_869,In_2196);
xnor U4374 (N_4374,In_311,In_840);
nand U4375 (N_4375,In_1995,In_2223);
or U4376 (N_4376,In_1384,In_2470);
or U4377 (N_4377,In_1480,In_1963);
nand U4378 (N_4378,In_111,In_1480);
or U4379 (N_4379,In_1986,In_2153);
or U4380 (N_4380,In_1525,In_731);
nor U4381 (N_4381,In_8,In_677);
or U4382 (N_4382,In_2037,In_261);
nand U4383 (N_4383,In_1920,In_2203);
nand U4384 (N_4384,In_1998,In_1889);
xor U4385 (N_4385,In_1390,In_1708);
and U4386 (N_4386,In_1616,In_1774);
xor U4387 (N_4387,In_709,In_513);
and U4388 (N_4388,In_2045,In_326);
or U4389 (N_4389,In_1739,In_2421);
xor U4390 (N_4390,In_723,In_575);
nand U4391 (N_4391,In_2478,In_99);
and U4392 (N_4392,In_746,In_241);
and U4393 (N_4393,In_494,In_845);
and U4394 (N_4394,In_668,In_157);
nand U4395 (N_4395,In_816,In_1547);
nand U4396 (N_4396,In_433,In_2094);
and U4397 (N_4397,In_802,In_286);
or U4398 (N_4398,In_1557,In_443);
xor U4399 (N_4399,In_2087,In_749);
or U4400 (N_4400,In_1706,In_476);
xor U4401 (N_4401,In_1001,In_784);
xor U4402 (N_4402,In_1498,In_2056);
and U4403 (N_4403,In_532,In_173);
nor U4404 (N_4404,In_1957,In_615);
nor U4405 (N_4405,In_1994,In_2179);
and U4406 (N_4406,In_74,In_781);
and U4407 (N_4407,In_2006,In_1086);
and U4408 (N_4408,In_2350,In_1046);
and U4409 (N_4409,In_1223,In_2376);
nand U4410 (N_4410,In_959,In_180);
nor U4411 (N_4411,In_1195,In_2385);
and U4412 (N_4412,In_564,In_1480);
nand U4413 (N_4413,In_22,In_2391);
nand U4414 (N_4414,In_998,In_633);
and U4415 (N_4415,In_2444,In_296);
nor U4416 (N_4416,In_1782,In_1970);
nor U4417 (N_4417,In_1562,In_1349);
xor U4418 (N_4418,In_2180,In_301);
nand U4419 (N_4419,In_559,In_2425);
nand U4420 (N_4420,In_2354,In_386);
nand U4421 (N_4421,In_2340,In_1674);
or U4422 (N_4422,In_2422,In_1031);
or U4423 (N_4423,In_470,In_748);
xnor U4424 (N_4424,In_995,In_1478);
nand U4425 (N_4425,In_2425,In_2270);
nor U4426 (N_4426,In_1852,In_1618);
nand U4427 (N_4427,In_629,In_1914);
xnor U4428 (N_4428,In_1633,In_69);
nor U4429 (N_4429,In_995,In_1132);
and U4430 (N_4430,In_1286,In_1899);
nor U4431 (N_4431,In_2318,In_2397);
and U4432 (N_4432,In_1123,In_711);
nor U4433 (N_4433,In_434,In_623);
or U4434 (N_4434,In_310,In_122);
nor U4435 (N_4435,In_335,In_1702);
and U4436 (N_4436,In_2465,In_1713);
nor U4437 (N_4437,In_221,In_2209);
xnor U4438 (N_4438,In_1628,In_1394);
or U4439 (N_4439,In_1796,In_1571);
or U4440 (N_4440,In_1598,In_2438);
xor U4441 (N_4441,In_1803,In_1757);
nand U4442 (N_4442,In_1469,In_1970);
and U4443 (N_4443,In_530,In_182);
nor U4444 (N_4444,In_804,In_1994);
nor U4445 (N_4445,In_1630,In_1912);
and U4446 (N_4446,In_1934,In_793);
xnor U4447 (N_4447,In_991,In_1699);
or U4448 (N_4448,In_1371,In_654);
or U4449 (N_4449,In_2458,In_103);
or U4450 (N_4450,In_567,In_1331);
xnor U4451 (N_4451,In_1723,In_1202);
and U4452 (N_4452,In_550,In_1385);
xnor U4453 (N_4453,In_179,In_2473);
and U4454 (N_4454,In_1152,In_459);
xnor U4455 (N_4455,In_1722,In_1868);
and U4456 (N_4456,In_1957,In_1805);
nor U4457 (N_4457,In_1373,In_1490);
xnor U4458 (N_4458,In_344,In_661);
xnor U4459 (N_4459,In_1380,In_256);
or U4460 (N_4460,In_174,In_2110);
or U4461 (N_4461,In_961,In_2398);
nand U4462 (N_4462,In_1899,In_479);
or U4463 (N_4463,In_325,In_273);
nand U4464 (N_4464,In_1867,In_1321);
nand U4465 (N_4465,In_1736,In_1138);
xor U4466 (N_4466,In_649,In_2116);
nand U4467 (N_4467,In_1864,In_2181);
or U4468 (N_4468,In_2107,In_2157);
xor U4469 (N_4469,In_1574,In_1198);
nor U4470 (N_4470,In_456,In_823);
nand U4471 (N_4471,In_1433,In_1640);
nor U4472 (N_4472,In_259,In_110);
or U4473 (N_4473,In_514,In_1504);
xor U4474 (N_4474,In_757,In_2249);
and U4475 (N_4475,In_1716,In_1118);
and U4476 (N_4476,In_57,In_736);
nand U4477 (N_4477,In_658,In_2285);
xnor U4478 (N_4478,In_2293,In_1418);
or U4479 (N_4479,In_691,In_165);
xnor U4480 (N_4480,In_891,In_1221);
xor U4481 (N_4481,In_226,In_2386);
and U4482 (N_4482,In_2210,In_530);
nor U4483 (N_4483,In_272,In_747);
nor U4484 (N_4484,In_1656,In_1860);
nand U4485 (N_4485,In_2379,In_333);
and U4486 (N_4486,In_2115,In_2005);
nand U4487 (N_4487,In_1180,In_2042);
nor U4488 (N_4488,In_351,In_1589);
nand U4489 (N_4489,In_1081,In_1728);
nor U4490 (N_4490,In_1919,In_2063);
nand U4491 (N_4491,In_2268,In_1928);
or U4492 (N_4492,In_2173,In_2474);
xor U4493 (N_4493,In_2190,In_166);
nor U4494 (N_4494,In_2096,In_1818);
and U4495 (N_4495,In_124,In_2112);
and U4496 (N_4496,In_2126,In_1882);
or U4497 (N_4497,In_1886,In_372);
nor U4498 (N_4498,In_2142,In_586);
nor U4499 (N_4499,In_534,In_1028);
nand U4500 (N_4500,In_1798,In_2100);
and U4501 (N_4501,In_2201,In_182);
and U4502 (N_4502,In_1227,In_2422);
nor U4503 (N_4503,In_2476,In_435);
nand U4504 (N_4504,In_96,In_2278);
xnor U4505 (N_4505,In_204,In_240);
xnor U4506 (N_4506,In_1786,In_1161);
and U4507 (N_4507,In_2329,In_831);
or U4508 (N_4508,In_2118,In_2064);
or U4509 (N_4509,In_1342,In_370);
or U4510 (N_4510,In_2490,In_1160);
and U4511 (N_4511,In_1973,In_2196);
nor U4512 (N_4512,In_1894,In_1714);
xor U4513 (N_4513,In_359,In_2127);
xor U4514 (N_4514,In_377,In_202);
or U4515 (N_4515,In_1631,In_1982);
xnor U4516 (N_4516,In_987,In_1681);
nand U4517 (N_4517,In_358,In_200);
nand U4518 (N_4518,In_1073,In_378);
nand U4519 (N_4519,In_472,In_831);
and U4520 (N_4520,In_2334,In_296);
xnor U4521 (N_4521,In_545,In_2055);
and U4522 (N_4522,In_900,In_679);
nor U4523 (N_4523,In_93,In_1413);
or U4524 (N_4524,In_2021,In_1687);
or U4525 (N_4525,In_1944,In_2370);
and U4526 (N_4526,In_1247,In_1747);
nand U4527 (N_4527,In_1598,In_780);
or U4528 (N_4528,In_1732,In_1655);
and U4529 (N_4529,In_468,In_1530);
and U4530 (N_4530,In_1543,In_2064);
nand U4531 (N_4531,In_2178,In_23);
nand U4532 (N_4532,In_1569,In_325);
nor U4533 (N_4533,In_1530,In_1668);
or U4534 (N_4534,In_429,In_995);
and U4535 (N_4535,In_327,In_167);
or U4536 (N_4536,In_326,In_26);
or U4537 (N_4537,In_906,In_888);
nor U4538 (N_4538,In_266,In_1400);
or U4539 (N_4539,In_1187,In_1491);
nor U4540 (N_4540,In_1526,In_1414);
or U4541 (N_4541,In_1951,In_1955);
or U4542 (N_4542,In_169,In_502);
and U4543 (N_4543,In_829,In_2077);
nor U4544 (N_4544,In_2270,In_1525);
nor U4545 (N_4545,In_2149,In_2398);
xor U4546 (N_4546,In_1314,In_2081);
nand U4547 (N_4547,In_1815,In_591);
xnor U4548 (N_4548,In_1003,In_1746);
xnor U4549 (N_4549,In_1112,In_2374);
or U4550 (N_4550,In_2328,In_636);
nor U4551 (N_4551,In_1166,In_1390);
or U4552 (N_4552,In_488,In_2318);
or U4553 (N_4553,In_2357,In_264);
nand U4554 (N_4554,In_309,In_1412);
nand U4555 (N_4555,In_974,In_704);
nand U4556 (N_4556,In_2292,In_1192);
xnor U4557 (N_4557,In_631,In_1983);
xor U4558 (N_4558,In_301,In_1620);
or U4559 (N_4559,In_868,In_1123);
xor U4560 (N_4560,In_2172,In_986);
nor U4561 (N_4561,In_1029,In_1987);
and U4562 (N_4562,In_325,In_6);
nand U4563 (N_4563,In_2321,In_1793);
nor U4564 (N_4564,In_266,In_108);
nor U4565 (N_4565,In_92,In_774);
nor U4566 (N_4566,In_2134,In_25);
and U4567 (N_4567,In_616,In_1268);
or U4568 (N_4568,In_1076,In_1530);
or U4569 (N_4569,In_33,In_2138);
xnor U4570 (N_4570,In_1486,In_669);
xor U4571 (N_4571,In_1988,In_1580);
and U4572 (N_4572,In_1852,In_2117);
or U4573 (N_4573,In_954,In_791);
or U4574 (N_4574,In_638,In_348);
xor U4575 (N_4575,In_34,In_1365);
or U4576 (N_4576,In_1819,In_518);
and U4577 (N_4577,In_305,In_1268);
xnor U4578 (N_4578,In_1014,In_1293);
nor U4579 (N_4579,In_2040,In_2218);
nor U4580 (N_4580,In_516,In_666);
and U4581 (N_4581,In_106,In_99);
or U4582 (N_4582,In_2263,In_1146);
or U4583 (N_4583,In_2246,In_908);
and U4584 (N_4584,In_1711,In_792);
xor U4585 (N_4585,In_34,In_1190);
or U4586 (N_4586,In_640,In_2064);
xor U4587 (N_4587,In_377,In_643);
and U4588 (N_4588,In_36,In_784);
xor U4589 (N_4589,In_1166,In_652);
or U4590 (N_4590,In_507,In_310);
nor U4591 (N_4591,In_729,In_2177);
nor U4592 (N_4592,In_1306,In_345);
nor U4593 (N_4593,In_2426,In_1742);
nor U4594 (N_4594,In_1826,In_173);
nor U4595 (N_4595,In_1324,In_2190);
nand U4596 (N_4596,In_1931,In_1194);
xnor U4597 (N_4597,In_1231,In_1852);
nand U4598 (N_4598,In_239,In_827);
xor U4599 (N_4599,In_432,In_487);
or U4600 (N_4600,In_874,In_1494);
xnor U4601 (N_4601,In_1448,In_1754);
nand U4602 (N_4602,In_951,In_1282);
nor U4603 (N_4603,In_1602,In_1724);
nand U4604 (N_4604,In_2278,In_1746);
and U4605 (N_4605,In_1764,In_1717);
xor U4606 (N_4606,In_2431,In_266);
xor U4607 (N_4607,In_1560,In_180);
or U4608 (N_4608,In_181,In_31);
nand U4609 (N_4609,In_343,In_465);
nand U4610 (N_4610,In_1269,In_1569);
and U4611 (N_4611,In_1632,In_2174);
nor U4612 (N_4612,In_497,In_1907);
xnor U4613 (N_4613,In_154,In_1622);
and U4614 (N_4614,In_1393,In_2029);
xor U4615 (N_4615,In_1397,In_1377);
or U4616 (N_4616,In_1999,In_610);
or U4617 (N_4617,In_1802,In_598);
or U4618 (N_4618,In_162,In_1469);
or U4619 (N_4619,In_753,In_579);
nor U4620 (N_4620,In_1648,In_1897);
xnor U4621 (N_4621,In_1817,In_1888);
or U4622 (N_4622,In_109,In_1815);
and U4623 (N_4623,In_926,In_2046);
xor U4624 (N_4624,In_21,In_1818);
nand U4625 (N_4625,In_1868,In_2018);
nand U4626 (N_4626,In_5,In_2162);
nor U4627 (N_4627,In_778,In_1818);
xor U4628 (N_4628,In_1518,In_300);
nor U4629 (N_4629,In_2484,In_2069);
and U4630 (N_4630,In_1295,In_1504);
or U4631 (N_4631,In_2423,In_1398);
nand U4632 (N_4632,In_1546,In_983);
nor U4633 (N_4633,In_2322,In_2292);
and U4634 (N_4634,In_733,In_1032);
xor U4635 (N_4635,In_303,In_214);
and U4636 (N_4636,In_199,In_1851);
nand U4637 (N_4637,In_603,In_1387);
xor U4638 (N_4638,In_2367,In_1230);
xnor U4639 (N_4639,In_453,In_1514);
nor U4640 (N_4640,In_1003,In_997);
nand U4641 (N_4641,In_134,In_28);
nand U4642 (N_4642,In_554,In_909);
xnor U4643 (N_4643,In_2086,In_1132);
or U4644 (N_4644,In_2125,In_1986);
nor U4645 (N_4645,In_1014,In_1610);
nor U4646 (N_4646,In_2277,In_1092);
xor U4647 (N_4647,In_2410,In_2468);
nor U4648 (N_4648,In_2430,In_396);
nor U4649 (N_4649,In_940,In_1203);
nor U4650 (N_4650,In_1399,In_921);
xnor U4651 (N_4651,In_848,In_720);
nor U4652 (N_4652,In_996,In_281);
and U4653 (N_4653,In_1384,In_294);
xnor U4654 (N_4654,In_1191,In_1490);
xnor U4655 (N_4655,In_39,In_299);
nor U4656 (N_4656,In_2033,In_1589);
nor U4657 (N_4657,In_2108,In_1281);
nor U4658 (N_4658,In_888,In_1952);
and U4659 (N_4659,In_1670,In_753);
or U4660 (N_4660,In_2067,In_2032);
xor U4661 (N_4661,In_1138,In_465);
xor U4662 (N_4662,In_510,In_2022);
xnor U4663 (N_4663,In_945,In_1716);
nor U4664 (N_4664,In_145,In_1170);
nand U4665 (N_4665,In_2194,In_223);
and U4666 (N_4666,In_2370,In_1953);
xnor U4667 (N_4667,In_1668,In_1848);
and U4668 (N_4668,In_933,In_1642);
and U4669 (N_4669,In_195,In_2242);
xnor U4670 (N_4670,In_277,In_357);
nand U4671 (N_4671,In_5,In_1764);
nor U4672 (N_4672,In_1339,In_740);
nand U4673 (N_4673,In_1941,In_1506);
nor U4674 (N_4674,In_1445,In_1259);
and U4675 (N_4675,In_2232,In_615);
or U4676 (N_4676,In_725,In_33);
or U4677 (N_4677,In_2094,In_568);
nand U4678 (N_4678,In_1725,In_1207);
xnor U4679 (N_4679,In_1241,In_1027);
nand U4680 (N_4680,In_10,In_2289);
nor U4681 (N_4681,In_2134,In_334);
and U4682 (N_4682,In_940,In_486);
xor U4683 (N_4683,In_18,In_207);
or U4684 (N_4684,In_2115,In_452);
and U4685 (N_4685,In_1049,In_1172);
xor U4686 (N_4686,In_2181,In_1887);
and U4687 (N_4687,In_317,In_1774);
nor U4688 (N_4688,In_2155,In_1373);
xor U4689 (N_4689,In_631,In_2195);
nand U4690 (N_4690,In_1652,In_1089);
and U4691 (N_4691,In_1548,In_1774);
and U4692 (N_4692,In_2481,In_292);
nand U4693 (N_4693,In_169,In_875);
nor U4694 (N_4694,In_1446,In_2422);
and U4695 (N_4695,In_446,In_1038);
and U4696 (N_4696,In_486,In_1666);
xor U4697 (N_4697,In_1223,In_1256);
nand U4698 (N_4698,In_1871,In_1929);
xnor U4699 (N_4699,In_373,In_840);
xnor U4700 (N_4700,In_577,In_1988);
nor U4701 (N_4701,In_554,In_229);
xnor U4702 (N_4702,In_1677,In_1294);
nor U4703 (N_4703,In_619,In_1978);
nor U4704 (N_4704,In_1346,In_2310);
nand U4705 (N_4705,In_608,In_1558);
and U4706 (N_4706,In_1076,In_252);
or U4707 (N_4707,In_2306,In_2056);
nand U4708 (N_4708,In_248,In_503);
and U4709 (N_4709,In_768,In_1994);
nand U4710 (N_4710,In_757,In_843);
or U4711 (N_4711,In_851,In_1738);
and U4712 (N_4712,In_811,In_716);
nand U4713 (N_4713,In_1284,In_597);
or U4714 (N_4714,In_2417,In_1175);
xor U4715 (N_4715,In_1790,In_2028);
or U4716 (N_4716,In_2109,In_677);
xnor U4717 (N_4717,In_332,In_1519);
or U4718 (N_4718,In_1854,In_2178);
nand U4719 (N_4719,In_2091,In_1757);
nor U4720 (N_4720,In_362,In_1919);
or U4721 (N_4721,In_2370,In_1633);
nand U4722 (N_4722,In_1693,In_1314);
and U4723 (N_4723,In_501,In_597);
nor U4724 (N_4724,In_1079,In_2382);
nor U4725 (N_4725,In_2106,In_1765);
nand U4726 (N_4726,In_1856,In_1790);
nand U4727 (N_4727,In_923,In_1344);
nor U4728 (N_4728,In_595,In_2124);
or U4729 (N_4729,In_2369,In_2424);
or U4730 (N_4730,In_257,In_1387);
xor U4731 (N_4731,In_2453,In_1728);
nor U4732 (N_4732,In_2173,In_1338);
nand U4733 (N_4733,In_2189,In_1565);
xnor U4734 (N_4734,In_548,In_365);
nand U4735 (N_4735,In_1634,In_2380);
nor U4736 (N_4736,In_809,In_2344);
xor U4737 (N_4737,In_529,In_944);
or U4738 (N_4738,In_43,In_1765);
nor U4739 (N_4739,In_1500,In_68);
or U4740 (N_4740,In_647,In_1584);
xor U4741 (N_4741,In_4,In_1657);
xnor U4742 (N_4742,In_2355,In_1132);
xor U4743 (N_4743,In_150,In_379);
xnor U4744 (N_4744,In_1233,In_1506);
nand U4745 (N_4745,In_2292,In_1829);
or U4746 (N_4746,In_1226,In_570);
nor U4747 (N_4747,In_1235,In_2110);
nor U4748 (N_4748,In_2037,In_2434);
and U4749 (N_4749,In_1649,In_2008);
and U4750 (N_4750,In_2428,In_501);
nand U4751 (N_4751,In_986,In_555);
and U4752 (N_4752,In_1671,In_1222);
nand U4753 (N_4753,In_2320,In_605);
or U4754 (N_4754,In_2052,In_2468);
and U4755 (N_4755,In_1919,In_2074);
nor U4756 (N_4756,In_67,In_1334);
nor U4757 (N_4757,In_1389,In_1782);
or U4758 (N_4758,In_200,In_1397);
xor U4759 (N_4759,In_1390,In_116);
nor U4760 (N_4760,In_1405,In_1723);
nand U4761 (N_4761,In_633,In_1506);
and U4762 (N_4762,In_1932,In_2389);
nand U4763 (N_4763,In_144,In_2485);
nand U4764 (N_4764,In_1836,In_550);
xor U4765 (N_4765,In_309,In_793);
and U4766 (N_4766,In_833,In_929);
xor U4767 (N_4767,In_1711,In_1231);
or U4768 (N_4768,In_1224,In_866);
nand U4769 (N_4769,In_722,In_1421);
nand U4770 (N_4770,In_2438,In_737);
or U4771 (N_4771,In_1466,In_1448);
xnor U4772 (N_4772,In_1844,In_2060);
or U4773 (N_4773,In_2022,In_2284);
nor U4774 (N_4774,In_1128,In_1015);
nand U4775 (N_4775,In_2390,In_1491);
nor U4776 (N_4776,In_2090,In_1566);
xor U4777 (N_4777,In_580,In_521);
or U4778 (N_4778,In_2080,In_1691);
nor U4779 (N_4779,In_379,In_168);
nand U4780 (N_4780,In_1202,In_363);
and U4781 (N_4781,In_590,In_1692);
nand U4782 (N_4782,In_506,In_1326);
or U4783 (N_4783,In_467,In_1989);
or U4784 (N_4784,In_1583,In_862);
xnor U4785 (N_4785,In_2165,In_684);
or U4786 (N_4786,In_1105,In_718);
nor U4787 (N_4787,In_764,In_132);
nand U4788 (N_4788,In_2256,In_997);
nor U4789 (N_4789,In_1826,In_2407);
or U4790 (N_4790,In_551,In_1033);
xnor U4791 (N_4791,In_1932,In_960);
and U4792 (N_4792,In_1235,In_2238);
nand U4793 (N_4793,In_1297,In_2179);
nor U4794 (N_4794,In_55,In_1532);
nor U4795 (N_4795,In_2318,In_302);
xnor U4796 (N_4796,In_1912,In_527);
or U4797 (N_4797,In_1134,In_0);
nand U4798 (N_4798,In_1455,In_1309);
nand U4799 (N_4799,In_285,In_527);
and U4800 (N_4800,In_1497,In_1578);
nand U4801 (N_4801,In_1887,In_208);
or U4802 (N_4802,In_265,In_1073);
nor U4803 (N_4803,In_995,In_351);
nor U4804 (N_4804,In_2035,In_1355);
nor U4805 (N_4805,In_1426,In_88);
or U4806 (N_4806,In_1349,In_1960);
xnor U4807 (N_4807,In_1355,In_2136);
or U4808 (N_4808,In_1839,In_1636);
or U4809 (N_4809,In_2042,In_74);
and U4810 (N_4810,In_200,In_651);
nor U4811 (N_4811,In_2370,In_1585);
and U4812 (N_4812,In_1516,In_408);
nand U4813 (N_4813,In_1322,In_728);
xnor U4814 (N_4814,In_826,In_1121);
and U4815 (N_4815,In_2477,In_1832);
xor U4816 (N_4816,In_1822,In_174);
xor U4817 (N_4817,In_2026,In_1185);
or U4818 (N_4818,In_1137,In_1711);
and U4819 (N_4819,In_429,In_2018);
or U4820 (N_4820,In_1700,In_1590);
and U4821 (N_4821,In_1479,In_2313);
nor U4822 (N_4822,In_1064,In_1447);
nand U4823 (N_4823,In_2010,In_535);
nand U4824 (N_4824,In_1418,In_1388);
or U4825 (N_4825,In_771,In_10);
or U4826 (N_4826,In_1581,In_1602);
or U4827 (N_4827,In_2489,In_2352);
and U4828 (N_4828,In_1603,In_2490);
or U4829 (N_4829,In_2262,In_1631);
or U4830 (N_4830,In_544,In_2281);
or U4831 (N_4831,In_1820,In_1929);
nor U4832 (N_4832,In_1660,In_559);
nor U4833 (N_4833,In_902,In_322);
or U4834 (N_4834,In_82,In_1753);
nand U4835 (N_4835,In_1796,In_1443);
xnor U4836 (N_4836,In_17,In_2182);
nor U4837 (N_4837,In_2307,In_968);
nor U4838 (N_4838,In_2051,In_206);
nand U4839 (N_4839,In_2135,In_629);
nor U4840 (N_4840,In_550,In_1821);
or U4841 (N_4841,In_1915,In_811);
nor U4842 (N_4842,In_1597,In_1596);
nor U4843 (N_4843,In_1465,In_678);
or U4844 (N_4844,In_1327,In_1613);
xor U4845 (N_4845,In_333,In_940);
nand U4846 (N_4846,In_978,In_2274);
or U4847 (N_4847,In_900,In_858);
nand U4848 (N_4848,In_387,In_1226);
xnor U4849 (N_4849,In_361,In_2311);
or U4850 (N_4850,In_1390,In_83);
nand U4851 (N_4851,In_1567,In_24);
nor U4852 (N_4852,In_2041,In_1834);
xnor U4853 (N_4853,In_1571,In_1178);
or U4854 (N_4854,In_2206,In_824);
or U4855 (N_4855,In_2471,In_1452);
xnor U4856 (N_4856,In_918,In_1791);
nand U4857 (N_4857,In_2027,In_1884);
nand U4858 (N_4858,In_119,In_1765);
nand U4859 (N_4859,In_1405,In_849);
nand U4860 (N_4860,In_1745,In_230);
xnor U4861 (N_4861,In_967,In_2423);
nor U4862 (N_4862,In_2113,In_1912);
and U4863 (N_4863,In_2464,In_2496);
xnor U4864 (N_4864,In_1372,In_1151);
xnor U4865 (N_4865,In_1088,In_139);
xor U4866 (N_4866,In_856,In_905);
nor U4867 (N_4867,In_2095,In_1026);
nand U4868 (N_4868,In_2203,In_1616);
xnor U4869 (N_4869,In_815,In_1453);
nor U4870 (N_4870,In_830,In_671);
nor U4871 (N_4871,In_855,In_1526);
nor U4872 (N_4872,In_1822,In_1762);
xor U4873 (N_4873,In_1032,In_1715);
and U4874 (N_4874,In_1880,In_2365);
xnor U4875 (N_4875,In_124,In_2153);
xor U4876 (N_4876,In_301,In_2080);
nand U4877 (N_4877,In_2022,In_1957);
xor U4878 (N_4878,In_1207,In_158);
nor U4879 (N_4879,In_1488,In_64);
nand U4880 (N_4880,In_2226,In_1194);
and U4881 (N_4881,In_1165,In_2451);
or U4882 (N_4882,In_718,In_2286);
xor U4883 (N_4883,In_1080,In_2031);
and U4884 (N_4884,In_1824,In_1053);
xnor U4885 (N_4885,In_994,In_1517);
nor U4886 (N_4886,In_1695,In_19);
nor U4887 (N_4887,In_1165,In_1648);
or U4888 (N_4888,In_2342,In_1723);
nor U4889 (N_4889,In_294,In_305);
or U4890 (N_4890,In_676,In_1638);
nor U4891 (N_4891,In_774,In_451);
xor U4892 (N_4892,In_2379,In_586);
and U4893 (N_4893,In_621,In_2140);
xor U4894 (N_4894,In_578,In_1637);
and U4895 (N_4895,In_1132,In_396);
nand U4896 (N_4896,In_1353,In_2340);
or U4897 (N_4897,In_31,In_1490);
nand U4898 (N_4898,In_409,In_1186);
or U4899 (N_4899,In_325,In_1900);
and U4900 (N_4900,In_348,In_2166);
nor U4901 (N_4901,In_1101,In_1177);
or U4902 (N_4902,In_1394,In_778);
xnor U4903 (N_4903,In_412,In_1015);
or U4904 (N_4904,In_1146,In_1469);
xor U4905 (N_4905,In_1772,In_1842);
nor U4906 (N_4906,In_736,In_520);
nor U4907 (N_4907,In_820,In_189);
and U4908 (N_4908,In_594,In_15);
and U4909 (N_4909,In_150,In_1798);
xnor U4910 (N_4910,In_240,In_1792);
xnor U4911 (N_4911,In_981,In_915);
and U4912 (N_4912,In_1564,In_387);
xnor U4913 (N_4913,In_1612,In_1410);
xor U4914 (N_4914,In_2369,In_447);
or U4915 (N_4915,In_410,In_1040);
nor U4916 (N_4916,In_2017,In_564);
nor U4917 (N_4917,In_1933,In_817);
xor U4918 (N_4918,In_2439,In_1419);
xnor U4919 (N_4919,In_980,In_2365);
and U4920 (N_4920,In_1156,In_2404);
xor U4921 (N_4921,In_170,In_692);
nand U4922 (N_4922,In_1277,In_1275);
nor U4923 (N_4923,In_1859,In_716);
nand U4924 (N_4924,In_863,In_438);
or U4925 (N_4925,In_908,In_918);
and U4926 (N_4926,In_2350,In_709);
xnor U4927 (N_4927,In_428,In_481);
nor U4928 (N_4928,In_1716,In_192);
xor U4929 (N_4929,In_32,In_2249);
nand U4930 (N_4930,In_1140,In_817);
xor U4931 (N_4931,In_2022,In_2244);
xor U4932 (N_4932,In_1690,In_1147);
and U4933 (N_4933,In_276,In_1558);
nor U4934 (N_4934,In_968,In_556);
or U4935 (N_4935,In_2106,In_1641);
nand U4936 (N_4936,In_612,In_2328);
xor U4937 (N_4937,In_1309,In_281);
nand U4938 (N_4938,In_663,In_1443);
nor U4939 (N_4939,In_1096,In_658);
nor U4940 (N_4940,In_1216,In_1238);
nand U4941 (N_4941,In_1641,In_1783);
nand U4942 (N_4942,In_819,In_666);
or U4943 (N_4943,In_1998,In_1882);
or U4944 (N_4944,In_442,In_2124);
nand U4945 (N_4945,In_495,In_2153);
and U4946 (N_4946,In_2349,In_99);
nand U4947 (N_4947,In_615,In_2302);
nor U4948 (N_4948,In_179,In_686);
or U4949 (N_4949,In_822,In_2005);
xor U4950 (N_4950,In_931,In_1070);
nor U4951 (N_4951,In_2309,In_116);
nor U4952 (N_4952,In_2223,In_1713);
xnor U4953 (N_4953,In_929,In_2352);
or U4954 (N_4954,In_1560,In_2344);
and U4955 (N_4955,In_1779,In_1975);
or U4956 (N_4956,In_1251,In_695);
xor U4957 (N_4957,In_504,In_509);
and U4958 (N_4958,In_2138,In_1211);
and U4959 (N_4959,In_86,In_2001);
xor U4960 (N_4960,In_279,In_1293);
nand U4961 (N_4961,In_2036,In_1539);
or U4962 (N_4962,In_2112,In_315);
and U4963 (N_4963,In_967,In_1924);
nand U4964 (N_4964,In_152,In_816);
or U4965 (N_4965,In_1348,In_1506);
xor U4966 (N_4966,In_403,In_1074);
xnor U4967 (N_4967,In_1904,In_324);
xnor U4968 (N_4968,In_1826,In_1568);
or U4969 (N_4969,In_445,In_1694);
nor U4970 (N_4970,In_645,In_1277);
xor U4971 (N_4971,In_1724,In_883);
nand U4972 (N_4972,In_2192,In_799);
xnor U4973 (N_4973,In_2263,In_2407);
or U4974 (N_4974,In_1060,In_2417);
nand U4975 (N_4975,In_1053,In_461);
or U4976 (N_4976,In_877,In_1082);
and U4977 (N_4977,In_1310,In_157);
nor U4978 (N_4978,In_186,In_1320);
nor U4979 (N_4979,In_72,In_205);
or U4980 (N_4980,In_383,In_2236);
xnor U4981 (N_4981,In_764,In_1635);
and U4982 (N_4982,In_216,In_1969);
or U4983 (N_4983,In_916,In_1501);
nor U4984 (N_4984,In_1822,In_577);
nand U4985 (N_4985,In_606,In_298);
nand U4986 (N_4986,In_882,In_390);
nand U4987 (N_4987,In_964,In_527);
and U4988 (N_4988,In_832,In_1912);
nand U4989 (N_4989,In_2433,In_232);
nand U4990 (N_4990,In_2438,In_999);
xor U4991 (N_4991,In_2184,In_2236);
or U4992 (N_4992,In_1574,In_908);
xnor U4993 (N_4993,In_1450,In_2482);
and U4994 (N_4994,In_1869,In_1069);
nor U4995 (N_4995,In_1798,In_1806);
and U4996 (N_4996,In_337,In_1508);
nor U4997 (N_4997,In_2452,In_183);
and U4998 (N_4998,In_817,In_1436);
nand U4999 (N_4999,In_2467,In_999);
xor U5000 (N_5000,In_835,In_1703);
nor U5001 (N_5001,In_911,In_1614);
and U5002 (N_5002,In_1060,In_1771);
and U5003 (N_5003,In_1806,In_1963);
nand U5004 (N_5004,In_104,In_938);
nor U5005 (N_5005,In_1341,In_1099);
xnor U5006 (N_5006,In_1951,In_1211);
nand U5007 (N_5007,In_1105,In_1390);
or U5008 (N_5008,In_2465,In_2188);
or U5009 (N_5009,In_731,In_2292);
xor U5010 (N_5010,In_2497,In_768);
xor U5011 (N_5011,In_605,In_57);
nor U5012 (N_5012,In_634,In_790);
or U5013 (N_5013,In_2413,In_2027);
nand U5014 (N_5014,In_662,In_618);
nor U5015 (N_5015,In_1612,In_2036);
xor U5016 (N_5016,In_346,In_594);
nand U5017 (N_5017,In_530,In_848);
and U5018 (N_5018,In_995,In_607);
xor U5019 (N_5019,In_1927,In_1677);
nand U5020 (N_5020,In_656,In_2292);
and U5021 (N_5021,In_1842,In_15);
nand U5022 (N_5022,In_716,In_1384);
or U5023 (N_5023,In_2251,In_2022);
xor U5024 (N_5024,In_666,In_1687);
nand U5025 (N_5025,In_569,In_416);
xnor U5026 (N_5026,In_2449,In_2448);
nand U5027 (N_5027,In_2293,In_1890);
nor U5028 (N_5028,In_2427,In_221);
nor U5029 (N_5029,In_1450,In_684);
xnor U5030 (N_5030,In_310,In_1438);
nand U5031 (N_5031,In_251,In_2135);
or U5032 (N_5032,In_1668,In_930);
nor U5033 (N_5033,In_1196,In_1165);
and U5034 (N_5034,In_1675,In_2201);
xor U5035 (N_5035,In_144,In_2355);
xnor U5036 (N_5036,In_2111,In_537);
nand U5037 (N_5037,In_1522,In_1414);
and U5038 (N_5038,In_1294,In_1039);
xor U5039 (N_5039,In_349,In_84);
nor U5040 (N_5040,In_221,In_1311);
xnor U5041 (N_5041,In_584,In_211);
nor U5042 (N_5042,In_2096,In_750);
nand U5043 (N_5043,In_1823,In_1084);
and U5044 (N_5044,In_272,In_1134);
or U5045 (N_5045,In_867,In_1756);
nand U5046 (N_5046,In_1626,In_271);
or U5047 (N_5047,In_629,In_1460);
and U5048 (N_5048,In_507,In_2168);
nand U5049 (N_5049,In_1870,In_795);
nand U5050 (N_5050,In_2363,In_1141);
and U5051 (N_5051,In_1320,In_1218);
nor U5052 (N_5052,In_667,In_1220);
nor U5053 (N_5053,In_441,In_1534);
and U5054 (N_5054,In_2475,In_1834);
or U5055 (N_5055,In_1602,In_2385);
and U5056 (N_5056,In_984,In_1334);
nor U5057 (N_5057,In_2109,In_2330);
nor U5058 (N_5058,In_523,In_2159);
nor U5059 (N_5059,In_1889,In_2119);
nand U5060 (N_5060,In_1580,In_110);
nand U5061 (N_5061,In_835,In_1188);
xnor U5062 (N_5062,In_1170,In_374);
and U5063 (N_5063,In_1814,In_2254);
nand U5064 (N_5064,In_508,In_2498);
nand U5065 (N_5065,In_1782,In_1895);
and U5066 (N_5066,In_375,In_1825);
nor U5067 (N_5067,In_1689,In_859);
and U5068 (N_5068,In_1360,In_1531);
xor U5069 (N_5069,In_30,In_1134);
and U5070 (N_5070,In_1714,In_1603);
or U5071 (N_5071,In_1332,In_228);
nand U5072 (N_5072,In_1454,In_1298);
xnor U5073 (N_5073,In_1027,In_511);
or U5074 (N_5074,In_1842,In_1722);
nand U5075 (N_5075,In_522,In_2259);
xnor U5076 (N_5076,In_1999,In_2169);
nand U5077 (N_5077,In_1010,In_982);
nor U5078 (N_5078,In_2318,In_2316);
or U5079 (N_5079,In_2031,In_1542);
and U5080 (N_5080,In_1191,In_1477);
and U5081 (N_5081,In_1522,In_537);
xnor U5082 (N_5082,In_774,In_569);
nand U5083 (N_5083,In_2243,In_19);
and U5084 (N_5084,In_396,In_1115);
and U5085 (N_5085,In_573,In_16);
or U5086 (N_5086,In_2408,In_1854);
nand U5087 (N_5087,In_1220,In_1541);
and U5088 (N_5088,In_1493,In_372);
xor U5089 (N_5089,In_880,In_998);
nor U5090 (N_5090,In_2095,In_29);
nor U5091 (N_5091,In_1531,In_2473);
or U5092 (N_5092,In_149,In_2268);
or U5093 (N_5093,In_2255,In_625);
xnor U5094 (N_5094,In_1539,In_93);
nor U5095 (N_5095,In_375,In_956);
nor U5096 (N_5096,In_521,In_1693);
xnor U5097 (N_5097,In_2040,In_2123);
nor U5098 (N_5098,In_346,In_1614);
and U5099 (N_5099,In_888,In_496);
or U5100 (N_5100,In_489,In_1840);
xor U5101 (N_5101,In_433,In_1242);
or U5102 (N_5102,In_360,In_67);
or U5103 (N_5103,In_1865,In_922);
xor U5104 (N_5104,In_1549,In_319);
or U5105 (N_5105,In_1090,In_370);
xor U5106 (N_5106,In_361,In_1064);
nor U5107 (N_5107,In_2476,In_2461);
xor U5108 (N_5108,In_2089,In_1010);
xnor U5109 (N_5109,In_890,In_1993);
and U5110 (N_5110,In_711,In_1098);
nor U5111 (N_5111,In_2483,In_726);
or U5112 (N_5112,In_124,In_2350);
nand U5113 (N_5113,In_481,In_1248);
and U5114 (N_5114,In_233,In_651);
xnor U5115 (N_5115,In_338,In_271);
nand U5116 (N_5116,In_948,In_142);
nand U5117 (N_5117,In_75,In_1832);
nor U5118 (N_5118,In_397,In_2016);
and U5119 (N_5119,In_1294,In_195);
and U5120 (N_5120,In_358,In_2250);
or U5121 (N_5121,In_852,In_729);
nand U5122 (N_5122,In_1067,In_635);
nand U5123 (N_5123,In_2455,In_1082);
and U5124 (N_5124,In_1383,In_1187);
or U5125 (N_5125,In_118,In_155);
and U5126 (N_5126,In_1539,In_1726);
or U5127 (N_5127,In_1155,In_2362);
nor U5128 (N_5128,In_110,In_2302);
nor U5129 (N_5129,In_26,In_757);
nand U5130 (N_5130,In_581,In_904);
nor U5131 (N_5131,In_1492,In_1887);
nor U5132 (N_5132,In_2256,In_2037);
or U5133 (N_5133,In_1592,In_863);
nand U5134 (N_5134,In_480,In_1619);
xor U5135 (N_5135,In_2443,In_2447);
xor U5136 (N_5136,In_635,In_69);
nand U5137 (N_5137,In_2330,In_24);
nor U5138 (N_5138,In_2114,In_1);
or U5139 (N_5139,In_301,In_147);
xor U5140 (N_5140,In_106,In_386);
xnor U5141 (N_5141,In_1353,In_926);
and U5142 (N_5142,In_445,In_307);
xnor U5143 (N_5143,In_1786,In_1958);
nor U5144 (N_5144,In_639,In_331);
and U5145 (N_5145,In_945,In_1590);
xnor U5146 (N_5146,In_773,In_2389);
and U5147 (N_5147,In_582,In_2403);
nand U5148 (N_5148,In_23,In_1325);
or U5149 (N_5149,In_142,In_2216);
xor U5150 (N_5150,In_1314,In_2145);
nor U5151 (N_5151,In_967,In_1213);
nor U5152 (N_5152,In_856,In_319);
and U5153 (N_5153,In_1296,In_1385);
nand U5154 (N_5154,In_2099,In_1384);
xnor U5155 (N_5155,In_6,In_1791);
or U5156 (N_5156,In_14,In_595);
nor U5157 (N_5157,In_2341,In_522);
nor U5158 (N_5158,In_1201,In_2300);
or U5159 (N_5159,In_110,In_1029);
or U5160 (N_5160,In_2306,In_1091);
nand U5161 (N_5161,In_518,In_32);
xnor U5162 (N_5162,In_1604,In_2423);
nand U5163 (N_5163,In_2222,In_1503);
nor U5164 (N_5164,In_2180,In_2241);
and U5165 (N_5165,In_1421,In_2158);
nand U5166 (N_5166,In_1764,In_2188);
nor U5167 (N_5167,In_1817,In_334);
or U5168 (N_5168,In_257,In_1805);
nor U5169 (N_5169,In_1020,In_2081);
nand U5170 (N_5170,In_323,In_1286);
nor U5171 (N_5171,In_712,In_1786);
nor U5172 (N_5172,In_1283,In_645);
or U5173 (N_5173,In_1310,In_1358);
xnor U5174 (N_5174,In_303,In_995);
and U5175 (N_5175,In_683,In_201);
or U5176 (N_5176,In_2016,In_294);
and U5177 (N_5177,In_1058,In_2492);
or U5178 (N_5178,In_1441,In_1733);
or U5179 (N_5179,In_542,In_1217);
or U5180 (N_5180,In_1944,In_904);
or U5181 (N_5181,In_1391,In_1515);
and U5182 (N_5182,In_1045,In_293);
xnor U5183 (N_5183,In_2385,In_342);
and U5184 (N_5184,In_1408,In_1409);
xnor U5185 (N_5185,In_1989,In_259);
or U5186 (N_5186,In_950,In_2344);
xnor U5187 (N_5187,In_2030,In_1034);
xnor U5188 (N_5188,In_1781,In_1770);
nor U5189 (N_5189,In_650,In_1766);
xnor U5190 (N_5190,In_1081,In_312);
nand U5191 (N_5191,In_505,In_1004);
nor U5192 (N_5192,In_2133,In_661);
and U5193 (N_5193,In_1779,In_51);
nor U5194 (N_5194,In_546,In_1798);
xor U5195 (N_5195,In_139,In_909);
nand U5196 (N_5196,In_1529,In_1447);
nand U5197 (N_5197,In_1221,In_2350);
nand U5198 (N_5198,In_1872,In_749);
or U5199 (N_5199,In_408,In_2419);
nand U5200 (N_5200,In_276,In_1467);
or U5201 (N_5201,In_1932,In_594);
and U5202 (N_5202,In_2459,In_1597);
and U5203 (N_5203,In_1217,In_735);
and U5204 (N_5204,In_1924,In_703);
nand U5205 (N_5205,In_91,In_1494);
nand U5206 (N_5206,In_438,In_1380);
xnor U5207 (N_5207,In_521,In_953);
xnor U5208 (N_5208,In_256,In_2151);
nand U5209 (N_5209,In_1519,In_536);
or U5210 (N_5210,In_360,In_1423);
nor U5211 (N_5211,In_1589,In_911);
or U5212 (N_5212,In_1327,In_2124);
or U5213 (N_5213,In_1222,In_1106);
nand U5214 (N_5214,In_338,In_545);
nor U5215 (N_5215,In_2039,In_609);
or U5216 (N_5216,In_654,In_672);
nor U5217 (N_5217,In_1716,In_1108);
xnor U5218 (N_5218,In_1660,In_735);
xor U5219 (N_5219,In_882,In_1431);
nor U5220 (N_5220,In_2347,In_1507);
xor U5221 (N_5221,In_1225,In_923);
and U5222 (N_5222,In_1372,In_1699);
xor U5223 (N_5223,In_1756,In_1472);
nor U5224 (N_5224,In_1519,In_1677);
and U5225 (N_5225,In_777,In_924);
and U5226 (N_5226,In_1205,In_51);
xnor U5227 (N_5227,In_1884,In_382);
nand U5228 (N_5228,In_93,In_442);
or U5229 (N_5229,In_1049,In_2469);
xnor U5230 (N_5230,In_2075,In_1092);
or U5231 (N_5231,In_1023,In_1795);
nor U5232 (N_5232,In_2168,In_797);
or U5233 (N_5233,In_94,In_1976);
xor U5234 (N_5234,In_2245,In_2106);
or U5235 (N_5235,In_1806,In_721);
and U5236 (N_5236,In_666,In_2287);
and U5237 (N_5237,In_1530,In_839);
or U5238 (N_5238,In_2197,In_1346);
nand U5239 (N_5239,In_1755,In_1126);
xor U5240 (N_5240,In_1205,In_1642);
nand U5241 (N_5241,In_1566,In_240);
nand U5242 (N_5242,In_305,In_885);
or U5243 (N_5243,In_1158,In_127);
and U5244 (N_5244,In_1265,In_1078);
nand U5245 (N_5245,In_612,In_56);
nor U5246 (N_5246,In_51,In_1960);
or U5247 (N_5247,In_899,In_1793);
and U5248 (N_5248,In_792,In_1521);
or U5249 (N_5249,In_2487,In_1490);
xor U5250 (N_5250,In_8,In_261);
nor U5251 (N_5251,In_2075,In_433);
nand U5252 (N_5252,In_1041,In_2408);
xnor U5253 (N_5253,In_2482,In_300);
nand U5254 (N_5254,In_1493,In_427);
nand U5255 (N_5255,In_1641,In_1873);
and U5256 (N_5256,In_1333,In_2071);
xnor U5257 (N_5257,In_2042,In_1193);
and U5258 (N_5258,In_1133,In_1679);
or U5259 (N_5259,In_2180,In_197);
nor U5260 (N_5260,In_2331,In_1025);
nand U5261 (N_5261,In_1454,In_2139);
or U5262 (N_5262,In_18,In_1641);
and U5263 (N_5263,In_68,In_651);
xor U5264 (N_5264,In_2147,In_1699);
nor U5265 (N_5265,In_400,In_67);
or U5266 (N_5266,In_1571,In_1937);
and U5267 (N_5267,In_53,In_1345);
or U5268 (N_5268,In_1668,In_2342);
or U5269 (N_5269,In_1801,In_1874);
nand U5270 (N_5270,In_1406,In_1909);
nor U5271 (N_5271,In_173,In_2466);
or U5272 (N_5272,In_1606,In_1802);
nand U5273 (N_5273,In_1126,In_1897);
nor U5274 (N_5274,In_146,In_1991);
xnor U5275 (N_5275,In_1120,In_1865);
or U5276 (N_5276,In_656,In_1470);
xnor U5277 (N_5277,In_397,In_1318);
nand U5278 (N_5278,In_219,In_160);
or U5279 (N_5279,In_1643,In_2013);
and U5280 (N_5280,In_77,In_1644);
nor U5281 (N_5281,In_951,In_2261);
nor U5282 (N_5282,In_2223,In_852);
or U5283 (N_5283,In_1728,In_1148);
or U5284 (N_5284,In_801,In_654);
nand U5285 (N_5285,In_1717,In_2263);
xnor U5286 (N_5286,In_738,In_213);
nor U5287 (N_5287,In_93,In_2374);
xor U5288 (N_5288,In_1732,In_2326);
xor U5289 (N_5289,In_2175,In_1469);
nor U5290 (N_5290,In_202,In_414);
or U5291 (N_5291,In_912,In_358);
nand U5292 (N_5292,In_2473,In_1013);
or U5293 (N_5293,In_1725,In_2250);
and U5294 (N_5294,In_1565,In_163);
nor U5295 (N_5295,In_1423,In_1980);
or U5296 (N_5296,In_16,In_1650);
xnor U5297 (N_5297,In_43,In_583);
xnor U5298 (N_5298,In_1909,In_822);
nand U5299 (N_5299,In_690,In_533);
and U5300 (N_5300,In_1862,In_1873);
and U5301 (N_5301,In_2244,In_972);
nor U5302 (N_5302,In_1640,In_2206);
and U5303 (N_5303,In_1037,In_15);
nand U5304 (N_5304,In_450,In_761);
nor U5305 (N_5305,In_1309,In_2419);
nor U5306 (N_5306,In_229,In_766);
nand U5307 (N_5307,In_1723,In_2288);
xnor U5308 (N_5308,In_872,In_1758);
and U5309 (N_5309,In_981,In_526);
xor U5310 (N_5310,In_1242,In_1608);
nand U5311 (N_5311,In_204,In_937);
xnor U5312 (N_5312,In_2028,In_1529);
and U5313 (N_5313,In_975,In_2410);
xnor U5314 (N_5314,In_221,In_1691);
or U5315 (N_5315,In_1328,In_2139);
xnor U5316 (N_5316,In_1037,In_590);
nand U5317 (N_5317,In_919,In_2040);
and U5318 (N_5318,In_2399,In_459);
nor U5319 (N_5319,In_976,In_181);
and U5320 (N_5320,In_676,In_1980);
nand U5321 (N_5321,In_1697,In_1951);
nor U5322 (N_5322,In_34,In_273);
and U5323 (N_5323,In_2089,In_1541);
and U5324 (N_5324,In_1697,In_122);
nand U5325 (N_5325,In_1926,In_1745);
or U5326 (N_5326,In_617,In_70);
or U5327 (N_5327,In_1081,In_541);
and U5328 (N_5328,In_899,In_1208);
nand U5329 (N_5329,In_1424,In_985);
nor U5330 (N_5330,In_431,In_1285);
nor U5331 (N_5331,In_2133,In_1817);
or U5332 (N_5332,In_116,In_559);
nand U5333 (N_5333,In_974,In_163);
or U5334 (N_5334,In_1148,In_2172);
nand U5335 (N_5335,In_2302,In_2024);
xor U5336 (N_5336,In_2492,In_2423);
xor U5337 (N_5337,In_1301,In_1862);
xnor U5338 (N_5338,In_448,In_1829);
nand U5339 (N_5339,In_238,In_1738);
nand U5340 (N_5340,In_1778,In_1173);
nand U5341 (N_5341,In_1118,In_1134);
and U5342 (N_5342,In_1570,In_819);
nor U5343 (N_5343,In_128,In_2215);
or U5344 (N_5344,In_1062,In_762);
xor U5345 (N_5345,In_2404,In_727);
xnor U5346 (N_5346,In_1993,In_2489);
xor U5347 (N_5347,In_2441,In_1050);
nor U5348 (N_5348,In_1716,In_1810);
nor U5349 (N_5349,In_1318,In_1528);
and U5350 (N_5350,In_1677,In_1081);
or U5351 (N_5351,In_1156,In_919);
nor U5352 (N_5352,In_747,In_651);
xor U5353 (N_5353,In_268,In_17);
and U5354 (N_5354,In_241,In_1467);
xnor U5355 (N_5355,In_1252,In_1311);
and U5356 (N_5356,In_2231,In_462);
nand U5357 (N_5357,In_704,In_1278);
and U5358 (N_5358,In_2244,In_110);
nor U5359 (N_5359,In_701,In_2422);
nand U5360 (N_5360,In_364,In_1290);
and U5361 (N_5361,In_2393,In_1259);
xnor U5362 (N_5362,In_197,In_1614);
nor U5363 (N_5363,In_3,In_2137);
nor U5364 (N_5364,In_15,In_414);
xnor U5365 (N_5365,In_1566,In_1431);
nor U5366 (N_5366,In_1061,In_956);
nor U5367 (N_5367,In_1493,In_926);
xnor U5368 (N_5368,In_2344,In_1602);
and U5369 (N_5369,In_2350,In_1005);
nor U5370 (N_5370,In_492,In_2416);
nor U5371 (N_5371,In_2023,In_1243);
and U5372 (N_5372,In_1341,In_924);
xor U5373 (N_5373,In_1636,In_2305);
and U5374 (N_5374,In_1098,In_1572);
nand U5375 (N_5375,In_1998,In_2058);
nand U5376 (N_5376,In_2435,In_2419);
xor U5377 (N_5377,In_1048,In_2316);
nor U5378 (N_5378,In_371,In_1436);
xor U5379 (N_5379,In_2202,In_347);
nor U5380 (N_5380,In_2462,In_476);
nand U5381 (N_5381,In_134,In_1529);
and U5382 (N_5382,In_1528,In_1305);
or U5383 (N_5383,In_2287,In_1196);
xor U5384 (N_5384,In_763,In_2199);
or U5385 (N_5385,In_719,In_1110);
nand U5386 (N_5386,In_1636,In_1524);
nor U5387 (N_5387,In_2385,In_1019);
and U5388 (N_5388,In_1017,In_1894);
or U5389 (N_5389,In_2010,In_1333);
nor U5390 (N_5390,In_1619,In_1002);
nand U5391 (N_5391,In_1785,In_445);
nand U5392 (N_5392,In_159,In_862);
xnor U5393 (N_5393,In_958,In_1567);
nand U5394 (N_5394,In_2358,In_1293);
nand U5395 (N_5395,In_1974,In_2073);
xor U5396 (N_5396,In_361,In_749);
and U5397 (N_5397,In_288,In_1439);
and U5398 (N_5398,In_1167,In_1188);
xnor U5399 (N_5399,In_561,In_1882);
and U5400 (N_5400,In_482,In_2444);
or U5401 (N_5401,In_1036,In_760);
and U5402 (N_5402,In_1878,In_356);
xnor U5403 (N_5403,In_2190,In_633);
and U5404 (N_5404,In_952,In_1024);
or U5405 (N_5405,In_1304,In_939);
nor U5406 (N_5406,In_1347,In_2108);
nor U5407 (N_5407,In_1906,In_1843);
nand U5408 (N_5408,In_1477,In_255);
or U5409 (N_5409,In_2267,In_792);
and U5410 (N_5410,In_970,In_1784);
nor U5411 (N_5411,In_1886,In_907);
nor U5412 (N_5412,In_949,In_1253);
and U5413 (N_5413,In_1241,In_1494);
xor U5414 (N_5414,In_2463,In_2136);
xor U5415 (N_5415,In_1596,In_2126);
xnor U5416 (N_5416,In_1981,In_314);
and U5417 (N_5417,In_433,In_678);
xor U5418 (N_5418,In_1997,In_43);
and U5419 (N_5419,In_546,In_2201);
xor U5420 (N_5420,In_2454,In_1388);
xor U5421 (N_5421,In_1250,In_1764);
nor U5422 (N_5422,In_2270,In_1894);
or U5423 (N_5423,In_2341,In_923);
xnor U5424 (N_5424,In_1526,In_786);
xor U5425 (N_5425,In_1458,In_639);
nor U5426 (N_5426,In_2375,In_908);
nand U5427 (N_5427,In_1717,In_2045);
and U5428 (N_5428,In_1626,In_837);
and U5429 (N_5429,In_2382,In_128);
or U5430 (N_5430,In_1031,In_441);
xor U5431 (N_5431,In_2396,In_2479);
nor U5432 (N_5432,In_2491,In_2293);
or U5433 (N_5433,In_291,In_1610);
xnor U5434 (N_5434,In_1729,In_1057);
or U5435 (N_5435,In_539,In_729);
xor U5436 (N_5436,In_2309,In_54);
xor U5437 (N_5437,In_1763,In_236);
nand U5438 (N_5438,In_503,In_1805);
xnor U5439 (N_5439,In_427,In_439);
nand U5440 (N_5440,In_2482,In_2259);
nand U5441 (N_5441,In_973,In_338);
or U5442 (N_5442,In_367,In_2133);
and U5443 (N_5443,In_1998,In_2180);
or U5444 (N_5444,In_2260,In_2154);
or U5445 (N_5445,In_569,In_1287);
nor U5446 (N_5446,In_270,In_411);
xor U5447 (N_5447,In_1874,In_1843);
nand U5448 (N_5448,In_665,In_2484);
and U5449 (N_5449,In_1213,In_2471);
nand U5450 (N_5450,In_1713,In_1393);
nor U5451 (N_5451,In_208,In_621);
or U5452 (N_5452,In_443,In_992);
nor U5453 (N_5453,In_623,In_1962);
nand U5454 (N_5454,In_1725,In_582);
and U5455 (N_5455,In_658,In_52);
xnor U5456 (N_5456,In_244,In_1485);
or U5457 (N_5457,In_245,In_463);
nor U5458 (N_5458,In_1696,In_43);
xnor U5459 (N_5459,In_1584,In_104);
or U5460 (N_5460,In_298,In_1325);
or U5461 (N_5461,In_1643,In_928);
nor U5462 (N_5462,In_821,In_818);
nor U5463 (N_5463,In_1664,In_1852);
nand U5464 (N_5464,In_1783,In_1850);
nor U5465 (N_5465,In_155,In_263);
nand U5466 (N_5466,In_2115,In_1239);
nand U5467 (N_5467,In_244,In_1758);
xnor U5468 (N_5468,In_798,In_2097);
xnor U5469 (N_5469,In_2161,In_324);
nand U5470 (N_5470,In_938,In_2350);
and U5471 (N_5471,In_1572,In_896);
or U5472 (N_5472,In_688,In_1317);
nor U5473 (N_5473,In_2235,In_1527);
and U5474 (N_5474,In_2068,In_1372);
nor U5475 (N_5475,In_1953,In_2185);
and U5476 (N_5476,In_1086,In_1459);
xor U5477 (N_5477,In_1336,In_1897);
and U5478 (N_5478,In_1843,In_2378);
nor U5479 (N_5479,In_1989,In_831);
xnor U5480 (N_5480,In_163,In_1426);
nand U5481 (N_5481,In_1291,In_119);
or U5482 (N_5482,In_2417,In_78);
xor U5483 (N_5483,In_478,In_964);
and U5484 (N_5484,In_1788,In_1931);
or U5485 (N_5485,In_815,In_388);
nor U5486 (N_5486,In_1736,In_372);
xnor U5487 (N_5487,In_1139,In_244);
or U5488 (N_5488,In_2,In_1836);
nand U5489 (N_5489,In_487,In_2154);
xor U5490 (N_5490,In_2328,In_2044);
nor U5491 (N_5491,In_535,In_1400);
or U5492 (N_5492,In_1206,In_488);
and U5493 (N_5493,In_1764,In_1772);
nor U5494 (N_5494,In_1988,In_1540);
nor U5495 (N_5495,In_1710,In_977);
or U5496 (N_5496,In_2460,In_811);
nand U5497 (N_5497,In_1718,In_2113);
nor U5498 (N_5498,In_248,In_75);
or U5499 (N_5499,In_766,In_668);
or U5500 (N_5500,In_1737,In_1996);
nor U5501 (N_5501,In_1997,In_1627);
xor U5502 (N_5502,In_676,In_922);
nand U5503 (N_5503,In_1490,In_959);
nand U5504 (N_5504,In_174,In_902);
and U5505 (N_5505,In_1886,In_2268);
or U5506 (N_5506,In_1641,In_386);
xnor U5507 (N_5507,In_1312,In_1199);
nand U5508 (N_5508,In_782,In_1740);
nand U5509 (N_5509,In_2346,In_268);
nand U5510 (N_5510,In_2425,In_2294);
or U5511 (N_5511,In_1303,In_1067);
nand U5512 (N_5512,In_2451,In_1449);
or U5513 (N_5513,In_2426,In_817);
nand U5514 (N_5514,In_90,In_1835);
and U5515 (N_5515,In_1798,In_559);
nor U5516 (N_5516,In_297,In_1717);
xor U5517 (N_5517,In_267,In_1518);
nand U5518 (N_5518,In_853,In_106);
or U5519 (N_5519,In_2232,In_83);
or U5520 (N_5520,In_23,In_232);
and U5521 (N_5521,In_1219,In_1567);
nor U5522 (N_5522,In_2113,In_1186);
nor U5523 (N_5523,In_658,In_454);
nand U5524 (N_5524,In_1167,In_2414);
xnor U5525 (N_5525,In_1879,In_1287);
nor U5526 (N_5526,In_1627,In_528);
xnor U5527 (N_5527,In_1782,In_464);
and U5528 (N_5528,In_1672,In_86);
or U5529 (N_5529,In_1914,In_2471);
and U5530 (N_5530,In_2493,In_970);
nand U5531 (N_5531,In_1364,In_1507);
nor U5532 (N_5532,In_1714,In_1819);
nand U5533 (N_5533,In_703,In_401);
nor U5534 (N_5534,In_1038,In_1234);
xnor U5535 (N_5535,In_1386,In_445);
or U5536 (N_5536,In_2399,In_718);
or U5537 (N_5537,In_1800,In_2073);
xor U5538 (N_5538,In_1992,In_2284);
nand U5539 (N_5539,In_960,In_612);
or U5540 (N_5540,In_1985,In_1480);
nand U5541 (N_5541,In_299,In_1240);
or U5542 (N_5542,In_844,In_2348);
or U5543 (N_5543,In_818,In_52);
and U5544 (N_5544,In_1399,In_1065);
and U5545 (N_5545,In_966,In_1661);
nor U5546 (N_5546,In_1845,In_1039);
nand U5547 (N_5547,In_2311,In_1367);
and U5548 (N_5548,In_375,In_1154);
nand U5549 (N_5549,In_1118,In_2030);
and U5550 (N_5550,In_2075,In_2378);
and U5551 (N_5551,In_2228,In_970);
nand U5552 (N_5552,In_1352,In_2349);
nor U5553 (N_5553,In_1713,In_1002);
nor U5554 (N_5554,In_2075,In_199);
xor U5555 (N_5555,In_609,In_842);
or U5556 (N_5556,In_1384,In_1783);
or U5557 (N_5557,In_1452,In_1557);
nor U5558 (N_5558,In_372,In_668);
nand U5559 (N_5559,In_534,In_1598);
nand U5560 (N_5560,In_144,In_2409);
or U5561 (N_5561,In_2147,In_517);
nand U5562 (N_5562,In_1231,In_88);
xnor U5563 (N_5563,In_2019,In_1037);
nor U5564 (N_5564,In_1807,In_1450);
or U5565 (N_5565,In_1066,In_944);
or U5566 (N_5566,In_2052,In_44);
nand U5567 (N_5567,In_305,In_1362);
xnor U5568 (N_5568,In_1463,In_405);
nand U5569 (N_5569,In_1487,In_1406);
and U5570 (N_5570,In_1739,In_310);
xor U5571 (N_5571,In_114,In_265);
xnor U5572 (N_5572,In_91,In_519);
nor U5573 (N_5573,In_1036,In_2310);
xor U5574 (N_5574,In_2113,In_1685);
xnor U5575 (N_5575,In_618,In_596);
nor U5576 (N_5576,In_975,In_1354);
nand U5577 (N_5577,In_1300,In_940);
nor U5578 (N_5578,In_1627,In_1827);
xnor U5579 (N_5579,In_420,In_274);
xor U5580 (N_5580,In_1924,In_741);
or U5581 (N_5581,In_780,In_2077);
xor U5582 (N_5582,In_2177,In_318);
nor U5583 (N_5583,In_876,In_709);
and U5584 (N_5584,In_934,In_188);
xor U5585 (N_5585,In_884,In_198);
or U5586 (N_5586,In_82,In_1047);
nand U5587 (N_5587,In_1994,In_302);
and U5588 (N_5588,In_317,In_2445);
or U5589 (N_5589,In_2376,In_703);
or U5590 (N_5590,In_988,In_287);
nor U5591 (N_5591,In_520,In_1477);
xnor U5592 (N_5592,In_1150,In_2169);
or U5593 (N_5593,In_2299,In_1975);
or U5594 (N_5594,In_1526,In_1914);
or U5595 (N_5595,In_1414,In_160);
and U5596 (N_5596,In_491,In_1252);
or U5597 (N_5597,In_1739,In_2377);
nand U5598 (N_5598,In_702,In_1087);
and U5599 (N_5599,In_2352,In_2311);
or U5600 (N_5600,In_47,In_1541);
and U5601 (N_5601,In_1054,In_933);
and U5602 (N_5602,In_2394,In_2281);
and U5603 (N_5603,In_589,In_2251);
nor U5604 (N_5604,In_2151,In_1805);
or U5605 (N_5605,In_652,In_362);
xnor U5606 (N_5606,In_2372,In_646);
xor U5607 (N_5607,In_194,In_2424);
nor U5608 (N_5608,In_697,In_1569);
nand U5609 (N_5609,In_963,In_1870);
nand U5610 (N_5610,In_1194,In_1565);
or U5611 (N_5611,In_1311,In_174);
xnor U5612 (N_5612,In_1816,In_1920);
nor U5613 (N_5613,In_1120,In_1038);
or U5614 (N_5614,In_71,In_647);
and U5615 (N_5615,In_289,In_499);
xor U5616 (N_5616,In_1862,In_766);
xnor U5617 (N_5617,In_1970,In_1297);
or U5618 (N_5618,In_13,In_1747);
or U5619 (N_5619,In_2286,In_998);
xnor U5620 (N_5620,In_1844,In_1958);
xnor U5621 (N_5621,In_508,In_2042);
or U5622 (N_5622,In_1221,In_1964);
nand U5623 (N_5623,In_1097,In_2212);
xor U5624 (N_5624,In_1502,In_2229);
nand U5625 (N_5625,In_126,In_2292);
xnor U5626 (N_5626,In_1187,In_1924);
nor U5627 (N_5627,In_67,In_2011);
nor U5628 (N_5628,In_1094,In_872);
nand U5629 (N_5629,In_480,In_814);
nor U5630 (N_5630,In_2118,In_1077);
and U5631 (N_5631,In_382,In_1990);
nor U5632 (N_5632,In_2488,In_1642);
nor U5633 (N_5633,In_1416,In_1984);
nor U5634 (N_5634,In_814,In_2185);
nor U5635 (N_5635,In_412,In_2112);
and U5636 (N_5636,In_1481,In_1879);
nor U5637 (N_5637,In_1245,In_1446);
xnor U5638 (N_5638,In_341,In_33);
nand U5639 (N_5639,In_662,In_2299);
xnor U5640 (N_5640,In_760,In_2296);
or U5641 (N_5641,In_2222,In_2189);
xnor U5642 (N_5642,In_149,In_996);
nor U5643 (N_5643,In_1573,In_672);
xor U5644 (N_5644,In_2079,In_554);
nor U5645 (N_5645,In_430,In_1912);
nand U5646 (N_5646,In_579,In_2295);
nand U5647 (N_5647,In_2192,In_842);
nor U5648 (N_5648,In_879,In_496);
xnor U5649 (N_5649,In_1141,In_407);
nor U5650 (N_5650,In_515,In_1342);
or U5651 (N_5651,In_1198,In_1825);
nor U5652 (N_5652,In_2374,In_2195);
nand U5653 (N_5653,In_1156,In_1675);
nand U5654 (N_5654,In_2300,In_1925);
nand U5655 (N_5655,In_1106,In_1771);
nand U5656 (N_5656,In_1331,In_2341);
nor U5657 (N_5657,In_1345,In_1119);
nand U5658 (N_5658,In_1986,In_1999);
xor U5659 (N_5659,In_270,In_1497);
and U5660 (N_5660,In_230,In_25);
nand U5661 (N_5661,In_2293,In_1915);
xnor U5662 (N_5662,In_2089,In_364);
nor U5663 (N_5663,In_1309,In_1966);
xnor U5664 (N_5664,In_383,In_300);
and U5665 (N_5665,In_1699,In_1082);
or U5666 (N_5666,In_868,In_2389);
nand U5667 (N_5667,In_547,In_2108);
nand U5668 (N_5668,In_1351,In_458);
and U5669 (N_5669,In_1011,In_996);
nor U5670 (N_5670,In_1888,In_1766);
and U5671 (N_5671,In_2405,In_971);
xnor U5672 (N_5672,In_1955,In_2040);
nand U5673 (N_5673,In_1342,In_1994);
xnor U5674 (N_5674,In_1782,In_1515);
and U5675 (N_5675,In_1349,In_815);
or U5676 (N_5676,In_1996,In_1645);
xor U5677 (N_5677,In_958,In_1672);
nor U5678 (N_5678,In_1881,In_2077);
nor U5679 (N_5679,In_2232,In_876);
nor U5680 (N_5680,In_1352,In_2486);
xnor U5681 (N_5681,In_2145,In_542);
and U5682 (N_5682,In_875,In_63);
nor U5683 (N_5683,In_2273,In_1933);
or U5684 (N_5684,In_2214,In_2430);
and U5685 (N_5685,In_133,In_789);
and U5686 (N_5686,In_1918,In_1320);
xnor U5687 (N_5687,In_928,In_1838);
and U5688 (N_5688,In_1120,In_1221);
nand U5689 (N_5689,In_2083,In_2375);
or U5690 (N_5690,In_1466,In_897);
nand U5691 (N_5691,In_582,In_1443);
xor U5692 (N_5692,In_884,In_488);
nand U5693 (N_5693,In_199,In_1967);
nor U5694 (N_5694,In_83,In_2133);
or U5695 (N_5695,In_2479,In_998);
and U5696 (N_5696,In_2256,In_399);
or U5697 (N_5697,In_2078,In_1003);
nor U5698 (N_5698,In_2240,In_1587);
nand U5699 (N_5699,In_245,In_319);
nor U5700 (N_5700,In_2116,In_1602);
or U5701 (N_5701,In_1171,In_2316);
or U5702 (N_5702,In_732,In_759);
xor U5703 (N_5703,In_1672,In_2025);
xnor U5704 (N_5704,In_263,In_2388);
xor U5705 (N_5705,In_961,In_421);
and U5706 (N_5706,In_1287,In_1718);
or U5707 (N_5707,In_1631,In_119);
nand U5708 (N_5708,In_199,In_1161);
xnor U5709 (N_5709,In_500,In_468);
or U5710 (N_5710,In_237,In_2162);
and U5711 (N_5711,In_2064,In_2198);
nor U5712 (N_5712,In_2094,In_767);
xnor U5713 (N_5713,In_129,In_2022);
nand U5714 (N_5714,In_917,In_1603);
nor U5715 (N_5715,In_1363,In_1516);
nor U5716 (N_5716,In_662,In_1380);
xor U5717 (N_5717,In_2203,In_2444);
nand U5718 (N_5718,In_1087,In_190);
or U5719 (N_5719,In_1829,In_1080);
nand U5720 (N_5720,In_1618,In_1917);
or U5721 (N_5721,In_1413,In_1241);
nor U5722 (N_5722,In_2332,In_1319);
nor U5723 (N_5723,In_551,In_736);
and U5724 (N_5724,In_2387,In_590);
nor U5725 (N_5725,In_228,In_680);
nor U5726 (N_5726,In_953,In_2409);
nor U5727 (N_5727,In_560,In_1451);
nand U5728 (N_5728,In_8,In_607);
or U5729 (N_5729,In_1486,In_918);
nand U5730 (N_5730,In_454,In_971);
xnor U5731 (N_5731,In_1906,In_1760);
nand U5732 (N_5732,In_1040,In_323);
nand U5733 (N_5733,In_1958,In_923);
nand U5734 (N_5734,In_1927,In_823);
nand U5735 (N_5735,In_2252,In_908);
xnor U5736 (N_5736,In_1296,In_536);
nor U5737 (N_5737,In_2149,In_1427);
and U5738 (N_5738,In_2228,In_559);
nand U5739 (N_5739,In_1656,In_1928);
and U5740 (N_5740,In_1766,In_1141);
nand U5741 (N_5741,In_1318,In_34);
or U5742 (N_5742,In_2388,In_434);
nand U5743 (N_5743,In_1996,In_505);
nand U5744 (N_5744,In_1608,In_2016);
nor U5745 (N_5745,In_553,In_328);
and U5746 (N_5746,In_1733,In_159);
or U5747 (N_5747,In_937,In_135);
nand U5748 (N_5748,In_910,In_265);
nor U5749 (N_5749,In_1961,In_367);
and U5750 (N_5750,In_520,In_1918);
nor U5751 (N_5751,In_616,In_505);
nor U5752 (N_5752,In_815,In_2287);
and U5753 (N_5753,In_724,In_2116);
nand U5754 (N_5754,In_96,In_2280);
or U5755 (N_5755,In_123,In_2443);
xnor U5756 (N_5756,In_232,In_622);
or U5757 (N_5757,In_2312,In_702);
or U5758 (N_5758,In_461,In_362);
or U5759 (N_5759,In_163,In_172);
nor U5760 (N_5760,In_409,In_2151);
and U5761 (N_5761,In_2218,In_1798);
and U5762 (N_5762,In_1657,In_1464);
nand U5763 (N_5763,In_781,In_2334);
nor U5764 (N_5764,In_1831,In_2378);
or U5765 (N_5765,In_1926,In_2280);
or U5766 (N_5766,In_887,In_174);
xnor U5767 (N_5767,In_1698,In_2247);
nor U5768 (N_5768,In_2365,In_598);
xor U5769 (N_5769,In_638,In_1007);
or U5770 (N_5770,In_1314,In_1697);
xor U5771 (N_5771,In_2318,In_2428);
xor U5772 (N_5772,In_1282,In_638);
xor U5773 (N_5773,In_1281,In_832);
or U5774 (N_5774,In_483,In_673);
nor U5775 (N_5775,In_409,In_2429);
nand U5776 (N_5776,In_897,In_977);
and U5777 (N_5777,In_2121,In_1339);
nand U5778 (N_5778,In_895,In_2177);
and U5779 (N_5779,In_1575,In_2267);
or U5780 (N_5780,In_1926,In_1357);
nor U5781 (N_5781,In_2263,In_771);
nand U5782 (N_5782,In_504,In_331);
xnor U5783 (N_5783,In_1204,In_1078);
and U5784 (N_5784,In_2171,In_283);
nand U5785 (N_5785,In_1944,In_1075);
and U5786 (N_5786,In_2218,In_2455);
and U5787 (N_5787,In_848,In_1638);
nand U5788 (N_5788,In_1933,In_2235);
nor U5789 (N_5789,In_871,In_1214);
nor U5790 (N_5790,In_2220,In_487);
and U5791 (N_5791,In_1919,In_1727);
xnor U5792 (N_5792,In_2062,In_498);
nor U5793 (N_5793,In_1509,In_134);
nand U5794 (N_5794,In_781,In_1152);
xor U5795 (N_5795,In_1051,In_1993);
or U5796 (N_5796,In_2437,In_1152);
xnor U5797 (N_5797,In_21,In_337);
nor U5798 (N_5798,In_1310,In_1630);
xor U5799 (N_5799,In_557,In_1557);
or U5800 (N_5800,In_1027,In_460);
and U5801 (N_5801,In_1177,In_2446);
or U5802 (N_5802,In_2255,In_1937);
or U5803 (N_5803,In_2217,In_2328);
or U5804 (N_5804,In_93,In_2345);
or U5805 (N_5805,In_734,In_947);
and U5806 (N_5806,In_977,In_2338);
nand U5807 (N_5807,In_998,In_1676);
or U5808 (N_5808,In_1969,In_203);
nand U5809 (N_5809,In_1512,In_2255);
nor U5810 (N_5810,In_2117,In_1032);
nand U5811 (N_5811,In_1762,In_1704);
and U5812 (N_5812,In_1322,In_657);
and U5813 (N_5813,In_921,In_909);
xor U5814 (N_5814,In_500,In_2170);
and U5815 (N_5815,In_1582,In_1115);
nand U5816 (N_5816,In_1535,In_1283);
or U5817 (N_5817,In_1221,In_1202);
nor U5818 (N_5818,In_587,In_906);
nand U5819 (N_5819,In_1792,In_163);
xnor U5820 (N_5820,In_967,In_406);
and U5821 (N_5821,In_1949,In_2315);
and U5822 (N_5822,In_639,In_1014);
and U5823 (N_5823,In_386,In_2457);
xnor U5824 (N_5824,In_1932,In_1950);
and U5825 (N_5825,In_2100,In_1606);
xnor U5826 (N_5826,In_2128,In_870);
nor U5827 (N_5827,In_1836,In_1282);
xnor U5828 (N_5828,In_103,In_1552);
xor U5829 (N_5829,In_2325,In_729);
nor U5830 (N_5830,In_756,In_2096);
and U5831 (N_5831,In_1831,In_2169);
xor U5832 (N_5832,In_2029,In_99);
or U5833 (N_5833,In_170,In_1943);
nor U5834 (N_5834,In_985,In_681);
nor U5835 (N_5835,In_842,In_2344);
and U5836 (N_5836,In_779,In_138);
nand U5837 (N_5837,In_407,In_740);
xor U5838 (N_5838,In_1517,In_40);
xor U5839 (N_5839,In_2030,In_1906);
xnor U5840 (N_5840,In_1429,In_1582);
nor U5841 (N_5841,In_823,In_932);
nor U5842 (N_5842,In_103,In_1112);
nor U5843 (N_5843,In_986,In_1831);
or U5844 (N_5844,In_951,In_79);
nand U5845 (N_5845,In_396,In_358);
and U5846 (N_5846,In_2316,In_760);
and U5847 (N_5847,In_1607,In_753);
nor U5848 (N_5848,In_2471,In_2146);
xnor U5849 (N_5849,In_1053,In_782);
and U5850 (N_5850,In_1466,In_1268);
nand U5851 (N_5851,In_1269,In_211);
xor U5852 (N_5852,In_607,In_1945);
nor U5853 (N_5853,In_375,In_2272);
and U5854 (N_5854,In_1303,In_76);
or U5855 (N_5855,In_2169,In_1553);
nand U5856 (N_5856,In_994,In_986);
nand U5857 (N_5857,In_2406,In_2328);
and U5858 (N_5858,In_2206,In_635);
or U5859 (N_5859,In_364,In_1334);
and U5860 (N_5860,In_2444,In_151);
nand U5861 (N_5861,In_116,In_1399);
nand U5862 (N_5862,In_894,In_340);
and U5863 (N_5863,In_151,In_2098);
nand U5864 (N_5864,In_358,In_1863);
and U5865 (N_5865,In_2432,In_2126);
nor U5866 (N_5866,In_571,In_1457);
nor U5867 (N_5867,In_1748,In_1342);
nor U5868 (N_5868,In_2333,In_449);
xor U5869 (N_5869,In_1042,In_496);
or U5870 (N_5870,In_2361,In_380);
xor U5871 (N_5871,In_145,In_349);
nor U5872 (N_5872,In_72,In_1248);
xor U5873 (N_5873,In_1502,In_1379);
xor U5874 (N_5874,In_1602,In_556);
nand U5875 (N_5875,In_2178,In_824);
nor U5876 (N_5876,In_1803,In_958);
or U5877 (N_5877,In_403,In_1278);
or U5878 (N_5878,In_1816,In_518);
and U5879 (N_5879,In_1496,In_1993);
and U5880 (N_5880,In_1711,In_1592);
nor U5881 (N_5881,In_1192,In_1692);
xor U5882 (N_5882,In_2253,In_914);
xnor U5883 (N_5883,In_1797,In_1450);
nor U5884 (N_5884,In_801,In_1690);
xor U5885 (N_5885,In_2103,In_1875);
and U5886 (N_5886,In_2198,In_594);
xnor U5887 (N_5887,In_2350,In_773);
xor U5888 (N_5888,In_2318,In_1490);
and U5889 (N_5889,In_1181,In_1116);
xor U5890 (N_5890,In_2347,In_1587);
or U5891 (N_5891,In_247,In_2203);
nand U5892 (N_5892,In_1924,In_1587);
or U5893 (N_5893,In_1222,In_2118);
nand U5894 (N_5894,In_933,In_1868);
nor U5895 (N_5895,In_1174,In_88);
nand U5896 (N_5896,In_1618,In_687);
and U5897 (N_5897,In_2047,In_2331);
nand U5898 (N_5898,In_297,In_193);
or U5899 (N_5899,In_827,In_486);
nor U5900 (N_5900,In_1428,In_2323);
and U5901 (N_5901,In_2275,In_1938);
or U5902 (N_5902,In_1752,In_1061);
or U5903 (N_5903,In_125,In_544);
nor U5904 (N_5904,In_1392,In_1856);
nor U5905 (N_5905,In_209,In_1170);
or U5906 (N_5906,In_955,In_1611);
xor U5907 (N_5907,In_399,In_2291);
or U5908 (N_5908,In_1928,In_1786);
xnor U5909 (N_5909,In_517,In_1880);
nor U5910 (N_5910,In_121,In_581);
or U5911 (N_5911,In_879,In_1664);
nor U5912 (N_5912,In_1244,In_33);
or U5913 (N_5913,In_2174,In_1544);
xor U5914 (N_5914,In_1372,In_885);
xor U5915 (N_5915,In_2003,In_1243);
xor U5916 (N_5916,In_1095,In_856);
or U5917 (N_5917,In_1824,In_1605);
nor U5918 (N_5918,In_89,In_1209);
xor U5919 (N_5919,In_2396,In_600);
or U5920 (N_5920,In_110,In_2036);
nor U5921 (N_5921,In_1250,In_1935);
xor U5922 (N_5922,In_862,In_797);
and U5923 (N_5923,In_1808,In_54);
or U5924 (N_5924,In_2274,In_719);
or U5925 (N_5925,In_987,In_1193);
xor U5926 (N_5926,In_500,In_240);
and U5927 (N_5927,In_1075,In_1309);
and U5928 (N_5928,In_349,In_1293);
nand U5929 (N_5929,In_1761,In_2462);
nor U5930 (N_5930,In_730,In_551);
and U5931 (N_5931,In_831,In_352);
or U5932 (N_5932,In_1235,In_2184);
nand U5933 (N_5933,In_193,In_1160);
nand U5934 (N_5934,In_2016,In_1309);
or U5935 (N_5935,In_142,In_1165);
xor U5936 (N_5936,In_130,In_2463);
xor U5937 (N_5937,In_230,In_2455);
nor U5938 (N_5938,In_1271,In_2224);
xor U5939 (N_5939,In_2332,In_1364);
and U5940 (N_5940,In_1394,In_1377);
or U5941 (N_5941,In_1242,In_2091);
or U5942 (N_5942,In_2475,In_2082);
nor U5943 (N_5943,In_1278,In_2238);
nor U5944 (N_5944,In_1958,In_2340);
or U5945 (N_5945,In_2183,In_2445);
and U5946 (N_5946,In_643,In_685);
or U5947 (N_5947,In_219,In_1450);
nor U5948 (N_5948,In_2400,In_951);
nor U5949 (N_5949,In_2254,In_243);
nor U5950 (N_5950,In_1612,In_1867);
or U5951 (N_5951,In_2032,In_1828);
nand U5952 (N_5952,In_361,In_1867);
xnor U5953 (N_5953,In_151,In_705);
or U5954 (N_5954,In_1894,In_1360);
xnor U5955 (N_5955,In_1899,In_2270);
nand U5956 (N_5956,In_372,In_280);
or U5957 (N_5957,In_1407,In_2351);
xnor U5958 (N_5958,In_1939,In_342);
and U5959 (N_5959,In_593,In_1256);
xnor U5960 (N_5960,In_1149,In_574);
nand U5961 (N_5961,In_1646,In_1202);
nand U5962 (N_5962,In_305,In_1912);
or U5963 (N_5963,In_387,In_284);
nand U5964 (N_5964,In_2196,In_2026);
nand U5965 (N_5965,In_1364,In_2180);
or U5966 (N_5966,In_1717,In_28);
xnor U5967 (N_5967,In_1749,In_202);
nor U5968 (N_5968,In_592,In_1506);
nand U5969 (N_5969,In_183,In_697);
nor U5970 (N_5970,In_2245,In_1672);
nor U5971 (N_5971,In_60,In_980);
or U5972 (N_5972,In_1784,In_119);
or U5973 (N_5973,In_908,In_1352);
xnor U5974 (N_5974,In_441,In_196);
nor U5975 (N_5975,In_1023,In_1829);
xor U5976 (N_5976,In_2346,In_1698);
nand U5977 (N_5977,In_2318,In_1234);
and U5978 (N_5978,In_2192,In_1480);
nor U5979 (N_5979,In_1252,In_110);
and U5980 (N_5980,In_1282,In_2292);
nand U5981 (N_5981,In_943,In_347);
and U5982 (N_5982,In_2450,In_935);
and U5983 (N_5983,In_921,In_263);
and U5984 (N_5984,In_1661,In_566);
nand U5985 (N_5985,In_1696,In_95);
nor U5986 (N_5986,In_2460,In_42);
nand U5987 (N_5987,In_2476,In_656);
and U5988 (N_5988,In_916,In_897);
nor U5989 (N_5989,In_73,In_177);
xnor U5990 (N_5990,In_2090,In_1942);
or U5991 (N_5991,In_1333,In_1740);
nor U5992 (N_5992,In_1869,In_1343);
and U5993 (N_5993,In_1022,In_1423);
nor U5994 (N_5994,In_1120,In_368);
and U5995 (N_5995,In_228,In_1937);
xor U5996 (N_5996,In_1385,In_1533);
xnor U5997 (N_5997,In_1360,In_314);
or U5998 (N_5998,In_2189,In_1874);
nor U5999 (N_5999,In_79,In_2241);
nand U6000 (N_6000,In_93,In_613);
or U6001 (N_6001,In_1397,In_1799);
nor U6002 (N_6002,In_1456,In_2277);
nand U6003 (N_6003,In_154,In_754);
and U6004 (N_6004,In_1215,In_1508);
and U6005 (N_6005,In_130,In_1167);
and U6006 (N_6006,In_856,In_897);
xnor U6007 (N_6007,In_2416,In_1970);
xnor U6008 (N_6008,In_1697,In_2240);
and U6009 (N_6009,In_647,In_2251);
and U6010 (N_6010,In_1304,In_1961);
nor U6011 (N_6011,In_1459,In_2287);
or U6012 (N_6012,In_2238,In_1202);
and U6013 (N_6013,In_1049,In_688);
nand U6014 (N_6014,In_2056,In_596);
and U6015 (N_6015,In_1837,In_1346);
xnor U6016 (N_6016,In_2282,In_2054);
and U6017 (N_6017,In_213,In_916);
xnor U6018 (N_6018,In_2085,In_1571);
and U6019 (N_6019,In_2193,In_850);
and U6020 (N_6020,In_301,In_543);
xor U6021 (N_6021,In_1808,In_1743);
and U6022 (N_6022,In_1289,In_403);
nand U6023 (N_6023,In_1674,In_1145);
nor U6024 (N_6024,In_2058,In_1290);
and U6025 (N_6025,In_2454,In_1635);
nor U6026 (N_6026,In_2347,In_76);
nor U6027 (N_6027,In_12,In_1538);
xnor U6028 (N_6028,In_1327,In_2389);
and U6029 (N_6029,In_1008,In_1779);
xnor U6030 (N_6030,In_1614,In_1542);
nor U6031 (N_6031,In_444,In_233);
nand U6032 (N_6032,In_1668,In_38);
nand U6033 (N_6033,In_705,In_539);
xnor U6034 (N_6034,In_2483,In_513);
nand U6035 (N_6035,In_2031,In_813);
nor U6036 (N_6036,In_1517,In_143);
and U6037 (N_6037,In_1281,In_52);
nor U6038 (N_6038,In_1952,In_1601);
xor U6039 (N_6039,In_2119,In_168);
and U6040 (N_6040,In_2498,In_2310);
and U6041 (N_6041,In_150,In_686);
and U6042 (N_6042,In_920,In_116);
nor U6043 (N_6043,In_2455,In_1077);
xor U6044 (N_6044,In_1830,In_2358);
and U6045 (N_6045,In_724,In_115);
and U6046 (N_6046,In_553,In_922);
nor U6047 (N_6047,In_2160,In_140);
or U6048 (N_6048,In_1429,In_1444);
xor U6049 (N_6049,In_1273,In_115);
or U6050 (N_6050,In_6,In_251);
and U6051 (N_6051,In_2394,In_1026);
nand U6052 (N_6052,In_274,In_2050);
and U6053 (N_6053,In_1290,In_721);
or U6054 (N_6054,In_2361,In_554);
xor U6055 (N_6055,In_754,In_330);
nor U6056 (N_6056,In_1514,In_666);
and U6057 (N_6057,In_2058,In_746);
and U6058 (N_6058,In_902,In_71);
and U6059 (N_6059,In_2332,In_2330);
or U6060 (N_6060,In_2454,In_724);
nand U6061 (N_6061,In_807,In_363);
nor U6062 (N_6062,In_204,In_1421);
and U6063 (N_6063,In_238,In_2249);
xor U6064 (N_6064,In_411,In_320);
xnor U6065 (N_6065,In_1673,In_558);
xor U6066 (N_6066,In_1256,In_1846);
or U6067 (N_6067,In_2316,In_1392);
and U6068 (N_6068,In_84,In_655);
nor U6069 (N_6069,In_282,In_1874);
and U6070 (N_6070,In_515,In_2404);
xor U6071 (N_6071,In_390,In_1447);
xnor U6072 (N_6072,In_2092,In_1171);
nor U6073 (N_6073,In_341,In_859);
and U6074 (N_6074,In_562,In_1130);
xnor U6075 (N_6075,In_248,In_1282);
or U6076 (N_6076,In_898,In_1884);
and U6077 (N_6077,In_274,In_1197);
nand U6078 (N_6078,In_2204,In_952);
or U6079 (N_6079,In_67,In_57);
nor U6080 (N_6080,In_1763,In_1963);
xor U6081 (N_6081,In_846,In_1945);
xnor U6082 (N_6082,In_1280,In_334);
or U6083 (N_6083,In_2118,In_396);
or U6084 (N_6084,In_2264,In_2093);
and U6085 (N_6085,In_2381,In_1381);
or U6086 (N_6086,In_1776,In_2481);
xor U6087 (N_6087,In_2113,In_2379);
nor U6088 (N_6088,In_1541,In_186);
nor U6089 (N_6089,In_1957,In_1700);
or U6090 (N_6090,In_779,In_970);
nor U6091 (N_6091,In_1859,In_897);
nand U6092 (N_6092,In_926,In_1381);
nand U6093 (N_6093,In_726,In_1917);
nor U6094 (N_6094,In_1781,In_1554);
nand U6095 (N_6095,In_2012,In_1594);
nor U6096 (N_6096,In_2190,In_276);
or U6097 (N_6097,In_823,In_1750);
nor U6098 (N_6098,In_760,In_1859);
nand U6099 (N_6099,In_604,In_629);
nor U6100 (N_6100,In_1840,In_1166);
nor U6101 (N_6101,In_781,In_391);
nand U6102 (N_6102,In_2245,In_1674);
xnor U6103 (N_6103,In_1522,In_2337);
or U6104 (N_6104,In_2380,In_845);
or U6105 (N_6105,In_298,In_866);
and U6106 (N_6106,In_560,In_902);
and U6107 (N_6107,In_483,In_803);
and U6108 (N_6108,In_1952,In_492);
nand U6109 (N_6109,In_1971,In_514);
xor U6110 (N_6110,In_5,In_956);
or U6111 (N_6111,In_564,In_776);
and U6112 (N_6112,In_1025,In_1542);
nor U6113 (N_6113,In_261,In_1590);
and U6114 (N_6114,In_1362,In_325);
nand U6115 (N_6115,In_437,In_913);
or U6116 (N_6116,In_980,In_777);
xor U6117 (N_6117,In_1191,In_424);
nand U6118 (N_6118,In_833,In_666);
and U6119 (N_6119,In_881,In_371);
or U6120 (N_6120,In_1884,In_948);
xnor U6121 (N_6121,In_158,In_1661);
and U6122 (N_6122,In_1878,In_1953);
or U6123 (N_6123,In_1285,In_1313);
xor U6124 (N_6124,In_2225,In_2367);
nor U6125 (N_6125,In_1905,In_358);
nor U6126 (N_6126,In_1051,In_1035);
nand U6127 (N_6127,In_706,In_795);
nand U6128 (N_6128,In_1020,In_1302);
xor U6129 (N_6129,In_1483,In_2187);
and U6130 (N_6130,In_2299,In_136);
nand U6131 (N_6131,In_1854,In_1386);
and U6132 (N_6132,In_733,In_1487);
or U6133 (N_6133,In_2074,In_969);
and U6134 (N_6134,In_519,In_2220);
xor U6135 (N_6135,In_2361,In_730);
xnor U6136 (N_6136,In_1335,In_864);
and U6137 (N_6137,In_1611,In_1516);
xnor U6138 (N_6138,In_191,In_129);
xnor U6139 (N_6139,In_113,In_849);
or U6140 (N_6140,In_818,In_1571);
nor U6141 (N_6141,In_222,In_1683);
xnor U6142 (N_6142,In_2137,In_1023);
or U6143 (N_6143,In_1118,In_1890);
or U6144 (N_6144,In_2086,In_1068);
or U6145 (N_6145,In_2106,In_18);
xor U6146 (N_6146,In_1118,In_1160);
or U6147 (N_6147,In_1186,In_894);
nand U6148 (N_6148,In_891,In_1399);
and U6149 (N_6149,In_581,In_1469);
or U6150 (N_6150,In_1558,In_1933);
nor U6151 (N_6151,In_1651,In_977);
or U6152 (N_6152,In_2209,In_666);
nor U6153 (N_6153,In_1479,In_1612);
nor U6154 (N_6154,In_638,In_1006);
nor U6155 (N_6155,In_1618,In_938);
nor U6156 (N_6156,In_340,In_65);
nor U6157 (N_6157,In_1694,In_1354);
xor U6158 (N_6158,In_654,In_1240);
nor U6159 (N_6159,In_1732,In_1553);
nand U6160 (N_6160,In_948,In_1277);
and U6161 (N_6161,In_2184,In_1290);
or U6162 (N_6162,In_1431,In_2115);
nor U6163 (N_6163,In_2427,In_1701);
xnor U6164 (N_6164,In_1549,In_502);
nand U6165 (N_6165,In_1798,In_1496);
nor U6166 (N_6166,In_425,In_1836);
or U6167 (N_6167,In_1658,In_2201);
and U6168 (N_6168,In_1668,In_353);
xnor U6169 (N_6169,In_2420,In_342);
and U6170 (N_6170,In_416,In_575);
nor U6171 (N_6171,In_2026,In_1263);
or U6172 (N_6172,In_1514,In_1351);
and U6173 (N_6173,In_653,In_1595);
and U6174 (N_6174,In_775,In_1339);
and U6175 (N_6175,In_782,In_750);
and U6176 (N_6176,In_283,In_1037);
or U6177 (N_6177,In_1202,In_1190);
and U6178 (N_6178,In_1504,In_111);
or U6179 (N_6179,In_268,In_1775);
and U6180 (N_6180,In_2007,In_1208);
nand U6181 (N_6181,In_1886,In_1649);
and U6182 (N_6182,In_1000,In_2265);
nand U6183 (N_6183,In_1099,In_919);
nand U6184 (N_6184,In_2277,In_1396);
or U6185 (N_6185,In_1920,In_767);
nand U6186 (N_6186,In_1555,In_2180);
nand U6187 (N_6187,In_1602,In_2332);
and U6188 (N_6188,In_2243,In_2417);
or U6189 (N_6189,In_944,In_653);
nand U6190 (N_6190,In_1058,In_665);
xnor U6191 (N_6191,In_664,In_2499);
xnor U6192 (N_6192,In_348,In_1507);
and U6193 (N_6193,In_1594,In_732);
nand U6194 (N_6194,In_625,In_599);
xnor U6195 (N_6195,In_358,In_887);
and U6196 (N_6196,In_1966,In_881);
nor U6197 (N_6197,In_445,In_763);
nor U6198 (N_6198,In_1266,In_1265);
nand U6199 (N_6199,In_1818,In_916);
and U6200 (N_6200,In_1373,In_112);
nand U6201 (N_6201,In_2382,In_1348);
and U6202 (N_6202,In_1623,In_1030);
nor U6203 (N_6203,In_1480,In_1640);
nand U6204 (N_6204,In_2361,In_1461);
nand U6205 (N_6205,In_930,In_1546);
and U6206 (N_6206,In_2361,In_1146);
xnor U6207 (N_6207,In_720,In_550);
nor U6208 (N_6208,In_478,In_403);
nand U6209 (N_6209,In_610,In_522);
or U6210 (N_6210,In_2179,In_78);
nand U6211 (N_6211,In_278,In_1132);
nand U6212 (N_6212,In_1273,In_1008);
nand U6213 (N_6213,In_1854,In_1001);
xnor U6214 (N_6214,In_1702,In_1508);
nor U6215 (N_6215,In_1946,In_2444);
xnor U6216 (N_6216,In_980,In_2285);
and U6217 (N_6217,In_2286,In_1167);
xor U6218 (N_6218,In_1757,In_5);
nand U6219 (N_6219,In_2408,In_252);
and U6220 (N_6220,In_1776,In_601);
xor U6221 (N_6221,In_1638,In_322);
xor U6222 (N_6222,In_1076,In_423);
nand U6223 (N_6223,In_1948,In_1940);
or U6224 (N_6224,In_735,In_747);
xor U6225 (N_6225,In_192,In_1033);
xor U6226 (N_6226,In_1969,In_2254);
nor U6227 (N_6227,In_727,In_1694);
xor U6228 (N_6228,In_55,In_1402);
and U6229 (N_6229,In_1851,In_1462);
nand U6230 (N_6230,In_220,In_493);
nor U6231 (N_6231,In_1408,In_2115);
or U6232 (N_6232,In_1098,In_2203);
nand U6233 (N_6233,In_1831,In_1845);
nor U6234 (N_6234,In_1086,In_1263);
and U6235 (N_6235,In_75,In_818);
nor U6236 (N_6236,In_54,In_933);
or U6237 (N_6237,In_1173,In_7);
nor U6238 (N_6238,In_1013,In_1960);
xor U6239 (N_6239,In_1952,In_5);
xnor U6240 (N_6240,In_478,In_60);
nor U6241 (N_6241,In_591,In_71);
xor U6242 (N_6242,In_891,In_1284);
nand U6243 (N_6243,In_133,In_971);
nand U6244 (N_6244,In_1490,In_1869);
and U6245 (N_6245,In_22,In_1866);
nor U6246 (N_6246,In_2490,In_1172);
xor U6247 (N_6247,In_2254,In_1223);
nand U6248 (N_6248,In_1044,In_217);
or U6249 (N_6249,In_618,In_1772);
xnor U6250 (N_6250,N_5682,N_2080);
or U6251 (N_6251,N_4629,N_5382);
and U6252 (N_6252,N_3111,N_2569);
nor U6253 (N_6253,N_3781,N_227);
xnor U6254 (N_6254,N_5509,N_4018);
xnor U6255 (N_6255,N_5997,N_1828);
nor U6256 (N_6256,N_5319,N_5920);
or U6257 (N_6257,N_3123,N_1253);
xor U6258 (N_6258,N_5246,N_4370);
xor U6259 (N_6259,N_5392,N_2617);
or U6260 (N_6260,N_4570,N_4012);
and U6261 (N_6261,N_431,N_504);
or U6262 (N_6262,N_6201,N_3203);
nand U6263 (N_6263,N_4666,N_3462);
nand U6264 (N_6264,N_363,N_5328);
nor U6265 (N_6265,N_4619,N_3972);
nand U6266 (N_6266,N_144,N_966);
and U6267 (N_6267,N_1975,N_6081);
xor U6268 (N_6268,N_5119,N_4016);
nor U6269 (N_6269,N_2973,N_4186);
nand U6270 (N_6270,N_5092,N_1643);
nor U6271 (N_6271,N_1297,N_2361);
and U6272 (N_6272,N_890,N_5015);
or U6273 (N_6273,N_2280,N_2657);
or U6274 (N_6274,N_5551,N_1562);
or U6275 (N_6275,N_5209,N_52);
or U6276 (N_6276,N_4234,N_168);
nor U6277 (N_6277,N_1158,N_2220);
nand U6278 (N_6278,N_2188,N_3929);
nor U6279 (N_6279,N_4882,N_2134);
nand U6280 (N_6280,N_661,N_725);
nor U6281 (N_6281,N_4854,N_5419);
xnor U6282 (N_6282,N_3580,N_627);
nor U6283 (N_6283,N_2349,N_2518);
nor U6284 (N_6284,N_2020,N_1872);
nand U6285 (N_6285,N_1395,N_2417);
and U6286 (N_6286,N_5527,N_2311);
xnor U6287 (N_6287,N_2607,N_189);
and U6288 (N_6288,N_1084,N_3371);
nor U6289 (N_6289,N_5884,N_4161);
and U6290 (N_6290,N_2189,N_503);
nor U6291 (N_6291,N_2771,N_270);
or U6292 (N_6292,N_2181,N_479);
and U6293 (N_6293,N_1368,N_1560);
or U6294 (N_6294,N_3512,N_4167);
nand U6295 (N_6295,N_5008,N_3387);
and U6296 (N_6296,N_4057,N_4308);
and U6297 (N_6297,N_6212,N_493);
xnor U6298 (N_6298,N_6046,N_2309);
nor U6299 (N_6299,N_170,N_1342);
nand U6300 (N_6300,N_6061,N_461);
nand U6301 (N_6301,N_3966,N_6202);
nor U6302 (N_6302,N_1539,N_38);
xnor U6303 (N_6303,N_5240,N_3602);
nand U6304 (N_6304,N_5722,N_1908);
and U6305 (N_6305,N_4336,N_6032);
or U6306 (N_6306,N_2158,N_1119);
nand U6307 (N_6307,N_5348,N_4302);
xnor U6308 (N_6308,N_1548,N_4246);
and U6309 (N_6309,N_5309,N_5981);
and U6310 (N_6310,N_3098,N_762);
xnor U6311 (N_6311,N_4711,N_1061);
nor U6312 (N_6312,N_2039,N_4038);
or U6313 (N_6313,N_1407,N_951);
or U6314 (N_6314,N_1673,N_822);
nor U6315 (N_6315,N_585,N_5408);
nand U6316 (N_6316,N_2946,N_2094);
or U6317 (N_6317,N_5790,N_5116);
xor U6318 (N_6318,N_4696,N_3311);
nor U6319 (N_6319,N_324,N_2301);
nor U6320 (N_6320,N_3663,N_1277);
xor U6321 (N_6321,N_837,N_4853);
xnor U6322 (N_6322,N_5118,N_5534);
nor U6323 (N_6323,N_5315,N_3686);
and U6324 (N_6324,N_1893,N_2979);
and U6325 (N_6325,N_1477,N_5476);
nor U6326 (N_6326,N_5168,N_1517);
nand U6327 (N_6327,N_2252,N_5034);
nor U6328 (N_6328,N_3285,N_2376);
and U6329 (N_6329,N_4596,N_5656);
and U6330 (N_6330,N_570,N_2886);
or U6331 (N_6331,N_1419,N_3600);
xor U6332 (N_6332,N_6111,N_4777);
nor U6333 (N_6333,N_1612,N_380);
xor U6334 (N_6334,N_4996,N_4738);
nand U6335 (N_6335,N_2776,N_1162);
nor U6336 (N_6336,N_5342,N_3169);
nand U6337 (N_6337,N_1139,N_6205);
xor U6338 (N_6338,N_1155,N_1646);
nand U6339 (N_6339,N_5074,N_5125);
or U6340 (N_6340,N_2131,N_5291);
or U6341 (N_6341,N_3012,N_2701);
or U6342 (N_6342,N_1465,N_5373);
or U6343 (N_6343,N_2648,N_5128);
nand U6344 (N_6344,N_2185,N_1718);
xnor U6345 (N_6345,N_4683,N_197);
and U6346 (N_6346,N_2924,N_5735);
xnor U6347 (N_6347,N_2370,N_4367);
xnor U6348 (N_6348,N_542,N_2618);
and U6349 (N_6349,N_2026,N_1727);
nor U6350 (N_6350,N_4764,N_375);
xor U6351 (N_6351,N_1732,N_3644);
nand U6352 (N_6352,N_5212,N_4475);
or U6353 (N_6353,N_2705,N_1046);
and U6354 (N_6354,N_3397,N_3131);
nand U6355 (N_6355,N_4869,N_4735);
or U6356 (N_6356,N_124,N_3734);
nor U6357 (N_6357,N_2741,N_6213);
or U6358 (N_6358,N_2918,N_3087);
nand U6359 (N_6359,N_5570,N_2982);
or U6360 (N_6360,N_3040,N_738);
nor U6361 (N_6361,N_509,N_4624);
nand U6362 (N_6362,N_3857,N_1603);
xnor U6363 (N_6363,N_492,N_3838);
xor U6364 (N_6364,N_5395,N_3172);
nand U6365 (N_6365,N_1042,N_2631);
or U6366 (N_6366,N_4219,N_4140);
xnor U6367 (N_6367,N_348,N_5208);
or U6368 (N_6368,N_1399,N_5117);
and U6369 (N_6369,N_1627,N_5266);
or U6370 (N_6370,N_6054,N_1945);
nand U6371 (N_6371,N_4344,N_2251);
and U6372 (N_6372,N_5102,N_3078);
or U6373 (N_6373,N_4914,N_2344);
nor U6374 (N_6374,N_1642,N_2229);
nand U6375 (N_6375,N_895,N_1495);
nor U6376 (N_6376,N_1705,N_2327);
nand U6377 (N_6377,N_2294,N_5635);
nor U6378 (N_6378,N_3220,N_4254);
or U6379 (N_6379,N_2849,N_6165);
nand U6380 (N_6380,N_5367,N_1271);
or U6381 (N_6381,N_1207,N_3354);
or U6382 (N_6382,N_4223,N_2580);
nand U6383 (N_6383,N_21,N_1039);
and U6384 (N_6384,N_89,N_4413);
xor U6385 (N_6385,N_3628,N_5148);
or U6386 (N_6386,N_1756,N_1807);
and U6387 (N_6387,N_524,N_5202);
nor U6388 (N_6388,N_460,N_5082);
xor U6389 (N_6389,N_5751,N_5178);
xor U6390 (N_6390,N_1009,N_5417);
nand U6391 (N_6391,N_3180,N_3676);
xnor U6392 (N_6392,N_2422,N_548);
and U6393 (N_6393,N_5917,N_2642);
nor U6394 (N_6394,N_3035,N_845);
and U6395 (N_6395,N_5312,N_3719);
or U6396 (N_6396,N_3369,N_1510);
or U6397 (N_6397,N_3213,N_3992);
nand U6398 (N_6398,N_710,N_5127);
and U6399 (N_6399,N_217,N_3708);
nand U6400 (N_6400,N_2471,N_5085);
xnor U6401 (N_6401,N_2822,N_861);
xnor U6402 (N_6402,N_3652,N_5457);
and U6403 (N_6403,N_1634,N_833);
xor U6404 (N_6404,N_2775,N_1473);
or U6405 (N_6405,N_5965,N_150);
nor U6406 (N_6406,N_4540,N_5329);
nand U6407 (N_6407,N_6185,N_6123);
xnor U6408 (N_6408,N_4287,N_3445);
nand U6409 (N_6409,N_4887,N_5716);
nor U6410 (N_6410,N_112,N_5556);
nand U6411 (N_6411,N_1026,N_490);
nand U6412 (N_6412,N_2572,N_2183);
and U6413 (N_6413,N_582,N_15);
nand U6414 (N_6414,N_1187,N_2655);
nand U6415 (N_6415,N_3244,N_4159);
or U6416 (N_6416,N_667,N_2792);
nand U6417 (N_6417,N_429,N_3709);
xnor U6418 (N_6418,N_2842,N_462);
or U6419 (N_6419,N_2854,N_3878);
and U6420 (N_6420,N_1757,N_2747);
nor U6421 (N_6421,N_893,N_422);
xor U6422 (N_6422,N_1946,N_5577);
or U6423 (N_6423,N_6156,N_1497);
nor U6424 (N_6424,N_278,N_3245);
nand U6425 (N_6425,N_1645,N_476);
nand U6426 (N_6426,N_4637,N_5520);
xnor U6427 (N_6427,N_3845,N_612);
xnor U6428 (N_6428,N_5169,N_3233);
xor U6429 (N_6429,N_4640,N_5779);
nor U6430 (N_6430,N_2351,N_79);
nor U6431 (N_6431,N_5054,N_4249);
or U6432 (N_6432,N_3687,N_4689);
xnor U6433 (N_6433,N_5278,N_4794);
xnor U6434 (N_6434,N_2009,N_5606);
xnor U6435 (N_6435,N_987,N_4305);
or U6436 (N_6436,N_3474,N_3269);
xor U6437 (N_6437,N_6215,N_1607);
nand U6438 (N_6438,N_4950,N_1886);
or U6439 (N_6439,N_2509,N_5404);
or U6440 (N_6440,N_37,N_4512);
xnor U6441 (N_6441,N_4210,N_3112);
nor U6442 (N_6442,N_415,N_247);
nand U6443 (N_6443,N_322,N_434);
nand U6444 (N_6444,N_1408,N_2820);
xnor U6445 (N_6445,N_2388,N_2332);
nor U6446 (N_6446,N_779,N_5177);
xnor U6447 (N_6447,N_2780,N_834);
nand U6448 (N_6448,N_3711,N_1597);
nand U6449 (N_6449,N_3818,N_5040);
nor U6450 (N_6450,N_697,N_2060);
and U6451 (N_6451,N_5619,N_1781);
xnor U6452 (N_6452,N_4388,N_2041);
nand U6453 (N_6453,N_2708,N_6070);
or U6454 (N_6454,N_942,N_654);
xor U6455 (N_6455,N_723,N_4100);
and U6456 (N_6456,N_2016,N_5925);
nand U6457 (N_6457,N_899,N_6225);
nor U6458 (N_6458,N_4417,N_2787);
and U6459 (N_6459,N_2192,N_5327);
nand U6460 (N_6460,N_4991,N_4829);
xor U6461 (N_6461,N_67,N_2983);
nor U6462 (N_6462,N_940,N_647);
or U6463 (N_6463,N_865,N_2940);
or U6464 (N_6464,N_440,N_3858);
nand U6465 (N_6465,N_5306,N_4929);
and U6466 (N_6466,N_4430,N_3359);
xnor U6467 (N_6467,N_742,N_2857);
or U6468 (N_6468,N_949,N_5699);
nor U6469 (N_6469,N_849,N_4313);
or U6470 (N_6470,N_2481,N_4438);
nor U6471 (N_6471,N_2706,N_3433);
nand U6472 (N_6472,N_2646,N_4114);
and U6473 (N_6473,N_1697,N_3258);
and U6474 (N_6474,N_3331,N_1197);
and U6475 (N_6475,N_5603,N_5032);
nor U6476 (N_6476,N_3034,N_3473);
xor U6477 (N_6477,N_1972,N_229);
xor U6478 (N_6478,N_3978,N_2152);
nor U6479 (N_6479,N_4421,N_4058);
xnor U6480 (N_6480,N_3262,N_3437);
and U6481 (N_6481,N_4300,N_1348);
xnor U6482 (N_6482,N_2906,N_1030);
or U6483 (N_6483,N_2413,N_6011);
nor U6484 (N_6484,N_3215,N_2879);
nor U6485 (N_6485,N_5614,N_5004);
nor U6486 (N_6486,N_4048,N_3316);
nor U6487 (N_6487,N_1710,N_4208);
nand U6488 (N_6488,N_2625,N_382);
and U6489 (N_6489,N_2904,N_4995);
nand U6490 (N_6490,N_3116,N_922);
nor U6491 (N_6491,N_523,N_5597);
xnor U6492 (N_6492,N_5160,N_1296);
or U6493 (N_6493,N_4986,N_471);
and U6494 (N_6494,N_5241,N_4897);
or U6495 (N_6495,N_2695,N_4549);
xor U6496 (N_6496,N_1104,N_4509);
and U6497 (N_6497,N_5953,N_3242);
nor U6498 (N_6498,N_2210,N_3015);
or U6499 (N_6499,N_4552,N_86);
nor U6500 (N_6500,N_675,N_3277);
nand U6501 (N_6501,N_4221,N_4976);
xor U6502 (N_6502,N_1987,N_5604);
xnor U6503 (N_6503,N_4977,N_555);
and U6504 (N_6504,N_464,N_5391);
and U6505 (N_6505,N_3063,N_1555);
nor U6506 (N_6506,N_409,N_1778);
nand U6507 (N_6507,N_2608,N_1879);
and U6508 (N_6508,N_2440,N_6040);
nand U6509 (N_6509,N_4027,N_5299);
or U6510 (N_6510,N_5446,N_3052);
and U6511 (N_6511,N_3140,N_5296);
and U6512 (N_6512,N_452,N_73);
and U6513 (N_6513,N_412,N_1907);
nand U6514 (N_6514,N_298,N_2851);
xor U6515 (N_6515,N_2750,N_2584);
nor U6516 (N_6516,N_4635,N_695);
and U6517 (N_6517,N_2389,N_317);
xnor U6518 (N_6518,N_130,N_3450);
nand U6519 (N_6519,N_5146,N_4880);
xor U6520 (N_6520,N_3486,N_4303);
or U6521 (N_6521,N_637,N_3617);
or U6522 (N_6522,N_5558,N_271);
or U6523 (N_6523,N_5625,N_2847);
or U6524 (N_6524,N_4754,N_3256);
and U6525 (N_6525,N_5647,N_6162);
and U6526 (N_6526,N_1801,N_3234);
and U6527 (N_6527,N_4983,N_5484);
nor U6528 (N_6528,N_3248,N_2406);
or U6529 (N_6529,N_780,N_5752);
nor U6530 (N_6530,N_3780,N_4056);
or U6531 (N_6531,N_5176,N_5811);
or U6532 (N_6532,N_2520,N_2670);
xnor U6533 (N_6533,N_5711,N_1052);
or U6534 (N_6534,N_3693,N_2279);
nor U6535 (N_6535,N_2169,N_3436);
nand U6536 (N_6536,N_181,N_3839);
and U6537 (N_6537,N_4973,N_5494);
xnor U6538 (N_6538,N_4989,N_5239);
or U6539 (N_6539,N_1926,N_1684);
xnor U6540 (N_6540,N_4377,N_2742);
nand U6541 (N_6541,N_4252,N_5448);
nor U6542 (N_6542,N_4604,N_4828);
xor U6543 (N_6543,N_1346,N_4442);
and U6544 (N_6544,N_4454,N_3683);
nand U6545 (N_6545,N_2155,N_6089);
or U6546 (N_6546,N_2304,N_512);
xor U6547 (N_6547,N_5502,N_3848);
and U6548 (N_6548,N_2385,N_1733);
or U6549 (N_6549,N_2687,N_1775);
nand U6550 (N_6550,N_283,N_5863);
and U6551 (N_6551,N_4803,N_5989);
and U6552 (N_6552,N_6073,N_5563);
or U6553 (N_6553,N_6195,N_4326);
or U6554 (N_6554,N_225,N_5836);
and U6555 (N_6555,N_4107,N_3353);
nand U6556 (N_6556,N_239,N_3575);
nand U6557 (N_6557,N_1923,N_765);
or U6558 (N_6558,N_4631,N_909);
nor U6559 (N_6559,N_1243,N_4726);
or U6560 (N_6560,N_2023,N_1029);
nand U6561 (N_6561,N_1004,N_2707);
nand U6562 (N_6562,N_2876,N_2285);
and U6563 (N_6563,N_1239,N_5380);
xnor U6564 (N_6564,N_3342,N_2613);
or U6565 (N_6565,N_280,N_5586);
and U6566 (N_6566,N_5005,N_592);
nand U6567 (N_6567,N_359,N_4724);
xor U6568 (N_6568,N_3951,N_4023);
xor U6569 (N_6569,N_4993,N_884);
and U6570 (N_6570,N_256,N_5261);
and U6571 (N_6571,N_1769,N_8);
and U6572 (N_6572,N_4518,N_3096);
xor U6573 (N_6573,N_1869,N_3967);
or U6574 (N_6574,N_5010,N_4704);
and U6575 (N_6575,N_3301,N_3044);
or U6576 (N_6576,N_2645,N_5056);
nand U6577 (N_6577,N_2084,N_4063);
xnor U6578 (N_6578,N_2844,N_6000);
xnor U6579 (N_6579,N_2383,N_3292);
or U6580 (N_6580,N_907,N_5636);
nor U6581 (N_6581,N_6221,N_3753);
xnor U6582 (N_6582,N_4690,N_1723);
nand U6583 (N_6583,N_5557,N_3415);
and U6584 (N_6584,N_5517,N_6025);
nand U6585 (N_6585,N_5445,N_5064);
nand U6586 (N_6586,N_6247,N_5564);
or U6587 (N_6587,N_2187,N_3906);
xnor U6588 (N_6588,N_2689,N_1859);
nand U6589 (N_6589,N_3950,N_5634);
and U6590 (N_6590,N_5999,N_4646);
nor U6591 (N_6591,N_4730,N_3612);
xor U6592 (N_6592,N_5284,N_2452);
nand U6593 (N_6593,N_5753,N_5662);
nor U6594 (N_6594,N_2395,N_2337);
or U6595 (N_6595,N_757,N_1527);
and U6596 (N_6596,N_474,N_2235);
nor U6597 (N_6597,N_3811,N_831);
and U6598 (N_6598,N_2265,N_897);
nand U6599 (N_6599,N_2615,N_1865);
xnor U6600 (N_6600,N_991,N_5621);
or U6601 (N_6601,N_6034,N_3005);
nor U6602 (N_6602,N_3304,N_6050);
nor U6603 (N_6603,N_2396,N_5120);
xnor U6604 (N_6604,N_4216,N_2791);
and U6605 (N_6605,N_952,N_5946);
nand U6606 (N_6606,N_3526,N_5803);
xnor U6607 (N_6607,N_5288,N_4801);
and U6608 (N_6608,N_1471,N_3358);
and U6609 (N_6609,N_1280,N_2401);
or U6610 (N_6610,N_1803,N_6134);
or U6611 (N_6611,N_515,N_6079);
nor U6612 (N_6612,N_4536,N_2516);
nand U6613 (N_6613,N_3247,N_141);
or U6614 (N_6614,N_2270,N_1345);
nand U6615 (N_6615,N_5043,N_5985);
or U6616 (N_6616,N_3980,N_6088);
and U6617 (N_6617,N_291,N_994);
nor U6618 (N_6618,N_5822,N_4407);
and U6619 (N_6619,N_2425,N_3902);
xor U6620 (N_6620,N_5472,N_968);
nor U6621 (N_6621,N_402,N_2863);
nand U6622 (N_6622,N_5479,N_3389);
or U6623 (N_6623,N_1501,N_5456);
nor U6624 (N_6624,N_473,N_5921);
and U6625 (N_6625,N_3901,N_3808);
xnor U6626 (N_6626,N_4296,N_163);
or U6627 (N_6627,N_336,N_2457);
xnor U6628 (N_6628,N_339,N_1429);
or U6629 (N_6629,N_3283,N_4931);
xor U6630 (N_6630,N_569,N_5990);
or U6631 (N_6631,N_3625,N_3658);
and U6632 (N_6632,N_3551,N_4386);
xnor U6633 (N_6633,N_3998,N_1719);
or U6634 (N_6634,N_1000,N_2164);
or U6635 (N_6635,N_126,N_4104);
nand U6636 (N_6636,N_1467,N_5891);
xnor U6637 (N_6637,N_5966,N_26);
nor U6638 (N_6638,N_5272,N_3372);
and U6639 (N_6639,N_5455,N_4797);
or U6640 (N_6640,N_2275,N_3797);
nor U6641 (N_6641,N_3201,N_1750);
nor U6642 (N_6642,N_1785,N_1092);
xor U6643 (N_6643,N_6096,N_3804);
or U6644 (N_6644,N_634,N_2394);
xor U6645 (N_6645,N_4395,N_5063);
nand U6646 (N_6646,N_3150,N_3241);
or U6647 (N_6647,N_4510,N_1797);
nand U6648 (N_6648,N_3491,N_1241);
or U6649 (N_6649,N_1482,N_3975);
or U6650 (N_6650,N_361,N_728);
or U6651 (N_6651,N_5856,N_1564);
nand U6652 (N_6652,N_4678,N_2365);
and U6653 (N_6653,N_2911,N_977);
nor U6654 (N_6654,N_5066,N_5366);
nand U6655 (N_6655,N_4691,N_5349);
nor U6656 (N_6656,N_1659,N_4196);
nand U6657 (N_6657,N_1861,N_4707);
xor U6658 (N_6658,N_1649,N_852);
xor U6659 (N_6659,N_2159,N_4831);
xnor U6660 (N_6660,N_5781,N_4187);
and U6661 (N_6661,N_2773,N_3318);
nand U6662 (N_6662,N_88,N_2709);
nor U6663 (N_6663,N_4815,N_3019);
xor U6664 (N_6664,N_2543,N_1380);
or U6665 (N_6665,N_2078,N_486);
nor U6666 (N_6666,N_1773,N_2952);
nand U6667 (N_6667,N_4598,N_2935);
or U6668 (N_6668,N_5858,N_1126);
nor U6669 (N_6669,N_6168,N_1500);
nor U6670 (N_6670,N_3882,N_1322);
or U6671 (N_6671,N_2660,N_4930);
and U6672 (N_6672,N_3046,N_3497);
nand U6673 (N_6673,N_5029,N_4125);
xor U6674 (N_6674,N_1057,N_1711);
xor U6675 (N_6675,N_3458,N_581);
or U6676 (N_6676,N_4019,N_1456);
or U6677 (N_6677,N_4889,N_2524);
and U6678 (N_6678,N_936,N_5215);
nor U6679 (N_6679,N_265,N_2355);
or U6680 (N_6680,N_1842,N_5036);
and U6681 (N_6681,N_636,N_3671);
xnor U6682 (N_6682,N_5251,N_3468);
and U6683 (N_6683,N_2928,N_5474);
or U6684 (N_6684,N_820,N_5050);
and U6685 (N_6685,N_5573,N_3995);
or U6686 (N_6686,N_1034,N_4410);
and U6687 (N_6687,N_1024,N_6214);
and U6688 (N_6688,N_1466,N_793);
nand U6689 (N_6689,N_4581,N_3231);
or U6690 (N_6690,N_1240,N_3051);
nand U6691 (N_6691,N_4886,N_4111);
nand U6692 (N_6692,N_1752,N_3057);
or U6693 (N_6693,N_2932,N_5844);
and U6694 (N_6694,N_1311,N_2323);
and U6695 (N_6695,N_6,N_3273);
and U6696 (N_6696,N_2745,N_5095);
and U6697 (N_6697,N_514,N_1613);
nor U6698 (N_6698,N_2259,N_676);
xnor U6699 (N_6699,N_3236,N_4933);
nor U6700 (N_6700,N_3717,N_2907);
or U6701 (N_6701,N_827,N_811);
nor U6702 (N_6702,N_4584,N_6237);
nor U6703 (N_6703,N_5041,N_4699);
xnor U6704 (N_6704,N_3528,N_4335);
nand U6705 (N_6705,N_2167,N_6208);
xnor U6706 (N_6706,N_132,N_2168);
or U6707 (N_6707,N_2082,N_2433);
nor U6708 (N_6708,N_943,N_4207);
nand U6709 (N_6709,N_5869,N_1929);
or U6710 (N_6710,N_5956,N_5812);
or U6711 (N_6711,N_2800,N_4906);
or U6712 (N_6712,N_1783,N_3640);
nand U6713 (N_6713,N_5220,N_3689);
or U6714 (N_6714,N_1333,N_4999);
and U6715 (N_6715,N_3076,N_5326);
xor U6716 (N_6716,N_3518,N_5231);
or U6717 (N_6717,N_1663,N_5919);
and U6718 (N_6718,N_997,N_5207);
xnor U6719 (N_6719,N_1763,N_4713);
xor U6720 (N_6720,N_2154,N_2531);
nor U6721 (N_6721,N_4486,N_748);
and U6722 (N_6722,N_346,N_3508);
xor U6723 (N_6723,N_3315,N_3505);
nor U6724 (N_6724,N_3250,N_4163);
and U6725 (N_6725,N_5524,N_1720);
and U6726 (N_6726,N_5607,N_1850);
nand U6727 (N_6727,N_3280,N_1248);
nand U6728 (N_6728,N_2825,N_6190);
nand U6729 (N_6729,N_962,N_307);
or U6730 (N_6730,N_6138,N_1263);
and U6731 (N_6731,N_5554,N_1236);
or U6732 (N_6732,N_4376,N_2179);
nand U6733 (N_6733,N_1290,N_2566);
and U6734 (N_6734,N_3144,N_1606);
nand U6735 (N_6735,N_1986,N_1999);
xnor U6736 (N_6736,N_2011,N_1261);
xnor U6737 (N_6737,N_3441,N_2393);
and U6738 (N_6738,N_2117,N_4118);
or U6739 (N_6739,N_4505,N_212);
nand U6740 (N_6740,N_1141,N_944);
nand U6741 (N_6741,N_2049,N_1505);
xnor U6742 (N_6742,N_3598,N_4155);
xor U6743 (N_6743,N_1635,N_4002);
xor U6744 (N_6744,N_4390,N_1567);
nor U6745 (N_6745,N_2557,N_3830);
and U6746 (N_6746,N_2338,N_249);
or U6747 (N_6747,N_454,N_1381);
xnor U6748 (N_6748,N_252,N_1679);
nor U6749 (N_6749,N_1192,N_5394);
xnor U6750 (N_6750,N_4564,N_411);
xor U6751 (N_6751,N_5470,N_2635);
nand U6752 (N_6752,N_5370,N_2203);
or U6753 (N_6753,N_2925,N_5866);
xnor U6754 (N_6754,N_3743,N_3635);
or U6755 (N_6755,N_4142,N_5998);
or U6756 (N_6756,N_1725,N_2106);
and U6757 (N_6757,N_1164,N_1938);
nand U6758 (N_6758,N_4881,N_74);
nand U6759 (N_6759,N_587,N_4403);
nand U6760 (N_6760,N_5491,N_5787);
or U6761 (N_6761,N_1117,N_1810);
and U6762 (N_6762,N_3667,N_1382);
and U6763 (N_6763,N_5764,N_290);
or U6764 (N_6764,N_4759,N_1526);
nand U6765 (N_6765,N_4013,N_1087);
or U6766 (N_6766,N_625,N_4820);
and U6767 (N_6767,N_3209,N_1109);
or U6768 (N_6768,N_5121,N_732);
or U6769 (N_6769,N_4270,N_1817);
nand U6770 (N_6770,N_1058,N_2130);
and U6771 (N_6771,N_2075,N_709);
xnor U6772 (N_6772,N_1588,N_4595);
and U6773 (N_6773,N_3573,N_744);
nand U6774 (N_6774,N_46,N_2447);
or U6775 (N_6775,N_6005,N_3194);
nor U6776 (N_6776,N_828,N_3478);
xnor U6777 (N_6777,N_3681,N_5644);
nand U6778 (N_6778,N_378,N_5519);
or U6779 (N_6779,N_802,N_1312);
or U6780 (N_6780,N_1328,N_5704);
or U6781 (N_6781,N_1270,N_2898);
nor U6782 (N_6782,N_1626,N_2721);
and U6783 (N_6783,N_726,N_3089);
nor U6784 (N_6784,N_5761,N_3604);
nand U6785 (N_6785,N_3442,N_756);
xor U6786 (N_6786,N_584,N_841);
and U6787 (N_6787,N_673,N_5599);
xnor U6788 (N_6788,N_3737,N_6242);
xor U6789 (N_6789,N_65,N_5281);
nor U6790 (N_6790,N_4841,N_3517);
or U6791 (N_6791,N_3707,N_5794);
nor U6792 (N_6792,N_4873,N_2120);
nor U6793 (N_6793,N_2418,N_238);
xor U6794 (N_6794,N_2867,N_5185);
xor U6795 (N_6795,N_1955,N_208);
or U6796 (N_6796,N_595,N_3293);
nand U6797 (N_6797,N_2624,N_3523);
xnor U6798 (N_6798,N_2544,N_4381);
nor U6799 (N_6799,N_3989,N_879);
nand U6800 (N_6800,N_4960,N_136);
nand U6801 (N_6801,N_1305,N_6052);
and U6802 (N_6802,N_3515,N_2170);
xor U6803 (N_6803,N_3464,N_1849);
or U6804 (N_6804,N_5561,N_2838);
nand U6805 (N_6805,N_5295,N_2665);
xnor U6806 (N_6806,N_2255,N_874);
nand U6807 (N_6807,N_2718,N_3591);
nor U6808 (N_6808,N_3179,N_1580);
nor U6809 (N_6809,N_543,N_3261);
or U6810 (N_6810,N_3321,N_1949);
or U6811 (N_6811,N_4682,N_795);
nor U6812 (N_6812,N_2953,N_955);
xnor U6813 (N_6813,N_2916,N_2410);
xor U6814 (N_6814,N_4768,N_3653);
xnor U6815 (N_6815,N_1877,N_158);
or U6816 (N_6816,N_2331,N_1871);
or U6817 (N_6817,N_4761,N_2470);
nand U6818 (N_6818,N_792,N_2128);
and U6819 (N_6819,N_818,N_2057);
xnor U6820 (N_6820,N_3917,N_6157);
nor U6821 (N_6821,N_173,N_1377);
xor U6822 (N_6822,N_385,N_5831);
nand U6823 (N_6823,N_3739,N_3428);
and U6824 (N_6824,N_4687,N_6108);
nand U6825 (N_6825,N_58,N_1165);
nand U6826 (N_6826,N_3988,N_2125);
xnor U6827 (N_6827,N_3350,N_644);
nor U6828 (N_6828,N_3119,N_1316);
and U6829 (N_6829,N_4623,N_1005);
or U6830 (N_6830,N_2784,N_755);
xnor U6831 (N_6831,N_374,N_2416);
xnor U6832 (N_6832,N_6174,N_1105);
nand U6833 (N_6833,N_1904,N_2748);
nand U6834 (N_6834,N_1385,N_1425);
xnor U6835 (N_6835,N_4171,N_387);
and U6836 (N_6836,N_4843,N_3206);
nand U6837 (N_6837,N_3759,N_1836);
xnor U6838 (N_6838,N_5141,N_1461);
nor U6839 (N_6839,N_4069,N_6042);
nor U6840 (N_6840,N_830,N_1128);
or U6841 (N_6841,N_3100,N_2633);
and U6842 (N_6842,N_1532,N_5842);
xor U6843 (N_6843,N_981,N_4408);
or U6844 (N_6844,N_5247,N_3160);
or U6845 (N_6845,N_20,N_2515);
nand U6846 (N_6846,N_5708,N_6072);
nor U6847 (N_6847,N_1294,N_3937);
nand U6848 (N_6848,N_3335,N_5642);
nand U6849 (N_6849,N_5007,N_663);
and U6850 (N_6850,N_2943,N_4545);
or U6851 (N_6851,N_4992,N_1541);
nor U6852 (N_6852,N_3716,N_3164);
nand U6853 (N_6853,N_1304,N_2673);
nand U6854 (N_6854,N_4784,N_1677);
xnor U6855 (N_6855,N_2363,N_4636);
and U6856 (N_6856,N_4130,N_5897);
nand U6857 (N_6857,N_875,N_5450);
nand U6858 (N_6858,N_986,N_1011);
nor U6859 (N_6859,N_254,N_3403);
nor U6860 (N_6860,N_2793,N_835);
nor U6861 (N_6861,N_4182,N_2348);
or U6862 (N_6862,N_2602,N_804);
and U6863 (N_6863,N_4416,N_5814);
and U6864 (N_6864,N_5437,N_4520);
nand U6865 (N_6865,N_3770,N_30);
nor U6866 (N_6866,N_3897,N_6105);
xor U6867 (N_6867,N_4258,N_4043);
nand U6868 (N_6868,N_3572,N_1257);
xor U6869 (N_6869,N_2286,N_2367);
and U6870 (N_6870,N_5645,N_4401);
nor U6871 (N_6871,N_5567,N_263);
and U6872 (N_6872,N_1214,N_2474);
nor U6873 (N_6873,N_3694,N_2215);
xor U6874 (N_6874,N_1813,N_2242);
xnor U6875 (N_6875,N_177,N_1088);
nor U6876 (N_6876,N_3161,N_1708);
nor U6877 (N_6877,N_1168,N_1596);
xor U6878 (N_6878,N_2977,N_5238);
nor U6879 (N_6879,N_2195,N_4608);
or U6880 (N_6880,N_1360,N_4345);
xor U6881 (N_6881,N_478,N_2209);
or U6882 (N_6882,N_1894,N_1232);
nor U6883 (N_6883,N_5249,N_4045);
or U6884 (N_6884,N_5789,N_3402);
xor U6885 (N_6885,N_5667,N_5531);
and U6886 (N_6886,N_2336,N_2579);
and U6887 (N_6887,N_3306,N_1244);
nand U6888 (N_6888,N_2988,N_988);
and U6889 (N_6889,N_4668,N_1854);
nand U6890 (N_6890,N_2243,N_1041);
or U6891 (N_6891,N_2223,N_301);
xor U6892 (N_6892,N_99,N_1549);
xnor U6893 (N_6893,N_960,N_396);
xnor U6894 (N_6894,N_5489,N_6244);
nor U6895 (N_6895,N_4651,N_917);
or U6896 (N_6896,N_1740,N_853);
nor U6897 (N_6897,N_5357,N_2102);
nor U6898 (N_6898,N_1636,N_5055);
nor U6899 (N_6899,N_5685,N_5413);
nor U6900 (N_6900,N_3944,N_3873);
xnor U6901 (N_6901,N_4015,N_3724);
nand U6902 (N_6902,N_180,N_3840);
or U6903 (N_6903,N_5726,N_398);
or U6904 (N_6904,N_1398,N_5444);
nor U6905 (N_6905,N_223,N_1930);
and U6906 (N_6906,N_809,N_3991);
or U6907 (N_6907,N_698,N_5313);
and U6908 (N_6908,N_741,N_1354);
nand U6909 (N_6909,N_699,N_4814);
xor U6910 (N_6910,N_437,N_6177);
xor U6911 (N_6911,N_2600,N_4215);
nand U6912 (N_6912,N_5903,N_355);
nor U6913 (N_6913,N_1737,N_4127);
or U6914 (N_6914,N_1423,N_3363);
or U6915 (N_6915,N_3487,N_4077);
xor U6916 (N_6916,N_5195,N_2813);
or U6917 (N_6917,N_975,N_1669);
or U6918 (N_6918,N_925,N_160);
nand U6919 (N_6919,N_4031,N_2710);
nand U6920 (N_6920,N_6230,N_5975);
nand U6921 (N_6921,N_2431,N_159);
or U6922 (N_6922,N_5739,N_2420);
and U6923 (N_6923,N_1330,N_631);
xor U6924 (N_6924,N_6233,N_2029);
or U6925 (N_6925,N_4474,N_3120);
xor U6926 (N_6926,N_1210,N_1958);
or U6927 (N_6927,N_3018,N_3356);
nand U6928 (N_6928,N_6140,N_6068);
and U6929 (N_6929,N_3132,N_930);
and U6930 (N_6930,N_696,N_3977);
and U6931 (N_6931,N_3888,N_2138);
xor U6932 (N_6932,N_530,N_4354);
or U6933 (N_6933,N_5521,N_5780);
nor U6934 (N_6934,N_4298,N_5905);
xnor U6935 (N_6935,N_2554,N_2957);
or U6936 (N_6936,N_1619,N_565);
nand U6937 (N_6937,N_685,N_312);
nor U6938 (N_6938,N_5734,N_2573);
nor U6939 (N_6939,N_2208,N_887);
nand U6940 (N_6940,N_3411,N_5432);
or U6941 (N_6941,N_4740,N_2240);
nor U6942 (N_6942,N_2779,N_3167);
xnor U6943 (N_6943,N_3567,N_5201);
nand U6944 (N_6944,N_5971,N_3863);
nand U6945 (N_6945,N_5047,N_3633);
and U6946 (N_6946,N_2503,N_1479);
nand U6947 (N_6947,N_1145,N_5454);
and U6948 (N_6948,N_2658,N_3843);
nand U6949 (N_6949,N_666,N_3507);
nand U6950 (N_6950,N_1918,N_2939);
nor U6951 (N_6951,N_4846,N_749);
xnor U6952 (N_6952,N_3143,N_1157);
xnor U6953 (N_6953,N_5129,N_3986);
xnor U6954 (N_6954,N_345,N_3802);
nor U6955 (N_6955,N_2409,N_2292);
and U6956 (N_6956,N_2593,N_2885);
nor U6957 (N_6957,N_3570,N_2291);
nor U6958 (N_6958,N_2437,N_5383);
xor U6959 (N_6959,N_4097,N_1375);
xnor U6960 (N_6960,N_5626,N_5114);
xor U6961 (N_6961,N_4200,N_4492);
xnor U6962 (N_6962,N_786,N_5600);
nor U6963 (N_6963,N_4628,N_483);
and U6964 (N_6964,N_3963,N_5019);
xnor U6965 (N_6965,N_5581,N_2941);
xnor U6966 (N_6966,N_4137,N_4934);
and U6967 (N_6967,N_3855,N_3422);
nor U6968 (N_6968,N_2180,N_2832);
nand U6969 (N_6969,N_4561,N_5837);
nand U6970 (N_6970,N_1115,N_4212);
xnor U6971 (N_6971,N_2501,N_2671);
or U6972 (N_6972,N_2722,N_3495);
or U6973 (N_6973,N_3158,N_444);
nor U6974 (N_6974,N_4263,N_5853);
and U6975 (N_6975,N_5820,N_776);
nor U6976 (N_6976,N_2881,N_1881);
nand U6977 (N_6977,N_4918,N_4538);
nand U6978 (N_6978,N_6055,N_5952);
and U6979 (N_6979,N_751,N_5828);
and U6980 (N_6980,N_2497,N_4387);
or U6981 (N_6981,N_4034,N_2111);
and U6982 (N_6982,N_3482,N_2092);
nand U6983 (N_6983,N_3920,N_2998);
nand U6984 (N_6984,N_3336,N_2528);
and U6985 (N_6985,N_583,N_4415);
nor U6986 (N_6986,N_3004,N_2731);
nand U6987 (N_6987,N_2369,N_898);
nor U6988 (N_6988,N_2521,N_854);
or U6989 (N_6989,N_451,N_4009);
nand U6990 (N_6990,N_2306,N_655);
or U6991 (N_6991,N_4493,N_3023);
nor U6992 (N_6992,N_3713,N_2205);
xnor U6993 (N_6993,N_1131,N_4790);
or U6994 (N_6994,N_4323,N_4819);
or U6995 (N_6995,N_652,N_3747);
or U6996 (N_6996,N_185,N_1478);
nor U6997 (N_6997,N_4149,N_564);
nor U6998 (N_6998,N_2017,N_3361);
nor U6999 (N_6999,N_5827,N_1457);
nand U7000 (N_7000,N_2693,N_2271);
and U7001 (N_7001,N_1362,N_4627);
and U7002 (N_7002,N_6131,N_2392);
nand U7003 (N_7003,N_1943,N_1488);
nor U7004 (N_7004,N_6056,N_5826);
xor U7005 (N_7005,N_6144,N_5659);
and U7006 (N_7006,N_2065,N_5878);
and U7007 (N_7007,N_4280,N_790);
and U7008 (N_7008,N_5609,N_4062);
nand U7009 (N_7009,N_5311,N_4022);
nor U7010 (N_7010,N_5829,N_5506);
or U7011 (N_7011,N_5935,N_3800);
and U7012 (N_7012,N_1199,N_5525);
xor U7013 (N_7013,N_4423,N_2599);
nor U7014 (N_7014,N_1644,N_4642);
nand U7015 (N_7015,N_1055,N_149);
and U7016 (N_7016,N_1786,N_3268);
nand U7017 (N_7017,N_1887,N_1313);
nor U7018 (N_7018,N_6194,N_368);
and U7019 (N_7019,N_3068,N_1386);
xnor U7020 (N_7020,N_1950,N_3235);
nor U7021 (N_7021,N_2987,N_554);
xnor U7022 (N_7022,N_2031,N_466);
nor U7023 (N_7023,N_3786,N_3896);
xnor U7024 (N_7024,N_4476,N_6113);
nor U7025 (N_7025,N_3844,N_499);
and U7026 (N_7026,N_3395,N_6047);
nor U7027 (N_7027,N_4990,N_3174);
and U7028 (N_7028,N_277,N_3548);
or U7029 (N_7029,N_1279,N_1866);
nand U7030 (N_7030,N_203,N_4667);
and U7031 (N_7031,N_4141,N_2353);
xor U7032 (N_7032,N_1043,N_519);
nand U7033 (N_7033,N_2864,N_560);
xnor U7034 (N_7034,N_5052,N_3065);
nand U7035 (N_7035,N_6186,N_4741);
nand U7036 (N_7036,N_1508,N_101);
and U7037 (N_7037,N_2715,N_5515);
or U7038 (N_7038,N_2048,N_1132);
nand U7039 (N_7039,N_4449,N_4020);
or U7040 (N_7040,N_3,N_4098);
nand U7041 (N_7041,N_5977,N_5399);
nor U7042 (N_7042,N_605,N_5723);
and U7043 (N_7043,N_3776,N_5379);
nand U7044 (N_7044,N_3574,N_6095);
and U7045 (N_7045,N_2414,N_4088);
nand U7046 (N_7046,N_6059,N_905);
nand U7047 (N_7047,N_5166,N_2828);
nor U7048 (N_7048,N_3381,N_2088);
nor U7049 (N_7049,N_3083,N_3494);
nand U7050 (N_7050,N_3409,N_3646);
nand U7051 (N_7051,N_3155,N_5660);
and U7052 (N_7052,N_6076,N_3380);
xnor U7053 (N_7053,N_2144,N_1489);
nor U7054 (N_7054,N_430,N_5818);
xnor U7055 (N_7055,N_2556,N_1651);
nor U7056 (N_7056,N_596,N_5617);
and U7057 (N_7057,N_2264,N_2761);
and U7058 (N_7058,N_4923,N_902);
xor U7059 (N_7059,N_2354,N_912);
nor U7060 (N_7060,N_2415,N_669);
nand U7061 (N_7061,N_4714,N_123);
or U7062 (N_7062,N_335,N_4237);
xnor U7063 (N_7063,N_6051,N_2561);
and U7064 (N_7064,N_964,N_4494);
or U7065 (N_7065,N_5629,N_4542);
and U7066 (N_7066,N_933,N_913);
nor U7067 (N_7067,N_540,N_3463);
or U7068 (N_7068,N_4330,N_3946);
nand U7069 (N_7069,N_4117,N_2590);
nor U7070 (N_7070,N_4152,N_5083);
nand U7071 (N_7071,N_3479,N_1161);
nand U7072 (N_7072,N_4364,N_1442);
nand U7073 (N_7073,N_1231,N_4025);
nor U7074 (N_7074,N_4269,N_498);
nor U7075 (N_7075,N_3421,N_4592);
and U7076 (N_7076,N_1324,N_3278);
nand U7077 (N_7077,N_6175,N_3714);
and U7078 (N_7078,N_152,N_3327);
xor U7079 (N_7079,N_1978,N_63);
or U7080 (N_7080,N_4213,N_4896);
or U7081 (N_7081,N_1018,N_4081);
and U7082 (N_7082,N_4400,N_672);
and U7083 (N_7083,N_7,N_2127);
and U7084 (N_7084,N_5158,N_2606);
nand U7085 (N_7085,N_2663,N_1933);
nand U7086 (N_7086,N_740,N_1432);
xnor U7087 (N_7087,N_5799,N_1873);
nand U7088 (N_7088,N_2342,N_5886);
or U7089 (N_7089,N_5944,N_2880);
or U7090 (N_7090,N_730,N_6159);
nor U7091 (N_7091,N_3357,N_3943);
xnor U7092 (N_7092,N_5256,N_3303);
xor U7093 (N_7093,N_117,N_5947);
nor U7094 (N_7094,N_2958,N_708);
nand U7095 (N_7095,N_3601,N_5732);
nand U7096 (N_7096,N_4673,N_1700);
and U7097 (N_7097,N_3037,N_198);
nor U7098 (N_7098,N_5738,N_4734);
xnor U7099 (N_7099,N_5268,N_4122);
nor U7100 (N_7100,N_4644,N_5200);
and U7101 (N_7101,N_5139,N_3349);
and U7102 (N_7102,N_5931,N_2989);
nand U7103 (N_7103,N_1019,N_6062);
or U7104 (N_7104,N_3490,N_1401);
nand U7105 (N_7105,N_179,N_64);
or U7106 (N_7106,N_1755,N_3024);
and U7107 (N_7107,N_1695,N_358);
nand U7108 (N_7108,N_752,N_1083);
xor U7109 (N_7109,N_862,N_5104);
nor U7110 (N_7110,N_294,N_164);
and U7111 (N_7111,N_985,N_3071);
and U7112 (N_7112,N_1997,N_683);
or U7113 (N_7113,N_3915,N_3386);
xor U7114 (N_7114,N_1762,N_5942);
nor U7115 (N_7115,N_3824,N_4793);
nand U7116 (N_7116,N_5805,N_1864);
or U7117 (N_7117,N_4365,N_2830);
nor U7118 (N_7118,N_3659,N_6003);
nand U7119 (N_7119,N_5967,N_4404);
nand U7120 (N_7120,N_4342,N_2686);
nand U7121 (N_7121,N_1184,N_2668);
and U7122 (N_7122,N_5002,N_1793);
nor U7123 (N_7123,N_3025,N_1438);
nand U7124 (N_7124,N_2104,N_2000);
nor U7125 (N_7125,N_1195,N_113);
nand U7126 (N_7126,N_5164,N_344);
xnor U7127 (N_7127,N_3513,N_6248);
nor U7128 (N_7128,N_747,N_2268);
xor U7129 (N_7129,N_3212,N_735);
nor U7130 (N_7130,N_200,N_5894);
or U7131 (N_7131,N_2448,N_4425);
xor U7132 (N_7132,N_3549,N_5363);
xor U7133 (N_7133,N_1583,N_6164);
nor U7134 (N_7134,N_5681,N_5286);
or U7135 (N_7135,N_4962,N_25);
xnor U7136 (N_7136,N_2453,N_4360);
or U7137 (N_7137,N_1256,N_2173);
nand U7138 (N_7138,N_972,N_1841);
and U7139 (N_7139,N_2499,N_2767);
nor U7140 (N_7140,N_2614,N_4647);
and U7141 (N_7141,N_800,N_459);
and U7142 (N_7142,N_4888,N_69);
xnor U7143 (N_7143,N_2035,N_4134);
nand U7144 (N_7144,N_243,N_4870);
nand U7145 (N_7145,N_4460,N_2491);
and U7146 (N_7146,N_1995,N_5611);
and U7147 (N_7147,N_2797,N_1899);
and U7148 (N_7148,N_5108,N_2214);
or U7149 (N_7149,N_4921,N_289);
and U7150 (N_7150,N_2045,N_1545);
nor U7151 (N_7151,N_216,N_606);
xnor U7152 (N_7152,N_2545,N_2489);
nor U7153 (N_7153,N_1100,N_4597);
nand U7154 (N_7154,N_5301,N_140);
nor U7155 (N_7155,N_3657,N_4733);
or U7156 (N_7156,N_2654,N_481);
nand U7157 (N_7157,N_1506,N_693);
nor U7158 (N_7158,N_4334,N_4328);
nor U7159 (N_7159,N_4284,N_1935);
or U7160 (N_7160,N_5124,N_5934);
nand U7161 (N_7161,N_165,N_4185);
and U7162 (N_7162,N_5463,N_2696);
nand U7163 (N_7163,N_108,N_3529);
nand U7164 (N_7164,N_1255,N_832);
and U7165 (N_7165,N_1736,N_3705);
xnor U7166 (N_7166,N_4705,N_4337);
xnor U7167 (N_7167,N_717,N_527);
and U7168 (N_7168,N_2917,N_839);
nand U7169 (N_7169,N_2766,N_4206);
and U7170 (N_7170,N_2372,N_1080);
nor U7171 (N_7171,N_1135,N_1601);
nand U7172 (N_7172,N_4902,N_1153);
or U7173 (N_7173,N_5098,N_2135);
nor U7174 (N_7174,N_5616,N_5641);
nand U7175 (N_7175,N_5012,N_253);
nor U7176 (N_7176,N_4708,N_360);
nand U7177 (N_7177,N_1130,N_2692);
nand U7178 (N_7178,N_6037,N_4003);
nand U7179 (N_7179,N_4363,N_4103);
nor U7180 (N_7180,N_880,N_2853);
nor U7181 (N_7181,N_2476,N_2870);
and U7182 (N_7182,N_1140,N_3021);
xnor U7183 (N_7183,N_4554,N_4685);
and U7184 (N_7184,N_3255,N_337);
or U7185 (N_7185,N_4656,N_2581);
nor U7186 (N_7186,N_3214,N_674);
and U7187 (N_7187,N_2032,N_5698);
or U7188 (N_7188,N_6171,N_2013);
or U7189 (N_7189,N_1287,N_963);
nand U7190 (N_7190,N_3775,N_648);
nand U7191 (N_7191,N_4198,N_1334);
and U7192 (N_7192,N_147,N_3305);
nand U7193 (N_7193,N_715,N_3594);
xor U7194 (N_7194,N_1956,N_2061);
nor U7195 (N_7195,N_3095,N_3524);
and U7196 (N_7196,N_684,N_3377);
or U7197 (N_7197,N_3769,N_2230);
or U7198 (N_7198,N_3320,N_670);
xnor U7199 (N_7199,N_4719,N_156);
nand U7200 (N_7200,N_505,N_3832);
nand U7201 (N_7201,N_1310,N_5154);
or U7202 (N_7202,N_3627,N_174);
and U7203 (N_7203,N_2166,N_1625);
nand U7204 (N_7204,N_1543,N_5255);
nor U7205 (N_7205,N_5320,N_5961);
nor U7206 (N_7206,N_6193,N_1211);
and U7207 (N_7207,N_3861,N_5318);
and U7208 (N_7208,N_5666,N_4725);
and U7209 (N_7209,N_2882,N_3251);
nand U7210 (N_7210,N_1383,N_4649);
nor U7211 (N_7211,N_589,N_81);
nor U7212 (N_7212,N_4080,N_3726);
xor U7213 (N_7213,N_4822,N_1538);
xnor U7214 (N_7214,N_274,N_1040);
xnor U7215 (N_7215,N_4382,N_677);
xnor U7216 (N_7216,N_3569,N_2836);
xnor U7217 (N_7217,N_642,N_5544);
and U7218 (N_7218,N_5907,N_1565);
nor U7219 (N_7219,N_3639,N_4925);
xor U7220 (N_7220,N_2373,N_729);
nor U7221 (N_7221,N_4679,N_3289);
or U7222 (N_7222,N_4052,N_3001);
nand U7223 (N_7223,N_3376,N_4614);
xor U7224 (N_7224,N_3779,N_1185);
xor U7225 (N_7225,N_4972,N_5279);
and U7226 (N_7226,N_3695,N_6211);
nand U7227 (N_7227,N_3533,N_5864);
or U7228 (N_7228,N_6152,N_633);
and U7229 (N_7229,N_4857,N_5543);
and U7230 (N_7230,N_1091,N_1503);
xnor U7231 (N_7231,N_266,N_2729);
or U7232 (N_7232,N_1373,N_3771);
nand U7233 (N_7233,N_5387,N_5758);
xnor U7234 (N_7234,N_6010,N_4044);
nand U7235 (N_7235,N_3352,N_2623);
or U7236 (N_7236,N_1855,N_2076);
nand U7237 (N_7237,N_547,N_6148);
nor U7238 (N_7238,N_660,N_3267);
nand U7239 (N_7239,N_3355,N_4650);
and U7240 (N_7240,N_6077,N_362);
xor U7241 (N_7241,N_941,N_3565);
xor U7242 (N_7242,N_183,N_1858);
or U7243 (N_7243,N_4301,N_2955);
nand U7244 (N_7244,N_3347,N_143);
nor U7245 (N_7245,N_3831,N_1616);
or U7246 (N_7246,N_6243,N_2788);
nand U7247 (N_7247,N_4271,N_5073);
nor U7248 (N_7248,N_2429,N_5217);
nor U7249 (N_7249,N_4499,N_5501);
and U7250 (N_7250,N_6120,N_1730);
nor U7251 (N_7251,N_2172,N_3718);
and U7252 (N_7252,N_3332,N_1965);
nand U7253 (N_7253,N_5857,N_488);
nand U7254 (N_7254,N_6013,N_193);
nand U7255 (N_7255,N_1982,N_128);
nor U7256 (N_7256,N_2737,N_4643);
or U7257 (N_7257,N_1747,N_4795);
or U7258 (N_7258,N_5890,N_594);
nand U7259 (N_7259,N_6058,N_2669);
nor U7260 (N_7260,N_341,N_2398);
and U7261 (N_7261,N_2612,N_4478);
nand U7262 (N_7262,N_4059,N_5742);
nor U7263 (N_7263,N_855,N_5653);
xor U7264 (N_7264,N_6012,N_2177);
nor U7265 (N_7265,N_3066,N_1566);
or U7266 (N_7266,N_3862,N_2400);
xnor U7267 (N_7267,N_3879,N_255);
and U7268 (N_7268,N_5677,N_4261);
xnor U7269 (N_7269,N_1509,N_1205);
xnor U7270 (N_7270,N_1202,N_1002);
and U7271 (N_7271,N_5507,N_2043);
nor U7272 (N_7272,N_2176,N_967);
nor U7273 (N_7273,N_3124,N_3432);
xnor U7274 (N_7274,N_4837,N_357);
nand U7275 (N_7275,N_1366,N_5223);
nand U7276 (N_7276,N_2644,N_3162);
xor U7277 (N_7277,N_3026,N_3701);
xor U7278 (N_7278,N_1306,N_3141);
and U7279 (N_7279,N_1654,N_3007);
nand U7280 (N_7280,N_3401,N_3557);
nand U7281 (N_7281,N_381,N_1143);
xnor U7282 (N_7282,N_1909,N_4503);
nand U7283 (N_7283,N_2523,N_300);
nand U7284 (N_7284,N_1487,N_2469);
xnor U7285 (N_7285,N_2384,N_1474);
nor U7286 (N_7286,N_1726,N_3762);
or U7287 (N_7287,N_5895,N_5331);
and U7288 (N_7288,N_3603,N_4230);
xor U7289 (N_7289,N_3566,N_1796);
nand U7290 (N_7290,N_586,N_736);
nand U7291 (N_7291,N_2472,N_245);
nor U7292 (N_7292,N_1670,N_1927);
nand U7293 (N_7293,N_1554,N_2295);
nor U7294 (N_7294,N_75,N_1078);
or U7295 (N_7295,N_2364,N_2576);
nand U7296 (N_7296,N_5571,N_2679);
xnor U7297 (N_7297,N_5583,N_5700);
and U7298 (N_7298,N_3735,N_338);
xnor U7299 (N_7299,N_5173,N_4522);
nor U7300 (N_7300,N_5523,N_4698);
nor U7301 (N_7301,N_4411,N_1824);
xnor U7302 (N_7302,N_470,N_3221);
nor U7303 (N_7303,N_176,N_6142);
or U7304 (N_7304,N_3393,N_3296);
and U7305 (N_7305,N_4633,N_767);
and U7306 (N_7306,N_1764,N_4266);
and U7307 (N_7307,N_1917,N_3545);
nor U7308 (N_7308,N_501,N_3097);
nand U7309 (N_7309,N_3469,N_104);
xnor U7310 (N_7310,N_658,N_3204);
xnor U7311 (N_7311,N_6030,N_5297);
nor U7312 (N_7312,N_4236,N_2869);
xor U7313 (N_7313,N_3622,N_6085);
nor U7314 (N_7314,N_4767,N_4565);
nand U7315 (N_7315,N_495,N_5362);
nand U7316 (N_7316,N_5912,N_3279);
and U7317 (N_7317,N_5443,N_3360);
or U7318 (N_7318,N_1133,N_2443);
and U7319 (N_7319,N_4176,N_297);
nand U7320 (N_7320,N_2992,N_4654);
nand U7321 (N_7321,N_3334,N_4177);
or U7322 (N_7322,N_4010,N_1598);
nand U7323 (N_7323,N_3597,N_1882);
xor U7324 (N_7324,N_5750,N_1671);
and U7325 (N_7325,N_3941,N_4630);
nand U7326 (N_7326,N_2053,N_918);
and U7327 (N_7327,N_3485,N_1661);
nor U7328 (N_7328,N_1496,N_6125);
or U7329 (N_7329,N_370,N_3792);
or U7330 (N_7330,N_4359,N_2677);
and U7331 (N_7331,N_5070,N_5377);
nand U7332 (N_7332,N_6075,N_1738);
and U7333 (N_7333,N_5590,N_3313);
xor U7334 (N_7334,N_2834,N_856);
and U7335 (N_7335,N_1082,N_2449);
xor U7336 (N_7336,N_2539,N_2839);
and U7337 (N_7337,N_4594,N_4245);
or U7338 (N_7338,N_3823,N_5233);
and U7339 (N_7339,N_3092,N_3733);
or U7340 (N_7340,N_3287,N_3562);
nor U7341 (N_7341,N_5060,N_745);
nand U7342 (N_7342,N_2391,N_1144);
xnor U7343 (N_7343,N_4927,N_1523);
xor U7344 (N_7344,N_6115,N_5982);
or U7345 (N_7345,N_134,N_1352);
or U7346 (N_7346,N_2837,N_5436);
xnor U7347 (N_7347,N_5134,N_4046);
and U7348 (N_7348,N_4179,N_3138);
nor U7349 (N_7349,N_864,N_1681);
and U7350 (N_7350,N_3431,N_553);
xnor U7351 (N_7351,N_2274,N_3029);
or U7352 (N_7352,N_195,N_2362);
nor U7353 (N_7353,N_3300,N_2700);
or U7354 (N_7354,N_4153,N_4504);
xor U7355 (N_7355,N_3419,N_2931);
nor U7356 (N_7356,N_5593,N_5596);
and U7357 (N_7357,N_4086,N_2627);
and U7358 (N_7358,N_3017,N_3677);
and U7359 (N_7359,N_2740,N_1447);
nor U7360 (N_7360,N_2293,N_3827);
or U7361 (N_7361,N_1667,N_6071);
xor U7362 (N_7362,N_1966,N_3767);
and U7363 (N_7363,N_4414,N_4047);
or U7364 (N_7364,N_4456,N_4321);
nor U7365 (N_7365,N_3238,N_2126);
nor U7366 (N_7366,N_6092,N_5289);
xor U7367 (N_7367,N_1099,N_2577);
and U7368 (N_7368,N_5307,N_4575);
nand U7369 (N_7369,N_4468,N_2206);
xnor U7370 (N_7370,N_1402,N_1338);
xor U7371 (N_7371,N_1766,N_5550);
xnor U7372 (N_7372,N_3006,N_5926);
nor U7373 (N_7373,N_5987,N_3553);
and U7374 (N_7374,N_235,N_5592);
or U7375 (N_7375,N_4168,N_3157);
and U7376 (N_7376,N_6207,N_3675);
nor U7377 (N_7377,N_4129,N_5462);
xor U7378 (N_7378,N_3429,N_2136);
and U7379 (N_7379,N_4297,N_4079);
nand U7380 (N_7380,N_611,N_2921);
xor U7381 (N_7381,N_2892,N_3543);
and U7382 (N_7382,N_1851,N_4798);
and U7383 (N_7383,N_5516,N_2754);
and U7384 (N_7384,N_1839,N_5615);
nand U7385 (N_7385,N_1919,N_3199);
and U7386 (N_7386,N_3809,N_2307);
xnor U7387 (N_7387,N_5579,N_6172);
or U7388 (N_7388,N_3211,N_2359);
and U7389 (N_7389,N_4602,N_320);
nand U7390 (N_7390,N_3893,N_4974);
nor U7391 (N_7391,N_1594,N_4235);
nor U7392 (N_7392,N_4380,N_1259);
or U7393 (N_7393,N_731,N_1410);
nand U7394 (N_7394,N_2010,N_4418);
nor U7395 (N_7395,N_1533,N_5813);
or U7396 (N_7396,N_4247,N_19);
nand U7397 (N_7397,N_2909,N_2062);
nand U7398 (N_7398,N_1300,N_3254);
xor U7399 (N_7399,N_1070,N_2310);
and U7400 (N_7400,N_566,N_983);
nor U7401 (N_7401,N_646,N_2278);
nand U7402 (N_7402,N_5763,N_1664);
xor U7403 (N_7403,N_4856,N_3822);
nor U7404 (N_7404,N_2,N_4903);
and U7405 (N_7405,N_1431,N_2643);
nand U7406 (N_7406,N_4277,N_3014);
or U7407 (N_7407,N_4802,N_3128);
nand U7408 (N_7408,N_6023,N_6121);
or U7409 (N_7409,N_4558,N_2439);
xor U7410 (N_7410,N_536,N_4420);
or U7411 (N_7411,N_939,N_5757);
or U7412 (N_7412,N_1595,N_5321);
and U7413 (N_7413,N_1822,N_4222);
xnor U7414 (N_7414,N_3763,N_2162);
nor U7415 (N_7415,N_4481,N_4955);
nand U7416 (N_7416,N_3889,N_85);
and U7417 (N_7417,N_1191,N_1863);
nand U7418 (N_7418,N_4288,N_6245);
or U7419 (N_7419,N_5672,N_5566);
and U7420 (N_7420,N_5441,N_4306);
xor U7421 (N_7421,N_3999,N_1156);
or U7422 (N_7422,N_1237,N_2450);
or U7423 (N_7423,N_783,N_4170);
and U7424 (N_7424,N_2419,N_3645);
or U7425 (N_7425,N_3976,N_995);
xor U7426 (N_7426,N_999,N_2585);
and U7427 (N_7427,N_369,N_2568);
or U7428 (N_7428,N_3749,N_2358);
or U7429 (N_7429,N_3877,N_5721);
or U7430 (N_7430,N_1376,N_3821);
and U7431 (N_7431,N_770,N_3643);
and U7432 (N_7432,N_1921,N_2222);
nand U7433 (N_7433,N_3796,N_178);
and U7434 (N_7434,N_5719,N_3404);
nor U7435 (N_7435,N_2538,N_1693);
nor U7436 (N_7436,N_414,N_1844);
and U7437 (N_7437,N_4368,N_5694);
and U7438 (N_7438,N_3875,N_5883);
nand U7439 (N_7439,N_4242,N_5442);
and U7440 (N_7440,N_6187,N_5668);
and U7441 (N_7441,N_260,N_1038);
xor U7442 (N_7442,N_620,N_946);
xnor U7443 (N_7443,N_4736,N_2250);
or U7444 (N_7444,N_400,N_4551);
or U7445 (N_7445,N_1530,N_5847);
nand U7446 (N_7446,N_3731,N_54);
nor U7447 (N_7447,N_576,N_3193);
nor U7448 (N_7448,N_2257,N_4007);
and U7449 (N_7449,N_6020,N_601);
xor U7450 (N_7450,N_145,N_6160);
nor U7451 (N_7451,N_3765,N_4658);
xor U7452 (N_7452,N_4915,N_4101);
or U7453 (N_7453,N_1534,N_2378);
and U7454 (N_7454,N_426,N_840);
xnor U7455 (N_7455,N_2727,N_794);
nor U7456 (N_7456,N_3812,N_4578);
nor U7457 (N_7457,N_5316,N_5974);
xnor U7458 (N_7458,N_5774,N_1678);
and U7459 (N_7459,N_17,N_4700);
xnor U7460 (N_7460,N_2165,N_1761);
xor U7461 (N_7461,N_5765,N_3218);
xnor U7462 (N_7462,N_1378,N_3819);
nor U7463 (N_7463,N_5453,N_4959);
nor U7464 (N_7464,N_196,N_4506);
xor U7465 (N_7465,N_366,N_4998);
nand U7466 (N_7466,N_5069,N_282);
nand U7467 (N_7467,N_2790,N_5710);
xnor U7468 (N_7468,N_2506,N_6064);
xnor U7469 (N_7469,N_1416,N_2379);
nor U7470 (N_7470,N_2287,N_5473);
nand U7471 (N_7471,N_2428,N_5171);
and U7472 (N_7472,N_4556,N_1891);
and U7473 (N_7473,N_4599,N_4113);
or U7474 (N_7474,N_327,N_3379);
nor U7475 (N_7475,N_4978,N_2887);
nor U7476 (N_7476,N_1504,N_891);
nand U7477 (N_7477,N_5426,N_1056);
xor U7478 (N_7478,N_1059,N_2937);
nand U7479 (N_7479,N_5786,N_4457);
xor U7480 (N_7480,N_6150,N_334);
xor U7481 (N_7481,N_5924,N_5655);
and U7482 (N_7482,N_4491,N_1309);
or U7483 (N_7483,N_847,N_127);
nor U7484 (N_7484,N_1069,N_2866);
nor U7485 (N_7485,N_1968,N_721);
and U7486 (N_7486,N_2063,N_4464);
nand U7487 (N_7487,N_2005,N_5749);
nor U7488 (N_7488,N_937,N_824);
or U7489 (N_7489,N_5338,N_4982);
nand U7490 (N_7490,N_214,N_2334);
or U7491 (N_7491,N_2547,N_167);
or U7492 (N_7492,N_4760,N_3641);
nor U7493 (N_7493,N_4318,N_3197);
nand U7494 (N_7494,N_4537,N_1942);
or U7495 (N_7495,N_2335,N_3610);
nand U7496 (N_7496,N_5161,N_2621);
and U7497 (N_7497,N_484,N_1633);
or U7498 (N_7498,N_5254,N_2097);
and U7499 (N_7499,N_4274,N_979);
or U7500 (N_7500,N_6234,N_5405);
nand U7501 (N_7501,N_3869,N_5712);
nand U7502 (N_7502,N_5497,N_1295);
xor U7503 (N_7503,N_3139,N_5754);
and U7504 (N_7504,N_5933,N_5627);
nor U7505 (N_7505,N_1630,N_894);
xor U7506 (N_7506,N_2632,N_2247);
xnor U7507 (N_7507,N_2877,N_2121);
nand U7508 (N_7508,N_2194,N_1470);
nand U7509 (N_7509,N_279,N_3472);
xnor U7510 (N_7510,N_3751,N_5401);
nor U7511 (N_7511,N_6236,N_5358);
or U7512 (N_7512,N_383,N_1318);
nand U7513 (N_7513,N_1712,N_2025);
xor U7514 (N_7514,N_1267,N_3434);
or U7515 (N_7515,N_2914,N_5332);
nand U7516 (N_7516,N_6158,N_77);
nand U7517 (N_7517,N_5954,N_5715);
nor U7518 (N_7518,N_5778,N_5492);
nand U7519 (N_7519,N_4458,N_3514);
and U7520 (N_7520,N_4729,N_4783);
nand U7521 (N_7521,N_2810,N_5340);
xor U7522 (N_7522,N_978,N_4225);
and U7523 (N_7523,N_3647,N_1947);
xnor U7524 (N_7524,N_4479,N_1676);
nor U7525 (N_7525,N_5425,N_393);
nor U7526 (N_7526,N_4488,N_120);
and U7527 (N_7527,N_5939,N_2008);
or U7528 (N_7528,N_1838,N_4813);
xor U7529 (N_7529,N_137,N_3227);
and U7530 (N_7530,N_2899,N_1514);
or U7531 (N_7531,N_269,N_4073);
nand U7532 (N_7532,N_6102,N_5649);
or U7533 (N_7533,N_6031,N_1170);
nand U7534 (N_7534,N_4576,N_5270);
xor U7535 (N_7535,N_3930,N_5009);
or U7536 (N_7536,N_5988,N_157);
or U7537 (N_7537,N_4910,N_2374);
or U7538 (N_7538,N_5386,N_511);
nand U7539 (N_7539,N_5736,N_5679);
nand U7540 (N_7540,N_1575,N_574);
and U7541 (N_7541,N_1903,N_3521);
nor U7542 (N_7542,N_3286,N_2639);
or U7543 (N_7543,N_2829,N_4904);
xnor U7544 (N_7544,N_5287,N_5585);
or U7545 (N_7545,N_982,N_3820);
xor U7546 (N_7546,N_3414,N_5132);
or U7547 (N_7547,N_5819,N_3516);
nor U7548 (N_7548,N_4664,N_2653);
or U7549 (N_7549,N_3813,N_1574);
nand U7550 (N_7550,N_5259,N_2345);
and U7551 (N_7551,N_1953,N_3968);
xnor U7552 (N_7552,N_2683,N_5973);
nor U7553 (N_7553,N_3850,N_3341);
xnor U7554 (N_7554,N_4786,N_5755);
and U7555 (N_7555,N_5402,N_1806);
and U7556 (N_7556,N_2553,N_6039);
nor U7557 (N_7557,N_4435,N_4577);
and U7558 (N_7558,N_1351,N_1349);
or U7559 (N_7559,N_1463,N_4095);
or U7560 (N_7560,N_1315,N_6179);
nand U7561 (N_7561,N_395,N_1450);
nor U7562 (N_7562,N_1846,N_4618);
and U7563 (N_7563,N_5372,N_1845);
nand U7564 (N_7564,N_2077,N_264);
or U7565 (N_7565,N_4517,N_3682);
nand U7566 (N_7566,N_4739,N_2003);
nor U7567 (N_7567,N_3459,N_3502);
nor U7568 (N_7568,N_2302,N_2231);
nand U7569 (N_7569,N_1417,N_1152);
nand U7570 (N_7570,N_4138,N_2896);
or U7571 (N_7571,N_425,N_3654);
nor U7572 (N_7572,N_4842,N_5434);
nand U7573 (N_7573,N_2272,N_1827);
and U7574 (N_7574,N_5675,N_3723);
nand U7575 (N_7575,N_5706,N_5678);
and U7576 (N_7576,N_2438,N_4939);
and U7577 (N_7577,N_2047,N_3730);
xor U7578 (N_7578,N_5260,N_1392);
nor U7579 (N_7579,N_1230,N_2744);
and U7580 (N_7580,N_6015,N_4611);
xnor U7581 (N_7581,N_4966,N_4037);
or U7582 (N_7582,N_5623,N_5839);
or U7583 (N_7583,N_868,N_700);
nor U7584 (N_7584,N_4467,N_1167);
xor U7585 (N_7585,N_1320,N_3368);
or U7586 (N_7586,N_772,N_3461);
nor U7587 (N_7587,N_4737,N_4484);
nor U7588 (N_7588,N_4994,N_5771);
nor U7589 (N_7589,N_2772,N_1483);
or U7590 (N_7590,N_376,N_401);
nand U7591 (N_7591,N_4262,N_1485);
nand U7592 (N_7592,N_1789,N_497);
or U7593 (N_7593,N_4890,N_6029);
xnor U7594 (N_7594,N_3208,N_5276);
or U7595 (N_7595,N_4979,N_32);
and U7596 (N_7596,N_1286,N_3519);
xor U7597 (N_7597,N_4151,N_3440);
or U7598 (N_7598,N_6153,N_2451);
nand U7599 (N_7599,N_773,N_4920);
and U7600 (N_7600,N_186,N_5068);
and U7601 (N_7601,N_1116,N_4477);
or U7602 (N_7602,N_2096,N_2963);
nand U7603 (N_7603,N_5598,N_4429);
or U7604 (N_7604,N_4776,N_4894);
nor U7605 (N_7605,N_4958,N_4473);
or U7606 (N_7606,N_3715,N_4068);
or U7607 (N_7607,N_420,N_537);
xnor U7608 (N_7608,N_2862,N_1805);
nor U7609 (N_7609,N_4174,N_679);
nand U7610 (N_7610,N_4123,N_1758);
xor U7611 (N_7611,N_5851,N_801);
or U7612 (N_7612,N_4877,N_4541);
xor U7613 (N_7613,N_4371,N_998);
or U7614 (N_7614,N_599,N_3192);
xor U7615 (N_7615,N_2492,N_419);
nor U7616 (N_7616,N_5464,N_4393);
nor U7617 (N_7617,N_0,N_754);
nor U7618 (N_7618,N_1754,N_2743);
nor U7619 (N_7619,N_598,N_5356);
xnor U7620 (N_7620,N_4255,N_1529);
nand U7621 (N_7621,N_3805,N_4448);
xnor U7622 (N_7622,N_651,N_5870);
xor U7623 (N_7623,N_3925,N_2555);
nor U7624 (N_7624,N_4124,N_5344);
xnor U7625 (N_7625,N_228,N_3534);
or U7626 (N_7626,N_4087,N_1862);
xor U7627 (N_7627,N_2232,N_5868);
xnor U7628 (N_7628,N_4279,N_6044);
nor U7629 (N_7629,N_2610,N_965);
and U7630 (N_7630,N_2454,N_4655);
nor U7631 (N_7631,N_575,N_4833);
or U7632 (N_7632,N_1249,N_3895);
and U7633 (N_7633,N_1435,N_3787);
or U7634 (N_7634,N_5511,N_3854);
or U7635 (N_7635,N_5684,N_2114);
and U7636 (N_7636,N_1544,N_568);
xor U7637 (N_7637,N_4796,N_1561);
nor U7638 (N_7638,N_3971,N_2550);
xor U7639 (N_7639,N_3282,N_4327);
and U7640 (N_7640,N_352,N_3177);
nor U7641 (N_7641,N_2891,N_5396);
xnor U7642 (N_7642,N_1183,N_3298);
xor U7643 (N_7643,N_4482,N_881);
nand U7644 (N_7644,N_299,N_4826);
nor U7645 (N_7645,N_4373,N_4041);
xnor U7646 (N_7646,N_522,N_1053);
nor U7647 (N_7647,N_3632,N_1017);
or U7648 (N_7648,N_785,N_2326);
nor U7649 (N_7649,N_544,N_2072);
xnor U7650 (N_7650,N_5701,N_5807);
or U7651 (N_7651,N_6083,N_5084);
nand U7652 (N_7652,N_1093,N_1308);
xor U7653 (N_7653,N_3452,N_5051);
and U7654 (N_7654,N_2681,N_591);
xnor U7655 (N_7655,N_5613,N_1742);
nand U7656 (N_7656,N_5024,N_3423);
or U7657 (N_7657,N_6132,N_122);
nor U7658 (N_7658,N_5336,N_250);
xnor U7659 (N_7659,N_333,N_4817);
nor U7660 (N_7660,N_6198,N_4366);
and U7661 (N_7661,N_2207,N_545);
xor U7662 (N_7662,N_4652,N_3069);
nor U7663 (N_7663,N_2704,N_1010);
and U7664 (N_7664,N_5631,N_2565);
xor U7665 (N_7665,N_2140,N_2984);
nand U7666 (N_7666,N_1768,N_3010);
nor U7667 (N_7667,N_3232,N_2997);
nor U7668 (N_7668,N_1418,N_5428);
nor U7669 (N_7669,N_80,N_1227);
and U7670 (N_7670,N_3816,N_4516);
or U7671 (N_7671,N_4716,N_6122);
nor U7672 (N_7672,N_1120,N_4144);
or U7673 (N_7673,N_468,N_2151);
nand U7674 (N_7674,N_3841,N_1704);
nor U7675 (N_7675,N_1213,N_3696);
and U7676 (N_7676,N_4340,N_1820);
and U7677 (N_7677,N_4607,N_6188);
or U7678 (N_7678,N_162,N_1706);
or U7679 (N_7679,N_1073,N_3965);
xnor U7680 (N_7680,N_3899,N_5948);
or U7681 (N_7681,N_4472,N_2004);
xor U7682 (N_7682,N_1068,N_796);
xor U7683 (N_7683,N_2478,N_1674);
xnor U7684 (N_7684,N_5236,N_2583);
nor U7685 (N_7685,N_2249,N_5167);
or U7686 (N_7686,N_706,N_3661);
or U7687 (N_7687,N_516,N_3585);
nand U7688 (N_7688,N_2426,N_2770);
and U7689 (N_7689,N_3532,N_2860);
or U7690 (N_7690,N_2930,N_4665);
nand U7691 (N_7691,N_1006,N_5815);
or U7692 (N_7692,N_2283,N_5513);
or U7693 (N_7693,N_6006,N_6045);
xor U7694 (N_7694,N_1137,N_2074);
nand U7695 (N_7695,N_3849,N_1653);
xor U7696 (N_7696,N_4912,N_5528);
nand U7697 (N_7697,N_5096,N_2263);
or U7698 (N_7698,N_5713,N_3766);
and U7699 (N_7699,N_5488,N_3094);
or U7700 (N_7700,N_2339,N_5830);
nor U7701 (N_7701,N_1014,N_2001);
nand U7702 (N_7702,N_1585,N_5020);
nor U7703 (N_7703,N_4265,N_3655);
nor U7704 (N_7704,N_5039,N_871);
nand U7705 (N_7705,N_4106,N_5088);
or U7706 (N_7706,N_5992,N_2244);
and U7707 (N_7707,N_2929,N_1136);
nor U7708 (N_7708,N_2161,N_5490);
and U7709 (N_7709,N_3060,N_4099);
or U7710 (N_7710,N_2071,N_5062);
or U7711 (N_7711,N_49,N_4310);
nand U7712 (N_7712,N_5147,N_3009);
and U7713 (N_7713,N_3867,N_2200);
nand U7714 (N_7714,N_4661,N_1952);
or U7715 (N_7715,N_2801,N_5825);
and U7716 (N_7716,N_2216,N_556);
nand U7717 (N_7717,N_5219,N_43);
and U7718 (N_7718,N_4232,N_4748);
and U7719 (N_7719,N_205,N_5709);
or U7720 (N_7720,N_1618,N_3903);
and U7721 (N_7721,N_5729,N_4093);
nor U7722 (N_7722,N_2149,N_433);
nor U7723 (N_7723,N_258,N_993);
nand U7724 (N_7724,N_4434,N_1459);
nand U7725 (N_7725,N_3922,N_4946);
nand U7726 (N_7726,N_959,N_3362);
xor U7727 (N_7727,N_4957,N_5135);
and U7728 (N_7728,N_6176,N_5335);
and U7729 (N_7729,N_5744,N_924);
nand U7730 (N_7730,N_5835,N_5747);
xor U7731 (N_7731,N_5252,N_844);
xor U7732 (N_7732,N_190,N_3798);
and U7733 (N_7733,N_1065,N_970);
nand U7734 (N_7734,N_3761,N_3118);
and U7735 (N_7735,N_1683,N_3159);
xnor U7736 (N_7736,N_3489,N_3496);
nand U7737 (N_7737,N_1460,N_5978);
or U7738 (N_7738,N_5911,N_4585);
nor U7739 (N_7739,N_240,N_4441);
nand U7740 (N_7740,N_559,N_5773);
or U7741 (N_7741,N_5180,N_931);
nand U7742 (N_7742,N_5017,N_878);
or U7743 (N_7743,N_347,N_4752);
xnor U7744 (N_7744,N_230,N_4603);
and U7745 (N_7745,N_1944,N_3081);
nor U7746 (N_7746,N_3918,N_4913);
xor U7747 (N_7747,N_3240,N_2006);
nor U7748 (N_7748,N_2723,N_1206);
xnor U7749 (N_7749,N_5689,N_3249);
nand U7750 (N_7750,N_572,N_6082);
or U7751 (N_7751,N_4136,N_2604);
xnor U7752 (N_7752,N_1033,N_6200);
nor U7753 (N_7753,N_1472,N_3453);
nor U7754 (N_7754,N_3987,N_2603);
nor U7755 (N_7755,N_2728,N_10);
xnor U7756 (N_7756,N_3836,N_2267);
and U7757 (N_7757,N_4135,N_4971);
nand U7758 (N_7758,N_5334,N_552);
nand U7759 (N_7759,N_1134,N_1825);
xor U7760 (N_7760,N_284,N_5354);
nor U7761 (N_7761,N_5539,N_3801);
or U7762 (N_7762,N_231,N_1340);
nor U7763 (N_7763,N_4653,N_2423);
nor U7764 (N_7764,N_1200,N_2241);
nand U7765 (N_7765,N_3182,N_5406);
nand U7766 (N_7766,N_4322,N_3080);
xnor U7767 (N_7767,N_5133,N_4774);
nand U7768 (N_7768,N_2468,N_3994);
and U7769 (N_7769,N_3480,N_1658);
and U7770 (N_7770,N_4818,N_4956);
and U7771 (N_7771,N_2237,N_4780);
and U7772 (N_7772,N_5885,N_4094);
and U7773 (N_7773,N_1668,N_3375);
xor U7774 (N_7774,N_4102,N_2424);
nand U7775 (N_7775,N_4004,N_1707);
nor U7776 (N_7776,N_5292,N_4527);
or U7777 (N_7777,N_1776,N_3184);
or U7778 (N_7778,N_4534,N_4811);
xnor U7779 (N_7779,N_2893,N_1880);
or U7780 (N_7780,N_3427,N_3202);
xor U7781 (N_7781,N_3264,N_1902);
nand U7782 (N_7782,N_4375,N_3493);
and U7783 (N_7783,N_4951,N_3308);
and U7784 (N_7784,N_5214,N_2831);
or U7785 (N_7785,N_5165,N_3173);
or U7786 (N_7786,N_2191,N_1221);
nand U7787 (N_7787,N_5415,N_4943);
nor U7788 (N_7788,N_3291,N_4944);
nand U7789 (N_7789,N_4562,N_5481);
nor U7790 (N_7790,N_3670,N_5061);
and U7791 (N_7791,N_2823,N_5028);
or U7792 (N_7792,N_4286,N_1814);
xnor U7793 (N_7793,N_4501,N_4461);
xnor U7794 (N_7794,N_2594,N_5226);
and U7795 (N_7795,N_3237,N_5138);
nand U7796 (N_7796,N_3626,N_1811);
xor U7797 (N_7797,N_2178,N_1388);
and U7798 (N_7798,N_1246,N_4569);
and U7799 (N_7799,N_5602,N_3075);
or U7800 (N_7800,N_5816,N_2938);
nand U7801 (N_7801,N_1557,N_4357);
and U7802 (N_7802,N_619,N_47);
or U7803 (N_7803,N_1792,N_3062);
nand U7804 (N_7804,N_2051,N_5000);
nand U7805 (N_7805,N_2978,N_5136);
nand U7806 (N_7806,N_4257,N_935);
nor U7807 (N_7807,N_2652,N_3082);
and U7808 (N_7808,N_6091,N_5540);
nand U7809 (N_7809,N_3871,N_209);
xnor U7810 (N_7810,N_5664,N_2421);
nor U7811 (N_7811,N_4749,N_224);
nand U7812 (N_7812,N_3107,N_4051);
and U7813 (N_7813,N_102,N_4240);
and U7814 (N_7814,N_187,N_604);
nor U7815 (N_7815,N_5230,N_4273);
nor U7816 (N_7816,N_3942,N_2258);
xor U7817 (N_7817,N_1691,N_3413);
xnor U7818 (N_7818,N_6094,N_4372);
nand U7819 (N_7819,N_330,N_4278);
nand U7820 (N_7820,N_2487,N_4469);
nor U7821 (N_7821,N_4396,N_1743);
or U7822 (N_7822,N_3599,N_2526);
nor U7823 (N_7823,N_4126,N_787);
xnor U7824 (N_7824,N_3790,N_5250);
xor U7825 (N_7825,N_4299,N_5461);
nand U7826 (N_7826,N_1188,N_3746);
and U7827 (N_7827,N_4834,N_3500);
and U7828 (N_7828,N_4358,N_5184);
nand U7829 (N_7829,N_2567,N_377);
or U7830 (N_7830,N_2146,N_2575);
xnor U7831 (N_7831,N_2405,N_447);
nor U7832 (N_7832,N_5533,N_1576);
and U7833 (N_7833,N_5638,N_5143);
and U7834 (N_7834,N_87,N_5097);
nand U7835 (N_7835,N_5025,N_118);
or U7836 (N_7836,N_1973,N_16);
and U7837 (N_7837,N_4311,N_13);
nor U7838 (N_7838,N_6147,N_2562);
and U7839 (N_7839,N_4732,N_5651);
or U7840 (N_7840,N_954,N_4601);
nor U7841 (N_7841,N_3782,N_5079);
nand U7842 (N_7842,N_5503,N_455);
nand U7843 (N_7843,N_4502,N_1025);
nand U7844 (N_7844,N_1641,N_3391);
and U7845 (N_7845,N_1138,N_3027);
nand U7846 (N_7846,N_2777,N_5957);
xor U7847 (N_7847,N_3002,N_6124);
xor U7848 (N_7848,N_3086,N_5381);
xnor U7849 (N_7849,N_3420,N_5555);
nand U7850 (N_7850,N_1941,N_1201);
xor U7851 (N_7851,N_4128,N_2994);
nor U7852 (N_7852,N_3587,N_4409);
nor U7853 (N_7853,N_242,N_608);
or U7854 (N_7854,N_607,N_276);
and U7855 (N_7855,N_125,N_1498);
nor U7856 (N_7856,N_275,N_1353);
nor U7857 (N_7857,N_2542,N_2855);
or U7858 (N_7858,N_763,N_3036);
and U7859 (N_7859,N_5654,N_5059);
xnor U7860 (N_7860,N_4406,N_4907);
xor U7861 (N_7861,N_873,N_6191);
nor U7862 (N_7862,N_6007,N_4808);
or U7863 (N_7863,N_5465,N_5179);
nor U7864 (N_7864,N_27,N_1951);
and U7865 (N_7865,N_5414,N_3912);
nand U7866 (N_7866,N_1439,N_1421);
nor U7867 (N_7867,N_4529,N_5665);
nand U7868 (N_7868,N_1771,N_5768);
and U7869 (N_7869,N_1370,N_5731);
nand U7870 (N_7870,N_4947,N_4806);
and U7871 (N_7871,N_5575,N_664);
nand U7872 (N_7872,N_3927,N_2190);
or U7873 (N_7873,N_2786,N_281);
or U7874 (N_7874,N_1971,N_5963);
nand U7875 (N_7875,N_4747,N_533);
and U7876 (N_7876,N_2559,N_6004);
nand U7877 (N_7877,N_3928,N_4082);
and U7878 (N_7878,N_1883,N_681);
xor U7879 (N_7879,N_889,N_2811);
nand U7880 (N_7880,N_2730,N_4550);
nand U7881 (N_7881,N_6093,N_4905);
nor U7882 (N_7882,N_2044,N_5122);
nand U7883 (N_7883,N_5152,N_4285);
or U7884 (N_7884,N_5485,N_3614);
and U7885 (N_7885,N_4621,N_3539);
or U7886 (N_7886,N_2402,N_876);
nor U7887 (N_7887,N_2456,N_6220);
or U7888 (N_7888,N_44,N_657);
xor U7889 (N_7889,N_3000,N_1035);
nand U7890 (N_7890,N_927,N_4911);
xnor U7891 (N_7891,N_4662,N_2674);
nand U7892 (N_7892,N_4453,N_1957);
or U7893 (N_7893,N_1874,N_5892);
or U7894 (N_7894,N_630,N_5574);
and U7895 (N_7895,N_201,N_1302);
or U7896 (N_7896,N_4514,N_5591);
and U7897 (N_7897,N_3911,N_3997);
or U7898 (N_7898,N_1837,N_2965);
xnor U7899 (N_7899,N_5422,N_3908);
xnor U7900 (N_7900,N_825,N_1834);
xnor U7901 (N_7901,N_3791,N_5745);
nand U7902 (N_7902,N_4132,N_4451);
nand U7903 (N_7903,N_2375,N_1552);
nand U7904 (N_7904,N_3467,N_2314);
nor U7905 (N_7905,N_5793,N_1593);
or U7906 (N_7906,N_4029,N_1307);
nor U7907 (N_7907,N_3219,N_1175);
nand U7908 (N_7908,N_2108,N_760);
xor U7909 (N_7909,N_4121,N_5549);
nand U7910 (N_7910,N_4470,N_4392);
nand U7911 (N_7911,N_5469,N_4771);
xor U7912 (N_7912,N_1335,N_2002);
and U7913 (N_7913,N_1856,N_3535);
nand U7914 (N_7914,N_1452,N_4238);
and U7915 (N_7915,N_2697,N_2764);
and U7916 (N_7916,N_513,N_5730);
xnor U7917 (N_7917,N_1962,N_5845);
or U7918 (N_7918,N_969,N_5440);
xor U7919 (N_7919,N_5077,N_2124);
and U7920 (N_7920,N_1499,N_5996);
and U7921 (N_7921,N_1512,N_3195);
xnor U7922 (N_7922,N_2611,N_3814);
xor U7923 (N_7923,N_5804,N_1238);
nor U7924 (N_7924,N_2970,N_2548);
nor U7925 (N_7925,N_3135,N_4156);
nor U7926 (N_7926,N_1672,N_4590);
and U7927 (N_7927,N_4825,N_866);
nor U7928 (N_7928,N_546,N_1314);
and U7929 (N_7929,N_6240,N_1905);
nor U7930 (N_7930,N_5006,N_500);
xnor U7931 (N_7931,N_4524,N_5683);
or U7932 (N_7932,N_712,N_5510);
and U7933 (N_7933,N_5810,N_2629);
nand U7934 (N_7934,N_3642,N_1077);
nor U7935 (N_7935,N_5618,N_3067);
nand U7936 (N_7936,N_1251,N_3892);
nand U7937 (N_7937,N_5359,N_5285);
nor U7938 (N_7938,N_2019,N_6182);
nor U7939 (N_7939,N_3629,N_1112);
xor U7940 (N_7940,N_1085,N_3166);
nand U7941 (N_7941,N_1067,N_4855);
xnor U7942 (N_7942,N_904,N_3272);
and U7943 (N_7943,N_1709,N_1391);
and U7944 (N_7944,N_3056,N_3186);
nand U7945 (N_7945,N_3592,N_5824);
or U7946 (N_7946,N_5099,N_1111);
or U7947 (N_7947,N_4231,N_5112);
nor U7948 (N_7948,N_5248,N_3757);
and U7949 (N_7949,N_5467,N_2211);
xnor U7950 (N_7950,N_6109,N_2317);
or U7951 (N_7951,N_808,N_2319);
or U7952 (N_7952,N_5221,N_4049);
nand U7953 (N_7953,N_3470,N_5530);
xnor U7954 (N_7954,N_2083,N_4197);
and U7955 (N_7955,N_1437,N_4341);
or U7956 (N_7956,N_5915,N_4391);
and U7957 (N_7957,N_798,N_551);
and U7958 (N_7958,N_617,N_4419);
and U7959 (N_7959,N_325,N_714);
or U7960 (N_7960,N_4785,N_3126);
nor U7961 (N_7961,N_109,N_206);
or U7962 (N_7962,N_4823,N_3865);
nand U7963 (N_7963,N_4544,N_6184);
nand U7964 (N_7964,N_3673,N_1522);
and U7965 (N_7965,N_261,N_5187);
and U7966 (N_7966,N_4938,N_391);
xnor U7967 (N_7967,N_1688,N_2616);
nand U7968 (N_7968,N_4800,N_5071);
or U7969 (N_7969,N_2227,N_3106);
xor U7970 (N_7970,N_3190,N_3638);
xor U7971 (N_7971,N_2103,N_3740);
nor U7972 (N_7972,N_2923,N_246);
xor U7973 (N_7973,N_4204,N_623);
nor U7974 (N_7974,N_3721,N_508);
nor U7975 (N_7975,N_1223,N_309);
xor U7976 (N_7976,N_6228,N_600);
and U7977 (N_7977,N_121,N_2856);
nor U7978 (N_7978,N_1282,N_4712);
nor U7979 (N_7979,N_2504,N_2995);
nor U7980 (N_7980,N_1384,N_529);
xor U7981 (N_7981,N_919,N_1780);
nand U7982 (N_7982,N_4463,N_1652);
nand U7983 (N_7983,N_4507,N_3935);
or U7984 (N_7984,N_4932,N_5949);
nand U7985 (N_7985,N_774,N_3475);
xor U7986 (N_7986,N_5170,N_769);
xnor U7987 (N_7987,N_6063,N_4061);
or U7988 (N_7988,N_1974,N_221);
and U7989 (N_7989,N_453,N_5089);
and U7990 (N_7990,N_5514,N_4559);
or U7991 (N_7991,N_2184,N_2116);
xnor U7992 (N_7992,N_4119,N_5109);
or U7993 (N_7993,N_2256,N_2666);
and U7994 (N_7994,N_4727,N_4293);
xnor U7995 (N_7995,N_1621,N_42);
xor U7996 (N_7996,N_6112,N_4076);
xor U7997 (N_7997,N_5846,N_2684);
nor U7998 (N_7998,N_1744,N_3454);
or U7999 (N_7999,N_3520,N_4884);
or U8000 (N_8000,N_5352,N_2996);
xor U8001 (N_8001,N_4876,N_2537);
nor U8002 (N_8002,N_2656,N_1716);
xor U8003 (N_8003,N_6026,N_4332);
nand U8004 (N_8004,N_3881,N_3583);
and U8005 (N_8005,N_2490,N_5508);
xnor U8006 (N_8006,N_5423,N_2734);
nand U8007 (N_8007,N_34,N_1393);
and U8008 (N_8008,N_1149,N_4096);
nand U8009 (N_8009,N_4686,N_95);
or U8010 (N_8010,N_438,N_640);
nor U8011 (N_8011,N_3274,N_3547);
or U8012 (N_8012,N_3540,N_4591);
nor U8013 (N_8013,N_5930,N_3894);
nor U8014 (N_8014,N_5235,N_1224);
and U8015 (N_8015,N_6009,N_4462);
and U8016 (N_8016,N_4402,N_2479);
and U8017 (N_8017,N_5026,N_3079);
xor U8018 (N_8018,N_3637,N_57);
and U8019 (N_8019,N_2807,N_1114);
xor U8020 (N_8020,N_1367,N_2551);
nand U8021 (N_8021,N_6239,N_3530);
nor U8022 (N_8022,N_6232,N_3615);
or U8023 (N_8023,N_116,N_2636);
nand U8024 (N_8024,N_1409,N_480);
nor U8025 (N_8025,N_114,N_4530);
nor U8026 (N_8026,N_4053,N_3383);
xnor U8027 (N_8027,N_93,N_1269);
xnor U8028 (N_8028,N_990,N_3323);
and U8029 (N_8029,N_5459,N_4312);
and U8030 (N_8030,N_5937,N_3447);
nor U8031 (N_8031,N_487,N_5244);
and U8032 (N_8032,N_788,N_5772);
xnor U8033 (N_8033,N_4543,N_6218);
xor U8034 (N_8034,N_3226,N_4861);
xnor U8035 (N_8035,N_5687,N_1920);
nor U8036 (N_8036,N_1356,N_4731);
nand U8037 (N_8037,N_2477,N_5361);
xnor U8038 (N_8038,N_3061,N_1357);
or U8039 (N_8039,N_446,N_3806);
nand U8040 (N_8040,N_4532,N_810);
and U8041 (N_8041,N_4483,N_1363);
nand U8042 (N_8042,N_6216,N_823);
and U8043 (N_8043,N_3188,N_3618);
nand U8044 (N_8044,N_4175,N_5189);
or U8045 (N_8045,N_5717,N_5397);
nand U8046 (N_8046,N_1749,N_2281);
xor U8047 (N_8047,N_5861,N_5431);
and U8048 (N_8048,N_3329,N_6227);
xor U8049 (N_8049,N_5172,N_3388);
nand U8050 (N_8050,N_1913,N_771);
and U8051 (N_8051,N_4275,N_3322);
or U8052 (N_8052,N_3504,N_4055);
and U8053 (N_8053,N_5115,N_5887);
or U8054 (N_8054,N_635,N_4355);
nor U8055 (N_8055,N_4264,N_3926);
and U8056 (N_8056,N_4317,N_1390);
or U8057 (N_8057,N_5576,N_5535);
or U8058 (N_8058,N_5430,N_3055);
nand U8059 (N_8059,N_384,N_3990);
or U8060 (N_8060,N_3077,N_4612);
and U8061 (N_8061,N_1326,N_3181);
or U8062 (N_8062,N_5671,N_2760);
and U8063 (N_8063,N_2768,N_5498);
nor U8064 (N_8064,N_4645,N_1615);
nand U8065 (N_8065,N_850,N_2069);
or U8066 (N_8066,N_4580,N_6049);
or U8067 (N_8067,N_4849,N_2934);
nand U8068 (N_8068,N_1696,N_5480);
nand U8069 (N_8069,N_1179,N_5913);
nand U8070 (N_8070,N_4600,N_4928);
nand U8071 (N_8071,N_2662,N_4710);
nand U8072 (N_8072,N_1823,N_6154);
and U8073 (N_8073,N_5832,N_48);
nor U8074 (N_8074,N_5972,N_4224);
nand U8075 (N_8075,N_5206,N_6098);
and U8076 (N_8076,N_1843,N_1129);
nand U8077 (N_8077,N_4981,N_5955);
and U8078 (N_8078,N_2814,N_3955);
xnor U8079 (N_8079,N_2441,N_5403);
nand U8080 (N_8080,N_2445,N_4214);
nand U8081 (N_8081,N_3378,N_4715);
nor U8082 (N_8082,N_83,N_668);
or U8083 (N_8083,N_3110,N_467);
nand U8084 (N_8084,N_4487,N_4011);
nand U8085 (N_8085,N_1964,N_5595);
and U8086 (N_8086,N_6246,N_3742);
xnor U8087 (N_8087,N_3147,N_2672);
or U8088 (N_8088,N_1264,N_2850);
or U8089 (N_8089,N_5439,N_5280);
nor U8090 (N_8090,N_2826,N_1301);
and U8091 (N_8091,N_6204,N_910);
xor U8092 (N_8092,N_2408,N_207);
nand U8093 (N_8093,N_2858,N_5293);
nor U8094 (N_8094,N_1895,N_1151);
nand U8095 (N_8095,N_4398,N_2248);
xor U8096 (N_8096,N_2058,N_3113);
and U8097 (N_8097,N_4028,N_815);
or U8098 (N_8098,N_3712,N_2525);
and U8099 (N_8099,N_2514,N_1480);
and U8100 (N_8100,N_3448,N_2799);
nor U8101 (N_8101,N_1896,N_616);
nor U8102 (N_8102,N_2541,N_1072);
xor U8103 (N_8103,N_2042,N_2313);
or U8104 (N_8104,N_6041,N_2199);
nand U8105 (N_8105,N_5562,N_932);
xor U8106 (N_8106,N_3133,N_2522);
nand U8107 (N_8107,N_4405,N_5191);
nand U8108 (N_8108,N_5228,N_2253);
nand U8109 (N_8109,N_1934,N_3466);
nor U8110 (N_8110,N_4008,N_1998);
or U8111 (N_8111,N_713,N_3623);
nor U8112 (N_8112,N_6022,N_4535);
xor U8113 (N_8113,N_3443,N_5460);
and U8114 (N_8114,N_5610,N_4871);
nor U8115 (N_8115,N_3481,N_3033);
and U8116 (N_8116,N_5163,N_5565);
nand U8117 (N_8117,N_4139,N_3104);
nand U8118 (N_8118,N_3923,N_5929);
and U8119 (N_8119,N_2712,N_1815);
nor U8120 (N_8120,N_4816,N_539);
nor U8121 (N_8121,N_791,N_28);
or U8122 (N_8122,N_1840,N_6028);
and U8123 (N_8123,N_4229,N_2308);
or U8124 (N_8124,N_4762,N_5714);
nor U8125 (N_8125,N_328,N_3145);
nand U8126 (N_8126,N_5435,N_3405);
nand U8127 (N_8127,N_3105,N_3117);
xor U8128 (N_8128,N_4721,N_1193);
or U8129 (N_8129,N_4307,N_528);
nand U8130 (N_8130,N_4782,N_6170);
nand U8131 (N_8131,N_5412,N_3973);
and U8132 (N_8132,N_6084,N_5748);
nor U8133 (N_8133,N_2143,N_5048);
nand U8134 (N_8134,N_2900,N_1589);
and U8135 (N_8135,N_4194,N_403);
xor U8136 (N_8136,N_3163,N_2724);
nor U8137 (N_8137,N_768,N_1910);
nand U8138 (N_8138,N_1021,N_4697);
or U8139 (N_8139,N_3424,N_4480);
and U8140 (N_8140,N_5053,N_2444);
nor U8141 (N_8141,N_5608,N_326);
or U8142 (N_8142,N_5411,N_686);
and U8143 (N_8143,N_1685,N_1096);
or U8144 (N_8144,N_1829,N_4634);
nand U8145 (N_8145,N_1629,N_5204);
nor U8146 (N_8146,N_6166,N_3309);
xnor U8147 (N_8147,N_1050,N_4523);
xor U8148 (N_8148,N_4965,N_1443);
nand U8149 (N_8149,N_2664,N_417);
or U8150 (N_8150,N_4508,N_3439);
and U8151 (N_8151,N_1028,N_2746);
nor U8152 (N_8152,N_1121,N_1258);
nand U8153 (N_8153,N_3187,N_4201);
xor U8154 (N_8154,N_3945,N_3588);
nand U8155 (N_8155,N_2738,N_671);
nand U8156 (N_8156,N_4773,N_4742);
xor U8157 (N_8157,N_2620,N_2808);
and U8158 (N_8158,N_6008,N_489);
and U8159 (N_8159,N_6002,N_1611);
nor U8160 (N_8160,N_5265,N_3392);
xor U8161 (N_8161,N_82,N_3898);
or U8162 (N_8162,N_232,N_2110);
nand U8163 (N_8163,N_4893,N_3175);
xnor U8164 (N_8164,N_2628,N_4353);
nand U8165 (N_8165,N_2819,N_1502);
or U8166 (N_8166,N_1799,N_138);
and U8167 (N_8167,N_1586,N_2446);
or U8168 (N_8168,N_5733,N_5175);
nand U8169 (N_8169,N_56,N_1274);
and U8170 (N_8170,N_4005,N_107);
and U8171 (N_8171,N_5720,N_4948);
nor U8172 (N_8172,N_3940,N_1980);
and U8173 (N_8173,N_5718,N_1798);
or U8174 (N_8174,N_1404,N_2196);
nor U8175 (N_8175,N_1173,N_356);
and U8176 (N_8176,N_5225,N_5674);
nand U8177 (N_8177,N_1110,N_3860);
xnor U8178 (N_8178,N_2960,N_1835);
or U8179 (N_8179,N_4490,N_6219);
nor U8180 (N_8180,N_1125,N_5728);
and U8181 (N_8181,N_5945,N_5447);
xor U8182 (N_8182,N_1901,N_115);
nor U8183 (N_8183,N_3577,N_2912);
nor U8184 (N_8184,N_5727,N_4292);
nor U8185 (N_8185,N_2841,N_5916);
nor U8186 (N_8186,N_2289,N_4940);
nand U8187 (N_8187,N_989,N_682);
nand U8188 (N_8188,N_2266,N_4241);
xnor U8189 (N_8189,N_1163,N_1623);
xor U8190 (N_8190,N_5690,N_2638);
nand U8191 (N_8191,N_4519,N_5495);
nand U8192 (N_8192,N_6038,N_1492);
and U8193 (N_8193,N_3127,N_5458);
or U8194 (N_8194,N_2404,N_5901);
nand U8195 (N_8195,N_2933,N_4572);
nor U8196 (N_8196,N_3552,N_6145);
or U8197 (N_8197,N_2461,N_1071);
and U8198 (N_8198,N_5553,N_6127);
nor U8199 (N_8199,N_237,N_2455);
or U8200 (N_8200,N_2948,N_1397);
nand U8201 (N_8201,N_5630,N_3752);
and U8202 (N_8202,N_579,N_1970);
xnor U8203 (N_8203,N_3471,N_2833);
nand U8204 (N_8204,N_351,N_3931);
nand U8205 (N_8205,N_68,N_2647);
xnor U8206 (N_8206,N_1660,N_1892);
nor U8207 (N_8207,N_3883,N_4648);
or U8208 (N_8208,N_4244,N_5737);
and U8209 (N_8209,N_1454,N_4146);
and U8210 (N_8210,N_3134,N_2333);
and U8211 (N_8211,N_4573,N_1468);
or U8212 (N_8212,N_4963,N_55);
nor U8213 (N_8213,N_4084,N_5072);
xor U8214 (N_8214,N_2460,N_813);
nand U8215 (N_8215,N_3703,N_2073);
and U8216 (N_8216,N_3560,N_4838);
nor U8217 (N_8217,N_1016,N_2763);
xor U8218 (N_8218,N_5875,N_1222);
xnor U8219 (N_8219,N_2260,N_1103);
and U8220 (N_8220,N_4883,N_2089);
nor U8221 (N_8221,N_4295,N_4333);
xor U8222 (N_8222,N_5427,N_3114);
or U8223 (N_8223,N_906,N_1602);
and U8224 (N_8224,N_5,N_719);
xor U8225 (N_8225,N_1516,N_3294);
xnor U8226 (N_8226,N_5203,N_6196);
xnor U8227 (N_8227,N_18,N_78);
nor U8228 (N_8228,N_379,N_3880);
and U8229 (N_8229,N_233,N_3728);
and U8230 (N_8230,N_5155,N_5038);
nand U8231 (N_8231,N_1948,N_1870);
xnor U8232 (N_8232,N_3425,N_703);
nor U8233 (N_8233,N_4531,N_2366);
or U8234 (N_8234,N_24,N_2981);
and U8235 (N_8235,N_2852,N_1458);
nand U8236 (N_8236,N_3045,N_1520);
nand U8237 (N_8237,N_6043,N_2848);
or U8238 (N_8238,N_2473,N_5605);
xnor U8239 (N_8239,N_5775,N_1790);
xnor U8240 (N_8240,N_5854,N_877);
nand U8241 (N_8241,N_2115,N_2105);
nand U8242 (N_8242,N_2922,N_5183);
and U8243 (N_8243,N_1563,N_4452);
and U8244 (N_8244,N_2329,N_603);
and U8245 (N_8245,N_580,N_5126);
xnor U8246 (N_8246,N_5346,N_781);
xnor U8247 (N_8247,N_2762,N_4243);
or U8248 (N_8248,N_5283,N_525);
nor U8249 (N_8249,N_5282,N_373);
or U8250 (N_8250,N_2484,N_4799);
nand U8251 (N_8251,N_5314,N_4259);
xor U8252 (N_8252,N_4845,N_2070);
nand U8253 (N_8253,N_701,N_3936);
nor U8254 (N_8254,N_5049,N_3568);
xor U8255 (N_8255,N_3345,N_3171);
or U8256 (N_8256,N_5633,N_5680);
nand U8257 (N_8257,N_2667,N_3773);
nor U8258 (N_8258,N_5867,N_5707);
and U8259 (N_8259,N_4331,N_248);
nor U8260 (N_8260,N_4781,N_996);
xnor U8261 (N_8261,N_1662,N_4195);
xor U8262 (N_8262,N_3265,N_4835);
or U8263 (N_8263,N_5542,N_2589);
xnor U8264 (N_8264,N_2795,N_2147);
or U8265 (N_8265,N_4433,N_421);
nand U8266 (N_8266,N_1172,N_6126);
or U8267 (N_8267,N_3207,N_621);
nor U8268 (N_8268,N_6128,N_1051);
or U8269 (N_8269,N_2198,N_4791);
nor U8270 (N_8270,N_5848,N_1176);
xnor U8271 (N_8271,N_2843,N_1331);
or U8272 (N_8272,N_332,N_5552);
nor U8273 (N_8273,N_2685,N_5275);
or U8274 (N_8274,N_1430,N_3699);
or U8275 (N_8275,N_1066,N_5879);
xor U8276 (N_8276,N_992,N_3768);
nor U8277 (N_8277,N_5986,N_4671);
nor U8278 (N_8278,N_4546,N_2736);
and U8279 (N_8279,N_1150,N_4017);
nor U8280 (N_8280,N_4867,N_3276);
or U8281 (N_8281,N_2845,N_3465);
nand U8282 (N_8282,N_4158,N_3949);
and U8283 (N_8283,N_1446,N_1885);
or U8284 (N_8284,N_2971,N_5345);
or U8285 (N_8285,N_4253,N_5303);
xnor U8286 (N_8286,N_1494,N_2962);
nor U8287 (N_8287,N_4399,N_1180);
xnor U8288 (N_8288,N_1444,N_2346);
and U8289 (N_8289,N_1639,N_4385);
and U8290 (N_8290,N_5784,N_2883);
nand U8291 (N_8291,N_722,N_36);
and U8292 (N_8292,N_5496,N_5785);
and U8293 (N_8293,N_561,N_1177);
or U8294 (N_8294,N_2142,N_2046);
and U8295 (N_8295,N_3624,N_5308);
and U8296 (N_8296,N_1569,N_4489);
nand U8297 (N_8297,N_5850,N_3542);
xnor U8298 (N_8298,N_4557,N_4954);
nand U8299 (N_8299,N_2343,N_2381);
or U8300 (N_8300,N_161,N_2132);
nor U8301 (N_8301,N_5703,N_2678);
nand U8302 (N_8302,N_407,N_5876);
nand U8303 (N_8303,N_92,N_4397);
xor U8304 (N_8304,N_2079,N_1860);
xnor U8305 (N_8305,N_4447,N_1344);
and U8306 (N_8306,N_5378,N_4832);
nand U8307 (N_8307,N_427,N_2485);
nor U8308 (N_8308,N_3030,N_5263);
and U8309 (N_8309,N_1833,N_947);
nand U8310 (N_8310,N_3257,N_1572);
xnor U8311 (N_8311,N_302,N_1);
xnor U8312 (N_8312,N_662,N_5262);
or U8313 (N_8313,N_4804,N_916);
nand U8314 (N_8314,N_4745,N_1746);
xor U8315 (N_8315,N_5859,N_510);
and U8316 (N_8316,N_687,N_97);
xor U8317 (N_8317,N_1481,N_4949);
xnor U8318 (N_8318,N_310,N_1427);
or U8319 (N_8319,N_1878,N_2513);
xnor U8320 (N_8320,N_1518,N_3326);
nand U8321 (N_8321,N_3317,N_2888);
and U8322 (N_8322,N_1525,N_2944);
and U8323 (N_8323,N_3961,N_4347);
nor U8324 (N_8324,N_3444,N_5862);
xnor U8325 (N_8325,N_973,N_629);
nand U8326 (N_8326,N_1540,N_3200);
nor U8327 (N_8327,N_5769,N_2123);
or U8328 (N_8328,N_4108,N_4325);
xor U8329 (N_8329,N_3374,N_4879);
xnor U8330 (N_8330,N_3488,N_5841);
or U8331 (N_8331,N_1610,N_2148);
xnor U8332 (N_8332,N_3367,N_1609);
and U8333 (N_8333,N_3259,N_1283);
or U8334 (N_8334,N_5393,N_1812);
or U8335 (N_8335,N_921,N_2399);
and U8336 (N_8336,N_3476,N_2316);
or U8337 (N_8337,N_1573,N_1032);
nor U8338 (N_8338,N_3559,N_311);
and U8339 (N_8339,N_920,N_4526);
nand U8340 (N_8340,N_2066,N_1181);
or U8341 (N_8341,N_5927,N_3924);
or U8342 (N_8342,N_4919,N_934);
nor U8343 (N_8343,N_3477,N_4589);
nand U8344 (N_8344,N_4039,N_236);
and U8345 (N_8345,N_5657,N_3270);
and U8346 (N_8346,N_1108,N_2840);
or U8347 (N_8347,N_5658,N_1001);
or U8348 (N_8348,N_3783,N_4160);
and U8349 (N_8349,N_5759,N_1476);
nor U8350 (N_8350,N_2558,N_5560);
nor U8351 (N_8351,N_6104,N_191);
nor U8352 (N_8352,N_2564,N_1791);
nor U8353 (N_8353,N_3674,N_3668);
or U8354 (N_8354,N_1044,N_1713);
nor U8355 (N_8355,N_2153,N_2897);
nor U8356 (N_8356,N_5936,N_506);
and U8357 (N_8357,N_692,N_4329);
nor U8358 (N_8358,N_3913,N_1225);
xor U8359 (N_8359,N_5190,N_4975);
or U8360 (N_8360,N_5205,N_5541);
xnor U8361 (N_8361,N_3337,N_1079);
and U8362 (N_8362,N_6189,N_1889);
or U8363 (N_8363,N_1703,N_5783);
or U8364 (N_8364,N_3590,N_5640);
nand U8365 (N_8365,N_2022,N_2959);
nor U8366 (N_8366,N_1666,N_6249);
xor U8367 (N_8367,N_2872,N_6161);
xnor U8368 (N_8368,N_2815,N_2412);
xor U8369 (N_8369,N_1343,N_3297);
nand U8370 (N_8370,N_2889,N_520);
nand U8371 (N_8371,N_5661,N_3446);
and U8372 (N_8372,N_4154,N_2691);
and U8373 (N_8373,N_5388,N_4172);
nor U8374 (N_8374,N_3789,N_6033);
nor U8375 (N_8375,N_3042,N_4445);
nor U8376 (N_8376,N_958,N_4681);
nand U8377 (N_8377,N_5817,N_449);
and U8378 (N_8378,N_4694,N_3370);
or U8379 (N_8379,N_4571,N_4374);
xnor U8380 (N_8380,N_6149,N_2297);
or U8381 (N_8381,N_2570,N_3050);
and U8382 (N_8382,N_649,N_2702);
and U8383 (N_8383,N_3608,N_5865);
nand U8384 (N_8384,N_4935,N_4676);
nor U8385 (N_8385,N_448,N_4878);
nand U8386 (N_8386,N_2968,N_5065);
nand U8387 (N_8387,N_5798,N_3864);
xor U8388 (N_8388,N_5227,N_764);
or U8389 (N_8389,N_354,N_3607);
nor U8390 (N_8390,N_2972,N_4988);
and U8391 (N_8391,N_5323,N_4563);
or U8392 (N_8392,N_6210,N_4437);
nor U8393 (N_8393,N_1689,N_3310);
and U8394 (N_8394,N_2806,N_1531);
xor U8395 (N_8395,N_3136,N_5150);
nor U8396 (N_8396,N_4751,N_6133);
or U8397 (N_8397,N_5325,N_286);
nand U8398 (N_8398,N_5294,N_2467);
and U8399 (N_8399,N_3527,N_2488);
and U8400 (N_8400,N_1985,N_1198);
nand U8401 (N_8401,N_2086,N_1062);
xnor U8402 (N_8402,N_1327,N_442);
xnor U8403 (N_8403,N_665,N_6130);
or U8404 (N_8404,N_4706,N_1731);
nand U8405 (N_8405,N_4997,N_3859);
nand U8406 (N_8406,N_3909,N_5142);
nor U8407 (N_8407,N_974,N_6110);
xor U8408 (N_8408,N_2403,N_3108);
nor U8409 (N_8409,N_3554,N_3509);
nor U8410 (N_8410,N_5449,N_6097);
nor U8411 (N_8411,N_5505,N_2224);
and U8412 (N_8412,N_2024,N_4909);
nand U8413 (N_8413,N_2540,N_3581);
nor U8414 (N_8414,N_241,N_1599);
nor U8415 (N_8415,N_61,N_3634);
nand U8416 (N_8416,N_3281,N_2805);
and U8417 (N_8417,N_3544,N_4465);
xnor U8418 (N_8418,N_1008,N_4189);
nand U8419 (N_8419,N_3571,N_1319);
nand U8420 (N_8420,N_192,N_2574);
xnor U8421 (N_8421,N_4702,N_5888);
or U8422 (N_8422,N_3152,N_5196);
nand U8423 (N_8423,N_5537,N_364);
nand U8424 (N_8424,N_3408,N_615);
nand U8425 (N_8425,N_5242,N_5504);
and U8426 (N_8426,N_2174,N_5477);
nand U8427 (N_8427,N_4674,N_5923);
nand U8428 (N_8428,N_4941,N_1124);
or U8429 (N_8429,N_3016,N_3745);
nor U8430 (N_8430,N_4746,N_4228);
nand U8431 (N_8431,N_1767,N_2054);
nor U8432 (N_8432,N_4000,N_2634);
nand U8433 (N_8433,N_502,N_3702);
or U8434 (N_8434,N_1832,N_4267);
nor U8435 (N_8435,N_1007,N_5800);
nand U8436 (N_8436,N_549,N_2411);
nand U8437 (N_8437,N_6074,N_4583);
xor U8438 (N_8438,N_517,N_3536);
nand U8439 (N_8439,N_4339,N_4779);
and U8440 (N_8440,N_5310,N_5341);
and U8441 (N_8441,N_5253,N_1524);
nand U8442 (N_8442,N_526,N_639);
or U8443 (N_8443,N_2675,N_3088);
or U8444 (N_8444,N_1507,N_5483);
nand U8445 (N_8445,N_5045,N_3043);
and U8446 (N_8446,N_213,N_1582);
and U8447 (N_8447,N_4750,N_2719);
nor U8448 (N_8448,N_3947,N_3290);
nand U8449 (N_8449,N_3008,N_1989);
and U8450 (N_8450,N_4638,N_2592);
and U8451 (N_8451,N_5849,N_5792);
nor U8452 (N_8452,N_3722,N_323);
or U8453 (N_8453,N_6209,N_2859);
xnor U8454 (N_8454,N_4351,N_4744);
xor U8455 (N_8455,N_3621,N_4660);
xor U8456 (N_8456,N_3312,N_439);
nor U8457 (N_8457,N_896,N_557);
or U8458 (N_8458,N_5181,N_5486);
nor U8459 (N_8459,N_2967,N_4586);
nor U8460 (N_8460,N_5371,N_4193);
and U8461 (N_8461,N_9,N_5305);
and U8462 (N_8462,N_2322,N_3541);
xnor U8463 (N_8463,N_4720,N_428);
xor U8464 (N_8464,N_2782,N_148);
or U8465 (N_8465,N_2218,N_5622);
xnor U8466 (N_8466,N_2716,N_4859);
xnor U8467 (N_8467,N_5333,N_3828);
nor U8468 (N_8468,N_4770,N_6136);
and U8469 (N_8469,N_2785,N_797);
nor U8470 (N_8470,N_342,N_2236);
nor U8471 (N_8471,N_458,N_5264);
or U8472 (N_8472,N_1063,N_5995);
nor U8473 (N_8473,N_1022,N_5940);
xnor U8474 (N_8474,N_1414,N_12);
xnor U8475 (N_8475,N_6065,N_2269);
nand U8476 (N_8476,N_739,N_2091);
nor U8477 (N_8477,N_4840,N_5762);
or U8478 (N_8478,N_6086,N_1570);
or U8479 (N_8479,N_397,N_6223);
and U8480 (N_8480,N_2033,N_2276);
or U8481 (N_8481,N_2676,N_5044);
and U8482 (N_8482,N_5471,N_4824);
xnor U8483 (N_8483,N_3979,N_908);
and U8484 (N_8484,N_1690,N_5637);
xor U8485 (N_8485,N_2986,N_5188);
and U8486 (N_8486,N_1106,N_1203);
xnor U8487 (N_8487,N_1288,N_3847);
nand U8488 (N_8488,N_3983,N_3307);
nor U8489 (N_8489,N_1721,N_4089);
and U8490 (N_8490,N_4847,N_632);
nor U8491 (N_8491,N_2262,N_3777);
and U8492 (N_8492,N_3115,N_5149);
nand U8493 (N_8493,N_5224,N_5881);
and U8494 (N_8494,N_1218,N_6129);
and U8495 (N_8495,N_1960,N_4066);
and U8496 (N_8496,N_1632,N_5023);
nand U8497 (N_8497,N_2193,N_90);
nand U8498 (N_8498,N_883,N_5384);
xnor U8499 (N_8499,N_2494,N_1628);
and U8500 (N_8500,N_4294,N_980);
and U8501 (N_8501,N_2052,N_743);
xor U8502 (N_8502,N_4220,N_3691);
and U8503 (N_8503,N_3101,N_1559);
and U8504 (N_8504,N_2463,N_3185);
xor U8505 (N_8505,N_4024,N_3605);
or U8506 (N_8506,N_3829,N_4091);
or U8507 (N_8507,N_1961,N_1242);
nor U8508 (N_8508,N_2595,N_3698);
or U8509 (N_8509,N_618,N_367);
nand U8510 (N_8510,N_5153,N_1396);
xnor U8511 (N_8511,N_4620,N_753);
xor U8512 (N_8512,N_131,N_1890);
or U8513 (N_8513,N_4276,N_3596);
and U8514 (N_8514,N_6053,N_1003);
nor U8515 (N_8515,N_418,N_1372);
and U8516 (N_8516,N_3263,N_1788);
nor U8517 (N_8517,N_2305,N_3754);
xor U8518 (N_8518,N_5962,N_614);
nor U8519 (N_8519,N_3271,N_1015);
nand U8520 (N_8520,N_5776,N_4436);
nor U8521 (N_8521,N_5902,N_5014);
or U8522 (N_8522,N_4626,N_3032);
nand U8523 (N_8523,N_5559,N_948);
nand U8524 (N_8524,N_1655,N_2532);
or U8525 (N_8525,N_5343,N_1086);
xor U8526 (N_8526,N_3229,N_2758);
or U8527 (N_8527,N_6169,N_2510);
and U8528 (N_8528,N_2560,N_210);
nand U8529 (N_8529,N_2587,N_1347);
nor U8530 (N_8530,N_1469,N_3650);
and U8531 (N_8531,N_303,N_1513);
nor U8532 (N_8532,N_5692,N_4424);
nor U8533 (N_8533,N_2459,N_4178);
nand U8534 (N_8534,N_2688,N_5821);
xnor U8535 (N_8535,N_3168,N_3373);
nor U8536 (N_8536,N_4844,N_4984);
xnor U8537 (N_8537,N_5872,N_6106);
xor U8538 (N_8538,N_285,N_5910);
nor U8539 (N_8539,N_268,N_4809);
nor U8540 (N_8540,N_5908,N_3578);
and U8541 (N_8541,N_2122,N_2703);
nand U8542 (N_8542,N_1912,N_5390);
and U8543 (N_8543,N_1699,N_5691);
or U8544 (N_8544,N_475,N_1936);
xnor U8545 (N_8545,N_4432,N_4659);
nand U8546 (N_8546,N_1204,N_6067);
nor U8547 (N_8547,N_1284,N_171);
xnor U8548 (N_8548,N_2601,N_1990);
nand U8549 (N_8549,N_2901,N_1701);
and U8550 (N_8550,N_1090,N_872);
nor U8551 (N_8551,N_4763,N_2261);
nand U8552 (N_8552,N_1260,N_733);
nor U8553 (N_8553,N_151,N_5518);
or U8554 (N_8554,N_4547,N_3400);
nor U8555 (N_8555,N_5838,N_1759);
and U8556 (N_8556,N_2100,N_1939);
xnor U8557 (N_8557,N_5302,N_2619);
or U8558 (N_8558,N_3727,N_2037);
nor U8559 (N_8559,N_5964,N_4862);
nand U8560 (N_8560,N_3330,N_5686);
nor U8561 (N_8561,N_3885,N_541);
xor U8562 (N_8562,N_3794,N_5529);
xor U8563 (N_8563,N_2725,N_562);
and U8564 (N_8564,N_1687,N_5968);
or U8565 (N_8565,N_588,N_4937);
nand U8566 (N_8566,N_4868,N_1208);
nand U8567 (N_8567,N_4672,N_5075);
nand U8568 (N_8568,N_1455,N_1600);
xnor U8569 (N_8569,N_5466,N_2028);
nor U8570 (N_8570,N_5232,N_4428);
or U8571 (N_8571,N_3970,N_4064);
or U8572 (N_8572,N_5410,N_5174);
nand U8573 (N_8573,N_4239,N_2500);
nor U8574 (N_8574,N_5578,N_1445);
or U8575 (N_8575,N_2495,N_2527);
or U8576 (N_8576,N_1847,N_2915);
or U8577 (N_8577,N_2927,N_3680);
xor U8578 (N_8578,N_106,N_4394);
and U8579 (N_8579,N_2659,N_4606);
xnor U8580 (N_8580,N_1182,N_2596);
nor U8581 (N_8581,N_273,N_3343);
xor U8582 (N_8582,N_2238,N_4851);
or U8583 (N_8583,N_3576,N_4021);
or U8584 (N_8584,N_3456,N_1036);
and U8585 (N_8585,N_5130,N_2182);
and U8586 (N_8586,N_1424,N_314);
nand U8587 (N_8587,N_5330,N_5027);
and U8588 (N_8588,N_2605,N_1809);
xor U8589 (N_8589,N_1604,N_14);
nor U8590 (N_8590,N_799,N_914);
or U8591 (N_8591,N_5351,N_869);
nand U8592 (N_8592,N_4426,N_2432);
xor U8593 (N_8593,N_4980,N_306);
nand U8594 (N_8594,N_1729,N_3295);
and U8595 (N_8595,N_766,N_3156);
or U8596 (N_8596,N_1779,N_4605);
or U8597 (N_8597,N_6036,N_2090);
xor U8598 (N_8598,N_750,N_1148);
nand U8599 (N_8599,N_1212,N_1977);
nand U8600 (N_8600,N_4743,N_1924);
or U8601 (N_8601,N_1317,N_5620);
nand U8602 (N_8602,N_2650,N_4350);
or U8603 (N_8603,N_496,N_315);
nor U8604 (N_8604,N_1876,N_2894);
and U8605 (N_8605,N_4560,N_4444);
or U8606 (N_8606,N_1250,N_3396);
xnor U8607 (N_8607,N_4383,N_1853);
or U8608 (N_8608,N_4251,N_1760);
or U8609 (N_8609,N_3760,N_5416);
nor U8610 (N_8610,N_1262,N_169);
or U8611 (N_8611,N_316,N_2156);
xor U8612 (N_8612,N_234,N_5145);
xnor U8613 (N_8613,N_724,N_3678);
nand U8614 (N_8614,N_23,N_5140);
and U8615 (N_8615,N_4320,N_5113);
nor U8616 (N_8616,N_3072,N_5199);
nand U8617 (N_8617,N_4827,N_3074);
nor U8618 (N_8618,N_2757,N_2769);
nand U8619 (N_8619,N_3102,N_1900);
or U8620 (N_8620,N_929,N_3887);
nor U8621 (N_8621,N_2288,N_4319);
and U8622 (N_8622,N_3958,N_3921);
nor U8623 (N_8623,N_6103,N_5022);
xor U8624 (N_8624,N_1556,N_1620);
nor U8625 (N_8625,N_3692,N_2113);
or U8626 (N_8626,N_3365,N_392);
and U8627 (N_8627,N_2377,N_3648);
xnor U8628 (N_8628,N_5398,N_2277);
or U8629 (N_8629,N_1245,N_59);
nand U8630 (N_8630,N_1031,N_928);
nor U8631 (N_8631,N_1094,N_457);
and U8632 (N_8632,N_4684,N_5100);
and U8633 (N_8633,N_4582,N_4496);
xor U8634 (N_8634,N_5273,N_5003);
or U8635 (N_8635,N_534,N_3222);
nor U8636 (N_8636,N_3125,N_4006);
xor U8637 (N_8637,N_4891,N_4440);
and U8638 (N_8638,N_3196,N_5959);
or U8639 (N_8639,N_416,N_5090);
and U8640 (N_8640,N_4964,N_445);
or U8641 (N_8641,N_5976,N_2698);
and U8642 (N_8642,N_5809,N_2371);
and U8643 (N_8643,N_2951,N_5569);
nor U8644 (N_8644,N_6057,N_814);
xnor U8645 (N_8645,N_1571,N_638);
and U8646 (N_8646,N_4588,N_2961);
nor U8647 (N_8647,N_5245,N_806);
or U8648 (N_8648,N_2682,N_5093);
nand U8649 (N_8649,N_3435,N_1154);
and U8650 (N_8650,N_3664,N_4075);
and U8651 (N_8651,N_4625,N_5298);
and U8652 (N_8652,N_4343,N_1449);
nand U8653 (N_8653,N_3690,N_3616);
or U8654 (N_8654,N_3039,N_4001);
nor U8655 (N_8655,N_4112,N_5364);
nand U8656 (N_8656,N_340,N_1638);
xor U8657 (N_8657,N_1493,N_4693);
nand U8658 (N_8658,N_4291,N_5983);
nor U8659 (N_8659,N_1914,N_5833);
nor U8660 (N_8660,N_1922,N_1411);
xor U8661 (N_8661,N_1578,N_5594);
or U8662 (N_8662,N_2145,N_3666);
xnor U8663 (N_8663,N_331,N_2694);
nor U8664 (N_8664,N_2717,N_11);
nand U8665 (N_8665,N_5194,N_2341);
nand U8666 (N_8666,N_129,N_2622);
nand U8667 (N_8667,N_2036,N_211);
nand U8668 (N_8668,N_2890,N_4412);
xor U8669 (N_8669,N_5197,N_1171);
nand U8670 (N_8670,N_1486,N_923);
nor U8671 (N_8671,N_1994,N_1355);
xor U8672 (N_8672,N_319,N_1991);
nor U8673 (N_8673,N_5451,N_2038);
or U8674 (N_8674,N_1915,N_2739);
and U8675 (N_8675,N_465,N_6001);
xor U8676 (N_8676,N_4289,N_3364);
nand U8677 (N_8677,N_1631,N_5823);
and U8678 (N_8678,N_1916,N_5770);
nand U8679 (N_8679,N_3593,N_5182);
nand U8680 (N_8680,N_424,N_3886);
or U8681 (N_8681,N_4756,N_4466);
or U8682 (N_8682,N_5033,N_1728);
nor U8683 (N_8683,N_2356,N_6137);
xor U8684 (N_8684,N_5980,N_6017);
xor U8685 (N_8685,N_3684,N_2150);
xor U8686 (N_8686,N_1098,N_3153);
or U8687 (N_8687,N_3059,N_3744);
or U8688 (N_8688,N_5131,N_6107);
xor U8689 (N_8689,N_3417,N_3700);
or U8690 (N_8690,N_2290,N_1888);
nor U8691 (N_8691,N_3253,N_578);
and U8692 (N_8692,N_4775,N_1412);
and U8693 (N_8693,N_653,N_5368);
xor U8694 (N_8694,N_1940,N_805);
or U8695 (N_8695,N_3149,N_2868);
nand U8696 (N_8696,N_2067,N_5688);
and U8697 (N_8697,N_413,N_4515);
nand U8698 (N_8698,N_3216,N_222);
or U8699 (N_8699,N_2245,N_22);
nand U8700 (N_8700,N_1123,N_2752);
or U8701 (N_8701,N_1045,N_5418);
nand U8702 (N_8702,N_3835,N_2508);
and U8703 (N_8703,N_1228,N_6173);
or U8704 (N_8704,N_226,N_3669);
nor U8705 (N_8705,N_3563,N_2936);
xnor U8706 (N_8706,N_3874,N_2517);
and U8707 (N_8707,N_1782,N_1097);
nor U8708 (N_8708,N_188,N_2318);
and U8709 (N_8709,N_3058,N_1339);
xor U8710 (N_8710,N_2202,N_4211);
and U8711 (N_8711,N_1491,N_6197);
or U8712 (N_8712,N_2947,N_624);
and U8713 (N_8713,N_155,N_5852);
xnor U8714 (N_8714,N_1581,N_2756);
and U8715 (N_8715,N_4035,N_2969);
nor U8716 (N_8716,N_5970,N_6231);
and U8717 (N_8717,N_2380,N_2014);
and U8718 (N_8718,N_1897,N_1220);
or U8719 (N_8719,N_1741,N_1403);
xor U8720 (N_8720,N_3957,N_4872);
and U8721 (N_8721,N_3815,N_3704);
nand U8722 (N_8722,N_103,N_3070);
xor U8723 (N_8723,N_410,N_5873);
or U8724 (N_8724,N_4157,N_321);
or U8725 (N_8725,N_5087,N_5993);
nand U8726 (N_8726,N_1321,N_62);
and U8727 (N_8727,N_1303,N_532);
nor U8728 (N_8728,N_2475,N_71);
xor U8729 (N_8729,N_5526,N_1147);
and U8730 (N_8730,N_2204,N_1387);
xnor U8731 (N_8731,N_6183,N_3589);
and U8732 (N_8732,N_2778,N_4226);
nor U8733 (N_8733,N_3239,N_6060);
xnor U8734 (N_8734,N_2920,N_2018);
nand U8735 (N_8735,N_485,N_1122);
xor U8736 (N_8736,N_3868,N_1336);
nor U8737 (N_8737,N_2284,N_3890);
xnor U8738 (N_8738,N_1219,N_2027);
nor U8739 (N_8739,N_4316,N_3636);
nor U8740 (N_8740,N_3525,N_5589);
and U8741 (N_8741,N_3939,N_6078);
nor U8742 (N_8742,N_5374,N_2950);
nand U8743 (N_8743,N_390,N_690);
or U8744 (N_8744,N_2733,N_6090);
nand U8745 (N_8745,N_2821,N_4579);
xnor U8746 (N_8746,N_1521,N_5067);
nand U8747 (N_8747,N_3807,N_3662);
nand U8748 (N_8748,N_5046,N_2324);
xnor U8749 (N_8749,N_6181,N_135);
and U8750 (N_8750,N_5080,N_4942);
nand U8751 (N_8751,N_2427,N_4290);
and U8752 (N_8752,N_4092,N_3656);
nor U8753 (N_8753,N_2753,N_394);
xor U8754 (N_8754,N_3981,N_4533);
nand U8755 (N_8755,N_5475,N_3146);
xnor U8756 (N_8756,N_3660,N_1553);
or U8757 (N_8757,N_950,N_2711);
nand U8758 (N_8758,N_6226,N_5105);
and U8759 (N_8759,N_4528,N_2865);
nand U8760 (N_8760,N_4083,N_1102);
nor U8761 (N_8761,N_1448,N_6087);
and U8762 (N_8762,N_3129,N_1770);
or U8763 (N_8763,N_5648,N_5360);
and U8764 (N_8764,N_4166,N_2360);
xor U8765 (N_8765,N_2129,N_2690);
nor U8766 (N_8766,N_4553,N_5103);
nor U8767 (N_8767,N_5192,N_2529);
nand U8768 (N_8768,N_1194,N_4256);
xor U8769 (N_8769,N_4495,N_6224);
and U8770 (N_8770,N_3561,N_1648);
xor U8771 (N_8771,N_6163,N_5001);
nor U8772 (N_8772,N_3959,N_6222);
or U8773 (N_8773,N_3785,N_803);
or U8774 (N_8774,N_6021,N_4071);
and U8775 (N_8775,N_5304,N_3013);
nand U8776 (N_8776,N_3225,N_4369);
and U8777 (N_8777,N_816,N_2783);
nor U8778 (N_8778,N_6066,N_5695);
nand U8779 (N_8779,N_1558,N_5030);
or U8780 (N_8780,N_2435,N_2068);
or U8781 (N_8781,N_2902,N_1426);
nand U8782 (N_8782,N_1535,N_901);
or U8783 (N_8783,N_1884,N_2511);
or U8784 (N_8784,N_443,N_3205);
nor U8785 (N_8785,N_1537,N_3934);
nor U8786 (N_8786,N_2637,N_66);
xnor U8787 (N_8787,N_5243,N_5538);
xnor U8788 (N_8788,N_4065,N_2320);
or U8789 (N_8789,N_2732,N_3974);
and U8790 (N_8790,N_5612,N_6206);
xnor U8791 (N_8791,N_4863,N_851);
nor U8792 (N_8792,N_819,N_3778);
xnor U8793 (N_8793,N_5487,N_5855);
and U8794 (N_8794,N_5874,N_5950);
nand U8795 (N_8795,N_4755,N_1118);
xor U8796 (N_8796,N_1608,N_1337);
nor U8797 (N_8797,N_2254,N_2578);
and U8798 (N_8798,N_3904,N_5234);
and U8799 (N_8799,N_2794,N_5882);
and U8800 (N_8800,N_3910,N_720);
nor U8801 (N_8801,N_3810,N_2974);
or U8802 (N_8802,N_4917,N_259);
xnor U8803 (N_8803,N_650,N_3130);
and U8804 (N_8804,N_4688,N_5843);
nor U8805 (N_8805,N_6014,N_3872);
nor U8806 (N_8806,N_6151,N_1852);
nand U8807 (N_8807,N_5438,N_5499);
and U8808 (N_8808,N_4147,N_308);
xor U8809 (N_8809,N_3483,N_4969);
and U8810 (N_8810,N_3750,N_5669);
nand U8811 (N_8811,N_2512,N_6217);
nor U8812 (N_8812,N_39,N_4050);
and U8813 (N_8813,N_1159,N_3764);
or U8814 (N_8814,N_4821,N_1361);
and U8815 (N_8815,N_957,N_2571);
or U8816 (N_8816,N_1868,N_1420);
or U8817 (N_8817,N_1587,N_5806);
or U8818 (N_8818,N_3041,N_2798);
nand U8819 (N_8819,N_3837,N_5958);
and U8820 (N_8820,N_1490,N_3492);
nand U8821 (N_8821,N_482,N_3183);
and U8822 (N_8822,N_4362,N_3438);
nand U8823 (N_8823,N_4074,N_5984);
and U8824 (N_8824,N_711,N_3333);
and U8825 (N_8825,N_3584,N_5860);
xor U8826 (N_8826,N_4282,N_5904);
and U8827 (N_8827,N_1590,N_590);
nand U8828 (N_8828,N_1293,N_3501);
xor U8829 (N_8829,N_365,N_1622);
nor U8830 (N_8830,N_807,N_4);
nor U8831 (N_8831,N_142,N_4961);
and U8832 (N_8832,N_4670,N_5889);
nand U8833 (N_8833,N_1650,N_1983);
nand U8834 (N_8834,N_1434,N_6069);
or U8835 (N_8835,N_3319,N_2246);
or U8836 (N_8836,N_4766,N_602);
and U8837 (N_8837,N_3586,N_3048);
nand U8838 (N_8838,N_1107,N_2087);
xnor U8839 (N_8839,N_645,N_2299);
nor U8840 (N_8840,N_3720,N_3619);
or U8841 (N_8841,N_3366,N_2874);
or U8842 (N_8842,N_1406,N_926);
nor U8843 (N_8843,N_3953,N_4352);
xnor U8844 (N_8844,N_371,N_2465);
or U8845 (N_8845,N_31,N_1048);
or U8846 (N_8846,N_2056,N_2908);
nand U8847 (N_8847,N_1365,N_4217);
nor U8848 (N_8848,N_5106,N_3093);
and U8849 (N_8849,N_3884,N_5324);
xnor U8850 (N_8850,N_4109,N_5741);
or U8851 (N_8851,N_372,N_3932);
nand U8852 (N_8852,N_2875,N_3774);
xor U8853 (N_8853,N_3384,N_2219);
and U8854 (N_8854,N_1511,N_4723);
and U8855 (N_8855,N_4165,N_1830);
nor U8856 (N_8856,N_2350,N_2064);
or U8857 (N_8857,N_5650,N_5317);
or U8858 (N_8858,N_182,N_153);
or U8859 (N_8859,N_5376,N_1266);
or U8860 (N_8860,N_6155,N_4389);
nor U8861 (N_8861,N_5500,N_789);
nand U8862 (N_8862,N_4169,N_5938);
nand U8863 (N_8863,N_5743,N_2225);
nand U8864 (N_8864,N_3842,N_5186);
nor U8865 (N_8865,N_343,N_3531);
or U8866 (N_8866,N_1722,N_5587);
and U8867 (N_8867,N_4116,N_2530);
and U8868 (N_8868,N_2846,N_4248);
or U8869 (N_8869,N_2956,N_3788);
nand U8870 (N_8870,N_272,N_2464);
nand U8871 (N_8871,N_2015,N_1591);
nand U8872 (N_8872,N_4968,N_4807);
nand U8873 (N_8873,N_3579,N_1515);
nand U8874 (N_8874,N_1821,N_2496);
and U8875 (N_8875,N_3246,N_3620);
or U8876 (N_8876,N_5339,N_1675);
or U8877 (N_8877,N_5652,N_4675);
xor U8878 (N_8878,N_2030,N_1898);
and U8879 (N_8879,N_3938,N_836);
nand U8880 (N_8880,N_1637,N_4610);
xor U8881 (N_8881,N_1453,N_3154);
xor U8882 (N_8882,N_622,N_5740);
xor U8883 (N_8883,N_4348,N_1054);
nor U8884 (N_8884,N_4839,N_3996);
xnor U8885 (N_8885,N_3142,N_4908);
and U8886 (N_8886,N_4309,N_900);
and U8887 (N_8887,N_5385,N_4901);
nand U8888 (N_8888,N_4026,N_1276);
nor U8889 (N_8889,N_777,N_3210);
xnor U8890 (N_8890,N_1215,N_2816);
nor U8891 (N_8891,N_5409,N_2095);
xnor U8892 (N_8892,N_3914,N_1816);
or U8893 (N_8893,N_1074,N_3954);
nand U8894 (N_8894,N_3109,N_593);
nand U8895 (N_8895,N_1160,N_2357);
nor U8896 (N_8896,N_2640,N_3905);
xor U8897 (N_8897,N_2050,N_6199);
or U8898 (N_8898,N_5746,N_5365);
nor U8899 (N_8899,N_5375,N_4431);
xor U8900 (N_8900,N_2505,N_295);
and U8901 (N_8901,N_1359,N_6203);
and U8902 (N_8902,N_1329,N_842);
nand U8903 (N_8903,N_4188,N_3630);
or U8904 (N_8904,N_5760,N_2861);
nor U8905 (N_8905,N_1584,N_3558);
and U8906 (N_8906,N_782,N_5536);
or U8907 (N_8907,N_860,N_1963);
and U8908 (N_8908,N_4875,N_4769);
or U8909 (N_8909,N_1692,N_6178);
and U8910 (N_8910,N_4450,N_5198);
xnor U8911 (N_8911,N_863,N_2895);
and U8912 (N_8912,N_3054,N_1475);
nand U8913 (N_8913,N_51,N_4133);
nor U8914 (N_8914,N_2871,N_4162);
xor U8915 (N_8915,N_3964,N_1364);
or U8916 (N_8916,N_1379,N_5795);
nor U8917 (N_8917,N_3189,N_945);
and U8918 (N_8918,N_2563,N_5582);
nor U8919 (N_8919,N_2007,N_4145);
and U8920 (N_8920,N_3956,N_4616);
xor U8921 (N_8921,N_1988,N_1047);
nand U8922 (N_8922,N_2993,N_702);
or U8923 (N_8923,N_313,N_5424);
nand U8924 (N_8924,N_4250,N_1787);
and U8925 (N_8925,N_6101,N_4967);
nor U8926 (N_8926,N_408,N_3511);
nor U8927 (N_8927,N_2221,N_971);
or U8928 (N_8928,N_1196,N_4548);
xnor U8929 (N_8929,N_5899,N_1857);
nand U8930 (N_8930,N_1216,N_2713);
nor U8931 (N_8931,N_3416,N_704);
xor U8932 (N_8932,N_2296,N_4218);
and U8933 (N_8933,N_1400,N_705);
and U8934 (N_8934,N_3825,N_1724);
nor U8935 (N_8935,N_3856,N_5791);
or U8936 (N_8936,N_3706,N_5693);
and U8937 (N_8937,N_3038,N_610);
or U8938 (N_8938,N_1012,N_4924);
or U8939 (N_8939,N_45,N_2759);
nand U8940 (N_8940,N_6139,N_4874);
nand U8941 (N_8941,N_2835,N_4014);
xor U8942 (N_8942,N_3679,N_1209);
xnor U8943 (N_8943,N_6180,N_4164);
xor U8944 (N_8944,N_2954,N_4227);
and U8945 (N_8945,N_1984,N_40);
and U8946 (N_8946,N_4587,N_4033);
nor U8947 (N_8947,N_3176,N_3385);
and U8948 (N_8948,N_199,N_6018);
or U8949 (N_8949,N_2597,N_469);
nor U8950 (N_8950,N_1268,N_2507);
xnor U8951 (N_8951,N_886,N_1101);
or U8952 (N_8952,N_3430,N_399);
nand U8953 (N_8953,N_5237,N_1285);
and U8954 (N_8954,N_3498,N_5269);
nand U8955 (N_8955,N_3426,N_5350);
and U8956 (N_8956,N_305,N_1657);
and U8957 (N_8957,N_6118,N_2430);
or U8958 (N_8958,N_4427,N_4439);
nand U8959 (N_8959,N_3348,N_2137);
xor U8960 (N_8960,N_5808,N_1422);
nand U8961 (N_8961,N_2118,N_2582);
and U8962 (N_8962,N_4455,N_3049);
xor U8963 (N_8963,N_5322,N_3390);
or U8964 (N_8964,N_1932,N_2442);
or U8965 (N_8965,N_1415,N_1751);
nand U8966 (N_8966,N_4922,N_1217);
or U8967 (N_8967,N_2609,N_4110);
and U8968 (N_8968,N_2021,N_5016);
xnor U8969 (N_8969,N_3460,N_5900);
nor U8970 (N_8970,N_3394,N_2493);
and U8971 (N_8971,N_1075,N_3748);
nor U8972 (N_8972,N_5086,N_100);
and U8973 (N_8973,N_1614,N_5353);
or U8974 (N_8974,N_2328,N_3697);
xnor U8975 (N_8975,N_2586,N_4787);
xor U8976 (N_8976,N_1413,N_6167);
xor U8977 (N_8977,N_4810,N_3085);
and U8978 (N_8978,N_1519,N_3191);
nand U8979 (N_8979,N_5546,N_3672);
nand U8980 (N_8980,N_843,N_1928);
nor U8981 (N_8981,N_5229,N_1826);
xor U8982 (N_8982,N_4272,N_4078);
and U8983 (N_8983,N_2502,N_1624);
xor U8984 (N_8984,N_3793,N_1462);
and U8985 (N_8985,N_2720,N_4772);
nor U8986 (N_8986,N_5123,N_1060);
nor U8987 (N_8987,N_2789,N_2085);
and U8988 (N_8988,N_1169,N_2119);
nor U8989 (N_8989,N_405,N_218);
nor U8990 (N_8990,N_2055,N_1694);
xor U8991 (N_8991,N_2749,N_5011);
nand U8992 (N_8992,N_5840,N_1369);
and U8993 (N_8993,N_4792,N_4183);
or U8994 (N_8994,N_6119,N_494);
xnor U8995 (N_8995,N_350,N_4916);
or U8996 (N_8996,N_3412,N_1189);
nand U8997 (N_8997,N_6238,N_984);
and U8998 (N_8998,N_5076,N_1273);
xor U8999 (N_8999,N_727,N_641);
and U9000 (N_9000,N_2386,N_3178);
and U9001 (N_9001,N_5042,N_3451);
nor U9002 (N_9002,N_5091,N_3984);
xor U9003 (N_9003,N_4085,N_6027);
xor U9004 (N_9004,N_4090,N_139);
or U9005 (N_9005,N_5156,N_3710);
nor U9006 (N_9006,N_1332,N_3870);
nor U9007 (N_9007,N_643,N_2714);
nor U9008 (N_9008,N_5355,N_5545);
nor U9009 (N_9009,N_1959,N_1146);
or U9010 (N_9010,N_3230,N_4593);
nand U9011 (N_9011,N_4209,N_6235);
xnor U9012 (N_9012,N_1428,N_3755);
and U9013 (N_9013,N_389,N_72);
nor U9014 (N_9014,N_1717,N_5766);
and U9015 (N_9015,N_4765,N_1095);
xnor U9016 (N_9016,N_1702,N_2141);
and U9017 (N_9017,N_4864,N_4511);
xnor U9018 (N_9018,N_2273,N_2197);
and U9019 (N_9019,N_2774,N_3028);
xnor U9020 (N_9020,N_759,N_5277);
nor U9021 (N_9021,N_5111,N_1804);
nor U9022 (N_9022,N_3351,N_111);
nor U9023 (N_9023,N_5646,N_4173);
xnor U9024 (N_9024,N_2755,N_3252);
nor U9025 (N_9025,N_4378,N_1278);
and U9026 (N_9026,N_1680,N_2535);
or U9027 (N_9027,N_3732,N_567);
nand U9028 (N_9028,N_2699,N_2533);
xnor U9029 (N_9029,N_2387,N_5943);
or U9030 (N_9030,N_5420,N_911);
or U9031 (N_9031,N_2803,N_694);
xor U9032 (N_9032,N_219,N_2480);
nor U9033 (N_9033,N_5909,N_688);
or U9034 (N_9034,N_3165,N_3217);
xnor U9035 (N_9035,N_5159,N_2903);
nor U9036 (N_9036,N_1252,N_98);
xnor U9037 (N_9037,N_2661,N_689);
nor U9038 (N_9038,N_5960,N_3817);
and U9039 (N_9039,N_6099,N_2160);
or U9040 (N_9040,N_2966,N_3266);
xnor U9041 (N_9041,N_5267,N_775);
nand U9042 (N_9042,N_2626,N_3555);
xor U9043 (N_9043,N_3609,N_3900);
nand U9044 (N_9044,N_571,N_2817);
nand U9045 (N_9045,N_6024,N_2482);
nor U9046 (N_9046,N_220,N_563);
nand U9047 (N_9047,N_5210,N_2139);
nor U9048 (N_9048,N_3418,N_5696);
or U9049 (N_9049,N_5801,N_3410);
nand U9050 (N_9050,N_4315,N_870);
nor U9051 (N_9051,N_4143,N_531);
xor U9052 (N_9052,N_5478,N_329);
nand U9053 (N_9053,N_2552,N_3736);
nand U9054 (N_9054,N_4615,N_3484);
nand U9055 (N_9055,N_1993,N_1800);
xor U9056 (N_9056,N_1765,N_3556);
nand U9057 (N_9057,N_6241,N_5110);
xnor U9058 (N_9058,N_3228,N_3851);
and U9059 (N_9059,N_5216,N_3537);
xnor U9060 (N_9060,N_2368,N_4040);
nor U9061 (N_9061,N_2133,N_2282);
and U9062 (N_9062,N_1113,N_4260);
nand U9063 (N_9063,N_4865,N_1275);
nor U9064 (N_9064,N_2796,N_5797);
nand U9065 (N_9065,N_184,N_2186);
or U9066 (N_9066,N_5258,N_2942);
xnor U9067 (N_9067,N_2919,N_1289);
xnor U9068 (N_9068,N_2059,N_2436);
xor U9069 (N_9069,N_4718,N_3960);
or U9070 (N_9070,N_1049,N_5697);
and U9071 (N_9071,N_175,N_1568);
xnor U9072 (N_9072,N_3103,N_1969);
nor U9073 (N_9073,N_5389,N_3846);
nand U9074 (N_9074,N_3064,N_4663);
nor U9075 (N_9075,N_2651,N_1542);
xnor U9076 (N_9076,N_53,N_4936);
xnor U9077 (N_9077,N_1931,N_5777);
and U9078 (N_9078,N_4030,N_3099);
nand U9079 (N_9079,N_435,N_1665);
xor U9080 (N_9080,N_5057,N_4500);
nand U9081 (N_9081,N_1233,N_50);
or U9082 (N_9082,N_1142,N_915);
nand U9083 (N_9083,N_404,N_2347);
and U9084 (N_9084,N_3952,N_6019);
nor U9085 (N_9085,N_4692,N_3339);
xnor U9086 (N_9086,N_1605,N_2081);
and U9087 (N_9087,N_4281,N_3907);
nand U9088 (N_9088,N_3382,N_35);
xnor U9089 (N_9089,N_659,N_2802);
nor U9090 (N_9090,N_3962,N_3506);
xnor U9091 (N_9091,N_463,N_597);
nor U9092 (N_9092,N_5547,N_388);
nor U9093 (N_9093,N_4192,N_1818);
nand U9094 (N_9094,N_3328,N_888);
or U9095 (N_9095,N_1536,N_3314);
and U9096 (N_9096,N_882,N_1371);
and U9097 (N_9097,N_1178,N_3546);
or U9098 (N_9098,N_613,N_5941);
nand U9099 (N_9099,N_5918,N_2175);
nor U9100 (N_9100,N_2099,N_1734);
nand U9101 (N_9101,N_737,N_204);
nand U9102 (N_9102,N_2818,N_2352);
nand U9103 (N_9103,N_5643,N_4446);
nand U9104 (N_9104,N_2824,N_5724);
or U9105 (N_9105,N_172,N_2407);
nor U9106 (N_9106,N_5013,N_2630);
or U9107 (N_9107,N_5796,N_4361);
xor U9108 (N_9108,N_2462,N_1174);
xor U9109 (N_9109,N_318,N_3853);
or U9110 (N_9110,N_3299,N_4283);
and U9111 (N_9111,N_573,N_2975);
and U9112 (N_9112,N_3031,N_2991);
and U9113 (N_9113,N_1341,N_1777);
or U9114 (N_9114,N_3449,N_3550);
or U9115 (N_9115,N_194,N_76);
xnor U9116 (N_9116,N_1911,N_1027);
xor U9117 (N_9117,N_1405,N_5157);
or U9118 (N_9118,N_4190,N_4657);
xor U9119 (N_9119,N_3772,N_3084);
nand U9120 (N_9120,N_678,N_4521);
xor U9121 (N_9121,N_4205,N_5994);
and U9122 (N_9122,N_2233,N_2213);
and U9123 (N_9123,N_3982,N_4346);
nand U9124 (N_9124,N_1937,N_5580);
xnor U9125 (N_9125,N_41,N_2765);
nor U9126 (N_9126,N_3595,N_1081);
nor U9127 (N_9127,N_4356,N_1656);
and U9128 (N_9128,N_3993,N_3725);
nand U9129 (N_9129,N_5568,N_2098);
nand U9130 (N_9130,N_4622,N_4485);
nand U9131 (N_9131,N_4539,N_778);
and U9132 (N_9132,N_507,N_4985);
nand U9133 (N_9133,N_4203,N_84);
xor U9134 (N_9134,N_4042,N_406);
or U9135 (N_9135,N_293,N_5663);
or U9136 (N_9136,N_202,N_3122);
and U9137 (N_9137,N_4953,N_4836);
nor U9138 (N_9138,N_746,N_1577);
or U9139 (N_9139,N_5107,N_436);
xor U9140 (N_9140,N_5588,N_4202);
or U9141 (N_9141,N_4695,N_3399);
or U9142 (N_9142,N_4471,N_6143);
or U9143 (N_9143,N_5429,N_2157);
nand U9144 (N_9144,N_1753,N_5898);
xor U9145 (N_9145,N_4054,N_3834);
and U9146 (N_9146,N_2649,N_4852);
or U9147 (N_9147,N_2034,N_3170);
nor U9148 (N_9148,N_817,N_5670);
xnor U9149 (N_9149,N_1579,N_3685);
nor U9150 (N_9150,N_5639,N_2093);
xor U9151 (N_9151,N_3756,N_386);
xor U9152 (N_9152,N_859,N_5705);
xnor U9153 (N_9153,N_4701,N_1996);
xor U9154 (N_9154,N_3398,N_1234);
or U9155 (N_9155,N_4574,N_3003);
and U9156 (N_9156,N_2498,N_4926);
or U9157 (N_9157,N_4722,N_4525);
xnor U9158 (N_9158,N_3011,N_2112);
nand U9159 (N_9159,N_4778,N_1795);
nor U9160 (N_9160,N_5914,N_304);
or U9161 (N_9161,N_1976,N_4850);
nand U9162 (N_9162,N_4443,N_2315);
and U9163 (N_9163,N_3324,N_5290);
or U9164 (N_9164,N_3741,N_5922);
and U9165 (N_9165,N_4830,N_3288);
and U9166 (N_9166,N_3852,N_1592);
nor U9167 (N_9167,N_3795,N_3522);
nand U9168 (N_9168,N_857,N_1166);
xor U9169 (N_9169,N_4641,N_4067);
nand U9170 (N_9170,N_5018,N_3582);
and U9171 (N_9171,N_680,N_2234);
xor U9172 (N_9172,N_1925,N_2976);
nor U9173 (N_9173,N_577,N_2910);
nand U9174 (N_9174,N_1464,N_1698);
or U9175 (N_9175,N_3510,N_3784);
nand U9176 (N_9176,N_1867,N_3665);
xnor U9177 (N_9177,N_2884,N_718);
xnor U9178 (N_9178,N_3137,N_3738);
nand U9179 (N_9179,N_716,N_1291);
nor U9180 (N_9180,N_4459,N_1394);
nor U9181 (N_9181,N_812,N_5271);
nor U9182 (N_9182,N_518,N_3606);
nor U9183 (N_9183,N_1127,N_1440);
nor U9184 (N_9184,N_3325,N_4180);
nor U9185 (N_9185,N_5676,N_1906);
nor U9186 (N_9186,N_1298,N_6048);
and U9187 (N_9187,N_2999,N_4324);
xor U9188 (N_9188,N_5802,N_3243);
and U9189 (N_9189,N_2726,N_2591);
or U9190 (N_9190,N_6114,N_3799);
nor U9191 (N_9191,N_4379,N_1547);
xor U9192 (N_9192,N_3866,N_2905);
and U9193 (N_9193,N_4899,N_3457);
and U9194 (N_9194,N_349,N_2486);
and U9195 (N_9195,N_4131,N_5951);
nand U9196 (N_9196,N_1265,N_3538);
or U9197 (N_9197,N_6192,N_215);
nand U9198 (N_9198,N_5347,N_5081);
and U9199 (N_9199,N_4199,N_3803);
and U9200 (N_9200,N_5407,N_5400);
xor U9201 (N_9201,N_4497,N_609);
and U9202 (N_9202,N_441,N_5035);
and U9203 (N_9203,N_953,N_4120);
or U9204 (N_9204,N_5624,N_5979);
and U9205 (N_9205,N_5468,N_5274);
nand U9206 (N_9206,N_3919,N_91);
or U9207 (N_9207,N_691,N_2751);
and U9208 (N_9208,N_1808,N_2012);
and U9209 (N_9209,N_3073,N_472);
nand U9210 (N_9210,N_4758,N_4952);
nor U9211 (N_9211,N_838,N_288);
nor U9212 (N_9212,N_2300,N_867);
and U9213 (N_9213,N_846,N_4757);
nand U9214 (N_9214,N_2878,N_2312);
nand U9215 (N_9215,N_1235,N_3223);
and U9216 (N_9216,N_1350,N_4892);
or U9217 (N_9217,N_5218,N_826);
nor U9218 (N_9218,N_3758,N_5037);
nor U9219 (N_9219,N_33,N_2466);
nor U9220 (N_9220,N_2680,N_133);
nor U9221 (N_9221,N_5782,N_154);
nor U9222 (N_9222,N_5767,N_4568);
nand U9223 (N_9223,N_1819,N_1484);
nand U9224 (N_9224,N_3729,N_2735);
xor U9225 (N_9225,N_423,N_2519);
nor U9226 (N_9226,N_3284,N_4609);
and U9227 (N_9227,N_1272,N_707);
nor U9228 (N_9228,N_956,N_3891);
and U9229 (N_9229,N_477,N_2040);
or U9230 (N_9230,N_5532,N_2827);
or U9231 (N_9231,N_1433,N_5877);
and U9232 (N_9232,N_2588,N_4703);
nor U9233 (N_9233,N_1992,N_5058);
and U9234 (N_9234,N_4677,N_3346);
or U9235 (N_9235,N_4728,N_4498);
and U9236 (N_9236,N_5969,N_5144);
and U9237 (N_9237,N_2228,N_3826);
or U9238 (N_9238,N_5021,N_456);
or U9239 (N_9239,N_4349,N_2985);
xnor U9240 (N_9240,N_3022,N_4898);
or U9241 (N_9241,N_2980,N_2390);
and U9242 (N_9242,N_1226,N_287);
nor U9243 (N_9243,N_938,N_1323);
or U9244 (N_9244,N_2321,N_5928);
xor U9245 (N_9245,N_6141,N_5193);
or U9246 (N_9246,N_1802,N_1954);
xor U9247 (N_9247,N_4115,N_1281);
or U9248 (N_9248,N_1682,N_1745);
or U9249 (N_9249,N_267,N_292);
nor U9250 (N_9250,N_4848,N_1617);
or U9251 (N_9251,N_4970,N_1089);
or U9252 (N_9252,N_5257,N_262);
nand U9253 (N_9253,N_5222,N_5452);
or U9254 (N_9254,N_105,N_4513);
and U9255 (N_9255,N_4885,N_5031);
nand U9256 (N_9256,N_4788,N_4567);
nor U9257 (N_9257,N_4805,N_3020);
nand U9258 (N_9258,N_2534,N_4895);
nor U9259 (N_9259,N_1550,N_3344);
xor U9260 (N_9260,N_3406,N_1186);
and U9261 (N_9261,N_5493,N_4669);
nand U9262 (N_9262,N_656,N_2809);
or U9263 (N_9263,N_6117,N_5906);
nor U9264 (N_9264,N_2382,N_5433);
xnor U9265 (N_9265,N_6035,N_4617);
nand U9266 (N_9266,N_3338,N_4314);
nor U9267 (N_9267,N_3148,N_4555);
and U9268 (N_9268,N_4422,N_3302);
and U9269 (N_9269,N_4639,N_5300);
and U9270 (N_9270,N_3091,N_4060);
xnor U9271 (N_9271,N_6016,N_2212);
or U9272 (N_9272,N_244,N_6080);
or U9273 (N_9273,N_4150,N_2949);
nor U9274 (N_9274,N_3151,N_1714);
and U9275 (N_9275,N_1640,N_2536);
xnor U9276 (N_9276,N_296,N_1715);
xor U9277 (N_9277,N_5584,N_848);
nor U9278 (N_9278,N_1735,N_2217);
and U9279 (N_9279,N_1374,N_5137);
nor U9280 (N_9280,N_961,N_521);
and U9281 (N_9281,N_3340,N_3948);
and U9282 (N_9282,N_2101,N_976);
or U9283 (N_9283,N_1358,N_5369);
xor U9284 (N_9284,N_6229,N_4945);
xnor U9285 (N_9285,N_432,N_1528);
and U9286 (N_9286,N_110,N_3090);
nor U9287 (N_9287,N_1064,N_903);
nor U9288 (N_9288,N_2483,N_2873);
xor U9289 (N_9289,N_550,N_5893);
nand U9290 (N_9290,N_5337,N_2598);
xnor U9291 (N_9291,N_5756,N_3833);
or U9292 (N_9292,N_3631,N_1794);
nor U9293 (N_9293,N_1981,N_2990);
and U9294 (N_9294,N_4072,N_1247);
nor U9295 (N_9295,N_1299,N_5834);
xor U9296 (N_9296,N_5896,N_450);
and U9297 (N_9297,N_5628,N_3985);
and U9298 (N_9298,N_858,N_5421);
nand U9299 (N_9299,N_2171,N_1647);
or U9300 (N_9300,N_3649,N_4858);
xnor U9301 (N_9301,N_2239,N_4384);
or U9302 (N_9302,N_758,N_4613);
or U9303 (N_9303,N_3613,N_1739);
nor U9304 (N_9304,N_4680,N_3916);
nor U9305 (N_9305,N_5871,N_2434);
or U9306 (N_9306,N_1037,N_5880);
xnor U9307 (N_9307,N_4987,N_5482);
nor U9308 (N_9308,N_29,N_6116);
xor U9309 (N_9309,N_3933,N_1748);
or U9310 (N_9310,N_1076,N_2926);
xnor U9311 (N_9311,N_1451,N_821);
nor U9312 (N_9312,N_628,N_2964);
xor U9313 (N_9313,N_5601,N_1546);
nand U9314 (N_9314,N_2201,N_3224);
nor U9315 (N_9315,N_3651,N_2303);
nor U9316 (N_9316,N_3611,N_6135);
or U9317 (N_9317,N_1441,N_784);
and U9318 (N_9318,N_60,N_3564);
xor U9319 (N_9319,N_5101,N_3047);
or U9320 (N_9320,N_885,N_4268);
xnor U9321 (N_9321,N_5094,N_3198);
or U9322 (N_9322,N_3876,N_1784);
nor U9323 (N_9323,N_4900,N_2163);
nand U9324 (N_9324,N_5632,N_5702);
and U9325 (N_9325,N_1848,N_2325);
or U9326 (N_9326,N_2913,N_5213);
nand U9327 (N_9327,N_2109,N_3455);
nand U9328 (N_9328,N_1686,N_1325);
and U9329 (N_9329,N_5788,N_3053);
and U9330 (N_9330,N_257,N_5991);
nor U9331 (N_9331,N_1190,N_2546);
nor U9332 (N_9332,N_146,N_6146);
or U9333 (N_9333,N_1254,N_2340);
nand U9334 (N_9334,N_6100,N_2458);
xor U9335 (N_9335,N_5932,N_2298);
nand U9336 (N_9336,N_1967,N_2549);
nor U9337 (N_9337,N_353,N_1875);
nand U9338 (N_9338,N_4036,N_5078);
xor U9339 (N_9339,N_761,N_2945);
or U9340 (N_9340,N_535,N_1292);
nand U9341 (N_9341,N_1020,N_2812);
nor U9342 (N_9342,N_251,N_4070);
and U9343 (N_9343,N_3969,N_3503);
or U9344 (N_9344,N_4789,N_3407);
and U9345 (N_9345,N_3121,N_5162);
and U9346 (N_9346,N_4184,N_119);
nor U9347 (N_9347,N_2397,N_1229);
and U9348 (N_9348,N_1436,N_558);
or U9349 (N_9349,N_94,N_4812);
nor U9350 (N_9350,N_4632,N_1772);
nand U9351 (N_9351,N_4105,N_2781);
nor U9352 (N_9352,N_1389,N_1023);
xor U9353 (N_9353,N_5151,N_4032);
and U9354 (N_9354,N_5211,N_96);
or U9355 (N_9355,N_2804,N_5548);
nand U9356 (N_9356,N_734,N_3260);
nor U9357 (N_9357,N_4860,N_5572);
nor U9358 (N_9358,N_2226,N_1831);
xor U9359 (N_9359,N_4148,N_2641);
xor U9360 (N_9360,N_1774,N_2107);
nand U9361 (N_9361,N_4181,N_5725);
xnor U9362 (N_9362,N_5512,N_3275);
or U9363 (N_9363,N_2330,N_5522);
or U9364 (N_9364,N_491,N_892);
nor U9365 (N_9365,N_4717,N_4191);
nor U9366 (N_9366,N_70,N_4338);
xnor U9367 (N_9367,N_3688,N_1979);
or U9368 (N_9368,N_4709,N_4866);
and U9369 (N_9369,N_1551,N_1013);
xor U9370 (N_9370,N_166,N_626);
xnor U9371 (N_9371,N_4753,N_4304);
xor U9372 (N_9372,N_538,N_5673);
xnor U9373 (N_9373,N_829,N_4566);
xnor U9374 (N_9374,N_3499,N_4233);
nor U9375 (N_9375,N_1556,N_612);
nor U9376 (N_9376,N_1834,N_2674);
nand U9377 (N_9377,N_739,N_2360);
and U9378 (N_9378,N_1115,N_3790);
xnor U9379 (N_9379,N_4087,N_5659);
nor U9380 (N_9380,N_1308,N_1963);
or U9381 (N_9381,N_2075,N_67);
or U9382 (N_9382,N_4814,N_6021);
or U9383 (N_9383,N_2924,N_4932);
or U9384 (N_9384,N_4571,N_6060);
and U9385 (N_9385,N_1703,N_3369);
or U9386 (N_9386,N_3842,N_2335);
or U9387 (N_9387,N_467,N_2829);
or U9388 (N_9388,N_1589,N_5730);
xnor U9389 (N_9389,N_1425,N_2612);
nand U9390 (N_9390,N_2596,N_1097);
nor U9391 (N_9391,N_5421,N_5541);
nor U9392 (N_9392,N_4476,N_2352);
nor U9393 (N_9393,N_3884,N_4945);
or U9394 (N_9394,N_3209,N_213);
and U9395 (N_9395,N_4002,N_5694);
nand U9396 (N_9396,N_5780,N_5350);
xor U9397 (N_9397,N_720,N_275);
nor U9398 (N_9398,N_2863,N_2305);
or U9399 (N_9399,N_4912,N_5258);
xor U9400 (N_9400,N_5715,N_6008);
and U9401 (N_9401,N_3962,N_728);
or U9402 (N_9402,N_3258,N_3924);
and U9403 (N_9403,N_4889,N_2242);
nand U9404 (N_9404,N_3188,N_1080);
nor U9405 (N_9405,N_1764,N_336);
nor U9406 (N_9406,N_4147,N_2108);
nor U9407 (N_9407,N_4338,N_2562);
xor U9408 (N_9408,N_1100,N_716);
or U9409 (N_9409,N_1978,N_2588);
xnor U9410 (N_9410,N_3418,N_225);
and U9411 (N_9411,N_5808,N_4216);
nor U9412 (N_9412,N_2498,N_4601);
nand U9413 (N_9413,N_1396,N_5205);
and U9414 (N_9414,N_2067,N_2062);
nand U9415 (N_9415,N_374,N_1877);
nor U9416 (N_9416,N_6204,N_5877);
nor U9417 (N_9417,N_3753,N_966);
xnor U9418 (N_9418,N_3203,N_2131);
nor U9419 (N_9419,N_5618,N_4617);
xnor U9420 (N_9420,N_3678,N_5021);
nand U9421 (N_9421,N_4310,N_4789);
nand U9422 (N_9422,N_2834,N_6142);
or U9423 (N_9423,N_439,N_3700);
nand U9424 (N_9424,N_2414,N_4403);
nand U9425 (N_9425,N_5722,N_1028);
or U9426 (N_9426,N_4018,N_2197);
nor U9427 (N_9427,N_2734,N_3004);
nor U9428 (N_9428,N_3094,N_1251);
or U9429 (N_9429,N_1775,N_1763);
nand U9430 (N_9430,N_4409,N_1472);
nand U9431 (N_9431,N_801,N_3163);
nand U9432 (N_9432,N_2212,N_5870);
nand U9433 (N_9433,N_4915,N_4258);
nand U9434 (N_9434,N_1297,N_251);
and U9435 (N_9435,N_3426,N_495);
xor U9436 (N_9436,N_5874,N_3744);
nor U9437 (N_9437,N_2150,N_3625);
or U9438 (N_9438,N_2707,N_3990);
and U9439 (N_9439,N_374,N_264);
nand U9440 (N_9440,N_4024,N_3682);
xnor U9441 (N_9441,N_1922,N_3774);
nand U9442 (N_9442,N_197,N_3958);
and U9443 (N_9443,N_2878,N_5621);
xnor U9444 (N_9444,N_3721,N_6145);
xnor U9445 (N_9445,N_4433,N_880);
nor U9446 (N_9446,N_2968,N_3761);
nor U9447 (N_9447,N_3632,N_5141);
and U9448 (N_9448,N_3091,N_2441);
and U9449 (N_9449,N_1219,N_168);
or U9450 (N_9450,N_1955,N_5053);
and U9451 (N_9451,N_3938,N_2911);
or U9452 (N_9452,N_1492,N_3932);
nor U9453 (N_9453,N_657,N_4091);
xnor U9454 (N_9454,N_420,N_4148);
xnor U9455 (N_9455,N_5392,N_5767);
nand U9456 (N_9456,N_2040,N_5344);
nor U9457 (N_9457,N_91,N_4881);
nand U9458 (N_9458,N_1367,N_2452);
nand U9459 (N_9459,N_3191,N_4925);
nand U9460 (N_9460,N_2672,N_3893);
or U9461 (N_9461,N_2421,N_5358);
nand U9462 (N_9462,N_2802,N_692);
nor U9463 (N_9463,N_5414,N_3737);
xor U9464 (N_9464,N_2268,N_5797);
nor U9465 (N_9465,N_4151,N_2831);
nor U9466 (N_9466,N_4292,N_2067);
or U9467 (N_9467,N_3028,N_5063);
xor U9468 (N_9468,N_6168,N_4169);
or U9469 (N_9469,N_2069,N_4904);
or U9470 (N_9470,N_5038,N_2080);
nand U9471 (N_9471,N_3246,N_4072);
nand U9472 (N_9472,N_2194,N_4458);
nand U9473 (N_9473,N_4775,N_5572);
nor U9474 (N_9474,N_4994,N_4387);
xor U9475 (N_9475,N_1509,N_2657);
xnor U9476 (N_9476,N_1674,N_4479);
or U9477 (N_9477,N_3424,N_2803);
nor U9478 (N_9478,N_2146,N_349);
xor U9479 (N_9479,N_1191,N_5036);
or U9480 (N_9480,N_6179,N_893);
or U9481 (N_9481,N_3539,N_6146);
nor U9482 (N_9482,N_3254,N_3199);
nor U9483 (N_9483,N_5977,N_4753);
and U9484 (N_9484,N_1001,N_6116);
or U9485 (N_9485,N_5247,N_4094);
xor U9486 (N_9486,N_4174,N_1894);
and U9487 (N_9487,N_4021,N_6111);
and U9488 (N_9488,N_4414,N_4977);
xor U9489 (N_9489,N_6172,N_2681);
nor U9490 (N_9490,N_3021,N_3583);
or U9491 (N_9491,N_1834,N_3607);
nor U9492 (N_9492,N_5234,N_2381);
nor U9493 (N_9493,N_1489,N_3958);
nor U9494 (N_9494,N_494,N_1961);
nor U9495 (N_9495,N_3669,N_3941);
xor U9496 (N_9496,N_4033,N_4241);
or U9497 (N_9497,N_1218,N_446);
and U9498 (N_9498,N_4800,N_2124);
or U9499 (N_9499,N_5660,N_6119);
nand U9500 (N_9500,N_1390,N_4519);
or U9501 (N_9501,N_2743,N_912);
nand U9502 (N_9502,N_4505,N_4024);
nand U9503 (N_9503,N_1304,N_5779);
or U9504 (N_9504,N_5846,N_540);
nor U9505 (N_9505,N_3175,N_4399);
nor U9506 (N_9506,N_5311,N_189);
nand U9507 (N_9507,N_964,N_1202);
nand U9508 (N_9508,N_5223,N_4765);
nor U9509 (N_9509,N_1839,N_2382);
and U9510 (N_9510,N_4448,N_20);
or U9511 (N_9511,N_1978,N_2203);
or U9512 (N_9512,N_3053,N_1219);
nand U9513 (N_9513,N_3942,N_2280);
nor U9514 (N_9514,N_5304,N_5412);
nor U9515 (N_9515,N_4732,N_1012);
nor U9516 (N_9516,N_3088,N_5427);
or U9517 (N_9517,N_3808,N_749);
nor U9518 (N_9518,N_4071,N_1533);
and U9519 (N_9519,N_344,N_969);
nor U9520 (N_9520,N_1090,N_596);
nand U9521 (N_9521,N_4693,N_5226);
or U9522 (N_9522,N_5204,N_121);
or U9523 (N_9523,N_889,N_4502);
and U9524 (N_9524,N_3159,N_1036);
nor U9525 (N_9525,N_811,N_3260);
nor U9526 (N_9526,N_1811,N_2264);
nand U9527 (N_9527,N_1127,N_4881);
nand U9528 (N_9528,N_4117,N_4407);
nor U9529 (N_9529,N_5341,N_2728);
and U9530 (N_9530,N_6093,N_5037);
nor U9531 (N_9531,N_4037,N_6144);
and U9532 (N_9532,N_5300,N_2111);
nor U9533 (N_9533,N_3234,N_4977);
nand U9534 (N_9534,N_135,N_2078);
nand U9535 (N_9535,N_2796,N_3670);
nand U9536 (N_9536,N_3186,N_2676);
nor U9537 (N_9537,N_1264,N_2130);
and U9538 (N_9538,N_2411,N_4940);
xnor U9539 (N_9539,N_2932,N_246);
or U9540 (N_9540,N_5131,N_5616);
nand U9541 (N_9541,N_1122,N_540);
xnor U9542 (N_9542,N_3201,N_361);
nand U9543 (N_9543,N_6166,N_221);
nor U9544 (N_9544,N_4887,N_3288);
nand U9545 (N_9545,N_3138,N_5470);
or U9546 (N_9546,N_4644,N_2991);
and U9547 (N_9547,N_2738,N_5852);
nand U9548 (N_9548,N_1714,N_1835);
and U9549 (N_9549,N_211,N_3856);
and U9550 (N_9550,N_3427,N_3596);
or U9551 (N_9551,N_834,N_4829);
or U9552 (N_9552,N_864,N_3334);
xnor U9553 (N_9553,N_6121,N_4351);
nor U9554 (N_9554,N_5742,N_5921);
nor U9555 (N_9555,N_6009,N_2240);
nor U9556 (N_9556,N_5815,N_1560);
xnor U9557 (N_9557,N_1227,N_3151);
xnor U9558 (N_9558,N_5279,N_6233);
and U9559 (N_9559,N_1089,N_522);
and U9560 (N_9560,N_4410,N_1634);
or U9561 (N_9561,N_3962,N_1760);
nand U9562 (N_9562,N_5268,N_5117);
or U9563 (N_9563,N_4564,N_5133);
and U9564 (N_9564,N_5173,N_2324);
nand U9565 (N_9565,N_4209,N_2606);
and U9566 (N_9566,N_3158,N_65);
nor U9567 (N_9567,N_3373,N_2093);
xnor U9568 (N_9568,N_5624,N_2693);
nor U9569 (N_9569,N_5561,N_1823);
or U9570 (N_9570,N_4824,N_4987);
xnor U9571 (N_9571,N_3544,N_3887);
or U9572 (N_9572,N_1246,N_4125);
nor U9573 (N_9573,N_1047,N_1607);
and U9574 (N_9574,N_3555,N_2652);
or U9575 (N_9575,N_5314,N_2532);
nand U9576 (N_9576,N_5789,N_611);
nor U9577 (N_9577,N_3272,N_3130);
or U9578 (N_9578,N_656,N_4050);
or U9579 (N_9579,N_3531,N_2340);
or U9580 (N_9580,N_6174,N_4120);
and U9581 (N_9581,N_2261,N_2808);
or U9582 (N_9582,N_3238,N_862);
or U9583 (N_9583,N_5311,N_4579);
and U9584 (N_9584,N_276,N_4282);
nor U9585 (N_9585,N_870,N_4321);
and U9586 (N_9586,N_4887,N_3901);
or U9587 (N_9587,N_5249,N_1962);
nor U9588 (N_9588,N_2429,N_4513);
nand U9589 (N_9589,N_3397,N_2957);
nand U9590 (N_9590,N_327,N_5667);
nand U9591 (N_9591,N_4223,N_2651);
nor U9592 (N_9592,N_1991,N_2096);
xnor U9593 (N_9593,N_41,N_4657);
and U9594 (N_9594,N_1752,N_809);
or U9595 (N_9595,N_1246,N_2883);
nor U9596 (N_9596,N_4395,N_3376);
and U9597 (N_9597,N_3401,N_5773);
nor U9598 (N_9598,N_2100,N_463);
and U9599 (N_9599,N_5684,N_1095);
nor U9600 (N_9600,N_2436,N_2983);
nand U9601 (N_9601,N_697,N_5314);
nor U9602 (N_9602,N_4931,N_3992);
or U9603 (N_9603,N_781,N_1510);
and U9604 (N_9604,N_3512,N_2610);
nand U9605 (N_9605,N_2337,N_6119);
xnor U9606 (N_9606,N_201,N_6071);
or U9607 (N_9607,N_2215,N_6184);
nand U9608 (N_9608,N_5595,N_5139);
nand U9609 (N_9609,N_1898,N_1593);
nor U9610 (N_9610,N_5147,N_1423);
or U9611 (N_9611,N_3971,N_979);
nor U9612 (N_9612,N_1915,N_2059);
nand U9613 (N_9613,N_4371,N_5416);
xnor U9614 (N_9614,N_2520,N_3834);
or U9615 (N_9615,N_3003,N_540);
nand U9616 (N_9616,N_5094,N_5520);
xor U9617 (N_9617,N_2567,N_4214);
nor U9618 (N_9618,N_1314,N_417);
xnor U9619 (N_9619,N_5397,N_3755);
and U9620 (N_9620,N_5379,N_2414);
or U9621 (N_9621,N_3265,N_1434);
and U9622 (N_9622,N_2178,N_3020);
or U9623 (N_9623,N_2317,N_2526);
or U9624 (N_9624,N_4259,N_909);
or U9625 (N_9625,N_5598,N_5953);
or U9626 (N_9626,N_4008,N_384);
nand U9627 (N_9627,N_6124,N_304);
nand U9628 (N_9628,N_274,N_3845);
xor U9629 (N_9629,N_3849,N_4650);
and U9630 (N_9630,N_5965,N_2069);
or U9631 (N_9631,N_562,N_2077);
and U9632 (N_9632,N_5795,N_5530);
nor U9633 (N_9633,N_3651,N_5595);
nand U9634 (N_9634,N_2757,N_91);
xnor U9635 (N_9635,N_2000,N_5987);
and U9636 (N_9636,N_2801,N_3303);
xnor U9637 (N_9637,N_2832,N_3745);
xor U9638 (N_9638,N_1814,N_2465);
nand U9639 (N_9639,N_5172,N_4751);
and U9640 (N_9640,N_5254,N_2952);
nand U9641 (N_9641,N_1133,N_865);
xor U9642 (N_9642,N_375,N_4706);
and U9643 (N_9643,N_1622,N_6193);
nor U9644 (N_9644,N_875,N_5381);
nor U9645 (N_9645,N_5267,N_3908);
nand U9646 (N_9646,N_6232,N_4939);
xor U9647 (N_9647,N_4110,N_5492);
nor U9648 (N_9648,N_317,N_1509);
nand U9649 (N_9649,N_2543,N_5040);
xor U9650 (N_9650,N_4765,N_4784);
and U9651 (N_9651,N_5559,N_4041);
or U9652 (N_9652,N_4489,N_1198);
and U9653 (N_9653,N_5395,N_1373);
nand U9654 (N_9654,N_3772,N_2416);
or U9655 (N_9655,N_498,N_4102);
and U9656 (N_9656,N_5216,N_1666);
or U9657 (N_9657,N_369,N_4263);
nor U9658 (N_9658,N_2334,N_4408);
nand U9659 (N_9659,N_854,N_3221);
xnor U9660 (N_9660,N_531,N_1820);
xnor U9661 (N_9661,N_4559,N_2531);
xor U9662 (N_9662,N_6200,N_583);
or U9663 (N_9663,N_951,N_3952);
xor U9664 (N_9664,N_2950,N_3993);
xnor U9665 (N_9665,N_4845,N_5654);
or U9666 (N_9666,N_4771,N_1655);
xnor U9667 (N_9667,N_3639,N_3321);
xor U9668 (N_9668,N_4726,N_3865);
xor U9669 (N_9669,N_4420,N_4320);
xor U9670 (N_9670,N_2367,N_4481);
nor U9671 (N_9671,N_1811,N_710);
nor U9672 (N_9672,N_5861,N_6113);
or U9673 (N_9673,N_2258,N_3270);
and U9674 (N_9674,N_5163,N_2003);
or U9675 (N_9675,N_2122,N_3861);
xnor U9676 (N_9676,N_5092,N_3791);
nand U9677 (N_9677,N_823,N_4215);
nand U9678 (N_9678,N_4749,N_5366);
nand U9679 (N_9679,N_945,N_6023);
nand U9680 (N_9680,N_5273,N_2192);
nor U9681 (N_9681,N_5698,N_3767);
and U9682 (N_9682,N_3839,N_1604);
or U9683 (N_9683,N_4559,N_5379);
nor U9684 (N_9684,N_2239,N_5049);
or U9685 (N_9685,N_1106,N_4545);
and U9686 (N_9686,N_4934,N_3358);
and U9687 (N_9687,N_3849,N_6010);
nand U9688 (N_9688,N_5375,N_4591);
or U9689 (N_9689,N_1823,N_3931);
xor U9690 (N_9690,N_2010,N_626);
nand U9691 (N_9691,N_5921,N_3424);
nor U9692 (N_9692,N_5752,N_2484);
nand U9693 (N_9693,N_5498,N_5257);
and U9694 (N_9694,N_1294,N_3345);
nor U9695 (N_9695,N_5576,N_5245);
xnor U9696 (N_9696,N_5380,N_4501);
nor U9697 (N_9697,N_2709,N_3082);
nand U9698 (N_9698,N_4464,N_1808);
xnor U9699 (N_9699,N_1091,N_4311);
and U9700 (N_9700,N_5388,N_402);
xnor U9701 (N_9701,N_1786,N_3233);
nand U9702 (N_9702,N_1536,N_2228);
nor U9703 (N_9703,N_1152,N_1091);
or U9704 (N_9704,N_1272,N_1015);
xnor U9705 (N_9705,N_4319,N_4655);
nor U9706 (N_9706,N_28,N_3947);
nor U9707 (N_9707,N_1817,N_3279);
xor U9708 (N_9708,N_3181,N_6170);
xnor U9709 (N_9709,N_4493,N_729);
nand U9710 (N_9710,N_398,N_4369);
or U9711 (N_9711,N_1879,N_3106);
xor U9712 (N_9712,N_259,N_932);
or U9713 (N_9713,N_3681,N_2438);
or U9714 (N_9714,N_2913,N_1453);
nand U9715 (N_9715,N_3849,N_2697);
nor U9716 (N_9716,N_2818,N_2315);
or U9717 (N_9717,N_4991,N_4480);
xnor U9718 (N_9718,N_97,N_5394);
and U9719 (N_9719,N_2793,N_4712);
and U9720 (N_9720,N_4341,N_2869);
and U9721 (N_9721,N_2846,N_4545);
xnor U9722 (N_9722,N_4705,N_2733);
nand U9723 (N_9723,N_84,N_5646);
or U9724 (N_9724,N_2529,N_865);
xor U9725 (N_9725,N_6210,N_5194);
and U9726 (N_9726,N_1920,N_509);
nand U9727 (N_9727,N_2356,N_5133);
and U9728 (N_9728,N_1494,N_4532);
nor U9729 (N_9729,N_205,N_1052);
nand U9730 (N_9730,N_391,N_3355);
xnor U9731 (N_9731,N_2902,N_900);
nor U9732 (N_9732,N_5828,N_2913);
or U9733 (N_9733,N_1746,N_413);
xor U9734 (N_9734,N_5796,N_1347);
and U9735 (N_9735,N_3917,N_5310);
or U9736 (N_9736,N_6174,N_3891);
and U9737 (N_9737,N_3535,N_2366);
or U9738 (N_9738,N_2224,N_2426);
and U9739 (N_9739,N_4746,N_5304);
nand U9740 (N_9740,N_2357,N_5909);
nand U9741 (N_9741,N_5852,N_3324);
xnor U9742 (N_9742,N_1766,N_4010);
xor U9743 (N_9743,N_2890,N_2329);
nor U9744 (N_9744,N_526,N_3584);
nor U9745 (N_9745,N_4271,N_5234);
xnor U9746 (N_9746,N_879,N_3567);
xnor U9747 (N_9747,N_705,N_4601);
and U9748 (N_9748,N_1511,N_1077);
and U9749 (N_9749,N_1293,N_4428);
nor U9750 (N_9750,N_1550,N_5040);
xor U9751 (N_9751,N_5270,N_3852);
or U9752 (N_9752,N_3204,N_847);
or U9753 (N_9753,N_3702,N_1880);
nor U9754 (N_9754,N_2877,N_1171);
nor U9755 (N_9755,N_2711,N_933);
xor U9756 (N_9756,N_4678,N_2642);
and U9757 (N_9757,N_3556,N_4023);
nand U9758 (N_9758,N_1629,N_2551);
or U9759 (N_9759,N_5695,N_252);
or U9760 (N_9760,N_1151,N_1481);
nor U9761 (N_9761,N_2147,N_4231);
nand U9762 (N_9762,N_4300,N_756);
and U9763 (N_9763,N_3542,N_5044);
xor U9764 (N_9764,N_4865,N_4409);
xnor U9765 (N_9765,N_3526,N_2504);
nand U9766 (N_9766,N_4222,N_1782);
and U9767 (N_9767,N_2214,N_1129);
xnor U9768 (N_9768,N_5584,N_482);
nor U9769 (N_9769,N_4696,N_3246);
xnor U9770 (N_9770,N_3323,N_5786);
nor U9771 (N_9771,N_847,N_1603);
nor U9772 (N_9772,N_2610,N_6097);
nor U9773 (N_9773,N_1013,N_6055);
and U9774 (N_9774,N_4110,N_4461);
or U9775 (N_9775,N_981,N_1851);
xor U9776 (N_9776,N_1326,N_5923);
or U9777 (N_9777,N_2223,N_1701);
or U9778 (N_9778,N_2691,N_4731);
nand U9779 (N_9779,N_3320,N_2414);
nor U9780 (N_9780,N_434,N_2789);
nor U9781 (N_9781,N_3338,N_6113);
nor U9782 (N_9782,N_4609,N_5739);
and U9783 (N_9783,N_2366,N_3948);
nand U9784 (N_9784,N_5726,N_3093);
nand U9785 (N_9785,N_1368,N_4763);
nor U9786 (N_9786,N_5437,N_456);
and U9787 (N_9787,N_2553,N_131);
xor U9788 (N_9788,N_5332,N_4398);
nor U9789 (N_9789,N_4561,N_1350);
or U9790 (N_9790,N_499,N_5669);
and U9791 (N_9791,N_3618,N_6067);
or U9792 (N_9792,N_5716,N_5516);
or U9793 (N_9793,N_849,N_639);
xor U9794 (N_9794,N_2092,N_2313);
and U9795 (N_9795,N_1172,N_330);
or U9796 (N_9796,N_295,N_344);
or U9797 (N_9797,N_4457,N_3618);
or U9798 (N_9798,N_4431,N_2253);
or U9799 (N_9799,N_4462,N_6076);
xnor U9800 (N_9800,N_979,N_2348);
or U9801 (N_9801,N_5223,N_4369);
or U9802 (N_9802,N_1407,N_5939);
xor U9803 (N_9803,N_848,N_3292);
xor U9804 (N_9804,N_5917,N_1332);
nand U9805 (N_9805,N_2871,N_6249);
xor U9806 (N_9806,N_4041,N_3769);
and U9807 (N_9807,N_2796,N_6123);
and U9808 (N_9808,N_2759,N_5569);
and U9809 (N_9809,N_5477,N_1239);
and U9810 (N_9810,N_2326,N_869);
or U9811 (N_9811,N_1840,N_532);
and U9812 (N_9812,N_4732,N_5633);
xnor U9813 (N_9813,N_5403,N_2410);
nor U9814 (N_9814,N_483,N_1172);
xor U9815 (N_9815,N_485,N_1993);
nor U9816 (N_9816,N_4892,N_5505);
nand U9817 (N_9817,N_173,N_3065);
or U9818 (N_9818,N_534,N_5257);
nor U9819 (N_9819,N_5563,N_4632);
nand U9820 (N_9820,N_4895,N_1940);
nor U9821 (N_9821,N_5375,N_5525);
and U9822 (N_9822,N_3859,N_2519);
nor U9823 (N_9823,N_3234,N_1928);
or U9824 (N_9824,N_4453,N_3061);
nand U9825 (N_9825,N_4018,N_3358);
or U9826 (N_9826,N_863,N_5831);
nand U9827 (N_9827,N_1855,N_6118);
xor U9828 (N_9828,N_2800,N_2670);
nor U9829 (N_9829,N_3750,N_1147);
or U9830 (N_9830,N_5925,N_1393);
and U9831 (N_9831,N_3151,N_3655);
and U9832 (N_9832,N_1273,N_1353);
nor U9833 (N_9833,N_6019,N_1828);
or U9834 (N_9834,N_2835,N_3014);
or U9835 (N_9835,N_5788,N_3584);
nand U9836 (N_9836,N_75,N_4722);
or U9837 (N_9837,N_3308,N_3192);
xor U9838 (N_9838,N_1588,N_591);
or U9839 (N_9839,N_2869,N_4880);
or U9840 (N_9840,N_418,N_1724);
xnor U9841 (N_9841,N_1832,N_1818);
nor U9842 (N_9842,N_2126,N_2066);
or U9843 (N_9843,N_4111,N_5265);
or U9844 (N_9844,N_2769,N_6173);
xnor U9845 (N_9845,N_1419,N_3582);
and U9846 (N_9846,N_1080,N_3495);
or U9847 (N_9847,N_6007,N_4932);
or U9848 (N_9848,N_3552,N_6037);
xnor U9849 (N_9849,N_3323,N_3279);
nor U9850 (N_9850,N_1059,N_5867);
nand U9851 (N_9851,N_5272,N_4596);
nand U9852 (N_9852,N_814,N_5359);
nand U9853 (N_9853,N_2858,N_4530);
or U9854 (N_9854,N_635,N_5273);
or U9855 (N_9855,N_6110,N_5773);
and U9856 (N_9856,N_2961,N_2368);
or U9857 (N_9857,N_2903,N_0);
xor U9858 (N_9858,N_5341,N_3826);
nor U9859 (N_9859,N_4209,N_2645);
xor U9860 (N_9860,N_3446,N_3636);
and U9861 (N_9861,N_2565,N_3366);
xor U9862 (N_9862,N_5964,N_3851);
nor U9863 (N_9863,N_2856,N_2176);
nand U9864 (N_9864,N_568,N_4619);
and U9865 (N_9865,N_3441,N_5011);
xor U9866 (N_9866,N_337,N_5780);
and U9867 (N_9867,N_1093,N_3397);
or U9868 (N_9868,N_5804,N_4005);
and U9869 (N_9869,N_1671,N_4443);
xnor U9870 (N_9870,N_3330,N_4678);
or U9871 (N_9871,N_3925,N_3463);
nand U9872 (N_9872,N_3126,N_4540);
nor U9873 (N_9873,N_2571,N_3421);
and U9874 (N_9874,N_5918,N_3525);
xor U9875 (N_9875,N_4443,N_3514);
xor U9876 (N_9876,N_4243,N_4713);
nor U9877 (N_9877,N_4231,N_4885);
nand U9878 (N_9878,N_3938,N_3643);
nor U9879 (N_9879,N_5986,N_2280);
xor U9880 (N_9880,N_3905,N_5688);
and U9881 (N_9881,N_29,N_3040);
xor U9882 (N_9882,N_3205,N_2455);
and U9883 (N_9883,N_480,N_5118);
xnor U9884 (N_9884,N_5192,N_2414);
nor U9885 (N_9885,N_122,N_4227);
xor U9886 (N_9886,N_3650,N_923);
xor U9887 (N_9887,N_1540,N_4493);
or U9888 (N_9888,N_3884,N_4386);
nor U9889 (N_9889,N_4637,N_2577);
nor U9890 (N_9890,N_426,N_960);
or U9891 (N_9891,N_4676,N_5884);
nor U9892 (N_9892,N_3556,N_423);
xnor U9893 (N_9893,N_2519,N_3166);
nor U9894 (N_9894,N_5337,N_1550);
nor U9895 (N_9895,N_4152,N_3552);
nor U9896 (N_9896,N_4377,N_659);
or U9897 (N_9897,N_6051,N_1780);
or U9898 (N_9898,N_1928,N_2441);
or U9899 (N_9899,N_703,N_3486);
or U9900 (N_9900,N_5677,N_5239);
xor U9901 (N_9901,N_4282,N_4233);
and U9902 (N_9902,N_6186,N_238);
xnor U9903 (N_9903,N_184,N_6082);
nand U9904 (N_9904,N_1906,N_5166);
and U9905 (N_9905,N_5920,N_4544);
nand U9906 (N_9906,N_2920,N_5277);
or U9907 (N_9907,N_4951,N_5392);
and U9908 (N_9908,N_5738,N_1549);
nor U9909 (N_9909,N_5371,N_3008);
or U9910 (N_9910,N_5557,N_1772);
or U9911 (N_9911,N_934,N_5513);
nor U9912 (N_9912,N_1793,N_5478);
xnor U9913 (N_9913,N_208,N_3017);
nand U9914 (N_9914,N_2763,N_4728);
and U9915 (N_9915,N_4801,N_2404);
and U9916 (N_9916,N_1350,N_5391);
nor U9917 (N_9917,N_2533,N_3023);
or U9918 (N_9918,N_3872,N_5095);
xor U9919 (N_9919,N_5479,N_1169);
nor U9920 (N_9920,N_5547,N_3931);
nor U9921 (N_9921,N_5005,N_2051);
xnor U9922 (N_9922,N_16,N_363);
xor U9923 (N_9923,N_1336,N_3252);
or U9924 (N_9924,N_5993,N_5368);
xnor U9925 (N_9925,N_1707,N_546);
xnor U9926 (N_9926,N_4621,N_5291);
nand U9927 (N_9927,N_5499,N_1706);
or U9928 (N_9928,N_293,N_3084);
xor U9929 (N_9929,N_3894,N_1724);
and U9930 (N_9930,N_2808,N_5832);
and U9931 (N_9931,N_2403,N_5124);
and U9932 (N_9932,N_4486,N_3854);
nand U9933 (N_9933,N_5984,N_812);
xor U9934 (N_9934,N_3894,N_5545);
xor U9935 (N_9935,N_4486,N_1223);
or U9936 (N_9936,N_1037,N_3531);
and U9937 (N_9937,N_5387,N_2422);
xnor U9938 (N_9938,N_6213,N_5031);
xor U9939 (N_9939,N_5561,N_3969);
and U9940 (N_9940,N_3241,N_6182);
or U9941 (N_9941,N_1559,N_3783);
xor U9942 (N_9942,N_2144,N_3164);
nor U9943 (N_9943,N_1425,N_3716);
xnor U9944 (N_9944,N_2791,N_4320);
or U9945 (N_9945,N_2650,N_5254);
and U9946 (N_9946,N_3444,N_5688);
xor U9947 (N_9947,N_1808,N_2862);
or U9948 (N_9948,N_1830,N_1419);
or U9949 (N_9949,N_5532,N_1307);
or U9950 (N_9950,N_4994,N_4089);
xor U9951 (N_9951,N_108,N_991);
nand U9952 (N_9952,N_4442,N_3058);
nor U9953 (N_9953,N_4406,N_2361);
xor U9954 (N_9954,N_3358,N_5796);
nor U9955 (N_9955,N_2980,N_4579);
xnor U9956 (N_9956,N_2041,N_2955);
xnor U9957 (N_9957,N_4061,N_3133);
xnor U9958 (N_9958,N_1310,N_3020);
nand U9959 (N_9959,N_4014,N_2234);
xor U9960 (N_9960,N_1445,N_3971);
nand U9961 (N_9961,N_5190,N_3747);
and U9962 (N_9962,N_3364,N_1039);
or U9963 (N_9963,N_2688,N_4478);
xor U9964 (N_9964,N_5389,N_1111);
and U9965 (N_9965,N_5963,N_284);
or U9966 (N_9966,N_137,N_2082);
or U9967 (N_9967,N_1772,N_5944);
and U9968 (N_9968,N_4135,N_3837);
nor U9969 (N_9969,N_4381,N_1809);
nand U9970 (N_9970,N_5663,N_3446);
nand U9971 (N_9971,N_2281,N_2235);
and U9972 (N_9972,N_2916,N_1685);
nand U9973 (N_9973,N_1756,N_4524);
and U9974 (N_9974,N_939,N_1308);
xnor U9975 (N_9975,N_416,N_2588);
and U9976 (N_9976,N_854,N_5342);
nand U9977 (N_9977,N_713,N_5191);
or U9978 (N_9978,N_1912,N_4736);
nor U9979 (N_9979,N_5885,N_335);
xor U9980 (N_9980,N_5331,N_5385);
nand U9981 (N_9981,N_2934,N_5403);
or U9982 (N_9982,N_325,N_5454);
or U9983 (N_9983,N_6104,N_895);
nor U9984 (N_9984,N_2383,N_5198);
xnor U9985 (N_9985,N_4349,N_69);
xnor U9986 (N_9986,N_5552,N_633);
and U9987 (N_9987,N_5371,N_2742);
nor U9988 (N_9988,N_5720,N_2364);
nor U9989 (N_9989,N_1081,N_2294);
and U9990 (N_9990,N_3878,N_2571);
nor U9991 (N_9991,N_975,N_2413);
and U9992 (N_9992,N_859,N_1211);
nand U9993 (N_9993,N_438,N_3819);
xnor U9994 (N_9994,N_3098,N_3383);
or U9995 (N_9995,N_4705,N_4592);
or U9996 (N_9996,N_5123,N_3552);
nand U9997 (N_9997,N_904,N_3562);
nor U9998 (N_9998,N_2093,N_4828);
xor U9999 (N_9999,N_4174,N_4253);
xnor U10000 (N_10000,N_5415,N_5133);
and U10001 (N_10001,N_319,N_5425);
and U10002 (N_10002,N_1778,N_4606);
xor U10003 (N_10003,N_5257,N_2859);
nand U10004 (N_10004,N_5669,N_790);
and U10005 (N_10005,N_1197,N_964);
xnor U10006 (N_10006,N_490,N_1766);
xor U10007 (N_10007,N_548,N_4490);
nand U10008 (N_10008,N_5773,N_6244);
nor U10009 (N_10009,N_4611,N_5770);
nor U10010 (N_10010,N_1962,N_690);
or U10011 (N_10011,N_4319,N_6124);
or U10012 (N_10012,N_472,N_4046);
nor U10013 (N_10013,N_629,N_2163);
xor U10014 (N_10014,N_1510,N_5300);
or U10015 (N_10015,N_3489,N_985);
or U10016 (N_10016,N_1918,N_3621);
nand U10017 (N_10017,N_571,N_843);
and U10018 (N_10018,N_424,N_1663);
xnor U10019 (N_10019,N_2207,N_4906);
or U10020 (N_10020,N_4330,N_912);
xnor U10021 (N_10021,N_1113,N_2499);
or U10022 (N_10022,N_4872,N_1470);
nor U10023 (N_10023,N_1834,N_310);
and U10024 (N_10024,N_2812,N_4259);
xor U10025 (N_10025,N_4974,N_4191);
nand U10026 (N_10026,N_5129,N_4641);
and U10027 (N_10027,N_3532,N_5927);
and U10028 (N_10028,N_3112,N_1378);
xnor U10029 (N_10029,N_3453,N_2831);
nor U10030 (N_10030,N_4407,N_1423);
nand U10031 (N_10031,N_436,N_305);
or U10032 (N_10032,N_3580,N_1285);
or U10033 (N_10033,N_1537,N_5986);
nor U10034 (N_10034,N_977,N_4406);
nor U10035 (N_10035,N_5421,N_251);
and U10036 (N_10036,N_3103,N_4727);
nand U10037 (N_10037,N_3169,N_1765);
or U10038 (N_10038,N_273,N_5328);
xnor U10039 (N_10039,N_4909,N_2924);
nand U10040 (N_10040,N_6169,N_1391);
and U10041 (N_10041,N_2079,N_2803);
nand U10042 (N_10042,N_1655,N_2502);
xnor U10043 (N_10043,N_2450,N_1274);
xor U10044 (N_10044,N_2890,N_5866);
nand U10045 (N_10045,N_4865,N_182);
xor U10046 (N_10046,N_1848,N_1476);
or U10047 (N_10047,N_5569,N_543);
xnor U10048 (N_10048,N_1956,N_655);
or U10049 (N_10049,N_3804,N_3734);
xnor U10050 (N_10050,N_4285,N_4798);
nand U10051 (N_10051,N_5101,N_892);
or U10052 (N_10052,N_1050,N_4479);
nand U10053 (N_10053,N_1435,N_6021);
or U10054 (N_10054,N_4058,N_261);
and U10055 (N_10055,N_738,N_3930);
nor U10056 (N_10056,N_6077,N_5563);
nor U10057 (N_10057,N_5416,N_3877);
nand U10058 (N_10058,N_4793,N_5957);
or U10059 (N_10059,N_2293,N_72);
or U10060 (N_10060,N_3055,N_3639);
and U10061 (N_10061,N_4050,N_2186);
nor U10062 (N_10062,N_1801,N_3933);
and U10063 (N_10063,N_5011,N_834);
xnor U10064 (N_10064,N_1130,N_5905);
nor U10065 (N_10065,N_5971,N_3716);
xnor U10066 (N_10066,N_2899,N_479);
xor U10067 (N_10067,N_2684,N_2618);
nand U10068 (N_10068,N_3680,N_46);
nand U10069 (N_10069,N_1344,N_2783);
or U10070 (N_10070,N_4924,N_5113);
and U10071 (N_10071,N_1062,N_4920);
nor U10072 (N_10072,N_5102,N_2577);
or U10073 (N_10073,N_5586,N_3286);
and U10074 (N_10074,N_230,N_2093);
and U10075 (N_10075,N_5570,N_2069);
nor U10076 (N_10076,N_957,N_1831);
nor U10077 (N_10077,N_2120,N_1970);
nand U10078 (N_10078,N_4502,N_4900);
nand U10079 (N_10079,N_5053,N_6007);
xnor U10080 (N_10080,N_4876,N_3350);
xnor U10081 (N_10081,N_5163,N_4163);
nand U10082 (N_10082,N_1295,N_5049);
nor U10083 (N_10083,N_4192,N_5567);
and U10084 (N_10084,N_765,N_862);
or U10085 (N_10085,N_713,N_2039);
and U10086 (N_10086,N_5968,N_3259);
nor U10087 (N_10087,N_3727,N_791);
nand U10088 (N_10088,N_197,N_4604);
nand U10089 (N_10089,N_3261,N_4000);
nor U10090 (N_10090,N_4019,N_3687);
and U10091 (N_10091,N_1843,N_5134);
xnor U10092 (N_10092,N_1841,N_4795);
or U10093 (N_10093,N_3585,N_3991);
and U10094 (N_10094,N_5230,N_963);
nand U10095 (N_10095,N_3203,N_1585);
nand U10096 (N_10096,N_3187,N_1426);
or U10097 (N_10097,N_4822,N_3395);
or U10098 (N_10098,N_5649,N_3336);
and U10099 (N_10099,N_3809,N_2578);
xor U10100 (N_10100,N_5601,N_2674);
nand U10101 (N_10101,N_3854,N_1362);
xnor U10102 (N_10102,N_5735,N_1838);
and U10103 (N_10103,N_3649,N_5027);
and U10104 (N_10104,N_2384,N_5815);
and U10105 (N_10105,N_5656,N_3572);
xnor U10106 (N_10106,N_332,N_3525);
xor U10107 (N_10107,N_4652,N_402);
and U10108 (N_10108,N_1837,N_2464);
and U10109 (N_10109,N_1769,N_391);
or U10110 (N_10110,N_2556,N_4693);
xor U10111 (N_10111,N_3246,N_3852);
nand U10112 (N_10112,N_763,N_1894);
and U10113 (N_10113,N_5726,N_2513);
or U10114 (N_10114,N_4482,N_4916);
and U10115 (N_10115,N_3183,N_6070);
or U10116 (N_10116,N_1740,N_3858);
nand U10117 (N_10117,N_1057,N_5266);
xor U10118 (N_10118,N_6216,N_2119);
nor U10119 (N_10119,N_4381,N_3256);
nor U10120 (N_10120,N_1779,N_1088);
nor U10121 (N_10121,N_1460,N_3574);
nor U10122 (N_10122,N_3047,N_1813);
and U10123 (N_10123,N_7,N_5057);
nand U10124 (N_10124,N_1277,N_3856);
nand U10125 (N_10125,N_1801,N_3393);
nor U10126 (N_10126,N_1381,N_4667);
nand U10127 (N_10127,N_172,N_5579);
or U10128 (N_10128,N_3116,N_2962);
and U10129 (N_10129,N_1929,N_1863);
and U10130 (N_10130,N_6125,N_161);
nand U10131 (N_10131,N_2846,N_906);
and U10132 (N_10132,N_4539,N_82);
and U10133 (N_10133,N_4424,N_3044);
xnor U10134 (N_10134,N_5200,N_3528);
xor U10135 (N_10135,N_1005,N_5879);
nand U10136 (N_10136,N_6150,N_4300);
nand U10137 (N_10137,N_4515,N_661);
xnor U10138 (N_10138,N_5605,N_1103);
or U10139 (N_10139,N_200,N_5210);
and U10140 (N_10140,N_4970,N_3381);
nand U10141 (N_10141,N_4941,N_5014);
xor U10142 (N_10142,N_5670,N_3701);
nor U10143 (N_10143,N_1075,N_3197);
or U10144 (N_10144,N_5560,N_4716);
xnor U10145 (N_10145,N_402,N_1019);
or U10146 (N_10146,N_2758,N_1758);
xnor U10147 (N_10147,N_5301,N_1204);
nor U10148 (N_10148,N_1570,N_3611);
xnor U10149 (N_10149,N_1579,N_5513);
or U10150 (N_10150,N_1118,N_4940);
nor U10151 (N_10151,N_4533,N_5969);
or U10152 (N_10152,N_4717,N_1061);
nand U10153 (N_10153,N_1918,N_4640);
nand U10154 (N_10154,N_4738,N_4515);
and U10155 (N_10155,N_3145,N_3721);
or U10156 (N_10156,N_5175,N_295);
nand U10157 (N_10157,N_5697,N_564);
nor U10158 (N_10158,N_448,N_1246);
or U10159 (N_10159,N_706,N_5997);
nand U10160 (N_10160,N_3603,N_5631);
nor U10161 (N_10161,N_3334,N_148);
or U10162 (N_10162,N_5344,N_4862);
and U10163 (N_10163,N_5462,N_3401);
xnor U10164 (N_10164,N_4217,N_485);
or U10165 (N_10165,N_5024,N_2164);
xnor U10166 (N_10166,N_2851,N_3807);
nand U10167 (N_10167,N_2994,N_5981);
nand U10168 (N_10168,N_6228,N_314);
and U10169 (N_10169,N_6128,N_5821);
or U10170 (N_10170,N_3135,N_2552);
and U10171 (N_10171,N_4920,N_6058);
nand U10172 (N_10172,N_1214,N_3212);
and U10173 (N_10173,N_2769,N_2023);
nor U10174 (N_10174,N_5559,N_4544);
and U10175 (N_10175,N_1032,N_1687);
or U10176 (N_10176,N_1953,N_2904);
nor U10177 (N_10177,N_3339,N_3231);
and U10178 (N_10178,N_188,N_3905);
nand U10179 (N_10179,N_1873,N_3160);
and U10180 (N_10180,N_493,N_4637);
nand U10181 (N_10181,N_5121,N_5449);
nor U10182 (N_10182,N_1514,N_3544);
or U10183 (N_10183,N_320,N_5421);
nor U10184 (N_10184,N_5217,N_5576);
xor U10185 (N_10185,N_711,N_4159);
nand U10186 (N_10186,N_990,N_5486);
xnor U10187 (N_10187,N_1389,N_6100);
or U10188 (N_10188,N_2606,N_932);
or U10189 (N_10189,N_6057,N_3109);
and U10190 (N_10190,N_66,N_2627);
and U10191 (N_10191,N_5257,N_1732);
or U10192 (N_10192,N_2089,N_1164);
and U10193 (N_10193,N_5690,N_2413);
xor U10194 (N_10194,N_3382,N_2901);
xor U10195 (N_10195,N_5159,N_3810);
xnor U10196 (N_10196,N_1889,N_2143);
nand U10197 (N_10197,N_2549,N_271);
or U10198 (N_10198,N_4573,N_3446);
or U10199 (N_10199,N_6022,N_745);
or U10200 (N_10200,N_3378,N_1484);
xor U10201 (N_10201,N_6128,N_3990);
xnor U10202 (N_10202,N_450,N_3934);
xor U10203 (N_10203,N_2957,N_2674);
xor U10204 (N_10204,N_6099,N_4250);
nor U10205 (N_10205,N_4052,N_3612);
or U10206 (N_10206,N_6145,N_2476);
and U10207 (N_10207,N_2288,N_337);
xor U10208 (N_10208,N_2025,N_3608);
nand U10209 (N_10209,N_2523,N_3343);
nand U10210 (N_10210,N_4538,N_1827);
or U10211 (N_10211,N_5640,N_1684);
nor U10212 (N_10212,N_3830,N_4158);
xor U10213 (N_10213,N_2235,N_5439);
and U10214 (N_10214,N_1934,N_1039);
or U10215 (N_10215,N_5006,N_6224);
nor U10216 (N_10216,N_4282,N_1765);
or U10217 (N_10217,N_1409,N_1074);
nand U10218 (N_10218,N_4549,N_351);
nor U10219 (N_10219,N_5732,N_3031);
or U10220 (N_10220,N_357,N_5538);
nor U10221 (N_10221,N_5782,N_5883);
xnor U10222 (N_10222,N_5798,N_5759);
and U10223 (N_10223,N_4698,N_4468);
and U10224 (N_10224,N_357,N_3300);
and U10225 (N_10225,N_1740,N_3912);
nand U10226 (N_10226,N_6081,N_217);
nand U10227 (N_10227,N_1312,N_5557);
nand U10228 (N_10228,N_1838,N_5590);
and U10229 (N_10229,N_5984,N_4325);
and U10230 (N_10230,N_2691,N_4214);
or U10231 (N_10231,N_5736,N_3221);
or U10232 (N_10232,N_2405,N_5048);
and U10233 (N_10233,N_1350,N_2707);
xnor U10234 (N_10234,N_1805,N_2488);
or U10235 (N_10235,N_2201,N_6222);
xor U10236 (N_10236,N_2455,N_3868);
xnor U10237 (N_10237,N_2302,N_239);
nor U10238 (N_10238,N_3469,N_3547);
nand U10239 (N_10239,N_22,N_3356);
and U10240 (N_10240,N_4407,N_2260);
xnor U10241 (N_10241,N_916,N_3804);
nand U10242 (N_10242,N_9,N_4388);
nand U10243 (N_10243,N_3918,N_1067);
nor U10244 (N_10244,N_151,N_984);
or U10245 (N_10245,N_4953,N_1897);
and U10246 (N_10246,N_2946,N_1061);
and U10247 (N_10247,N_2108,N_355);
or U10248 (N_10248,N_2688,N_1765);
or U10249 (N_10249,N_1453,N_636);
or U10250 (N_10250,N_2629,N_2722);
and U10251 (N_10251,N_6051,N_3461);
or U10252 (N_10252,N_4796,N_813);
and U10253 (N_10253,N_3804,N_5221);
xnor U10254 (N_10254,N_3152,N_2078);
and U10255 (N_10255,N_3485,N_5909);
nor U10256 (N_10256,N_1828,N_3866);
and U10257 (N_10257,N_3624,N_4309);
nand U10258 (N_10258,N_5715,N_4792);
nand U10259 (N_10259,N_1811,N_3692);
xnor U10260 (N_10260,N_1135,N_5705);
nand U10261 (N_10261,N_950,N_4651);
nand U10262 (N_10262,N_5309,N_5522);
and U10263 (N_10263,N_1372,N_5577);
nand U10264 (N_10264,N_324,N_5882);
or U10265 (N_10265,N_5350,N_1413);
and U10266 (N_10266,N_4565,N_4325);
nand U10267 (N_10267,N_4657,N_3034);
xnor U10268 (N_10268,N_3135,N_2009);
nand U10269 (N_10269,N_5680,N_7);
xnor U10270 (N_10270,N_4178,N_5742);
nor U10271 (N_10271,N_3480,N_2625);
and U10272 (N_10272,N_2299,N_714);
nor U10273 (N_10273,N_1215,N_2931);
and U10274 (N_10274,N_4948,N_2149);
and U10275 (N_10275,N_5482,N_3098);
nand U10276 (N_10276,N_496,N_5233);
or U10277 (N_10277,N_3386,N_4031);
and U10278 (N_10278,N_1107,N_5550);
nand U10279 (N_10279,N_2398,N_2700);
xor U10280 (N_10280,N_1006,N_4087);
or U10281 (N_10281,N_3707,N_1054);
xnor U10282 (N_10282,N_938,N_920);
nand U10283 (N_10283,N_5427,N_1898);
and U10284 (N_10284,N_3510,N_5868);
nand U10285 (N_10285,N_5282,N_5528);
nand U10286 (N_10286,N_80,N_554);
nor U10287 (N_10287,N_1726,N_856);
nor U10288 (N_10288,N_1505,N_2382);
or U10289 (N_10289,N_692,N_909);
and U10290 (N_10290,N_2801,N_1322);
and U10291 (N_10291,N_2197,N_2563);
and U10292 (N_10292,N_1692,N_1232);
nand U10293 (N_10293,N_1480,N_3559);
or U10294 (N_10294,N_2756,N_4682);
and U10295 (N_10295,N_4375,N_1823);
and U10296 (N_10296,N_1669,N_946);
xnor U10297 (N_10297,N_2279,N_2305);
or U10298 (N_10298,N_5046,N_6008);
nor U10299 (N_10299,N_1635,N_5692);
or U10300 (N_10300,N_2281,N_476);
or U10301 (N_10301,N_1526,N_1096);
xnor U10302 (N_10302,N_4852,N_909);
xnor U10303 (N_10303,N_2883,N_368);
nand U10304 (N_10304,N_4314,N_2873);
nor U10305 (N_10305,N_3518,N_1353);
nand U10306 (N_10306,N_3844,N_2715);
xor U10307 (N_10307,N_1060,N_3723);
nor U10308 (N_10308,N_1341,N_5456);
nor U10309 (N_10309,N_3344,N_696);
and U10310 (N_10310,N_1621,N_141);
xnor U10311 (N_10311,N_604,N_643);
or U10312 (N_10312,N_2891,N_3489);
xnor U10313 (N_10313,N_5578,N_1565);
xor U10314 (N_10314,N_167,N_6116);
and U10315 (N_10315,N_3145,N_6033);
xnor U10316 (N_10316,N_251,N_3277);
xor U10317 (N_10317,N_1026,N_2638);
or U10318 (N_10318,N_3340,N_5262);
or U10319 (N_10319,N_1898,N_2328);
or U10320 (N_10320,N_4557,N_2540);
nand U10321 (N_10321,N_151,N_6132);
nand U10322 (N_10322,N_286,N_778);
or U10323 (N_10323,N_5595,N_127);
xnor U10324 (N_10324,N_2479,N_927);
xnor U10325 (N_10325,N_977,N_3709);
nand U10326 (N_10326,N_5136,N_1156);
and U10327 (N_10327,N_4584,N_3402);
xor U10328 (N_10328,N_3441,N_2456);
nor U10329 (N_10329,N_5398,N_3495);
xor U10330 (N_10330,N_2820,N_5665);
and U10331 (N_10331,N_1312,N_4);
or U10332 (N_10332,N_5662,N_1857);
nor U10333 (N_10333,N_2832,N_2520);
xnor U10334 (N_10334,N_5894,N_5379);
xor U10335 (N_10335,N_1628,N_1383);
nand U10336 (N_10336,N_5502,N_3003);
nand U10337 (N_10337,N_1208,N_2519);
xor U10338 (N_10338,N_2971,N_6012);
xnor U10339 (N_10339,N_217,N_1898);
xnor U10340 (N_10340,N_5219,N_6126);
nand U10341 (N_10341,N_4320,N_3637);
nor U10342 (N_10342,N_2780,N_2774);
xor U10343 (N_10343,N_4643,N_2253);
and U10344 (N_10344,N_277,N_3987);
nor U10345 (N_10345,N_3708,N_5674);
or U10346 (N_10346,N_5179,N_6130);
xor U10347 (N_10347,N_819,N_5532);
nand U10348 (N_10348,N_1919,N_3392);
and U10349 (N_10349,N_1196,N_2853);
nand U10350 (N_10350,N_68,N_3657);
xor U10351 (N_10351,N_3118,N_4666);
and U10352 (N_10352,N_4524,N_668);
nor U10353 (N_10353,N_5686,N_534);
nand U10354 (N_10354,N_5857,N_1271);
nand U10355 (N_10355,N_5257,N_4527);
or U10356 (N_10356,N_2108,N_2771);
or U10357 (N_10357,N_4029,N_1926);
nor U10358 (N_10358,N_4491,N_522);
xor U10359 (N_10359,N_3165,N_7);
nor U10360 (N_10360,N_3909,N_530);
or U10361 (N_10361,N_5520,N_941);
and U10362 (N_10362,N_146,N_385);
nor U10363 (N_10363,N_2525,N_6031);
or U10364 (N_10364,N_6083,N_5745);
nor U10365 (N_10365,N_2236,N_3743);
or U10366 (N_10366,N_2456,N_4080);
nor U10367 (N_10367,N_6153,N_679);
or U10368 (N_10368,N_5448,N_1886);
nor U10369 (N_10369,N_4694,N_6083);
or U10370 (N_10370,N_4796,N_2453);
nand U10371 (N_10371,N_6163,N_1844);
and U10372 (N_10372,N_2210,N_1446);
and U10373 (N_10373,N_407,N_3176);
xor U10374 (N_10374,N_2465,N_5730);
xor U10375 (N_10375,N_4365,N_4375);
xnor U10376 (N_10376,N_2891,N_5692);
xnor U10377 (N_10377,N_5645,N_5609);
nand U10378 (N_10378,N_5267,N_716);
or U10379 (N_10379,N_1943,N_6189);
nor U10380 (N_10380,N_2003,N_67);
nand U10381 (N_10381,N_559,N_980);
nand U10382 (N_10382,N_1033,N_5464);
nor U10383 (N_10383,N_6239,N_1835);
nand U10384 (N_10384,N_5350,N_3946);
xnor U10385 (N_10385,N_3981,N_5639);
and U10386 (N_10386,N_2007,N_2650);
nor U10387 (N_10387,N_2619,N_4379);
or U10388 (N_10388,N_542,N_3293);
nor U10389 (N_10389,N_4941,N_325);
or U10390 (N_10390,N_3635,N_4755);
nand U10391 (N_10391,N_5443,N_2383);
xor U10392 (N_10392,N_2818,N_5176);
nor U10393 (N_10393,N_5414,N_6158);
or U10394 (N_10394,N_1414,N_6087);
nor U10395 (N_10395,N_3673,N_6201);
and U10396 (N_10396,N_5303,N_3165);
and U10397 (N_10397,N_6090,N_5281);
xor U10398 (N_10398,N_2492,N_4074);
nor U10399 (N_10399,N_4678,N_4690);
xnor U10400 (N_10400,N_2575,N_3785);
nand U10401 (N_10401,N_5474,N_1719);
and U10402 (N_10402,N_857,N_5138);
xnor U10403 (N_10403,N_601,N_444);
nand U10404 (N_10404,N_4500,N_103);
or U10405 (N_10405,N_3762,N_2208);
and U10406 (N_10406,N_5785,N_4294);
and U10407 (N_10407,N_441,N_4887);
nor U10408 (N_10408,N_3472,N_3271);
or U10409 (N_10409,N_6248,N_529);
or U10410 (N_10410,N_1637,N_3540);
nor U10411 (N_10411,N_5833,N_100);
xnor U10412 (N_10412,N_5776,N_5729);
nor U10413 (N_10413,N_5755,N_4593);
and U10414 (N_10414,N_2178,N_2891);
and U10415 (N_10415,N_4872,N_2810);
nor U10416 (N_10416,N_2365,N_3892);
xnor U10417 (N_10417,N_1171,N_5867);
nand U10418 (N_10418,N_4953,N_3181);
xor U10419 (N_10419,N_3041,N_2496);
nand U10420 (N_10420,N_4860,N_3436);
and U10421 (N_10421,N_5596,N_616);
nor U10422 (N_10422,N_237,N_599);
or U10423 (N_10423,N_6229,N_3356);
xor U10424 (N_10424,N_2685,N_1359);
xnor U10425 (N_10425,N_1736,N_649);
and U10426 (N_10426,N_3863,N_2383);
nand U10427 (N_10427,N_2084,N_4764);
nand U10428 (N_10428,N_5934,N_3871);
xor U10429 (N_10429,N_3952,N_3924);
and U10430 (N_10430,N_5539,N_2946);
or U10431 (N_10431,N_1915,N_4310);
and U10432 (N_10432,N_3482,N_96);
nor U10433 (N_10433,N_4889,N_5745);
xor U10434 (N_10434,N_4329,N_1383);
and U10435 (N_10435,N_176,N_1432);
nand U10436 (N_10436,N_2305,N_5617);
nor U10437 (N_10437,N_5611,N_722);
and U10438 (N_10438,N_5332,N_106);
or U10439 (N_10439,N_212,N_6007);
xnor U10440 (N_10440,N_4752,N_4618);
or U10441 (N_10441,N_225,N_3900);
nand U10442 (N_10442,N_5383,N_3973);
or U10443 (N_10443,N_5869,N_4108);
and U10444 (N_10444,N_1931,N_3959);
xnor U10445 (N_10445,N_5064,N_4124);
and U10446 (N_10446,N_2496,N_2083);
nor U10447 (N_10447,N_5914,N_5017);
nor U10448 (N_10448,N_1105,N_4480);
nor U10449 (N_10449,N_4254,N_2461);
xnor U10450 (N_10450,N_3901,N_3772);
nand U10451 (N_10451,N_1628,N_4728);
or U10452 (N_10452,N_740,N_1363);
and U10453 (N_10453,N_624,N_2504);
or U10454 (N_10454,N_4928,N_3190);
nor U10455 (N_10455,N_34,N_5390);
and U10456 (N_10456,N_4128,N_544);
and U10457 (N_10457,N_4639,N_1842);
xnor U10458 (N_10458,N_3830,N_3112);
or U10459 (N_10459,N_4071,N_649);
or U10460 (N_10460,N_2801,N_1647);
or U10461 (N_10461,N_1353,N_242);
nand U10462 (N_10462,N_4885,N_564);
or U10463 (N_10463,N_5964,N_5376);
nor U10464 (N_10464,N_1094,N_1178);
xnor U10465 (N_10465,N_3549,N_5267);
nor U10466 (N_10466,N_5850,N_1139);
nand U10467 (N_10467,N_3924,N_5965);
xor U10468 (N_10468,N_220,N_876);
nor U10469 (N_10469,N_3979,N_2889);
or U10470 (N_10470,N_2801,N_3141);
and U10471 (N_10471,N_1612,N_6132);
or U10472 (N_10472,N_6162,N_2051);
and U10473 (N_10473,N_4349,N_4877);
or U10474 (N_10474,N_4308,N_6167);
or U10475 (N_10475,N_6204,N_3957);
nand U10476 (N_10476,N_2459,N_4608);
or U10477 (N_10477,N_348,N_4184);
nand U10478 (N_10478,N_3488,N_4907);
nor U10479 (N_10479,N_5531,N_3063);
nor U10480 (N_10480,N_2130,N_1476);
or U10481 (N_10481,N_1450,N_5998);
nand U10482 (N_10482,N_5093,N_6224);
and U10483 (N_10483,N_667,N_4125);
or U10484 (N_10484,N_2301,N_4066);
xor U10485 (N_10485,N_1554,N_2236);
xor U10486 (N_10486,N_2750,N_362);
xor U10487 (N_10487,N_1915,N_26);
and U10488 (N_10488,N_3292,N_889);
xnor U10489 (N_10489,N_1917,N_4256);
nor U10490 (N_10490,N_693,N_2555);
nand U10491 (N_10491,N_4961,N_2220);
xor U10492 (N_10492,N_4725,N_3096);
xor U10493 (N_10493,N_1041,N_2863);
nor U10494 (N_10494,N_2783,N_1966);
or U10495 (N_10495,N_2188,N_1772);
nand U10496 (N_10496,N_4257,N_2887);
or U10497 (N_10497,N_5621,N_4603);
nor U10498 (N_10498,N_4578,N_3398);
nand U10499 (N_10499,N_4229,N_2444);
nand U10500 (N_10500,N_4321,N_3546);
or U10501 (N_10501,N_2793,N_936);
and U10502 (N_10502,N_2607,N_257);
nand U10503 (N_10503,N_5230,N_4306);
or U10504 (N_10504,N_5262,N_5147);
and U10505 (N_10505,N_3430,N_3836);
xor U10506 (N_10506,N_503,N_1299);
nand U10507 (N_10507,N_4753,N_4773);
or U10508 (N_10508,N_5908,N_3512);
and U10509 (N_10509,N_1004,N_2320);
xnor U10510 (N_10510,N_2817,N_3897);
nor U10511 (N_10511,N_5618,N_5668);
xnor U10512 (N_10512,N_3830,N_996);
nor U10513 (N_10513,N_3489,N_1113);
nand U10514 (N_10514,N_1858,N_4068);
and U10515 (N_10515,N_6112,N_5509);
nand U10516 (N_10516,N_3480,N_1777);
or U10517 (N_10517,N_4383,N_2801);
nand U10518 (N_10518,N_4997,N_2629);
or U10519 (N_10519,N_4300,N_5585);
or U10520 (N_10520,N_4689,N_1125);
nor U10521 (N_10521,N_3230,N_2213);
xnor U10522 (N_10522,N_5944,N_5641);
or U10523 (N_10523,N_3025,N_5747);
nand U10524 (N_10524,N_2528,N_2640);
and U10525 (N_10525,N_745,N_1843);
xor U10526 (N_10526,N_5914,N_1479);
nor U10527 (N_10527,N_2172,N_2792);
nor U10528 (N_10528,N_714,N_3202);
nand U10529 (N_10529,N_1776,N_2374);
nand U10530 (N_10530,N_1847,N_805);
xnor U10531 (N_10531,N_1388,N_620);
and U10532 (N_10532,N_4502,N_5514);
nor U10533 (N_10533,N_671,N_4197);
xnor U10534 (N_10534,N_2307,N_5974);
or U10535 (N_10535,N_4070,N_4506);
nor U10536 (N_10536,N_4788,N_3898);
nand U10537 (N_10537,N_599,N_466);
or U10538 (N_10538,N_4444,N_2100);
or U10539 (N_10539,N_6044,N_2588);
xor U10540 (N_10540,N_4000,N_1690);
nand U10541 (N_10541,N_2628,N_2508);
nand U10542 (N_10542,N_4110,N_4790);
nand U10543 (N_10543,N_6197,N_2606);
and U10544 (N_10544,N_3875,N_358);
nand U10545 (N_10545,N_4639,N_5038);
and U10546 (N_10546,N_5323,N_4638);
nor U10547 (N_10547,N_4606,N_5815);
and U10548 (N_10548,N_1938,N_2539);
and U10549 (N_10549,N_2486,N_4277);
nor U10550 (N_10550,N_4539,N_3027);
nor U10551 (N_10551,N_892,N_1685);
or U10552 (N_10552,N_2449,N_446);
nand U10553 (N_10553,N_4232,N_831);
nand U10554 (N_10554,N_6215,N_3873);
or U10555 (N_10555,N_833,N_4907);
xor U10556 (N_10556,N_262,N_4189);
nand U10557 (N_10557,N_3466,N_2483);
nand U10558 (N_10558,N_5233,N_5521);
or U10559 (N_10559,N_5696,N_5741);
or U10560 (N_10560,N_5402,N_6219);
and U10561 (N_10561,N_3753,N_49);
xnor U10562 (N_10562,N_1323,N_680);
and U10563 (N_10563,N_1286,N_3702);
xnor U10564 (N_10564,N_815,N_1099);
xnor U10565 (N_10565,N_288,N_1379);
and U10566 (N_10566,N_4400,N_1911);
or U10567 (N_10567,N_4026,N_2185);
xor U10568 (N_10568,N_5379,N_1721);
nor U10569 (N_10569,N_1960,N_2598);
or U10570 (N_10570,N_2654,N_323);
nand U10571 (N_10571,N_770,N_1848);
and U10572 (N_10572,N_798,N_4151);
nor U10573 (N_10573,N_69,N_197);
xor U10574 (N_10574,N_3070,N_1484);
and U10575 (N_10575,N_515,N_5682);
or U10576 (N_10576,N_5965,N_4158);
or U10577 (N_10577,N_1216,N_2304);
and U10578 (N_10578,N_6122,N_5854);
xor U10579 (N_10579,N_5403,N_1049);
xor U10580 (N_10580,N_384,N_2704);
xor U10581 (N_10581,N_515,N_5472);
nand U10582 (N_10582,N_5123,N_291);
xnor U10583 (N_10583,N_4103,N_720);
nor U10584 (N_10584,N_1727,N_499);
and U10585 (N_10585,N_2626,N_1548);
nor U10586 (N_10586,N_974,N_2431);
or U10587 (N_10587,N_3742,N_2742);
nand U10588 (N_10588,N_4461,N_2019);
and U10589 (N_10589,N_2362,N_1231);
or U10590 (N_10590,N_2693,N_6030);
xor U10591 (N_10591,N_2983,N_3837);
nor U10592 (N_10592,N_1300,N_250);
and U10593 (N_10593,N_5883,N_1347);
nand U10594 (N_10594,N_1770,N_408);
nor U10595 (N_10595,N_10,N_5212);
and U10596 (N_10596,N_5756,N_5291);
nor U10597 (N_10597,N_3467,N_4097);
nand U10598 (N_10598,N_2865,N_3221);
nor U10599 (N_10599,N_4151,N_5359);
and U10600 (N_10600,N_3212,N_1479);
xnor U10601 (N_10601,N_4277,N_5471);
or U10602 (N_10602,N_275,N_6010);
nor U10603 (N_10603,N_5654,N_4070);
and U10604 (N_10604,N_3892,N_4212);
nor U10605 (N_10605,N_5078,N_4924);
nand U10606 (N_10606,N_1764,N_1436);
xnor U10607 (N_10607,N_956,N_4762);
xnor U10608 (N_10608,N_1601,N_5504);
nor U10609 (N_10609,N_5108,N_1773);
or U10610 (N_10610,N_3122,N_6188);
or U10611 (N_10611,N_4790,N_5081);
nand U10612 (N_10612,N_6130,N_716);
or U10613 (N_10613,N_2320,N_40);
nand U10614 (N_10614,N_5298,N_5564);
nand U10615 (N_10615,N_4357,N_3847);
xnor U10616 (N_10616,N_4822,N_968);
or U10617 (N_10617,N_5408,N_2461);
and U10618 (N_10618,N_4709,N_309);
nand U10619 (N_10619,N_5480,N_2128);
or U10620 (N_10620,N_669,N_103);
xor U10621 (N_10621,N_2556,N_2630);
and U10622 (N_10622,N_6084,N_5448);
nor U10623 (N_10623,N_5244,N_1056);
nor U10624 (N_10624,N_129,N_4049);
xnor U10625 (N_10625,N_751,N_3425);
nor U10626 (N_10626,N_6246,N_1988);
nor U10627 (N_10627,N_989,N_436);
and U10628 (N_10628,N_3962,N_1618);
and U10629 (N_10629,N_8,N_4490);
nor U10630 (N_10630,N_299,N_4521);
nor U10631 (N_10631,N_3867,N_2880);
or U10632 (N_10632,N_1507,N_6194);
nor U10633 (N_10633,N_5956,N_2383);
and U10634 (N_10634,N_4201,N_388);
or U10635 (N_10635,N_1139,N_712);
or U10636 (N_10636,N_1184,N_3138);
xor U10637 (N_10637,N_1210,N_3593);
or U10638 (N_10638,N_2996,N_2593);
nor U10639 (N_10639,N_1903,N_4173);
and U10640 (N_10640,N_4676,N_2042);
nand U10641 (N_10641,N_1801,N_4641);
nand U10642 (N_10642,N_1971,N_647);
and U10643 (N_10643,N_986,N_2252);
and U10644 (N_10644,N_2259,N_3339);
or U10645 (N_10645,N_1707,N_4628);
nor U10646 (N_10646,N_1495,N_4248);
nor U10647 (N_10647,N_4376,N_2094);
nand U10648 (N_10648,N_1688,N_4629);
or U10649 (N_10649,N_2286,N_417);
xor U10650 (N_10650,N_1996,N_1244);
and U10651 (N_10651,N_5728,N_5385);
and U10652 (N_10652,N_256,N_1131);
and U10653 (N_10653,N_4972,N_1071);
nand U10654 (N_10654,N_634,N_3284);
nand U10655 (N_10655,N_2294,N_5555);
or U10656 (N_10656,N_5075,N_443);
and U10657 (N_10657,N_6031,N_3244);
or U10658 (N_10658,N_2696,N_4918);
nor U10659 (N_10659,N_2316,N_1765);
xnor U10660 (N_10660,N_4672,N_897);
nand U10661 (N_10661,N_2227,N_746);
xor U10662 (N_10662,N_2403,N_1805);
nor U10663 (N_10663,N_355,N_3988);
nand U10664 (N_10664,N_2474,N_1335);
nor U10665 (N_10665,N_4543,N_3883);
or U10666 (N_10666,N_5119,N_1474);
nor U10667 (N_10667,N_2577,N_4674);
xor U10668 (N_10668,N_4293,N_3603);
nand U10669 (N_10669,N_2175,N_3525);
nand U10670 (N_10670,N_2935,N_3748);
nand U10671 (N_10671,N_2498,N_510);
and U10672 (N_10672,N_4174,N_366);
nor U10673 (N_10673,N_2644,N_3745);
and U10674 (N_10674,N_1410,N_5163);
nor U10675 (N_10675,N_1377,N_5842);
nor U10676 (N_10676,N_890,N_5510);
and U10677 (N_10677,N_2366,N_1982);
nand U10678 (N_10678,N_3516,N_832);
xnor U10679 (N_10679,N_2629,N_1318);
nand U10680 (N_10680,N_5314,N_4736);
and U10681 (N_10681,N_6118,N_1591);
xor U10682 (N_10682,N_4360,N_2954);
or U10683 (N_10683,N_5553,N_2279);
or U10684 (N_10684,N_399,N_424);
or U10685 (N_10685,N_3801,N_4244);
nor U10686 (N_10686,N_1783,N_3150);
nand U10687 (N_10687,N_3721,N_4848);
and U10688 (N_10688,N_4377,N_5308);
nand U10689 (N_10689,N_4061,N_820);
xnor U10690 (N_10690,N_2275,N_4954);
xnor U10691 (N_10691,N_864,N_3122);
nand U10692 (N_10692,N_5581,N_1963);
and U10693 (N_10693,N_1050,N_2377);
nand U10694 (N_10694,N_5946,N_1215);
or U10695 (N_10695,N_271,N_1929);
xnor U10696 (N_10696,N_1350,N_3751);
nor U10697 (N_10697,N_3828,N_1055);
or U10698 (N_10698,N_1175,N_5295);
and U10699 (N_10699,N_5951,N_6155);
or U10700 (N_10700,N_2133,N_1901);
xor U10701 (N_10701,N_4739,N_1234);
nand U10702 (N_10702,N_2176,N_5828);
or U10703 (N_10703,N_6247,N_6073);
or U10704 (N_10704,N_6081,N_6016);
nand U10705 (N_10705,N_1031,N_232);
or U10706 (N_10706,N_4988,N_645);
nand U10707 (N_10707,N_3983,N_5045);
nor U10708 (N_10708,N_5132,N_4260);
nor U10709 (N_10709,N_3512,N_3407);
and U10710 (N_10710,N_4100,N_3928);
nand U10711 (N_10711,N_4305,N_756);
xor U10712 (N_10712,N_4345,N_1572);
nor U10713 (N_10713,N_2612,N_1113);
nand U10714 (N_10714,N_1759,N_3921);
nor U10715 (N_10715,N_2008,N_5255);
nor U10716 (N_10716,N_3883,N_2261);
nand U10717 (N_10717,N_3415,N_3551);
and U10718 (N_10718,N_1376,N_2331);
xnor U10719 (N_10719,N_1649,N_3563);
nor U10720 (N_10720,N_2362,N_3196);
nor U10721 (N_10721,N_2527,N_3885);
xor U10722 (N_10722,N_3391,N_3527);
or U10723 (N_10723,N_3697,N_5627);
nand U10724 (N_10724,N_2539,N_1288);
or U10725 (N_10725,N_5506,N_1175);
nand U10726 (N_10726,N_5879,N_158);
nand U10727 (N_10727,N_4159,N_4571);
xnor U10728 (N_10728,N_512,N_5882);
nand U10729 (N_10729,N_4481,N_2078);
and U10730 (N_10730,N_784,N_956);
xnor U10731 (N_10731,N_2793,N_1079);
and U10732 (N_10732,N_904,N_1930);
or U10733 (N_10733,N_799,N_1720);
nor U10734 (N_10734,N_170,N_2951);
and U10735 (N_10735,N_3947,N_5920);
or U10736 (N_10736,N_5088,N_5284);
nor U10737 (N_10737,N_3802,N_4812);
and U10738 (N_10738,N_2102,N_5838);
xor U10739 (N_10739,N_1542,N_3606);
nor U10740 (N_10740,N_3394,N_458);
and U10741 (N_10741,N_3741,N_2177);
and U10742 (N_10742,N_1274,N_1341);
xnor U10743 (N_10743,N_5876,N_2776);
nor U10744 (N_10744,N_4990,N_1087);
or U10745 (N_10745,N_5348,N_4800);
or U10746 (N_10746,N_3173,N_1226);
or U10747 (N_10747,N_4494,N_1021);
nand U10748 (N_10748,N_2404,N_2873);
xnor U10749 (N_10749,N_3238,N_631);
nor U10750 (N_10750,N_1913,N_4478);
nor U10751 (N_10751,N_1528,N_3985);
nor U10752 (N_10752,N_2917,N_1131);
nand U10753 (N_10753,N_5769,N_130);
and U10754 (N_10754,N_1782,N_5204);
nor U10755 (N_10755,N_182,N_4505);
or U10756 (N_10756,N_910,N_3939);
nand U10757 (N_10757,N_916,N_3635);
nand U10758 (N_10758,N_1668,N_4572);
and U10759 (N_10759,N_4522,N_4286);
xor U10760 (N_10760,N_6012,N_1559);
nand U10761 (N_10761,N_5495,N_2402);
xnor U10762 (N_10762,N_2439,N_188);
nand U10763 (N_10763,N_5565,N_1666);
nand U10764 (N_10764,N_5930,N_41);
or U10765 (N_10765,N_164,N_3342);
and U10766 (N_10766,N_4888,N_3683);
nand U10767 (N_10767,N_266,N_496);
xnor U10768 (N_10768,N_1381,N_1001);
or U10769 (N_10769,N_3485,N_978);
or U10770 (N_10770,N_663,N_2877);
xnor U10771 (N_10771,N_2297,N_4505);
and U10772 (N_10772,N_1369,N_41);
and U10773 (N_10773,N_987,N_4557);
nand U10774 (N_10774,N_1537,N_5589);
nor U10775 (N_10775,N_3521,N_5231);
nor U10776 (N_10776,N_4018,N_5396);
and U10777 (N_10777,N_5621,N_1876);
nor U10778 (N_10778,N_756,N_1265);
and U10779 (N_10779,N_3886,N_4476);
nand U10780 (N_10780,N_2971,N_4327);
or U10781 (N_10781,N_1492,N_4360);
xnor U10782 (N_10782,N_3915,N_5411);
or U10783 (N_10783,N_5608,N_5283);
and U10784 (N_10784,N_2723,N_37);
or U10785 (N_10785,N_24,N_2911);
nand U10786 (N_10786,N_5364,N_1043);
xor U10787 (N_10787,N_1643,N_2568);
or U10788 (N_10788,N_909,N_3686);
and U10789 (N_10789,N_1723,N_3957);
nand U10790 (N_10790,N_905,N_3536);
and U10791 (N_10791,N_4798,N_719);
nor U10792 (N_10792,N_4512,N_1398);
and U10793 (N_10793,N_686,N_2345);
nand U10794 (N_10794,N_425,N_302);
and U10795 (N_10795,N_983,N_3889);
xor U10796 (N_10796,N_2620,N_6231);
nor U10797 (N_10797,N_4204,N_2250);
xnor U10798 (N_10798,N_5282,N_3401);
and U10799 (N_10799,N_624,N_212);
xnor U10800 (N_10800,N_4929,N_4304);
nor U10801 (N_10801,N_408,N_4825);
nand U10802 (N_10802,N_1224,N_1019);
or U10803 (N_10803,N_4269,N_5145);
nand U10804 (N_10804,N_3663,N_5296);
nand U10805 (N_10805,N_3728,N_44);
or U10806 (N_10806,N_5325,N_3942);
and U10807 (N_10807,N_4979,N_1003);
nor U10808 (N_10808,N_308,N_4012);
xnor U10809 (N_10809,N_5315,N_3241);
or U10810 (N_10810,N_1471,N_2357);
and U10811 (N_10811,N_2026,N_908);
xor U10812 (N_10812,N_3030,N_2071);
or U10813 (N_10813,N_1160,N_4229);
and U10814 (N_10814,N_235,N_3621);
and U10815 (N_10815,N_5859,N_2592);
or U10816 (N_10816,N_2990,N_3378);
or U10817 (N_10817,N_1973,N_1442);
and U10818 (N_10818,N_4263,N_5293);
or U10819 (N_10819,N_1619,N_3566);
and U10820 (N_10820,N_3379,N_463);
or U10821 (N_10821,N_5420,N_1713);
and U10822 (N_10822,N_4228,N_490);
xor U10823 (N_10823,N_506,N_1177);
nand U10824 (N_10824,N_4080,N_3538);
and U10825 (N_10825,N_4475,N_695);
and U10826 (N_10826,N_5035,N_5890);
nand U10827 (N_10827,N_4160,N_5709);
nand U10828 (N_10828,N_6084,N_2192);
or U10829 (N_10829,N_3372,N_733);
and U10830 (N_10830,N_4770,N_49);
nor U10831 (N_10831,N_4688,N_2275);
xor U10832 (N_10832,N_3908,N_2008);
or U10833 (N_10833,N_2618,N_2548);
xnor U10834 (N_10834,N_5247,N_5457);
or U10835 (N_10835,N_1562,N_6106);
nor U10836 (N_10836,N_661,N_263);
nand U10837 (N_10837,N_5106,N_2430);
xnor U10838 (N_10838,N_1435,N_1482);
or U10839 (N_10839,N_2376,N_4690);
and U10840 (N_10840,N_4793,N_5998);
or U10841 (N_10841,N_3000,N_3502);
and U10842 (N_10842,N_5657,N_3977);
nand U10843 (N_10843,N_667,N_3370);
and U10844 (N_10844,N_1929,N_4861);
and U10845 (N_10845,N_5107,N_4734);
nor U10846 (N_10846,N_4154,N_5864);
or U10847 (N_10847,N_1536,N_1253);
and U10848 (N_10848,N_1265,N_6203);
and U10849 (N_10849,N_838,N_5);
or U10850 (N_10850,N_1103,N_968);
and U10851 (N_10851,N_3141,N_4485);
nand U10852 (N_10852,N_942,N_867);
nor U10853 (N_10853,N_2444,N_3562);
xor U10854 (N_10854,N_3989,N_6013);
nand U10855 (N_10855,N_1285,N_3213);
or U10856 (N_10856,N_2787,N_418);
nand U10857 (N_10857,N_375,N_1935);
or U10858 (N_10858,N_5973,N_1861);
nor U10859 (N_10859,N_4266,N_3105);
xor U10860 (N_10860,N_4297,N_977);
or U10861 (N_10861,N_2501,N_831);
or U10862 (N_10862,N_2431,N_3249);
xor U10863 (N_10863,N_2073,N_2964);
xnor U10864 (N_10864,N_1914,N_2659);
nor U10865 (N_10865,N_5695,N_2190);
nand U10866 (N_10866,N_2342,N_1339);
or U10867 (N_10867,N_1604,N_3572);
xor U10868 (N_10868,N_3803,N_4100);
nand U10869 (N_10869,N_5517,N_5152);
and U10870 (N_10870,N_4939,N_5826);
nand U10871 (N_10871,N_4448,N_782);
nand U10872 (N_10872,N_953,N_1537);
nand U10873 (N_10873,N_5183,N_1619);
xor U10874 (N_10874,N_4858,N_5327);
xnor U10875 (N_10875,N_3460,N_4291);
and U10876 (N_10876,N_3103,N_2704);
nor U10877 (N_10877,N_4544,N_3921);
nand U10878 (N_10878,N_4393,N_43);
or U10879 (N_10879,N_4075,N_3496);
and U10880 (N_10880,N_1135,N_4108);
xor U10881 (N_10881,N_1221,N_287);
nor U10882 (N_10882,N_4495,N_4006);
nand U10883 (N_10883,N_3817,N_5902);
xnor U10884 (N_10884,N_2530,N_5741);
xnor U10885 (N_10885,N_4784,N_2555);
nor U10886 (N_10886,N_2130,N_6099);
nor U10887 (N_10887,N_5434,N_853);
nor U10888 (N_10888,N_2546,N_979);
nand U10889 (N_10889,N_867,N_5745);
xnor U10890 (N_10890,N_5884,N_1646);
xnor U10891 (N_10891,N_2401,N_1137);
xor U10892 (N_10892,N_3611,N_67);
nor U10893 (N_10893,N_5678,N_4988);
nor U10894 (N_10894,N_3405,N_6102);
nor U10895 (N_10895,N_5886,N_5183);
nor U10896 (N_10896,N_4618,N_1140);
xnor U10897 (N_10897,N_3226,N_2387);
or U10898 (N_10898,N_1735,N_5742);
and U10899 (N_10899,N_1294,N_4919);
and U10900 (N_10900,N_3218,N_927);
or U10901 (N_10901,N_4504,N_6077);
nor U10902 (N_10902,N_1952,N_504);
or U10903 (N_10903,N_1301,N_168);
nor U10904 (N_10904,N_2789,N_3388);
xnor U10905 (N_10905,N_4212,N_3008);
or U10906 (N_10906,N_1582,N_2734);
nor U10907 (N_10907,N_4092,N_5121);
nand U10908 (N_10908,N_1472,N_2502);
or U10909 (N_10909,N_4942,N_4830);
or U10910 (N_10910,N_5019,N_1017);
nor U10911 (N_10911,N_5706,N_5207);
and U10912 (N_10912,N_3658,N_2685);
nor U10913 (N_10913,N_1404,N_2325);
xor U10914 (N_10914,N_1869,N_2704);
nand U10915 (N_10915,N_2268,N_4325);
nand U10916 (N_10916,N_6246,N_5122);
or U10917 (N_10917,N_4797,N_3235);
nor U10918 (N_10918,N_5821,N_3569);
nand U10919 (N_10919,N_476,N_5076);
or U10920 (N_10920,N_1559,N_68);
xnor U10921 (N_10921,N_1981,N_2239);
xnor U10922 (N_10922,N_4701,N_5219);
or U10923 (N_10923,N_1116,N_600);
or U10924 (N_10924,N_5516,N_2523);
nand U10925 (N_10925,N_881,N_4455);
nand U10926 (N_10926,N_1353,N_1759);
or U10927 (N_10927,N_774,N_2511);
and U10928 (N_10928,N_5636,N_4905);
nor U10929 (N_10929,N_5806,N_5949);
and U10930 (N_10930,N_2873,N_3819);
nor U10931 (N_10931,N_446,N_5236);
xnor U10932 (N_10932,N_1642,N_4298);
and U10933 (N_10933,N_419,N_735);
or U10934 (N_10934,N_5925,N_2098);
nand U10935 (N_10935,N_3741,N_254);
xor U10936 (N_10936,N_700,N_4863);
nand U10937 (N_10937,N_1074,N_621);
xor U10938 (N_10938,N_3065,N_5794);
nand U10939 (N_10939,N_3718,N_636);
nor U10940 (N_10940,N_2848,N_1898);
xnor U10941 (N_10941,N_944,N_4026);
nand U10942 (N_10942,N_6132,N_3926);
xnor U10943 (N_10943,N_271,N_2049);
nand U10944 (N_10944,N_2361,N_524);
and U10945 (N_10945,N_2440,N_2566);
and U10946 (N_10946,N_65,N_3438);
and U10947 (N_10947,N_337,N_1764);
xnor U10948 (N_10948,N_4347,N_1767);
and U10949 (N_10949,N_3124,N_5713);
and U10950 (N_10950,N_6090,N_4521);
nand U10951 (N_10951,N_4827,N_96);
nand U10952 (N_10952,N_4440,N_742);
nor U10953 (N_10953,N_216,N_3673);
and U10954 (N_10954,N_4418,N_5215);
xnor U10955 (N_10955,N_2632,N_5617);
nor U10956 (N_10956,N_2323,N_5146);
nand U10957 (N_10957,N_3946,N_105);
nand U10958 (N_10958,N_1332,N_3531);
or U10959 (N_10959,N_98,N_6211);
nor U10960 (N_10960,N_2208,N_5866);
or U10961 (N_10961,N_1938,N_758);
or U10962 (N_10962,N_114,N_2589);
nand U10963 (N_10963,N_5381,N_5639);
and U10964 (N_10964,N_5811,N_3214);
nand U10965 (N_10965,N_5032,N_5732);
nor U10966 (N_10966,N_3905,N_3217);
xnor U10967 (N_10967,N_3327,N_3853);
xor U10968 (N_10968,N_691,N_4532);
or U10969 (N_10969,N_566,N_3856);
and U10970 (N_10970,N_583,N_3279);
or U10971 (N_10971,N_6100,N_4661);
nor U10972 (N_10972,N_4683,N_3891);
xor U10973 (N_10973,N_5813,N_4066);
xor U10974 (N_10974,N_5565,N_3425);
nor U10975 (N_10975,N_5591,N_5621);
xor U10976 (N_10976,N_3734,N_2013);
nor U10977 (N_10977,N_1360,N_2192);
or U10978 (N_10978,N_3251,N_1753);
or U10979 (N_10979,N_2749,N_4605);
or U10980 (N_10980,N_3219,N_1955);
nand U10981 (N_10981,N_1604,N_6205);
and U10982 (N_10982,N_5783,N_5320);
nand U10983 (N_10983,N_1673,N_5190);
or U10984 (N_10984,N_1605,N_4676);
and U10985 (N_10985,N_3434,N_4291);
nor U10986 (N_10986,N_750,N_133);
or U10987 (N_10987,N_1236,N_6067);
nand U10988 (N_10988,N_1595,N_853);
nand U10989 (N_10989,N_398,N_1948);
and U10990 (N_10990,N_5253,N_9);
xnor U10991 (N_10991,N_1605,N_91);
nor U10992 (N_10992,N_5500,N_5957);
nand U10993 (N_10993,N_5970,N_5988);
xor U10994 (N_10994,N_285,N_4112);
nand U10995 (N_10995,N_3313,N_1216);
nand U10996 (N_10996,N_468,N_2509);
nor U10997 (N_10997,N_4983,N_1270);
nor U10998 (N_10998,N_3521,N_4556);
and U10999 (N_10999,N_3739,N_332);
and U11000 (N_11000,N_2285,N_5656);
and U11001 (N_11001,N_2814,N_3366);
or U11002 (N_11002,N_3502,N_804);
xnor U11003 (N_11003,N_2404,N_1789);
and U11004 (N_11004,N_4382,N_2454);
nor U11005 (N_11005,N_5537,N_2219);
or U11006 (N_11006,N_1799,N_5554);
and U11007 (N_11007,N_277,N_1785);
xnor U11008 (N_11008,N_3558,N_5217);
nand U11009 (N_11009,N_1009,N_2064);
nand U11010 (N_11010,N_5705,N_5974);
nor U11011 (N_11011,N_2954,N_5390);
nor U11012 (N_11012,N_5548,N_4955);
or U11013 (N_11013,N_5915,N_2719);
xor U11014 (N_11014,N_4769,N_6197);
and U11015 (N_11015,N_2772,N_2508);
nand U11016 (N_11016,N_3824,N_5281);
and U11017 (N_11017,N_5573,N_5986);
nand U11018 (N_11018,N_312,N_3696);
nor U11019 (N_11019,N_68,N_5150);
and U11020 (N_11020,N_1607,N_5808);
nor U11021 (N_11021,N_700,N_5702);
nor U11022 (N_11022,N_387,N_3582);
nand U11023 (N_11023,N_1114,N_4799);
nor U11024 (N_11024,N_4101,N_1603);
xnor U11025 (N_11025,N_736,N_977);
nor U11026 (N_11026,N_3503,N_1005);
and U11027 (N_11027,N_2948,N_3620);
nand U11028 (N_11028,N_551,N_3570);
and U11029 (N_11029,N_3135,N_2025);
nor U11030 (N_11030,N_5254,N_3699);
or U11031 (N_11031,N_1549,N_2659);
or U11032 (N_11032,N_3701,N_4714);
and U11033 (N_11033,N_2639,N_4340);
nor U11034 (N_11034,N_5680,N_3432);
xnor U11035 (N_11035,N_1837,N_854);
or U11036 (N_11036,N_3315,N_1947);
xor U11037 (N_11037,N_1564,N_3214);
and U11038 (N_11038,N_1517,N_1962);
and U11039 (N_11039,N_5924,N_3653);
nand U11040 (N_11040,N_2591,N_111);
xor U11041 (N_11041,N_5526,N_4251);
or U11042 (N_11042,N_14,N_4035);
xor U11043 (N_11043,N_3517,N_1503);
and U11044 (N_11044,N_1427,N_3770);
xor U11045 (N_11045,N_2736,N_6139);
nand U11046 (N_11046,N_6223,N_6033);
xor U11047 (N_11047,N_4102,N_908);
nand U11048 (N_11048,N_1519,N_4260);
or U11049 (N_11049,N_4065,N_76);
xnor U11050 (N_11050,N_4293,N_3165);
nand U11051 (N_11051,N_1466,N_111);
and U11052 (N_11052,N_2347,N_2819);
nor U11053 (N_11053,N_4058,N_4672);
or U11054 (N_11054,N_5010,N_3460);
xnor U11055 (N_11055,N_2643,N_5312);
xnor U11056 (N_11056,N_2088,N_4652);
or U11057 (N_11057,N_4643,N_4043);
xor U11058 (N_11058,N_3259,N_1934);
nor U11059 (N_11059,N_469,N_3425);
nand U11060 (N_11060,N_5448,N_3851);
or U11061 (N_11061,N_2484,N_2483);
or U11062 (N_11062,N_2256,N_5734);
nor U11063 (N_11063,N_5125,N_4528);
nor U11064 (N_11064,N_4380,N_4855);
xnor U11065 (N_11065,N_5961,N_1109);
nand U11066 (N_11066,N_981,N_2553);
xnor U11067 (N_11067,N_167,N_5346);
nand U11068 (N_11068,N_3526,N_3848);
and U11069 (N_11069,N_1904,N_2096);
nand U11070 (N_11070,N_1753,N_25);
and U11071 (N_11071,N_338,N_5266);
or U11072 (N_11072,N_6151,N_5857);
and U11073 (N_11073,N_5201,N_1881);
or U11074 (N_11074,N_5841,N_5452);
or U11075 (N_11075,N_106,N_2510);
nor U11076 (N_11076,N_1652,N_3667);
xor U11077 (N_11077,N_1228,N_346);
nand U11078 (N_11078,N_5876,N_1616);
nand U11079 (N_11079,N_5135,N_4936);
xnor U11080 (N_11080,N_2259,N_5881);
xor U11081 (N_11081,N_4078,N_1998);
and U11082 (N_11082,N_620,N_6153);
and U11083 (N_11083,N_2680,N_3843);
nor U11084 (N_11084,N_904,N_4696);
nor U11085 (N_11085,N_5124,N_1992);
or U11086 (N_11086,N_826,N_3331);
nor U11087 (N_11087,N_954,N_5513);
nand U11088 (N_11088,N_855,N_5772);
and U11089 (N_11089,N_4555,N_5083);
nand U11090 (N_11090,N_5385,N_585);
and U11091 (N_11091,N_5583,N_3944);
nand U11092 (N_11092,N_5921,N_658);
xor U11093 (N_11093,N_2646,N_3275);
or U11094 (N_11094,N_5717,N_3749);
and U11095 (N_11095,N_4532,N_694);
or U11096 (N_11096,N_3380,N_5917);
xnor U11097 (N_11097,N_3200,N_4052);
and U11098 (N_11098,N_1060,N_5405);
xnor U11099 (N_11099,N_4678,N_5481);
and U11100 (N_11100,N_1842,N_2740);
and U11101 (N_11101,N_1961,N_3016);
nand U11102 (N_11102,N_3017,N_4402);
nor U11103 (N_11103,N_2395,N_329);
and U11104 (N_11104,N_646,N_4484);
nor U11105 (N_11105,N_1921,N_5983);
or U11106 (N_11106,N_1836,N_2166);
nand U11107 (N_11107,N_503,N_3866);
or U11108 (N_11108,N_3854,N_6079);
or U11109 (N_11109,N_16,N_227);
xor U11110 (N_11110,N_1593,N_4815);
or U11111 (N_11111,N_5642,N_1662);
nor U11112 (N_11112,N_1884,N_828);
or U11113 (N_11113,N_2293,N_1653);
xnor U11114 (N_11114,N_3082,N_5394);
or U11115 (N_11115,N_4267,N_5525);
and U11116 (N_11116,N_2812,N_3355);
and U11117 (N_11117,N_1646,N_6210);
nor U11118 (N_11118,N_216,N_4540);
or U11119 (N_11119,N_3845,N_1476);
and U11120 (N_11120,N_590,N_4218);
or U11121 (N_11121,N_5380,N_3683);
nand U11122 (N_11122,N_1037,N_5208);
xnor U11123 (N_11123,N_4469,N_3883);
and U11124 (N_11124,N_5745,N_5647);
xor U11125 (N_11125,N_654,N_4519);
nor U11126 (N_11126,N_6111,N_2504);
or U11127 (N_11127,N_1585,N_1968);
nand U11128 (N_11128,N_4927,N_913);
nand U11129 (N_11129,N_1611,N_3774);
xor U11130 (N_11130,N_5341,N_3848);
nand U11131 (N_11131,N_5918,N_443);
nand U11132 (N_11132,N_693,N_1184);
and U11133 (N_11133,N_2061,N_5627);
xor U11134 (N_11134,N_4239,N_6016);
xnor U11135 (N_11135,N_3845,N_6158);
xor U11136 (N_11136,N_3669,N_3827);
xor U11137 (N_11137,N_546,N_5887);
or U11138 (N_11138,N_1546,N_1416);
and U11139 (N_11139,N_5815,N_5454);
or U11140 (N_11140,N_316,N_963);
or U11141 (N_11141,N_4269,N_6194);
and U11142 (N_11142,N_5544,N_1562);
nor U11143 (N_11143,N_1445,N_2346);
or U11144 (N_11144,N_4038,N_6057);
nand U11145 (N_11145,N_2335,N_4125);
xor U11146 (N_11146,N_3003,N_704);
nand U11147 (N_11147,N_5154,N_3122);
nand U11148 (N_11148,N_4846,N_3656);
or U11149 (N_11149,N_4680,N_238);
xor U11150 (N_11150,N_2454,N_1060);
or U11151 (N_11151,N_3491,N_4854);
or U11152 (N_11152,N_4801,N_4724);
nor U11153 (N_11153,N_3303,N_5710);
or U11154 (N_11154,N_2908,N_3894);
nor U11155 (N_11155,N_4354,N_6013);
nor U11156 (N_11156,N_2559,N_51);
xnor U11157 (N_11157,N_264,N_5909);
and U11158 (N_11158,N_4596,N_2715);
nor U11159 (N_11159,N_2899,N_904);
xnor U11160 (N_11160,N_4061,N_5203);
xnor U11161 (N_11161,N_5967,N_1679);
nor U11162 (N_11162,N_5987,N_4221);
xor U11163 (N_11163,N_3836,N_5568);
or U11164 (N_11164,N_1281,N_1619);
xnor U11165 (N_11165,N_4422,N_5226);
xor U11166 (N_11166,N_4159,N_4381);
xnor U11167 (N_11167,N_2494,N_4017);
xnor U11168 (N_11168,N_4957,N_4182);
nor U11169 (N_11169,N_4640,N_76);
and U11170 (N_11170,N_5010,N_202);
nand U11171 (N_11171,N_5909,N_4192);
or U11172 (N_11172,N_3958,N_1325);
and U11173 (N_11173,N_3839,N_5937);
nor U11174 (N_11174,N_695,N_4704);
nor U11175 (N_11175,N_5729,N_1831);
nor U11176 (N_11176,N_1517,N_320);
xnor U11177 (N_11177,N_2813,N_2544);
xnor U11178 (N_11178,N_1832,N_5365);
nor U11179 (N_11179,N_6223,N_2588);
and U11180 (N_11180,N_3477,N_3000);
nand U11181 (N_11181,N_3192,N_4075);
and U11182 (N_11182,N_445,N_268);
xnor U11183 (N_11183,N_171,N_1758);
xnor U11184 (N_11184,N_5050,N_3258);
xnor U11185 (N_11185,N_4181,N_3699);
and U11186 (N_11186,N_4656,N_5087);
xnor U11187 (N_11187,N_5925,N_4158);
and U11188 (N_11188,N_4278,N_3833);
or U11189 (N_11189,N_3315,N_5804);
nor U11190 (N_11190,N_2345,N_4526);
or U11191 (N_11191,N_2221,N_1190);
xor U11192 (N_11192,N_3172,N_5850);
and U11193 (N_11193,N_3392,N_5636);
and U11194 (N_11194,N_1629,N_260);
nor U11195 (N_11195,N_2547,N_5344);
xnor U11196 (N_11196,N_913,N_1243);
nand U11197 (N_11197,N_382,N_3229);
nor U11198 (N_11198,N_528,N_1374);
or U11199 (N_11199,N_4751,N_2833);
xor U11200 (N_11200,N_5492,N_4683);
nand U11201 (N_11201,N_5968,N_5967);
and U11202 (N_11202,N_5051,N_3294);
and U11203 (N_11203,N_4329,N_2110);
nand U11204 (N_11204,N_1753,N_2152);
and U11205 (N_11205,N_5722,N_2928);
or U11206 (N_11206,N_6,N_2621);
and U11207 (N_11207,N_354,N_3378);
xnor U11208 (N_11208,N_4369,N_2710);
and U11209 (N_11209,N_2029,N_2447);
xor U11210 (N_11210,N_3410,N_1589);
xor U11211 (N_11211,N_2321,N_6155);
nor U11212 (N_11212,N_4310,N_607);
xor U11213 (N_11213,N_4698,N_4566);
nand U11214 (N_11214,N_1672,N_4269);
nor U11215 (N_11215,N_5627,N_684);
nor U11216 (N_11216,N_979,N_2843);
xor U11217 (N_11217,N_5909,N_1102);
xor U11218 (N_11218,N_4159,N_5908);
or U11219 (N_11219,N_3678,N_964);
or U11220 (N_11220,N_6140,N_4722);
nor U11221 (N_11221,N_5263,N_3922);
and U11222 (N_11222,N_6220,N_676);
and U11223 (N_11223,N_4835,N_2086);
nor U11224 (N_11224,N_4972,N_3014);
or U11225 (N_11225,N_4128,N_5009);
and U11226 (N_11226,N_4979,N_5268);
and U11227 (N_11227,N_1774,N_5940);
xnor U11228 (N_11228,N_3189,N_1626);
nand U11229 (N_11229,N_515,N_6176);
xnor U11230 (N_11230,N_1409,N_5315);
nor U11231 (N_11231,N_3055,N_5424);
or U11232 (N_11232,N_6133,N_1157);
and U11233 (N_11233,N_597,N_2787);
nand U11234 (N_11234,N_5220,N_1414);
nor U11235 (N_11235,N_975,N_3693);
nand U11236 (N_11236,N_5200,N_5988);
xnor U11237 (N_11237,N_1200,N_5903);
nor U11238 (N_11238,N_6101,N_844);
xor U11239 (N_11239,N_6137,N_1908);
or U11240 (N_11240,N_4980,N_626);
xnor U11241 (N_11241,N_480,N_5249);
nand U11242 (N_11242,N_1552,N_5543);
nor U11243 (N_11243,N_2625,N_3095);
or U11244 (N_11244,N_2177,N_607);
nand U11245 (N_11245,N_4549,N_4314);
nand U11246 (N_11246,N_6114,N_4270);
or U11247 (N_11247,N_1433,N_3365);
xor U11248 (N_11248,N_2155,N_4670);
or U11249 (N_11249,N_2032,N_2928);
nor U11250 (N_11250,N_2105,N_1605);
and U11251 (N_11251,N_3149,N_5326);
nand U11252 (N_11252,N_5754,N_5727);
nand U11253 (N_11253,N_3784,N_3155);
and U11254 (N_11254,N_3509,N_5094);
nor U11255 (N_11255,N_5459,N_412);
or U11256 (N_11256,N_2287,N_597);
nor U11257 (N_11257,N_2322,N_1990);
xnor U11258 (N_11258,N_3951,N_337);
and U11259 (N_11259,N_3216,N_664);
and U11260 (N_11260,N_714,N_5144);
nor U11261 (N_11261,N_2789,N_1864);
and U11262 (N_11262,N_5702,N_5090);
xor U11263 (N_11263,N_1601,N_3681);
and U11264 (N_11264,N_232,N_6235);
or U11265 (N_11265,N_884,N_2229);
and U11266 (N_11266,N_2873,N_1175);
and U11267 (N_11267,N_2093,N_4158);
nand U11268 (N_11268,N_4124,N_2912);
and U11269 (N_11269,N_4185,N_2581);
nand U11270 (N_11270,N_6149,N_3012);
nand U11271 (N_11271,N_178,N_5666);
xor U11272 (N_11272,N_5679,N_1145);
nor U11273 (N_11273,N_3191,N_1220);
nand U11274 (N_11274,N_1910,N_1720);
and U11275 (N_11275,N_4816,N_157);
xor U11276 (N_11276,N_4463,N_6033);
nand U11277 (N_11277,N_5818,N_6074);
nand U11278 (N_11278,N_2124,N_4479);
xor U11279 (N_11279,N_4133,N_3835);
nand U11280 (N_11280,N_2868,N_4830);
xor U11281 (N_11281,N_4659,N_2746);
or U11282 (N_11282,N_1439,N_2507);
or U11283 (N_11283,N_1152,N_116);
or U11284 (N_11284,N_5767,N_4710);
nand U11285 (N_11285,N_2573,N_696);
and U11286 (N_11286,N_2307,N_1521);
and U11287 (N_11287,N_6246,N_2399);
nor U11288 (N_11288,N_5965,N_2518);
xnor U11289 (N_11289,N_5918,N_2661);
nand U11290 (N_11290,N_854,N_4589);
nor U11291 (N_11291,N_3863,N_310);
or U11292 (N_11292,N_314,N_4585);
nand U11293 (N_11293,N_4866,N_1866);
nand U11294 (N_11294,N_4276,N_2016);
or U11295 (N_11295,N_5441,N_4652);
and U11296 (N_11296,N_1523,N_5480);
xnor U11297 (N_11297,N_2003,N_2132);
nor U11298 (N_11298,N_5925,N_3728);
nor U11299 (N_11299,N_1377,N_2449);
nor U11300 (N_11300,N_6148,N_1448);
nor U11301 (N_11301,N_5102,N_4124);
nor U11302 (N_11302,N_5233,N_3017);
or U11303 (N_11303,N_1432,N_6214);
nor U11304 (N_11304,N_3219,N_3139);
xor U11305 (N_11305,N_1363,N_5675);
nor U11306 (N_11306,N_3328,N_2668);
nand U11307 (N_11307,N_5481,N_2291);
and U11308 (N_11308,N_6076,N_1171);
xnor U11309 (N_11309,N_5753,N_1017);
xor U11310 (N_11310,N_2558,N_3994);
or U11311 (N_11311,N_1567,N_5836);
nor U11312 (N_11312,N_5913,N_468);
nor U11313 (N_11313,N_4785,N_6096);
xor U11314 (N_11314,N_4743,N_3534);
or U11315 (N_11315,N_2851,N_6214);
and U11316 (N_11316,N_5625,N_4702);
or U11317 (N_11317,N_4851,N_5414);
nand U11318 (N_11318,N_2366,N_3709);
nand U11319 (N_11319,N_5572,N_701);
and U11320 (N_11320,N_4663,N_6019);
nor U11321 (N_11321,N_5667,N_5652);
xnor U11322 (N_11322,N_418,N_341);
xor U11323 (N_11323,N_1288,N_1648);
xor U11324 (N_11324,N_4900,N_2816);
and U11325 (N_11325,N_2632,N_1358);
or U11326 (N_11326,N_2652,N_3563);
nand U11327 (N_11327,N_2232,N_3585);
nand U11328 (N_11328,N_2310,N_2433);
or U11329 (N_11329,N_2849,N_2373);
and U11330 (N_11330,N_4110,N_538);
nand U11331 (N_11331,N_1903,N_1178);
and U11332 (N_11332,N_4389,N_4056);
xnor U11333 (N_11333,N_5079,N_5035);
nor U11334 (N_11334,N_6015,N_954);
or U11335 (N_11335,N_139,N_4876);
nand U11336 (N_11336,N_282,N_1438);
xor U11337 (N_11337,N_43,N_5004);
or U11338 (N_11338,N_3891,N_5382);
xnor U11339 (N_11339,N_1708,N_6159);
nand U11340 (N_11340,N_2689,N_5307);
or U11341 (N_11341,N_4757,N_4175);
and U11342 (N_11342,N_4123,N_3941);
and U11343 (N_11343,N_6205,N_1669);
and U11344 (N_11344,N_449,N_3352);
nor U11345 (N_11345,N_455,N_6053);
xor U11346 (N_11346,N_4951,N_709);
or U11347 (N_11347,N_4415,N_2743);
xor U11348 (N_11348,N_1860,N_3209);
nor U11349 (N_11349,N_810,N_985);
nor U11350 (N_11350,N_6170,N_2460);
and U11351 (N_11351,N_1940,N_3533);
nor U11352 (N_11352,N_1978,N_4562);
or U11353 (N_11353,N_4041,N_2828);
nor U11354 (N_11354,N_5191,N_4953);
nand U11355 (N_11355,N_6175,N_780);
and U11356 (N_11356,N_212,N_4411);
nor U11357 (N_11357,N_5240,N_1901);
and U11358 (N_11358,N_4292,N_953);
xor U11359 (N_11359,N_3993,N_1625);
or U11360 (N_11360,N_224,N_5250);
and U11361 (N_11361,N_1860,N_3288);
nand U11362 (N_11362,N_1199,N_5969);
nand U11363 (N_11363,N_4094,N_4280);
nor U11364 (N_11364,N_1056,N_4203);
nand U11365 (N_11365,N_3660,N_5888);
nor U11366 (N_11366,N_3361,N_4474);
or U11367 (N_11367,N_5928,N_655);
xnor U11368 (N_11368,N_6007,N_5683);
nor U11369 (N_11369,N_5966,N_2194);
nand U11370 (N_11370,N_5794,N_523);
nand U11371 (N_11371,N_2829,N_4977);
nor U11372 (N_11372,N_4667,N_2383);
xnor U11373 (N_11373,N_5134,N_5769);
xnor U11374 (N_11374,N_3175,N_3285);
and U11375 (N_11375,N_5344,N_4254);
nand U11376 (N_11376,N_3781,N_5373);
nand U11377 (N_11377,N_1311,N_2404);
or U11378 (N_11378,N_3698,N_3213);
nor U11379 (N_11379,N_1009,N_4854);
and U11380 (N_11380,N_497,N_5965);
xnor U11381 (N_11381,N_392,N_1913);
or U11382 (N_11382,N_3286,N_5220);
nand U11383 (N_11383,N_4771,N_1757);
and U11384 (N_11384,N_3101,N_5490);
nand U11385 (N_11385,N_1460,N_1308);
xnor U11386 (N_11386,N_3595,N_2461);
and U11387 (N_11387,N_3609,N_4618);
nor U11388 (N_11388,N_5528,N_4742);
nand U11389 (N_11389,N_4884,N_2416);
and U11390 (N_11390,N_1705,N_6082);
nor U11391 (N_11391,N_4599,N_3554);
nand U11392 (N_11392,N_4326,N_4932);
nand U11393 (N_11393,N_751,N_5929);
nand U11394 (N_11394,N_5836,N_3191);
or U11395 (N_11395,N_5720,N_541);
or U11396 (N_11396,N_5550,N_4551);
xor U11397 (N_11397,N_3716,N_4381);
and U11398 (N_11398,N_4865,N_1364);
nand U11399 (N_11399,N_4976,N_77);
and U11400 (N_11400,N_5328,N_3408);
xor U11401 (N_11401,N_5555,N_1818);
or U11402 (N_11402,N_2434,N_4117);
nand U11403 (N_11403,N_1250,N_629);
xnor U11404 (N_11404,N_525,N_4886);
xor U11405 (N_11405,N_3462,N_3121);
or U11406 (N_11406,N_3912,N_3491);
nor U11407 (N_11407,N_4705,N_1341);
or U11408 (N_11408,N_5464,N_3866);
or U11409 (N_11409,N_2493,N_1061);
nor U11410 (N_11410,N_5672,N_5924);
xor U11411 (N_11411,N_2297,N_2341);
xor U11412 (N_11412,N_1280,N_42);
and U11413 (N_11413,N_4992,N_2221);
nor U11414 (N_11414,N_1686,N_3797);
xnor U11415 (N_11415,N_944,N_4135);
or U11416 (N_11416,N_6219,N_3484);
or U11417 (N_11417,N_1038,N_2685);
xor U11418 (N_11418,N_3397,N_1916);
and U11419 (N_11419,N_923,N_1341);
nand U11420 (N_11420,N_2767,N_4749);
or U11421 (N_11421,N_4449,N_3959);
and U11422 (N_11422,N_4613,N_5429);
nand U11423 (N_11423,N_2512,N_4338);
xnor U11424 (N_11424,N_4076,N_688);
and U11425 (N_11425,N_3580,N_295);
or U11426 (N_11426,N_5938,N_783);
nor U11427 (N_11427,N_2045,N_2312);
nand U11428 (N_11428,N_2773,N_5730);
nor U11429 (N_11429,N_2890,N_2352);
nand U11430 (N_11430,N_6100,N_4569);
nor U11431 (N_11431,N_1285,N_2129);
nand U11432 (N_11432,N_2198,N_2395);
xor U11433 (N_11433,N_4483,N_2306);
nand U11434 (N_11434,N_665,N_28);
nor U11435 (N_11435,N_1756,N_3012);
nand U11436 (N_11436,N_5147,N_811);
nand U11437 (N_11437,N_169,N_3907);
xnor U11438 (N_11438,N_1410,N_3955);
xor U11439 (N_11439,N_3482,N_4457);
and U11440 (N_11440,N_5602,N_3346);
nand U11441 (N_11441,N_235,N_2181);
xnor U11442 (N_11442,N_4977,N_3000);
nand U11443 (N_11443,N_6139,N_3849);
nand U11444 (N_11444,N_2929,N_3203);
nor U11445 (N_11445,N_5953,N_2140);
nor U11446 (N_11446,N_36,N_2878);
nor U11447 (N_11447,N_2420,N_5734);
or U11448 (N_11448,N_1818,N_534);
xnor U11449 (N_11449,N_166,N_361);
nand U11450 (N_11450,N_402,N_3572);
nor U11451 (N_11451,N_1402,N_5849);
and U11452 (N_11452,N_4499,N_5158);
and U11453 (N_11453,N_2345,N_4023);
or U11454 (N_11454,N_5324,N_1031);
or U11455 (N_11455,N_4959,N_2619);
nor U11456 (N_11456,N_2756,N_406);
or U11457 (N_11457,N_4783,N_2042);
or U11458 (N_11458,N_5132,N_5112);
and U11459 (N_11459,N_4249,N_2427);
xnor U11460 (N_11460,N_4454,N_3511);
or U11461 (N_11461,N_3683,N_4195);
or U11462 (N_11462,N_3140,N_4391);
nand U11463 (N_11463,N_4495,N_2244);
nand U11464 (N_11464,N_4676,N_1189);
nor U11465 (N_11465,N_1610,N_776);
or U11466 (N_11466,N_540,N_3732);
nor U11467 (N_11467,N_5980,N_2541);
nor U11468 (N_11468,N_3432,N_5348);
xor U11469 (N_11469,N_5501,N_2379);
xnor U11470 (N_11470,N_4136,N_4119);
or U11471 (N_11471,N_790,N_5123);
or U11472 (N_11472,N_2973,N_3586);
nor U11473 (N_11473,N_1015,N_3241);
or U11474 (N_11474,N_1747,N_6171);
nor U11475 (N_11475,N_1688,N_2883);
or U11476 (N_11476,N_3308,N_3722);
and U11477 (N_11477,N_690,N_1100);
nor U11478 (N_11478,N_1263,N_138);
nand U11479 (N_11479,N_253,N_4506);
xnor U11480 (N_11480,N_2146,N_1404);
and U11481 (N_11481,N_2433,N_245);
nand U11482 (N_11482,N_525,N_1532);
nor U11483 (N_11483,N_2022,N_1624);
and U11484 (N_11484,N_6197,N_1510);
nand U11485 (N_11485,N_5723,N_2045);
nor U11486 (N_11486,N_5886,N_164);
nand U11487 (N_11487,N_1696,N_2281);
nor U11488 (N_11488,N_3930,N_878);
nor U11489 (N_11489,N_2516,N_2429);
or U11490 (N_11490,N_5193,N_5956);
nand U11491 (N_11491,N_4853,N_647);
or U11492 (N_11492,N_213,N_5167);
nand U11493 (N_11493,N_2793,N_1590);
nand U11494 (N_11494,N_520,N_5942);
nor U11495 (N_11495,N_757,N_2551);
and U11496 (N_11496,N_3230,N_5197);
nor U11497 (N_11497,N_5747,N_5911);
nor U11498 (N_11498,N_377,N_3311);
nor U11499 (N_11499,N_5694,N_5206);
or U11500 (N_11500,N_5789,N_13);
and U11501 (N_11501,N_5213,N_5162);
nor U11502 (N_11502,N_2047,N_3585);
and U11503 (N_11503,N_4825,N_5476);
or U11504 (N_11504,N_3,N_645);
nand U11505 (N_11505,N_3560,N_1409);
xor U11506 (N_11506,N_5089,N_1412);
and U11507 (N_11507,N_2240,N_5241);
and U11508 (N_11508,N_340,N_2595);
xnor U11509 (N_11509,N_1708,N_2673);
or U11510 (N_11510,N_2217,N_3755);
xnor U11511 (N_11511,N_1012,N_3800);
or U11512 (N_11512,N_1365,N_5037);
xnor U11513 (N_11513,N_1178,N_5766);
nor U11514 (N_11514,N_2266,N_4699);
nand U11515 (N_11515,N_5813,N_1188);
nand U11516 (N_11516,N_4443,N_2376);
nand U11517 (N_11517,N_2096,N_6157);
nand U11518 (N_11518,N_4993,N_3427);
nand U11519 (N_11519,N_4913,N_3087);
xnor U11520 (N_11520,N_525,N_5769);
nor U11521 (N_11521,N_4750,N_4725);
nor U11522 (N_11522,N_4660,N_820);
and U11523 (N_11523,N_3928,N_2968);
and U11524 (N_11524,N_1087,N_5839);
nand U11525 (N_11525,N_141,N_2968);
xor U11526 (N_11526,N_943,N_2246);
nand U11527 (N_11527,N_5213,N_464);
xor U11528 (N_11528,N_1590,N_987);
and U11529 (N_11529,N_4831,N_6140);
nand U11530 (N_11530,N_5737,N_552);
nand U11531 (N_11531,N_4954,N_3236);
and U11532 (N_11532,N_633,N_5595);
nand U11533 (N_11533,N_215,N_5174);
nor U11534 (N_11534,N_1230,N_676);
nor U11535 (N_11535,N_5936,N_145);
and U11536 (N_11536,N_4260,N_2947);
nand U11537 (N_11537,N_1971,N_5293);
nor U11538 (N_11538,N_1721,N_2827);
or U11539 (N_11539,N_3973,N_2928);
nand U11540 (N_11540,N_6242,N_4094);
or U11541 (N_11541,N_2607,N_1372);
xor U11542 (N_11542,N_2647,N_5514);
or U11543 (N_11543,N_4981,N_3358);
nor U11544 (N_11544,N_397,N_104);
and U11545 (N_11545,N_95,N_5043);
or U11546 (N_11546,N_3554,N_1664);
xor U11547 (N_11547,N_778,N_2111);
nand U11548 (N_11548,N_2997,N_1172);
xor U11549 (N_11549,N_3451,N_4086);
nor U11550 (N_11550,N_1967,N_1738);
xnor U11551 (N_11551,N_654,N_5952);
or U11552 (N_11552,N_4712,N_1043);
nand U11553 (N_11553,N_3562,N_3937);
nor U11554 (N_11554,N_4631,N_3695);
and U11555 (N_11555,N_4515,N_4288);
nand U11556 (N_11556,N_5659,N_5045);
and U11557 (N_11557,N_131,N_2190);
or U11558 (N_11558,N_5375,N_3917);
nand U11559 (N_11559,N_4596,N_3012);
nor U11560 (N_11560,N_5747,N_1412);
or U11561 (N_11561,N_4847,N_178);
xnor U11562 (N_11562,N_5246,N_3583);
xor U11563 (N_11563,N_1582,N_2114);
or U11564 (N_11564,N_3178,N_248);
nand U11565 (N_11565,N_4038,N_2337);
nor U11566 (N_11566,N_4849,N_6103);
nand U11567 (N_11567,N_2974,N_6060);
nor U11568 (N_11568,N_676,N_1871);
nand U11569 (N_11569,N_3285,N_1990);
xnor U11570 (N_11570,N_4338,N_538);
nor U11571 (N_11571,N_456,N_1067);
xnor U11572 (N_11572,N_1820,N_5713);
or U11573 (N_11573,N_3210,N_3535);
and U11574 (N_11574,N_3538,N_6149);
xor U11575 (N_11575,N_5481,N_899);
nor U11576 (N_11576,N_4288,N_3995);
nand U11577 (N_11577,N_3752,N_67);
and U11578 (N_11578,N_4662,N_1520);
nand U11579 (N_11579,N_1008,N_2644);
nor U11580 (N_11580,N_6005,N_3838);
xor U11581 (N_11581,N_5384,N_586);
and U11582 (N_11582,N_1413,N_2946);
xnor U11583 (N_11583,N_1820,N_2041);
nor U11584 (N_11584,N_556,N_3745);
nand U11585 (N_11585,N_5367,N_54);
nor U11586 (N_11586,N_2076,N_4592);
nor U11587 (N_11587,N_1161,N_4121);
and U11588 (N_11588,N_2540,N_1453);
nor U11589 (N_11589,N_3007,N_1081);
or U11590 (N_11590,N_2128,N_3407);
or U11591 (N_11591,N_2130,N_2604);
xor U11592 (N_11592,N_3706,N_5112);
nand U11593 (N_11593,N_5102,N_187);
xor U11594 (N_11594,N_3973,N_4452);
xor U11595 (N_11595,N_3173,N_3599);
nand U11596 (N_11596,N_4270,N_803);
nor U11597 (N_11597,N_3855,N_3129);
nor U11598 (N_11598,N_5055,N_2737);
xnor U11599 (N_11599,N_2068,N_513);
and U11600 (N_11600,N_5487,N_5992);
xnor U11601 (N_11601,N_2736,N_1797);
xor U11602 (N_11602,N_5522,N_4896);
nor U11603 (N_11603,N_6243,N_5580);
xor U11604 (N_11604,N_672,N_2687);
or U11605 (N_11605,N_2179,N_2071);
nor U11606 (N_11606,N_3508,N_6211);
and U11607 (N_11607,N_5141,N_3465);
nor U11608 (N_11608,N_4556,N_2643);
nand U11609 (N_11609,N_711,N_5037);
nand U11610 (N_11610,N_1036,N_3274);
nand U11611 (N_11611,N_4517,N_5986);
xor U11612 (N_11612,N_4798,N_3646);
and U11613 (N_11613,N_1407,N_3503);
nand U11614 (N_11614,N_23,N_1986);
nor U11615 (N_11615,N_3543,N_3568);
nor U11616 (N_11616,N_5342,N_4648);
or U11617 (N_11617,N_4737,N_1636);
nor U11618 (N_11618,N_1833,N_3453);
nand U11619 (N_11619,N_2254,N_4365);
xor U11620 (N_11620,N_5011,N_165);
xnor U11621 (N_11621,N_1679,N_5425);
and U11622 (N_11622,N_906,N_170);
nand U11623 (N_11623,N_4646,N_6050);
xor U11624 (N_11624,N_1613,N_5093);
xnor U11625 (N_11625,N_3112,N_3003);
nor U11626 (N_11626,N_1482,N_5647);
or U11627 (N_11627,N_951,N_1229);
xnor U11628 (N_11628,N_3616,N_33);
or U11629 (N_11629,N_5616,N_3968);
xnor U11630 (N_11630,N_1738,N_2456);
nor U11631 (N_11631,N_70,N_4640);
nor U11632 (N_11632,N_4265,N_4343);
nand U11633 (N_11633,N_2047,N_1030);
or U11634 (N_11634,N_141,N_105);
xnor U11635 (N_11635,N_5446,N_2028);
nor U11636 (N_11636,N_1141,N_668);
xor U11637 (N_11637,N_6174,N_5366);
nor U11638 (N_11638,N_2418,N_2217);
nor U11639 (N_11639,N_3543,N_437);
or U11640 (N_11640,N_612,N_2035);
xnor U11641 (N_11641,N_3212,N_4054);
nand U11642 (N_11642,N_5954,N_2534);
xor U11643 (N_11643,N_4906,N_4303);
or U11644 (N_11644,N_4630,N_2615);
nor U11645 (N_11645,N_1828,N_5992);
nor U11646 (N_11646,N_2713,N_4927);
xnor U11647 (N_11647,N_5408,N_6118);
nor U11648 (N_11648,N_2540,N_4614);
xnor U11649 (N_11649,N_4848,N_3255);
nand U11650 (N_11650,N_3039,N_5895);
nor U11651 (N_11651,N_4456,N_4611);
nand U11652 (N_11652,N_323,N_5631);
nand U11653 (N_11653,N_1906,N_4904);
and U11654 (N_11654,N_5409,N_4221);
or U11655 (N_11655,N_3478,N_4143);
xnor U11656 (N_11656,N_1086,N_1265);
nor U11657 (N_11657,N_4408,N_658);
nor U11658 (N_11658,N_5524,N_5778);
nor U11659 (N_11659,N_19,N_6217);
and U11660 (N_11660,N_658,N_4115);
xor U11661 (N_11661,N_2893,N_4976);
nand U11662 (N_11662,N_2615,N_3535);
nand U11663 (N_11663,N_6084,N_1176);
nor U11664 (N_11664,N_3171,N_4768);
xor U11665 (N_11665,N_5462,N_2681);
nor U11666 (N_11666,N_3045,N_1932);
nand U11667 (N_11667,N_1024,N_1156);
and U11668 (N_11668,N_5031,N_2390);
or U11669 (N_11669,N_2273,N_2477);
nor U11670 (N_11670,N_494,N_2447);
xor U11671 (N_11671,N_6043,N_4605);
and U11672 (N_11672,N_1235,N_682);
or U11673 (N_11673,N_2447,N_4118);
xor U11674 (N_11674,N_3809,N_5041);
or U11675 (N_11675,N_312,N_5913);
and U11676 (N_11676,N_4854,N_2087);
nand U11677 (N_11677,N_3065,N_2678);
and U11678 (N_11678,N_1063,N_6018);
xnor U11679 (N_11679,N_977,N_2375);
nor U11680 (N_11680,N_873,N_358);
nand U11681 (N_11681,N_1808,N_727);
or U11682 (N_11682,N_5404,N_4557);
or U11683 (N_11683,N_2540,N_5893);
nor U11684 (N_11684,N_579,N_5619);
xor U11685 (N_11685,N_3869,N_1794);
nand U11686 (N_11686,N_3867,N_496);
nor U11687 (N_11687,N_1807,N_3609);
or U11688 (N_11688,N_5739,N_5756);
nor U11689 (N_11689,N_331,N_3270);
and U11690 (N_11690,N_5026,N_4597);
nand U11691 (N_11691,N_1863,N_5702);
nor U11692 (N_11692,N_6148,N_424);
or U11693 (N_11693,N_1301,N_1798);
nor U11694 (N_11694,N_4405,N_1362);
nand U11695 (N_11695,N_874,N_5630);
or U11696 (N_11696,N_4495,N_1012);
xor U11697 (N_11697,N_2121,N_1784);
xor U11698 (N_11698,N_2842,N_663);
nand U11699 (N_11699,N_4690,N_1209);
or U11700 (N_11700,N_3506,N_4249);
xnor U11701 (N_11701,N_4010,N_1129);
nand U11702 (N_11702,N_30,N_1175);
nand U11703 (N_11703,N_4691,N_4438);
or U11704 (N_11704,N_1740,N_5977);
nor U11705 (N_11705,N_1381,N_1549);
or U11706 (N_11706,N_5117,N_6116);
nand U11707 (N_11707,N_4753,N_4054);
or U11708 (N_11708,N_3599,N_1798);
nand U11709 (N_11709,N_1786,N_1216);
nor U11710 (N_11710,N_3226,N_4156);
nor U11711 (N_11711,N_3238,N_4516);
and U11712 (N_11712,N_4856,N_5248);
nand U11713 (N_11713,N_4481,N_1707);
or U11714 (N_11714,N_5165,N_2790);
nand U11715 (N_11715,N_3646,N_5899);
or U11716 (N_11716,N_259,N_3019);
nand U11717 (N_11717,N_2747,N_4330);
nand U11718 (N_11718,N_2614,N_374);
nor U11719 (N_11719,N_2089,N_1328);
xor U11720 (N_11720,N_3717,N_1860);
xnor U11721 (N_11721,N_2802,N_4584);
nor U11722 (N_11722,N_5631,N_4873);
or U11723 (N_11723,N_1085,N_5513);
or U11724 (N_11724,N_5644,N_1873);
nand U11725 (N_11725,N_5651,N_2121);
nand U11726 (N_11726,N_1774,N_165);
nor U11727 (N_11727,N_4589,N_4263);
and U11728 (N_11728,N_5941,N_5348);
nor U11729 (N_11729,N_729,N_2837);
or U11730 (N_11730,N_385,N_87);
or U11731 (N_11731,N_2140,N_5616);
nand U11732 (N_11732,N_2517,N_4891);
or U11733 (N_11733,N_3121,N_2892);
or U11734 (N_11734,N_2862,N_96);
nand U11735 (N_11735,N_1616,N_5566);
nand U11736 (N_11736,N_641,N_6190);
nand U11737 (N_11737,N_6113,N_4420);
nand U11738 (N_11738,N_238,N_850);
or U11739 (N_11739,N_1328,N_5302);
nand U11740 (N_11740,N_5542,N_3521);
xor U11741 (N_11741,N_6011,N_5233);
xor U11742 (N_11742,N_1035,N_2346);
nor U11743 (N_11743,N_6169,N_3332);
xor U11744 (N_11744,N_1162,N_4480);
and U11745 (N_11745,N_6074,N_4169);
or U11746 (N_11746,N_2386,N_3824);
and U11747 (N_11747,N_3101,N_4819);
or U11748 (N_11748,N_4856,N_2913);
and U11749 (N_11749,N_4287,N_4496);
or U11750 (N_11750,N_1649,N_5665);
xor U11751 (N_11751,N_3823,N_313);
nor U11752 (N_11752,N_4162,N_2171);
nand U11753 (N_11753,N_5424,N_3120);
and U11754 (N_11754,N_1238,N_5006);
and U11755 (N_11755,N_5394,N_653);
nand U11756 (N_11756,N_5672,N_4332);
nor U11757 (N_11757,N_3782,N_4684);
nor U11758 (N_11758,N_4791,N_5166);
xnor U11759 (N_11759,N_316,N_2282);
nor U11760 (N_11760,N_4733,N_4378);
xor U11761 (N_11761,N_2303,N_2282);
nand U11762 (N_11762,N_4885,N_2438);
xnor U11763 (N_11763,N_2058,N_2385);
xnor U11764 (N_11764,N_2791,N_1884);
nand U11765 (N_11765,N_1601,N_4405);
or U11766 (N_11766,N_1661,N_4883);
nor U11767 (N_11767,N_1068,N_5869);
nor U11768 (N_11768,N_114,N_1904);
xor U11769 (N_11769,N_4016,N_4050);
or U11770 (N_11770,N_475,N_284);
and U11771 (N_11771,N_3448,N_5251);
xor U11772 (N_11772,N_3565,N_3592);
or U11773 (N_11773,N_417,N_2176);
nand U11774 (N_11774,N_1327,N_2833);
nand U11775 (N_11775,N_1123,N_227);
nand U11776 (N_11776,N_3249,N_277);
nor U11777 (N_11777,N_2637,N_3814);
xnor U11778 (N_11778,N_332,N_4801);
xnor U11779 (N_11779,N_3711,N_3533);
nand U11780 (N_11780,N_4151,N_5895);
nor U11781 (N_11781,N_3882,N_6191);
xnor U11782 (N_11782,N_1237,N_47);
and U11783 (N_11783,N_416,N_236);
and U11784 (N_11784,N_3133,N_3209);
nor U11785 (N_11785,N_3589,N_4411);
nor U11786 (N_11786,N_388,N_798);
xor U11787 (N_11787,N_2064,N_2431);
or U11788 (N_11788,N_3946,N_4951);
nor U11789 (N_11789,N_1710,N_6169);
nand U11790 (N_11790,N_4496,N_1530);
or U11791 (N_11791,N_6112,N_4782);
xor U11792 (N_11792,N_3280,N_5918);
and U11793 (N_11793,N_5997,N_1637);
xnor U11794 (N_11794,N_351,N_5988);
and U11795 (N_11795,N_118,N_5614);
or U11796 (N_11796,N_796,N_4428);
nor U11797 (N_11797,N_4730,N_4153);
xnor U11798 (N_11798,N_5760,N_1412);
nor U11799 (N_11799,N_2599,N_5972);
nor U11800 (N_11800,N_5497,N_220);
nor U11801 (N_11801,N_2645,N_1581);
and U11802 (N_11802,N_5072,N_713);
nand U11803 (N_11803,N_6226,N_179);
and U11804 (N_11804,N_455,N_3368);
xor U11805 (N_11805,N_6053,N_1000);
xor U11806 (N_11806,N_6247,N_2118);
xnor U11807 (N_11807,N_1099,N_6148);
or U11808 (N_11808,N_6158,N_883);
nor U11809 (N_11809,N_435,N_1384);
and U11810 (N_11810,N_1667,N_727);
or U11811 (N_11811,N_4739,N_5053);
or U11812 (N_11812,N_78,N_1185);
nor U11813 (N_11813,N_3081,N_2376);
nand U11814 (N_11814,N_483,N_2439);
nand U11815 (N_11815,N_6238,N_2553);
nand U11816 (N_11816,N_1598,N_1605);
xor U11817 (N_11817,N_511,N_2862);
nand U11818 (N_11818,N_1035,N_1782);
and U11819 (N_11819,N_5876,N_4150);
nor U11820 (N_11820,N_3232,N_6231);
or U11821 (N_11821,N_1204,N_1858);
nor U11822 (N_11822,N_4230,N_4219);
or U11823 (N_11823,N_4336,N_2067);
or U11824 (N_11824,N_2297,N_5742);
or U11825 (N_11825,N_1319,N_5270);
xnor U11826 (N_11826,N_5364,N_3161);
and U11827 (N_11827,N_1207,N_5135);
nor U11828 (N_11828,N_5623,N_1480);
or U11829 (N_11829,N_1359,N_271);
xor U11830 (N_11830,N_347,N_3979);
or U11831 (N_11831,N_5034,N_694);
nand U11832 (N_11832,N_1896,N_103);
or U11833 (N_11833,N_5150,N_1403);
or U11834 (N_11834,N_1786,N_273);
and U11835 (N_11835,N_3546,N_4712);
and U11836 (N_11836,N_940,N_5461);
and U11837 (N_11837,N_3164,N_4481);
and U11838 (N_11838,N_1936,N_188);
xnor U11839 (N_11839,N_3903,N_4994);
xor U11840 (N_11840,N_2110,N_298);
nand U11841 (N_11841,N_173,N_1577);
xnor U11842 (N_11842,N_1283,N_5062);
and U11843 (N_11843,N_2648,N_1656);
and U11844 (N_11844,N_6204,N_3714);
nor U11845 (N_11845,N_3355,N_5705);
or U11846 (N_11846,N_2393,N_2656);
xor U11847 (N_11847,N_4785,N_5586);
xnor U11848 (N_11848,N_6196,N_4669);
xor U11849 (N_11849,N_3584,N_4982);
nor U11850 (N_11850,N_4944,N_3921);
and U11851 (N_11851,N_5716,N_2371);
nand U11852 (N_11852,N_2447,N_1354);
and U11853 (N_11853,N_3127,N_4586);
or U11854 (N_11854,N_2379,N_4073);
nand U11855 (N_11855,N_4808,N_2326);
and U11856 (N_11856,N_5574,N_3641);
or U11857 (N_11857,N_39,N_5821);
nor U11858 (N_11858,N_3768,N_2114);
nand U11859 (N_11859,N_1685,N_5162);
and U11860 (N_11860,N_2920,N_4614);
and U11861 (N_11861,N_2067,N_793);
nand U11862 (N_11862,N_577,N_1796);
nand U11863 (N_11863,N_2682,N_1336);
nor U11864 (N_11864,N_45,N_3581);
and U11865 (N_11865,N_3753,N_4717);
or U11866 (N_11866,N_2716,N_2671);
or U11867 (N_11867,N_4096,N_4889);
or U11868 (N_11868,N_1198,N_501);
xnor U11869 (N_11869,N_4573,N_1886);
nand U11870 (N_11870,N_291,N_3753);
nor U11871 (N_11871,N_3415,N_216);
xor U11872 (N_11872,N_2473,N_1190);
nor U11873 (N_11873,N_5722,N_3349);
nor U11874 (N_11874,N_3732,N_5941);
or U11875 (N_11875,N_3248,N_5746);
nand U11876 (N_11876,N_4951,N_1103);
nand U11877 (N_11877,N_5268,N_46);
nor U11878 (N_11878,N_358,N_333);
nor U11879 (N_11879,N_6033,N_1181);
and U11880 (N_11880,N_2132,N_3807);
xnor U11881 (N_11881,N_497,N_491);
and U11882 (N_11882,N_2517,N_1314);
nand U11883 (N_11883,N_3400,N_804);
xor U11884 (N_11884,N_4732,N_1641);
xor U11885 (N_11885,N_1217,N_303);
or U11886 (N_11886,N_163,N_643);
or U11887 (N_11887,N_3880,N_4295);
and U11888 (N_11888,N_4979,N_888);
nor U11889 (N_11889,N_4108,N_5228);
and U11890 (N_11890,N_5686,N_4437);
nand U11891 (N_11891,N_3686,N_241);
or U11892 (N_11892,N_5179,N_4290);
xor U11893 (N_11893,N_6243,N_363);
and U11894 (N_11894,N_1955,N_4320);
nand U11895 (N_11895,N_2608,N_4024);
nand U11896 (N_11896,N_875,N_3934);
xnor U11897 (N_11897,N_2730,N_2796);
xor U11898 (N_11898,N_3414,N_2631);
nand U11899 (N_11899,N_507,N_1243);
nand U11900 (N_11900,N_5949,N_2176);
and U11901 (N_11901,N_5804,N_3505);
or U11902 (N_11902,N_3452,N_3266);
xnor U11903 (N_11903,N_501,N_5247);
or U11904 (N_11904,N_4933,N_569);
xor U11905 (N_11905,N_5799,N_927);
or U11906 (N_11906,N_225,N_563);
or U11907 (N_11907,N_4072,N_14);
or U11908 (N_11908,N_3625,N_217);
xnor U11909 (N_11909,N_3808,N_4370);
nor U11910 (N_11910,N_4647,N_5375);
nor U11911 (N_11911,N_4979,N_4702);
or U11912 (N_11912,N_673,N_4802);
or U11913 (N_11913,N_2690,N_6181);
nand U11914 (N_11914,N_1815,N_1728);
nor U11915 (N_11915,N_236,N_3169);
xor U11916 (N_11916,N_4115,N_241);
nand U11917 (N_11917,N_4691,N_2667);
nor U11918 (N_11918,N_846,N_2688);
nand U11919 (N_11919,N_595,N_4441);
or U11920 (N_11920,N_1652,N_916);
nand U11921 (N_11921,N_1620,N_863);
nor U11922 (N_11922,N_2385,N_4878);
nor U11923 (N_11923,N_62,N_6213);
or U11924 (N_11924,N_3033,N_577);
nor U11925 (N_11925,N_1451,N_3551);
nor U11926 (N_11926,N_2211,N_421);
nor U11927 (N_11927,N_1999,N_2083);
or U11928 (N_11928,N_3831,N_1905);
or U11929 (N_11929,N_4766,N_6016);
nand U11930 (N_11930,N_3013,N_4995);
nor U11931 (N_11931,N_1282,N_4203);
or U11932 (N_11932,N_894,N_1641);
and U11933 (N_11933,N_5383,N_4045);
or U11934 (N_11934,N_4532,N_2341);
or U11935 (N_11935,N_5767,N_4301);
nor U11936 (N_11936,N_5599,N_1758);
nor U11937 (N_11937,N_3284,N_5768);
and U11938 (N_11938,N_220,N_5833);
xor U11939 (N_11939,N_2164,N_3615);
nor U11940 (N_11940,N_5354,N_1496);
nor U11941 (N_11941,N_3493,N_5735);
nor U11942 (N_11942,N_320,N_5633);
xnor U11943 (N_11943,N_5996,N_4173);
and U11944 (N_11944,N_4430,N_258);
or U11945 (N_11945,N_1487,N_200);
or U11946 (N_11946,N_6036,N_1709);
and U11947 (N_11947,N_3939,N_3038);
nor U11948 (N_11948,N_3812,N_328);
or U11949 (N_11949,N_4125,N_1999);
nand U11950 (N_11950,N_5868,N_4879);
xor U11951 (N_11951,N_4886,N_4416);
nor U11952 (N_11952,N_6143,N_2012);
nor U11953 (N_11953,N_3189,N_1723);
nand U11954 (N_11954,N_5680,N_4152);
nor U11955 (N_11955,N_2856,N_4141);
xnor U11956 (N_11956,N_5815,N_3360);
or U11957 (N_11957,N_1034,N_917);
or U11958 (N_11958,N_1282,N_1070);
nor U11959 (N_11959,N_4176,N_1575);
and U11960 (N_11960,N_789,N_5371);
or U11961 (N_11961,N_526,N_6093);
nor U11962 (N_11962,N_2644,N_5263);
and U11963 (N_11963,N_4554,N_3379);
nand U11964 (N_11964,N_4789,N_2621);
nand U11965 (N_11965,N_3921,N_731);
xnor U11966 (N_11966,N_4080,N_661);
or U11967 (N_11967,N_5441,N_2302);
and U11968 (N_11968,N_1397,N_5279);
nor U11969 (N_11969,N_4328,N_3563);
nand U11970 (N_11970,N_5657,N_5673);
or U11971 (N_11971,N_4720,N_1868);
nand U11972 (N_11972,N_2499,N_1631);
xnor U11973 (N_11973,N_3984,N_2776);
xnor U11974 (N_11974,N_5982,N_5391);
xnor U11975 (N_11975,N_1918,N_3214);
xnor U11976 (N_11976,N_4060,N_2615);
xnor U11977 (N_11977,N_1269,N_1060);
nor U11978 (N_11978,N_4865,N_5409);
and U11979 (N_11979,N_5458,N_2529);
nor U11980 (N_11980,N_3540,N_2784);
and U11981 (N_11981,N_3626,N_3768);
and U11982 (N_11982,N_5104,N_2345);
nand U11983 (N_11983,N_2028,N_4966);
nand U11984 (N_11984,N_6133,N_142);
nor U11985 (N_11985,N_879,N_4741);
xnor U11986 (N_11986,N_1416,N_4463);
nor U11987 (N_11987,N_362,N_458);
nor U11988 (N_11988,N_4326,N_2557);
and U11989 (N_11989,N_3614,N_5619);
and U11990 (N_11990,N_4719,N_318);
nand U11991 (N_11991,N_193,N_1932);
nor U11992 (N_11992,N_4571,N_689);
or U11993 (N_11993,N_5387,N_4481);
xor U11994 (N_11994,N_4098,N_4993);
and U11995 (N_11995,N_887,N_2202);
xnor U11996 (N_11996,N_4659,N_2955);
nand U11997 (N_11997,N_690,N_4485);
or U11998 (N_11998,N_6147,N_1024);
nand U11999 (N_11999,N_1604,N_5655);
or U12000 (N_12000,N_5457,N_1565);
xnor U12001 (N_12001,N_593,N_3483);
nand U12002 (N_12002,N_3106,N_2373);
nand U12003 (N_12003,N_1244,N_2479);
nor U12004 (N_12004,N_442,N_3216);
and U12005 (N_12005,N_5906,N_5568);
and U12006 (N_12006,N_3538,N_738);
and U12007 (N_12007,N_3465,N_6161);
xor U12008 (N_12008,N_3890,N_5028);
or U12009 (N_12009,N_3936,N_3293);
nand U12010 (N_12010,N_340,N_2557);
or U12011 (N_12011,N_3520,N_549);
nor U12012 (N_12012,N_470,N_6014);
nand U12013 (N_12013,N_1185,N_1095);
xnor U12014 (N_12014,N_746,N_2095);
or U12015 (N_12015,N_3788,N_1692);
and U12016 (N_12016,N_2538,N_887);
nand U12017 (N_12017,N_4222,N_6033);
xor U12018 (N_12018,N_5773,N_3254);
nor U12019 (N_12019,N_1036,N_5546);
and U12020 (N_12020,N_3651,N_5008);
and U12021 (N_12021,N_3232,N_5140);
or U12022 (N_12022,N_467,N_3980);
and U12023 (N_12023,N_5609,N_5256);
nor U12024 (N_12024,N_872,N_5305);
nand U12025 (N_12025,N_1244,N_2184);
and U12026 (N_12026,N_824,N_2857);
nand U12027 (N_12027,N_4977,N_3743);
nor U12028 (N_12028,N_4441,N_683);
and U12029 (N_12029,N_4867,N_3024);
and U12030 (N_12030,N_2580,N_1512);
xor U12031 (N_12031,N_4902,N_383);
nand U12032 (N_12032,N_2527,N_4087);
nor U12033 (N_12033,N_346,N_2561);
nand U12034 (N_12034,N_1365,N_4532);
nor U12035 (N_12035,N_1458,N_335);
nor U12036 (N_12036,N_3320,N_5580);
or U12037 (N_12037,N_1380,N_5641);
xnor U12038 (N_12038,N_3128,N_3612);
nand U12039 (N_12039,N_131,N_4932);
and U12040 (N_12040,N_1579,N_2238);
or U12041 (N_12041,N_2399,N_2263);
nor U12042 (N_12042,N_2996,N_3244);
nand U12043 (N_12043,N_3598,N_1778);
or U12044 (N_12044,N_2273,N_1304);
and U12045 (N_12045,N_4392,N_1998);
or U12046 (N_12046,N_1740,N_3338);
nand U12047 (N_12047,N_5706,N_2434);
nand U12048 (N_12048,N_4309,N_3511);
or U12049 (N_12049,N_2582,N_859);
and U12050 (N_12050,N_1221,N_5135);
and U12051 (N_12051,N_26,N_2372);
or U12052 (N_12052,N_4577,N_1469);
or U12053 (N_12053,N_5168,N_2253);
nand U12054 (N_12054,N_6169,N_1001);
nor U12055 (N_12055,N_6067,N_5811);
xor U12056 (N_12056,N_5573,N_1543);
or U12057 (N_12057,N_1096,N_5697);
and U12058 (N_12058,N_123,N_3215);
and U12059 (N_12059,N_4465,N_6006);
or U12060 (N_12060,N_3104,N_1662);
nand U12061 (N_12061,N_2871,N_4841);
and U12062 (N_12062,N_1271,N_4077);
xnor U12063 (N_12063,N_5041,N_155);
nand U12064 (N_12064,N_4102,N_3101);
nor U12065 (N_12065,N_6223,N_6017);
nand U12066 (N_12066,N_631,N_3638);
or U12067 (N_12067,N_3739,N_2497);
or U12068 (N_12068,N_3193,N_6045);
xnor U12069 (N_12069,N_3378,N_5487);
and U12070 (N_12070,N_5835,N_321);
or U12071 (N_12071,N_2388,N_5206);
or U12072 (N_12072,N_5977,N_5132);
xnor U12073 (N_12073,N_4727,N_2913);
nor U12074 (N_12074,N_74,N_6028);
nor U12075 (N_12075,N_1293,N_5214);
or U12076 (N_12076,N_5393,N_5996);
nor U12077 (N_12077,N_2297,N_1753);
and U12078 (N_12078,N_2535,N_5763);
xnor U12079 (N_12079,N_3745,N_5482);
and U12080 (N_12080,N_1300,N_4467);
nand U12081 (N_12081,N_4575,N_817);
or U12082 (N_12082,N_2142,N_3305);
nand U12083 (N_12083,N_4566,N_1855);
and U12084 (N_12084,N_3301,N_4917);
and U12085 (N_12085,N_4738,N_4906);
and U12086 (N_12086,N_6129,N_4509);
nor U12087 (N_12087,N_2865,N_6218);
or U12088 (N_12088,N_5894,N_4651);
and U12089 (N_12089,N_5416,N_2064);
nand U12090 (N_12090,N_3200,N_4145);
xor U12091 (N_12091,N_745,N_3085);
or U12092 (N_12092,N_4326,N_4235);
or U12093 (N_12093,N_5834,N_5202);
nand U12094 (N_12094,N_4134,N_5900);
or U12095 (N_12095,N_4902,N_1086);
or U12096 (N_12096,N_1771,N_1526);
and U12097 (N_12097,N_3913,N_3343);
xor U12098 (N_12098,N_1203,N_1263);
nor U12099 (N_12099,N_1910,N_1695);
or U12100 (N_12100,N_5996,N_5200);
nand U12101 (N_12101,N_5841,N_4103);
xnor U12102 (N_12102,N_2781,N_4409);
nor U12103 (N_12103,N_1049,N_503);
xnor U12104 (N_12104,N_122,N_2320);
xor U12105 (N_12105,N_62,N_6128);
nand U12106 (N_12106,N_263,N_3590);
nand U12107 (N_12107,N_1792,N_5783);
or U12108 (N_12108,N_4447,N_5432);
nor U12109 (N_12109,N_3929,N_3469);
xor U12110 (N_12110,N_4561,N_6214);
nor U12111 (N_12111,N_6140,N_1978);
or U12112 (N_12112,N_5096,N_267);
and U12113 (N_12113,N_2365,N_6122);
xnor U12114 (N_12114,N_648,N_1081);
and U12115 (N_12115,N_2998,N_2229);
nand U12116 (N_12116,N_4578,N_3146);
and U12117 (N_12117,N_5340,N_2767);
nand U12118 (N_12118,N_6049,N_1493);
nand U12119 (N_12119,N_5318,N_889);
or U12120 (N_12120,N_6136,N_5028);
xnor U12121 (N_12121,N_1644,N_4400);
and U12122 (N_12122,N_1045,N_1968);
xor U12123 (N_12123,N_6009,N_2393);
and U12124 (N_12124,N_1071,N_3556);
xnor U12125 (N_12125,N_1398,N_500);
and U12126 (N_12126,N_4128,N_1088);
xnor U12127 (N_12127,N_3418,N_2257);
or U12128 (N_12128,N_1084,N_5218);
xnor U12129 (N_12129,N_378,N_5964);
and U12130 (N_12130,N_5660,N_599);
or U12131 (N_12131,N_977,N_5772);
and U12132 (N_12132,N_3405,N_4735);
or U12133 (N_12133,N_6093,N_3484);
and U12134 (N_12134,N_4610,N_4741);
nor U12135 (N_12135,N_1220,N_4562);
nor U12136 (N_12136,N_1243,N_3651);
nor U12137 (N_12137,N_836,N_3831);
xor U12138 (N_12138,N_4418,N_1164);
nand U12139 (N_12139,N_3199,N_3324);
and U12140 (N_12140,N_4643,N_5906);
or U12141 (N_12141,N_1079,N_253);
nand U12142 (N_12142,N_5775,N_1549);
xor U12143 (N_12143,N_4872,N_2338);
and U12144 (N_12144,N_1940,N_813);
nand U12145 (N_12145,N_1438,N_4600);
or U12146 (N_12146,N_258,N_587);
nand U12147 (N_12147,N_5137,N_1989);
or U12148 (N_12148,N_2385,N_2729);
and U12149 (N_12149,N_369,N_5417);
nand U12150 (N_12150,N_2742,N_680);
nand U12151 (N_12151,N_5698,N_3853);
nand U12152 (N_12152,N_121,N_5215);
xnor U12153 (N_12153,N_2671,N_5667);
xor U12154 (N_12154,N_4480,N_260);
and U12155 (N_12155,N_2045,N_1021);
nor U12156 (N_12156,N_4310,N_3907);
or U12157 (N_12157,N_1071,N_2595);
nor U12158 (N_12158,N_2747,N_1972);
xor U12159 (N_12159,N_1095,N_1204);
and U12160 (N_12160,N_4727,N_1543);
or U12161 (N_12161,N_1889,N_1679);
nor U12162 (N_12162,N_2225,N_3190);
nand U12163 (N_12163,N_571,N_2570);
xor U12164 (N_12164,N_4859,N_826);
and U12165 (N_12165,N_1408,N_4734);
nand U12166 (N_12166,N_3760,N_199);
or U12167 (N_12167,N_4869,N_3028);
xor U12168 (N_12168,N_3884,N_5926);
or U12169 (N_12169,N_1806,N_4816);
and U12170 (N_12170,N_1624,N_5144);
xor U12171 (N_12171,N_4789,N_5137);
nand U12172 (N_12172,N_3895,N_880);
nand U12173 (N_12173,N_1668,N_4784);
or U12174 (N_12174,N_3133,N_6161);
xor U12175 (N_12175,N_5788,N_1233);
and U12176 (N_12176,N_5400,N_317);
and U12177 (N_12177,N_2844,N_3331);
nor U12178 (N_12178,N_1585,N_307);
or U12179 (N_12179,N_1183,N_668);
xnor U12180 (N_12180,N_3121,N_1165);
nand U12181 (N_12181,N_4371,N_478);
and U12182 (N_12182,N_4122,N_440);
or U12183 (N_12183,N_2659,N_1171);
nand U12184 (N_12184,N_3726,N_2467);
nor U12185 (N_12185,N_3047,N_2492);
or U12186 (N_12186,N_4093,N_3656);
nand U12187 (N_12187,N_953,N_3823);
or U12188 (N_12188,N_5900,N_6098);
xnor U12189 (N_12189,N_4987,N_1907);
or U12190 (N_12190,N_890,N_4457);
and U12191 (N_12191,N_1586,N_6217);
nor U12192 (N_12192,N_2398,N_2618);
xnor U12193 (N_12193,N_4577,N_4666);
xnor U12194 (N_12194,N_3252,N_2120);
or U12195 (N_12195,N_1894,N_4047);
nand U12196 (N_12196,N_2762,N_1085);
nor U12197 (N_12197,N_2117,N_2740);
or U12198 (N_12198,N_816,N_4302);
nor U12199 (N_12199,N_5553,N_5852);
nor U12200 (N_12200,N_965,N_5911);
or U12201 (N_12201,N_2966,N_3197);
and U12202 (N_12202,N_2254,N_892);
or U12203 (N_12203,N_248,N_4769);
or U12204 (N_12204,N_1140,N_2275);
nand U12205 (N_12205,N_2646,N_5983);
nor U12206 (N_12206,N_5338,N_4481);
nand U12207 (N_12207,N_1849,N_869);
nor U12208 (N_12208,N_2637,N_2201);
nor U12209 (N_12209,N_4683,N_2585);
and U12210 (N_12210,N_5288,N_4516);
xnor U12211 (N_12211,N_1635,N_2858);
nand U12212 (N_12212,N_895,N_5359);
nor U12213 (N_12213,N_4484,N_4279);
xor U12214 (N_12214,N_1903,N_1266);
or U12215 (N_12215,N_257,N_5589);
and U12216 (N_12216,N_444,N_5836);
nand U12217 (N_12217,N_5580,N_5197);
xor U12218 (N_12218,N_420,N_5146);
nor U12219 (N_12219,N_5758,N_3006);
xor U12220 (N_12220,N_4651,N_3258);
nor U12221 (N_12221,N_3129,N_1348);
xnor U12222 (N_12222,N_1400,N_1595);
and U12223 (N_12223,N_3876,N_3340);
and U12224 (N_12224,N_2547,N_4182);
nand U12225 (N_12225,N_1087,N_2407);
nor U12226 (N_12226,N_5939,N_2324);
nor U12227 (N_12227,N_5095,N_398);
or U12228 (N_12228,N_4812,N_5379);
nor U12229 (N_12229,N_1643,N_4377);
or U12230 (N_12230,N_2735,N_4538);
or U12231 (N_12231,N_1029,N_1903);
and U12232 (N_12232,N_5750,N_5646);
and U12233 (N_12233,N_487,N_3575);
and U12234 (N_12234,N_2212,N_2710);
or U12235 (N_12235,N_572,N_2954);
or U12236 (N_12236,N_6226,N_5466);
nor U12237 (N_12237,N_1815,N_296);
nand U12238 (N_12238,N_274,N_3826);
and U12239 (N_12239,N_1039,N_3871);
nor U12240 (N_12240,N_4483,N_1062);
nor U12241 (N_12241,N_1462,N_3952);
or U12242 (N_12242,N_5822,N_1603);
nand U12243 (N_12243,N_724,N_5802);
xor U12244 (N_12244,N_2001,N_775);
xor U12245 (N_12245,N_5753,N_3385);
xnor U12246 (N_12246,N_5460,N_1163);
xnor U12247 (N_12247,N_2797,N_4630);
xor U12248 (N_12248,N_3248,N_5666);
or U12249 (N_12249,N_5909,N_1941);
nand U12250 (N_12250,N_2281,N_4048);
nor U12251 (N_12251,N_330,N_1938);
nand U12252 (N_12252,N_4129,N_337);
nor U12253 (N_12253,N_1984,N_3289);
or U12254 (N_12254,N_4598,N_4196);
and U12255 (N_12255,N_6200,N_2130);
nor U12256 (N_12256,N_956,N_3465);
nand U12257 (N_12257,N_3593,N_2970);
xor U12258 (N_12258,N_2601,N_2248);
or U12259 (N_12259,N_1980,N_1510);
nand U12260 (N_12260,N_4672,N_3645);
and U12261 (N_12261,N_1994,N_1531);
nand U12262 (N_12262,N_581,N_3963);
xor U12263 (N_12263,N_1347,N_273);
xnor U12264 (N_12264,N_3545,N_4741);
nor U12265 (N_12265,N_5439,N_4349);
and U12266 (N_12266,N_2052,N_1549);
xor U12267 (N_12267,N_570,N_5529);
and U12268 (N_12268,N_154,N_2957);
or U12269 (N_12269,N_5055,N_1773);
nor U12270 (N_12270,N_1886,N_3211);
xnor U12271 (N_12271,N_888,N_5242);
nand U12272 (N_12272,N_1061,N_4994);
or U12273 (N_12273,N_1594,N_4905);
nand U12274 (N_12274,N_4897,N_5735);
nand U12275 (N_12275,N_4173,N_5125);
or U12276 (N_12276,N_4926,N_5629);
and U12277 (N_12277,N_3196,N_1005);
or U12278 (N_12278,N_2455,N_6070);
nor U12279 (N_12279,N_5898,N_6243);
or U12280 (N_12280,N_1834,N_3285);
nor U12281 (N_12281,N_939,N_5291);
nand U12282 (N_12282,N_6022,N_2075);
nand U12283 (N_12283,N_3684,N_254);
or U12284 (N_12284,N_4551,N_4638);
and U12285 (N_12285,N_1378,N_4863);
xnor U12286 (N_12286,N_6012,N_6223);
xnor U12287 (N_12287,N_1764,N_933);
and U12288 (N_12288,N_2000,N_1750);
nor U12289 (N_12289,N_5842,N_3789);
xnor U12290 (N_12290,N_580,N_361);
or U12291 (N_12291,N_2032,N_2414);
nor U12292 (N_12292,N_875,N_1023);
and U12293 (N_12293,N_3335,N_2021);
xor U12294 (N_12294,N_1795,N_264);
xnor U12295 (N_12295,N_1777,N_447);
nand U12296 (N_12296,N_1103,N_4968);
and U12297 (N_12297,N_5675,N_4012);
or U12298 (N_12298,N_251,N_5437);
or U12299 (N_12299,N_2477,N_5489);
nor U12300 (N_12300,N_251,N_2400);
or U12301 (N_12301,N_4929,N_539);
nor U12302 (N_12302,N_5187,N_5525);
nand U12303 (N_12303,N_3704,N_2220);
nand U12304 (N_12304,N_1034,N_3503);
nand U12305 (N_12305,N_5640,N_2428);
nor U12306 (N_12306,N_5702,N_4651);
nor U12307 (N_12307,N_63,N_2657);
nand U12308 (N_12308,N_2565,N_5237);
xor U12309 (N_12309,N_2612,N_2794);
nor U12310 (N_12310,N_5271,N_3139);
nor U12311 (N_12311,N_5918,N_2920);
xor U12312 (N_12312,N_623,N_1538);
and U12313 (N_12313,N_731,N_1146);
or U12314 (N_12314,N_6184,N_6119);
or U12315 (N_12315,N_1384,N_114);
or U12316 (N_12316,N_1891,N_6248);
or U12317 (N_12317,N_3631,N_1119);
xor U12318 (N_12318,N_4752,N_3095);
or U12319 (N_12319,N_3544,N_5107);
or U12320 (N_12320,N_1567,N_4124);
and U12321 (N_12321,N_4704,N_4008);
nand U12322 (N_12322,N_3817,N_2672);
and U12323 (N_12323,N_5950,N_4116);
xor U12324 (N_12324,N_4270,N_1094);
or U12325 (N_12325,N_1531,N_2651);
nor U12326 (N_12326,N_4738,N_2708);
xor U12327 (N_12327,N_3530,N_6129);
and U12328 (N_12328,N_2374,N_5083);
nor U12329 (N_12329,N_1638,N_3774);
nor U12330 (N_12330,N_4907,N_1808);
nor U12331 (N_12331,N_5474,N_23);
and U12332 (N_12332,N_3773,N_4058);
or U12333 (N_12333,N_1680,N_801);
xnor U12334 (N_12334,N_3943,N_4719);
and U12335 (N_12335,N_1342,N_5788);
and U12336 (N_12336,N_8,N_2518);
or U12337 (N_12337,N_1143,N_4866);
nor U12338 (N_12338,N_1182,N_856);
nor U12339 (N_12339,N_1273,N_3270);
nor U12340 (N_12340,N_5934,N_299);
nand U12341 (N_12341,N_4961,N_660);
nand U12342 (N_12342,N_2349,N_68);
or U12343 (N_12343,N_4458,N_2060);
and U12344 (N_12344,N_4183,N_4871);
nor U12345 (N_12345,N_6092,N_4432);
nor U12346 (N_12346,N_453,N_3257);
nand U12347 (N_12347,N_2341,N_1983);
and U12348 (N_12348,N_4456,N_3428);
xnor U12349 (N_12349,N_625,N_2201);
or U12350 (N_12350,N_5329,N_5493);
or U12351 (N_12351,N_5320,N_5022);
nand U12352 (N_12352,N_3326,N_3974);
or U12353 (N_12353,N_3356,N_2994);
xnor U12354 (N_12354,N_986,N_375);
or U12355 (N_12355,N_383,N_5611);
xor U12356 (N_12356,N_4631,N_694);
or U12357 (N_12357,N_5297,N_699);
and U12358 (N_12358,N_5050,N_2650);
and U12359 (N_12359,N_3620,N_1516);
nand U12360 (N_12360,N_4472,N_5984);
and U12361 (N_12361,N_5652,N_5291);
xor U12362 (N_12362,N_704,N_2391);
xor U12363 (N_12363,N_2651,N_4990);
nor U12364 (N_12364,N_1376,N_947);
or U12365 (N_12365,N_3406,N_3226);
and U12366 (N_12366,N_5224,N_696);
nor U12367 (N_12367,N_4367,N_5233);
nor U12368 (N_12368,N_4989,N_1083);
and U12369 (N_12369,N_265,N_5275);
xor U12370 (N_12370,N_4362,N_4331);
and U12371 (N_12371,N_3359,N_3656);
nor U12372 (N_12372,N_2060,N_2949);
xor U12373 (N_12373,N_5040,N_4809);
nor U12374 (N_12374,N_535,N_2767);
nor U12375 (N_12375,N_2869,N_5661);
nor U12376 (N_12376,N_5770,N_6097);
nor U12377 (N_12377,N_7,N_2145);
xnor U12378 (N_12378,N_1751,N_5106);
nor U12379 (N_12379,N_5160,N_5017);
nor U12380 (N_12380,N_4875,N_6077);
and U12381 (N_12381,N_372,N_2669);
xnor U12382 (N_12382,N_2504,N_2169);
or U12383 (N_12383,N_4867,N_1164);
nor U12384 (N_12384,N_2937,N_3005);
xor U12385 (N_12385,N_928,N_4226);
nor U12386 (N_12386,N_4732,N_4778);
nand U12387 (N_12387,N_2760,N_940);
xor U12388 (N_12388,N_4194,N_4730);
nor U12389 (N_12389,N_7,N_230);
nand U12390 (N_12390,N_5201,N_2994);
or U12391 (N_12391,N_4407,N_2081);
nor U12392 (N_12392,N_3995,N_1382);
nand U12393 (N_12393,N_4836,N_2206);
and U12394 (N_12394,N_3918,N_6027);
and U12395 (N_12395,N_5521,N_2636);
and U12396 (N_12396,N_2415,N_4669);
nor U12397 (N_12397,N_5667,N_4232);
or U12398 (N_12398,N_5197,N_1967);
nand U12399 (N_12399,N_6103,N_3938);
xnor U12400 (N_12400,N_2638,N_2096);
nor U12401 (N_12401,N_4453,N_2302);
nor U12402 (N_12402,N_1516,N_4603);
and U12403 (N_12403,N_2468,N_5207);
and U12404 (N_12404,N_2982,N_3696);
or U12405 (N_12405,N_3562,N_2924);
or U12406 (N_12406,N_5982,N_2241);
nand U12407 (N_12407,N_5974,N_4133);
and U12408 (N_12408,N_5332,N_4899);
nor U12409 (N_12409,N_3870,N_1017);
xnor U12410 (N_12410,N_5115,N_2263);
or U12411 (N_12411,N_2383,N_1248);
xnor U12412 (N_12412,N_332,N_1901);
xor U12413 (N_12413,N_5732,N_1885);
nand U12414 (N_12414,N_4209,N_201);
or U12415 (N_12415,N_4307,N_3061);
and U12416 (N_12416,N_5033,N_1386);
xor U12417 (N_12417,N_4596,N_3643);
or U12418 (N_12418,N_659,N_618);
nor U12419 (N_12419,N_1786,N_5222);
nor U12420 (N_12420,N_1631,N_113);
nand U12421 (N_12421,N_4274,N_4673);
nand U12422 (N_12422,N_14,N_2278);
nand U12423 (N_12423,N_4597,N_1443);
nor U12424 (N_12424,N_566,N_4384);
nor U12425 (N_12425,N_2184,N_1955);
xnor U12426 (N_12426,N_4691,N_276);
nand U12427 (N_12427,N_5133,N_1355);
or U12428 (N_12428,N_2461,N_4909);
and U12429 (N_12429,N_3676,N_1849);
nor U12430 (N_12430,N_4860,N_2272);
or U12431 (N_12431,N_1304,N_3049);
xor U12432 (N_12432,N_2380,N_2137);
or U12433 (N_12433,N_2177,N_4715);
nor U12434 (N_12434,N_5731,N_5684);
xor U12435 (N_12435,N_2888,N_2985);
nor U12436 (N_12436,N_5646,N_2724);
nand U12437 (N_12437,N_2584,N_4278);
nor U12438 (N_12438,N_2458,N_2935);
and U12439 (N_12439,N_264,N_3111);
nor U12440 (N_12440,N_1718,N_6016);
and U12441 (N_12441,N_2998,N_3415);
and U12442 (N_12442,N_5159,N_1776);
nand U12443 (N_12443,N_4197,N_4599);
or U12444 (N_12444,N_5631,N_3862);
nand U12445 (N_12445,N_3246,N_4977);
xnor U12446 (N_12446,N_214,N_482);
and U12447 (N_12447,N_3475,N_4660);
or U12448 (N_12448,N_3532,N_2971);
nor U12449 (N_12449,N_189,N_4382);
or U12450 (N_12450,N_1941,N_930);
nand U12451 (N_12451,N_1163,N_4181);
nor U12452 (N_12452,N_225,N_4492);
and U12453 (N_12453,N_2704,N_5710);
nand U12454 (N_12454,N_5093,N_4906);
nand U12455 (N_12455,N_2217,N_865);
or U12456 (N_12456,N_1770,N_1047);
xor U12457 (N_12457,N_4200,N_6185);
nor U12458 (N_12458,N_2163,N_3402);
and U12459 (N_12459,N_1993,N_4874);
nor U12460 (N_12460,N_6042,N_2237);
xor U12461 (N_12461,N_4281,N_3529);
and U12462 (N_12462,N_5194,N_4342);
or U12463 (N_12463,N_1029,N_1101);
nand U12464 (N_12464,N_3210,N_1412);
xor U12465 (N_12465,N_1142,N_2833);
nand U12466 (N_12466,N_5029,N_3036);
nand U12467 (N_12467,N_5437,N_2154);
xor U12468 (N_12468,N_6148,N_1754);
nand U12469 (N_12469,N_323,N_5720);
and U12470 (N_12470,N_4124,N_2234);
nor U12471 (N_12471,N_4695,N_1253);
and U12472 (N_12472,N_6167,N_3266);
or U12473 (N_12473,N_1187,N_235);
and U12474 (N_12474,N_4337,N_4500);
or U12475 (N_12475,N_5556,N_2650);
xnor U12476 (N_12476,N_3183,N_3317);
or U12477 (N_12477,N_3972,N_5442);
nor U12478 (N_12478,N_3768,N_5313);
xnor U12479 (N_12479,N_5998,N_2653);
or U12480 (N_12480,N_1857,N_1155);
nor U12481 (N_12481,N_4166,N_5241);
nor U12482 (N_12482,N_3109,N_1299);
or U12483 (N_12483,N_3328,N_4367);
xor U12484 (N_12484,N_6143,N_3490);
and U12485 (N_12485,N_391,N_5219);
or U12486 (N_12486,N_4313,N_3437);
or U12487 (N_12487,N_6072,N_787);
nand U12488 (N_12488,N_811,N_3024);
or U12489 (N_12489,N_5927,N_2608);
or U12490 (N_12490,N_1391,N_1963);
nor U12491 (N_12491,N_1510,N_6196);
nor U12492 (N_12492,N_2882,N_4327);
or U12493 (N_12493,N_3627,N_4995);
or U12494 (N_12494,N_3257,N_5123);
or U12495 (N_12495,N_1764,N_88);
and U12496 (N_12496,N_5830,N_4537);
xnor U12497 (N_12497,N_1980,N_3691);
xor U12498 (N_12498,N_6175,N_4154);
and U12499 (N_12499,N_2272,N_4229);
or U12500 (N_12500,N_7863,N_7903);
and U12501 (N_12501,N_9728,N_7161);
or U12502 (N_12502,N_8949,N_8134);
and U12503 (N_12503,N_7306,N_8273);
nor U12504 (N_12504,N_11888,N_7993);
nor U12505 (N_12505,N_8158,N_11996);
and U12506 (N_12506,N_9784,N_7788);
and U12507 (N_12507,N_7553,N_12180);
xor U12508 (N_12508,N_12326,N_10526);
or U12509 (N_12509,N_8796,N_9775);
or U12510 (N_12510,N_9703,N_6851);
nor U12511 (N_12511,N_9938,N_8027);
and U12512 (N_12512,N_7260,N_6555);
or U12513 (N_12513,N_12019,N_8636);
or U12514 (N_12514,N_6908,N_7873);
nor U12515 (N_12515,N_12241,N_11825);
nor U12516 (N_12516,N_8913,N_12108);
and U12517 (N_12517,N_10321,N_11165);
and U12518 (N_12518,N_10896,N_9425);
nor U12519 (N_12519,N_8190,N_7213);
or U12520 (N_12520,N_6865,N_6975);
and U12521 (N_12521,N_8309,N_11855);
and U12522 (N_12522,N_10612,N_6564);
nand U12523 (N_12523,N_8300,N_8264);
nor U12524 (N_12524,N_6658,N_11893);
nand U12525 (N_12525,N_10755,N_8645);
or U12526 (N_12526,N_11708,N_7732);
and U12527 (N_12527,N_9308,N_9674);
xor U12528 (N_12528,N_7527,N_7057);
nor U12529 (N_12529,N_8821,N_9699);
nand U12530 (N_12530,N_11842,N_8302);
nor U12531 (N_12531,N_8056,N_7678);
or U12532 (N_12532,N_9767,N_8472);
or U12533 (N_12533,N_7882,N_10318);
xor U12534 (N_12534,N_11523,N_6873);
or U12535 (N_12535,N_11617,N_10892);
and U12536 (N_12536,N_9087,N_8103);
nor U12537 (N_12537,N_11358,N_10508);
nor U12538 (N_12538,N_10699,N_8034);
xor U12539 (N_12539,N_9397,N_12018);
and U12540 (N_12540,N_12394,N_10846);
xor U12541 (N_12541,N_10197,N_8515);
or U12542 (N_12542,N_6271,N_11146);
and U12543 (N_12543,N_7190,N_11507);
and U12544 (N_12544,N_10930,N_12112);
xnor U12545 (N_12545,N_6956,N_7032);
nand U12546 (N_12546,N_8428,N_6938);
xor U12547 (N_12547,N_6573,N_7962);
and U12548 (N_12548,N_10009,N_8047);
or U12549 (N_12549,N_7270,N_9446);
nor U12550 (N_12550,N_12385,N_11900);
nand U12551 (N_12551,N_7567,N_6822);
or U12552 (N_12552,N_10064,N_11707);
xor U12553 (N_12553,N_11044,N_11001);
nand U12554 (N_12554,N_8492,N_10333);
xor U12555 (N_12555,N_6932,N_11593);
or U12556 (N_12556,N_11244,N_7243);
and U12557 (N_12557,N_6621,N_9141);
and U12558 (N_12558,N_8377,N_6713);
and U12559 (N_12559,N_9972,N_10817);
or U12560 (N_12560,N_11684,N_9891);
nor U12561 (N_12561,N_11154,N_10998);
and U12562 (N_12562,N_6628,N_7599);
nor U12563 (N_12563,N_12012,N_6878);
nand U12564 (N_12564,N_7214,N_11706);
or U12565 (N_12565,N_9478,N_10981);
xnor U12566 (N_12566,N_11841,N_7954);
nor U12567 (N_12567,N_7562,N_7172);
or U12568 (N_12568,N_8731,N_8261);
nor U12569 (N_12569,N_9820,N_6807);
or U12570 (N_12570,N_10608,N_12477);
nor U12571 (N_12571,N_6422,N_9762);
nand U12572 (N_12572,N_9244,N_7300);
and U12573 (N_12573,N_10701,N_11092);
nand U12574 (N_12574,N_11489,N_7807);
xnor U12575 (N_12575,N_6858,N_8125);
nand U12576 (N_12576,N_9963,N_11636);
xnor U12577 (N_12577,N_8280,N_9856);
nand U12578 (N_12578,N_10587,N_6836);
nand U12579 (N_12579,N_6425,N_7900);
nand U12580 (N_12580,N_12202,N_12115);
nand U12581 (N_12581,N_10779,N_7920);
or U12582 (N_12582,N_11347,N_6337);
or U12583 (N_12583,N_9804,N_12049);
xor U12584 (N_12584,N_11186,N_9682);
nand U12585 (N_12585,N_8298,N_11433);
nor U12586 (N_12586,N_9223,N_9509);
nand U12587 (N_12587,N_12045,N_7593);
nor U12588 (N_12588,N_11534,N_7842);
and U12589 (N_12589,N_6659,N_8849);
xor U12590 (N_12590,N_10213,N_10268);
and U12591 (N_12591,N_8421,N_10827);
nand U12592 (N_12592,N_9000,N_9603);
and U12593 (N_12593,N_11651,N_9324);
xor U12594 (N_12594,N_11149,N_8714);
and U12595 (N_12595,N_9677,N_6970);
and U12596 (N_12596,N_11206,N_11133);
or U12597 (N_12597,N_10121,N_9951);
and U12598 (N_12598,N_7649,N_8434);
nor U12599 (N_12599,N_12214,N_10852);
and U12600 (N_12600,N_8962,N_8170);
or U12601 (N_12601,N_8781,N_10055);
nand U12602 (N_12602,N_10799,N_7269);
nor U12603 (N_12603,N_7049,N_9095);
or U12604 (N_12604,N_10641,N_6579);
and U12605 (N_12605,N_6445,N_10254);
nor U12606 (N_12606,N_6281,N_7228);
xor U12607 (N_12607,N_12261,N_7196);
nand U12608 (N_12608,N_11387,N_7360);
or U12609 (N_12609,N_9633,N_12095);
nor U12610 (N_12610,N_6374,N_11025);
nor U12611 (N_12611,N_7240,N_11731);
xor U12612 (N_12612,N_7970,N_10617);
nand U12613 (N_12613,N_12316,N_7587);
nor U12614 (N_12614,N_9042,N_12175);
and U12615 (N_12615,N_9940,N_7852);
or U12616 (N_12616,N_8609,N_12395);
nor U12617 (N_12617,N_10992,N_6771);
nand U12618 (N_12618,N_10491,N_7054);
nand U12619 (N_12619,N_8892,N_10474);
or U12620 (N_12620,N_9165,N_11123);
nand U12621 (N_12621,N_10306,N_10730);
xor U12622 (N_12622,N_7722,N_8851);
or U12623 (N_12623,N_9368,N_7025);
nor U12624 (N_12624,N_12336,N_12472);
nand U12625 (N_12625,N_7639,N_10678);
nand U12626 (N_12626,N_6761,N_6663);
nand U12627 (N_12627,N_6400,N_7946);
nand U12628 (N_12628,N_9568,N_10842);
xor U12629 (N_12629,N_6845,N_9328);
nor U12630 (N_12630,N_11212,N_6636);
or U12631 (N_12631,N_7832,N_7891);
or U12632 (N_12632,N_7723,N_10910);
xor U12633 (N_12633,N_6720,N_11882);
or U12634 (N_12634,N_7089,N_9737);
and U12635 (N_12635,N_10336,N_11908);
or U12636 (N_12636,N_10780,N_11744);
or U12637 (N_12637,N_11267,N_10821);
or U12638 (N_12638,N_9730,N_7336);
xor U12639 (N_12639,N_9823,N_9024);
xnor U12640 (N_12640,N_6841,N_8551);
or U12641 (N_12641,N_12235,N_9011);
nor U12642 (N_12642,N_9203,N_11819);
and U12643 (N_12643,N_11868,N_11254);
nor U12644 (N_12644,N_7503,N_6256);
or U12645 (N_12645,N_7719,N_10300);
xnor U12646 (N_12646,N_7717,N_7795);
xnor U12647 (N_12647,N_12183,N_11571);
and U12648 (N_12648,N_11375,N_8409);
nor U12649 (N_12649,N_11549,N_10179);
or U12650 (N_12650,N_7850,N_7684);
or U12651 (N_12651,N_12403,N_10099);
xnor U12652 (N_12652,N_6984,N_10411);
nand U12653 (N_12653,N_8932,N_12133);
and U12654 (N_12654,N_10996,N_9378);
nor U12655 (N_12655,N_11453,N_10890);
nor U12656 (N_12656,N_6541,N_11561);
or U12657 (N_12657,N_7446,N_11366);
xnor U12658 (N_12658,N_12090,N_12460);
or U12659 (N_12659,N_12282,N_6995);
nor U12660 (N_12660,N_8358,N_8328);
and U12661 (N_12661,N_8585,N_8933);
and U12662 (N_12662,N_11746,N_11289);
nand U12663 (N_12663,N_6405,N_9510);
and U12664 (N_12664,N_12493,N_11880);
or U12665 (N_12665,N_10923,N_7944);
xnor U12666 (N_12666,N_7739,N_9104);
or U12667 (N_12667,N_8343,N_9101);
nand U12668 (N_12668,N_8805,N_7131);
nand U12669 (N_12669,N_7072,N_8099);
nand U12670 (N_12670,N_10223,N_9868);
nand U12671 (N_12671,N_6593,N_11396);
and U12672 (N_12672,N_7620,N_11851);
or U12673 (N_12673,N_10797,N_8133);
and U12674 (N_12674,N_10100,N_9233);
nand U12675 (N_12675,N_6892,N_12343);
or U12676 (N_12676,N_7514,N_12161);
and U12677 (N_12677,N_10758,N_8919);
or U12678 (N_12678,N_10997,N_7576);
or U12679 (N_12679,N_7708,N_10078);
and U12680 (N_12680,N_11365,N_8896);
nand U12681 (N_12681,N_11693,N_9648);
or U12682 (N_12682,N_11831,N_6904);
or U12683 (N_12683,N_10528,N_6302);
nand U12684 (N_12684,N_10177,N_8397);
or U12685 (N_12685,N_6429,N_7542);
and U12686 (N_12686,N_9110,N_9172);
or U12687 (N_12687,N_9157,N_7835);
or U12688 (N_12688,N_8172,N_10230);
and U12689 (N_12689,N_12266,N_7074);
nor U12690 (N_12690,N_8114,N_8242);
and U12691 (N_12691,N_7656,N_7860);
nand U12692 (N_12692,N_11427,N_7184);
and U12693 (N_12693,N_7893,N_9337);
xor U12694 (N_12694,N_8680,N_11100);
and U12695 (N_12695,N_8366,N_11596);
or U12696 (N_12696,N_9596,N_10976);
nor U12697 (N_12697,N_12197,N_8149);
nor U12698 (N_12698,N_7023,N_7353);
xor U12699 (N_12699,N_11095,N_8578);
xnor U12700 (N_12700,N_10548,N_10317);
nor U12701 (N_12701,N_7142,N_12066);
or U12702 (N_12702,N_10119,N_11160);
xnor U12703 (N_12703,N_11899,N_11995);
xnor U12704 (N_12704,N_11203,N_10215);
nor U12705 (N_12705,N_9017,N_12354);
xnor U12706 (N_12706,N_8840,N_8670);
nor U12707 (N_12707,N_10253,N_7346);
xnor U12708 (N_12708,N_9592,N_9558);
and U12709 (N_12709,N_8323,N_7486);
nor U12710 (N_12710,N_8425,N_8598);
nor U12711 (N_12711,N_10598,N_10171);
or U12712 (N_12712,N_12335,N_8610);
nand U12713 (N_12713,N_11268,N_11921);
and U12714 (N_12714,N_11760,N_6766);
and U12715 (N_12715,N_9598,N_8757);
nand U12716 (N_12716,N_9560,N_11306);
or U12717 (N_12717,N_9247,N_7153);
and U12718 (N_12718,N_6787,N_11530);
xnor U12719 (N_12719,N_6708,N_8723);
xnor U12720 (N_12720,N_9915,N_8649);
and U12721 (N_12721,N_8550,N_7417);
nand U12722 (N_12722,N_7868,N_10676);
and U12723 (N_12723,N_6987,N_11350);
nand U12724 (N_12724,N_11015,N_8930);
xnor U12725 (N_12725,N_10979,N_6947);
nand U12726 (N_12726,N_9107,N_8613);
and U12727 (N_12727,N_10822,N_11259);
nand U12728 (N_12728,N_9202,N_6307);
or U12729 (N_12729,N_9710,N_7851);
nor U12730 (N_12730,N_10515,N_12439);
and U12731 (N_12731,N_9577,N_8245);
xnor U12732 (N_12732,N_11055,N_9576);
nor U12733 (N_12733,N_6781,N_10594);
or U12734 (N_12734,N_7741,N_9372);
xnor U12735 (N_12735,N_8235,N_10949);
xor U12736 (N_12736,N_8712,N_8766);
nand U12737 (N_12737,N_10487,N_7932);
nand U12738 (N_12738,N_9082,N_9062);
nor U12739 (N_12739,N_8935,N_9160);
nand U12740 (N_12740,N_8909,N_11935);
or U12741 (N_12741,N_9222,N_11543);
or U12742 (N_12742,N_7472,N_9718);
nor U12743 (N_12743,N_11733,N_9206);
nand U12744 (N_12744,N_8478,N_12285);
and U12745 (N_12745,N_9459,N_9394);
or U12746 (N_12746,N_10742,N_11012);
or U12747 (N_12747,N_11270,N_12069);
and U12748 (N_12748,N_10689,N_7922);
xnor U12749 (N_12749,N_8316,N_7767);
or U12750 (N_12750,N_10109,N_7134);
nand U12751 (N_12751,N_7766,N_9620);
nor U12752 (N_12752,N_6389,N_8648);
xnor U12753 (N_12753,N_9252,N_7056);
nand U12754 (N_12754,N_10694,N_7523);
and U12755 (N_12755,N_8278,N_8406);
nand U12756 (N_12756,N_10589,N_8622);
nand U12757 (N_12757,N_8755,N_10621);
or U12758 (N_12758,N_8485,N_12089);
nor U12759 (N_12759,N_8600,N_6409);
and U12760 (N_12760,N_7864,N_7425);
or U12761 (N_12761,N_9574,N_7955);
and U12762 (N_12762,N_11950,N_9589);
nor U12763 (N_12763,N_7156,N_7249);
and U12764 (N_12764,N_6876,N_7068);
nor U12765 (N_12765,N_6538,N_9382);
nor U12766 (N_12766,N_9586,N_11579);
and U12767 (N_12767,N_9117,N_6731);
nand U12768 (N_12768,N_7121,N_7365);
and U12769 (N_12769,N_10952,N_10373);
nand U12770 (N_12770,N_11457,N_10565);
and U12771 (N_12771,N_12368,N_10244);
nand U12772 (N_12772,N_11713,N_6830);
nor U12773 (N_12773,N_8524,N_8038);
or U12774 (N_12774,N_6812,N_6714);
or U12775 (N_12775,N_12130,N_9119);
and U12776 (N_12776,N_11305,N_7244);
nand U12777 (N_12777,N_6755,N_12149);
nand U12778 (N_12778,N_9213,N_11009);
nor U12779 (N_12779,N_11937,N_9814);
xor U12780 (N_12780,N_6253,N_7980);
nor U12781 (N_12781,N_10756,N_7449);
nand U12782 (N_12782,N_8546,N_7536);
nand U12783 (N_12783,N_11526,N_11637);
nor U12784 (N_12784,N_6428,N_11456);
and U12785 (N_12785,N_9237,N_7433);
nor U12786 (N_12786,N_9068,N_6375);
xnor U12787 (N_12787,N_11262,N_9356);
xnor U12788 (N_12788,N_12111,N_10953);
and U12789 (N_12789,N_11284,N_11234);
xnor U12790 (N_12790,N_11797,N_8972);
and U12791 (N_12791,N_6292,N_8496);
or U12792 (N_12792,N_6997,N_9114);
and U12793 (N_12793,N_12377,N_9601);
nand U12794 (N_12794,N_9112,N_8393);
nand U12795 (N_12795,N_9754,N_10811);
and U12796 (N_12796,N_9961,N_7781);
nand U12797 (N_12797,N_9018,N_9014);
nand U12798 (N_12798,N_12390,N_12297);
and U12799 (N_12799,N_8816,N_7841);
or U12800 (N_12800,N_9216,N_7402);
nor U12801 (N_12801,N_9201,N_7742);
and U12802 (N_12802,N_6570,N_6924);
and U12803 (N_12803,N_11339,N_8918);
or U12804 (N_12804,N_8463,N_10163);
nand U12805 (N_12805,N_8016,N_9725);
nand U12806 (N_12806,N_10521,N_10299);
nand U12807 (N_12807,N_9281,N_6453);
nor U12808 (N_12808,N_8824,N_10691);
or U12809 (N_12809,N_11475,N_8642);
or U12810 (N_12810,N_10314,N_7694);
or U12811 (N_12811,N_12432,N_8846);
or U12812 (N_12812,N_7256,N_11418);
and U12813 (N_12813,N_9834,N_7927);
xor U12814 (N_12814,N_7798,N_10205);
or U12815 (N_12815,N_9531,N_8415);
nor U12816 (N_12816,N_7330,N_9264);
nor U12817 (N_12817,N_7203,N_11681);
and U12818 (N_12818,N_6928,N_9266);
nand U12819 (N_12819,N_10518,N_12032);
xor U12820 (N_12820,N_9918,N_10172);
nor U12821 (N_12821,N_8223,N_9713);
nand U12822 (N_12822,N_10147,N_7357);
xor U12823 (N_12823,N_8961,N_10486);
nand U12824 (N_12824,N_10227,N_7102);
nand U12825 (N_12825,N_7200,N_7125);
nor U12826 (N_12826,N_12370,N_8845);
or U12827 (N_12827,N_10900,N_10266);
or U12828 (N_12828,N_6383,N_9003);
or U12829 (N_12829,N_8355,N_10005);
xor U12830 (N_12830,N_7199,N_9414);
xor U12831 (N_12831,N_7122,N_10361);
nand U12832 (N_12832,N_9341,N_10828);
nand U12833 (N_12833,N_9276,N_10281);
and U12834 (N_12834,N_10395,N_12144);
nand U12835 (N_12835,N_7375,N_9608);
or U12836 (N_12836,N_11582,N_8043);
or U12837 (N_12837,N_9225,N_7460);
nor U12838 (N_12838,N_9240,N_12451);
nand U12839 (N_12839,N_11255,N_10184);
nand U12840 (N_12840,N_7379,N_7556);
nand U12841 (N_12841,N_10818,N_11553);
nand U12842 (N_12842,N_9518,N_9283);
or U12843 (N_12843,N_10960,N_11173);
nand U12844 (N_12844,N_11907,N_6614);
xor U12845 (N_12845,N_11739,N_7869);
xnor U12846 (N_12846,N_8122,N_7947);
xor U12847 (N_12847,N_12152,N_6419);
nor U12848 (N_12848,N_8959,N_7515);
or U12849 (N_12849,N_6915,N_8014);
or U12850 (N_12850,N_10697,N_11600);
xnor U12851 (N_12851,N_6486,N_10935);
or U12852 (N_12852,N_10804,N_6922);
xnor U12853 (N_12853,N_11291,N_11266);
xor U12854 (N_12854,N_11522,N_12492);
nand U12855 (N_12855,N_9884,N_10854);
nor U12856 (N_12856,N_8678,N_6828);
or U12857 (N_12857,N_11020,N_11410);
xor U12858 (N_12858,N_12084,N_9824);
and U12859 (N_12859,N_10315,N_9641);
xor U12860 (N_12860,N_10661,N_9005);
or U12861 (N_12861,N_9569,N_7394);
xnor U12862 (N_12862,N_10083,N_10127);
nand U12863 (N_12863,N_6349,N_8558);
or U12864 (N_12864,N_10012,N_6480);
and U12865 (N_12865,N_10036,N_10824);
nor U12866 (N_12866,N_7296,N_11506);
nor U12867 (N_12867,N_7288,N_9178);
xor U12868 (N_12868,N_8522,N_12396);
nor U12869 (N_12869,N_8336,N_8454);
or U12870 (N_12870,N_12038,N_11898);
nor U12871 (N_12871,N_11346,N_6276);
or U12872 (N_12872,N_11780,N_6844);
nor U12873 (N_12873,N_6441,N_8722);
or U12874 (N_12874,N_8468,N_12230);
xnor U12875 (N_12875,N_12470,N_12123);
xor U12876 (N_12876,N_10603,N_10313);
and U12877 (N_12877,N_10042,N_11927);
nand U12878 (N_12878,N_10543,N_9214);
or U12879 (N_12879,N_11791,N_6634);
nor U12880 (N_12880,N_11429,N_6916);
and U12881 (N_12881,N_10047,N_7912);
nand U12882 (N_12882,N_11918,N_12309);
nand U12883 (N_12883,N_12146,N_8071);
nand U12884 (N_12884,N_6682,N_11945);
and U12885 (N_12885,N_6305,N_10525);
xnor U12886 (N_12886,N_10035,N_7455);
xnor U12887 (N_12887,N_7761,N_7311);
and U12888 (N_12888,N_11784,N_8976);
or U12889 (N_12889,N_7176,N_7602);
nand U12890 (N_12890,N_10708,N_8052);
nand U12891 (N_12891,N_10681,N_9353);
xnor U12892 (N_12892,N_9670,N_7398);
xor U12893 (N_12893,N_12176,N_11499);
nand U12894 (N_12894,N_7933,N_11829);
nor U12895 (N_12895,N_6484,N_8254);
or U12896 (N_12896,N_12221,N_12365);
nor U12897 (N_12897,N_6958,N_11360);
xor U12898 (N_12898,N_6750,N_7401);
nand U12899 (N_12899,N_10483,N_12189);
xnor U12900 (N_12900,N_10798,N_9319);
and U12901 (N_12901,N_12359,N_10413);
xor U12902 (N_12902,N_9188,N_10229);
and U12903 (N_12903,N_7743,N_6291);
xnor U12904 (N_12904,N_7259,N_11675);
nand U12905 (N_12905,N_10938,N_9691);
nand U12906 (N_12906,N_10611,N_12314);
and U12907 (N_12907,N_11743,N_8605);
nand U12908 (N_12908,N_7528,N_6933);
and U12909 (N_12909,N_6393,N_7611);
nand U12910 (N_12910,N_12148,N_10941);
nand U12911 (N_12911,N_6816,N_9159);
xor U12912 (N_12912,N_10712,N_10914);
or U12913 (N_12913,N_10540,N_9155);
nand U12914 (N_12914,N_7726,N_8542);
nand U12915 (N_12915,N_9423,N_10680);
nand U12916 (N_12916,N_12209,N_11049);
and U12917 (N_12917,N_10123,N_8691);
nor U12918 (N_12918,N_8943,N_8807);
nand U12919 (N_12919,N_10027,N_11860);
nor U12920 (N_12920,N_7294,N_7356);
xnor U12921 (N_12921,N_9991,N_11913);
or U12922 (N_12922,N_9395,N_12005);
and U12923 (N_12923,N_7565,N_10326);
nand U12924 (N_12924,N_6369,N_8102);
or U12925 (N_12925,N_9563,N_7909);
nor U12926 (N_12926,N_9289,N_8958);
and U12927 (N_12927,N_10634,N_9241);
nor U12928 (N_12928,N_8012,N_11157);
nor U12929 (N_12929,N_9354,N_8387);
and U12930 (N_12930,N_10718,N_8954);
xor U12931 (N_12931,N_10416,N_10874);
and U12932 (N_12932,N_12070,N_9817);
and U12933 (N_12933,N_8437,N_9841);
xnor U12934 (N_12934,N_9452,N_7039);
nand U12935 (N_12935,N_10902,N_7079);
xor U12936 (N_12936,N_10125,N_11283);
and U12937 (N_12937,N_8775,N_8562);
xnor U12938 (N_12938,N_8720,N_6410);
xnor U12939 (N_12939,N_9664,N_6528);
and U12940 (N_12940,N_7283,N_9148);
nor U12941 (N_12941,N_9708,N_8509);
xor U12942 (N_12942,N_10692,N_8279);
or U12943 (N_12943,N_6454,N_11403);
and U12944 (N_12944,N_10011,N_8615);
and U12945 (N_12945,N_6540,N_9086);
nor U12946 (N_12946,N_8380,N_8684);
or U12947 (N_12947,N_10776,N_6358);
or U12948 (N_12948,N_10867,N_6834);
nor U12949 (N_12949,N_7448,N_12346);
or U12950 (N_12950,N_7818,N_11464);
or U12951 (N_12951,N_11090,N_11354);
xnor U12952 (N_12952,N_12433,N_11672);
nand U12953 (N_12953,N_9795,N_11144);
nor U12954 (N_12954,N_10145,N_11147);
nor U12955 (N_12955,N_8064,N_7555);
xnor U12956 (N_12956,N_6443,N_9876);
nand U12957 (N_12957,N_7670,N_10576);
nor U12958 (N_12958,N_10664,N_7114);
and U12959 (N_12959,N_9654,N_7445);
nand U12960 (N_12960,N_12356,N_9440);
xnor U12961 (N_12961,N_9719,N_7547);
nand U12962 (N_12962,N_11424,N_9275);
nor U12963 (N_12963,N_9984,N_11207);
xnor U12964 (N_12964,N_6638,N_8104);
and U12965 (N_12965,N_10559,N_8674);
xnor U12966 (N_12966,N_9389,N_8221);
and U12967 (N_12967,N_8140,N_12210);
and U12968 (N_12968,N_7790,N_7958);
nor U12969 (N_12969,N_10506,N_7277);
nor U12970 (N_12970,N_9567,N_11202);
and U12971 (N_12971,N_8743,N_8867);
xor U12972 (N_12972,N_12384,N_10522);
xor U12973 (N_12973,N_11053,N_9717);
nand U12974 (N_12974,N_6299,N_8639);
xnor U12975 (N_12975,N_9438,N_9959);
nand U12976 (N_12976,N_7453,N_11341);
and U12977 (N_12977,N_10016,N_10865);
xnor U12978 (N_12978,N_6567,N_10880);
xnor U12979 (N_12979,N_7118,N_9617);
and U12980 (N_12980,N_9367,N_11324);
nor U12981 (N_12981,N_11171,N_11963);
or U12982 (N_12982,N_7133,N_7227);
nand U12983 (N_12983,N_8009,N_8695);
or U12984 (N_12984,N_7917,N_8862);
nand U12985 (N_12985,N_6348,N_11795);
or U12986 (N_12986,N_8378,N_9538);
and U12987 (N_12987,N_7937,N_8017);
and U12988 (N_12988,N_8443,N_9547);
nor U12989 (N_12989,N_10248,N_8283);
or U12990 (N_12990,N_11348,N_10695);
or U12991 (N_12991,N_10320,N_8157);
and U12992 (N_12992,N_7221,N_8269);
nor U12993 (N_12993,N_7724,N_12061);
and U12994 (N_12994,N_6804,N_12497);
xor U12995 (N_12995,N_10499,N_10734);
or U12996 (N_12996,N_10717,N_6972);
xnor U12997 (N_12997,N_6371,N_10459);
nand U12998 (N_12998,N_6357,N_7299);
xnor U12999 (N_12999,N_11197,N_11849);
xnor U13000 (N_13000,N_10157,N_11537);
and U13001 (N_13001,N_9714,N_12388);
xnor U13002 (N_13002,N_9473,N_9655);
and U13003 (N_13003,N_9145,N_10872);
or U13004 (N_13004,N_10944,N_10106);
nor U13005 (N_13005,N_11872,N_12106);
nor U13006 (N_13006,N_6774,N_9236);
nand U13007 (N_13007,N_11441,N_7302);
or U13008 (N_13008,N_11071,N_10688);
or U13009 (N_13009,N_12179,N_9744);
or U13010 (N_13010,N_9849,N_8537);
nand U13011 (N_13011,N_11303,N_11492);
or U13012 (N_13012,N_12438,N_9445);
or U13013 (N_13013,N_10477,N_10294);
xor U13014 (N_13014,N_9712,N_8469);
nand U13015 (N_13015,N_7544,N_7837);
and U13016 (N_13016,N_12340,N_12236);
nand U13017 (N_13017,N_8422,N_6953);
nor U13018 (N_13018,N_6625,N_10017);
or U13019 (N_13019,N_9061,N_11225);
xnor U13020 (N_13020,N_9535,N_8597);
nand U13021 (N_13021,N_10861,N_10975);
nor U13022 (N_13022,N_9422,N_9773);
and U13023 (N_13023,N_7540,N_9702);
nand U13024 (N_13024,N_12273,N_9671);
xor U13025 (N_13025,N_8966,N_9537);
nand U13026 (N_13026,N_6402,N_11538);
nor U13027 (N_13027,N_8555,N_10242);
or U13028 (N_13028,N_9152,N_11968);
and U13029 (N_13029,N_9479,N_8385);
nand U13030 (N_13030,N_6961,N_10087);
xnor U13031 (N_13031,N_8771,N_12139);
or U13032 (N_13032,N_10803,N_11551);
and U13033 (N_13033,N_7672,N_10497);
and U13034 (N_13034,N_7006,N_10580);
xnor U13035 (N_13035,N_7451,N_11077);
xnor U13036 (N_13036,N_12348,N_9905);
or U13037 (N_13037,N_8595,N_9584);
xor U13038 (N_13038,N_9854,N_8718);
xnor U13039 (N_13039,N_6855,N_7895);
or U13040 (N_13040,N_6679,N_12469);
and U13041 (N_13041,N_11576,N_11897);
or U13042 (N_13042,N_6346,N_8220);
or U13043 (N_13043,N_8689,N_11714);
nand U13044 (N_13044,N_11550,N_6661);
xnor U13045 (N_13045,N_9182,N_7042);
nand U13046 (N_13046,N_9365,N_11905);
nand U13047 (N_13047,N_9821,N_8465);
nor U13048 (N_13048,N_8942,N_9630);
xor U13049 (N_13049,N_10563,N_7491);
or U13050 (N_13050,N_12042,N_7972);
and U13051 (N_13051,N_9629,N_11136);
nor U13052 (N_13052,N_7612,N_8814);
xnor U13053 (N_13053,N_11616,N_10725);
xor U13054 (N_13054,N_10810,N_8398);
nor U13055 (N_13055,N_12298,N_9889);
nand U13056 (N_13056,N_8590,N_7348);
and U13057 (N_13057,N_11926,N_7280);
nand U13058 (N_13058,N_7994,N_8521);
nor U13059 (N_13059,N_9698,N_12104);
nor U13060 (N_13060,N_10840,N_7193);
nand U13061 (N_13061,N_10120,N_9043);
and U13062 (N_13062,N_9983,N_6355);
or U13063 (N_13063,N_9830,N_7660);
and U13064 (N_13064,N_11639,N_6911);
and U13065 (N_13065,N_11686,N_9852);
nand U13066 (N_13066,N_8182,N_8480);
nand U13067 (N_13067,N_12416,N_10899);
nand U13068 (N_13068,N_8081,N_8889);
xnor U13069 (N_13069,N_8074,N_8878);
nand U13070 (N_13070,N_8395,N_9667);
nand U13071 (N_13071,N_11170,N_6427);
xor U13072 (N_13072,N_11749,N_9809);
nand U13073 (N_13073,N_8493,N_9621);
xnor U13074 (N_13074,N_6379,N_11299);
and U13075 (N_13075,N_9872,N_7151);
and U13076 (N_13076,N_8100,N_8487);
nor U13077 (N_13077,N_8643,N_11021);
or U13078 (N_13078,N_11485,N_6539);
nand U13079 (N_13079,N_9226,N_9907);
nor U13080 (N_13080,N_10370,N_10358);
or U13081 (N_13081,N_12260,N_10945);
nand U13082 (N_13082,N_8367,N_8621);
and U13083 (N_13083,N_6386,N_8523);
and U13084 (N_13084,N_11112,N_9035);
nand U13085 (N_13085,N_9517,N_11258);
or U13086 (N_13086,N_10637,N_10115);
or U13087 (N_13087,N_10597,N_8364);
or U13088 (N_13088,N_12268,N_11753);
or U13089 (N_13089,N_7710,N_6862);
nand U13090 (N_13090,N_9771,N_8682);
nor U13091 (N_13091,N_11114,N_6959);
and U13092 (N_13092,N_9683,N_11177);
or U13093 (N_13093,N_12328,N_10307);
or U13094 (N_13094,N_9858,N_11952);
nor U13095 (N_13095,N_10095,N_7019);
nor U13096 (N_13096,N_12047,N_11957);
xor U13097 (N_13097,N_12484,N_9839);
or U13098 (N_13098,N_9314,N_6993);
nor U13099 (N_13099,N_9595,N_8022);
xor U13100 (N_13100,N_11574,N_10156);
nand U13101 (N_13101,N_8784,N_6704);
and U13102 (N_13102,N_10330,N_11653);
nor U13103 (N_13103,N_11500,N_6336);
and U13104 (N_13104,N_10585,N_8508);
xnor U13105 (N_13105,N_12218,N_6387);
xnor U13106 (N_13106,N_6727,N_7885);
or U13107 (N_13107,N_9229,N_11246);
xnor U13108 (N_13108,N_10832,N_8113);
and U13109 (N_13109,N_10626,N_10409);
or U13110 (N_13110,N_6849,N_11452);
nor U13111 (N_13111,N_8864,N_10288);
nand U13112 (N_13112,N_7846,N_9638);
nor U13113 (N_13113,N_7906,N_10869);
and U13114 (N_13114,N_10607,N_6806);
or U13115 (N_13115,N_6974,N_11302);
xor U13116 (N_13116,N_9653,N_11910);
nand U13117 (N_13117,N_7709,N_6746);
and U13118 (N_13118,N_11712,N_11028);
nor U13119 (N_13119,N_10783,N_8737);
nand U13120 (N_13120,N_8618,N_8640);
xor U13121 (N_13121,N_12204,N_11236);
and U13122 (N_13122,N_8351,N_11877);
nand U13123 (N_13123,N_10124,N_6381);
and U13124 (N_13124,N_6606,N_9146);
nand U13125 (N_13125,N_7859,N_8068);
or U13126 (N_13126,N_11959,N_10329);
xor U13127 (N_13127,N_6986,N_7358);
nand U13128 (N_13128,N_8249,N_6697);
and U13129 (N_13129,N_9009,N_8710);
xor U13130 (N_13130,N_10829,N_6610);
nand U13131 (N_13131,N_8599,N_8817);
nand U13132 (N_13132,N_8356,N_11556);
xor U13133 (N_13133,N_6925,N_9065);
nor U13134 (N_13134,N_9588,N_11252);
nand U13135 (N_13135,N_9811,N_7136);
nor U13136 (N_13136,N_12475,N_10774);
nor U13137 (N_13137,N_11759,N_8810);
nor U13138 (N_13138,N_11085,N_10451);
xor U13139 (N_13139,N_9193,N_8654);
nand U13140 (N_13140,N_7194,N_9258);
xor U13141 (N_13141,N_9657,N_11230);
nor U13142 (N_13142,N_8083,N_7516);
nor U13143 (N_13143,N_11158,N_6937);
and U13144 (N_13144,N_11478,N_8899);
nand U13145 (N_13145,N_6251,N_11376);
nor U13146 (N_13146,N_8226,N_10424);
or U13147 (N_13147,N_7340,N_11717);
nor U13148 (N_13148,N_6740,N_11026);
or U13149 (N_13149,N_11181,N_10619);
nor U13150 (N_13150,N_8863,N_11139);
or U13151 (N_13151,N_12238,N_8130);
and U13152 (N_13152,N_11756,N_9282);
xnor U13153 (N_13153,N_11106,N_10399);
nand U13154 (N_13154,N_9516,N_11205);
nor U13155 (N_13155,N_6895,N_10539);
and U13156 (N_13156,N_11887,N_11994);
nand U13157 (N_13157,N_10238,N_6776);
xnor U13158 (N_13158,N_9556,N_11034);
nor U13159 (N_13159,N_7866,N_9038);
nand U13160 (N_13160,N_12292,N_9920);
nand U13161 (N_13161,N_9929,N_7816);
or U13162 (N_13162,N_7347,N_7480);
and U13163 (N_13163,N_6784,N_7812);
nand U13164 (N_13164,N_12031,N_8123);
nor U13165 (N_13165,N_7548,N_9257);
nor U13166 (N_13166,N_9694,N_10898);
and U13167 (N_13167,N_8266,N_10167);
xor U13168 (N_13168,N_9679,N_10995);
xnor U13169 (N_13169,N_11271,N_11175);
nor U13170 (N_13170,N_6852,N_9302);
or U13171 (N_13171,N_10081,N_6971);
nand U13172 (N_13172,N_9100,N_7648);
nor U13173 (N_13173,N_8531,N_12002);
and U13174 (N_13174,N_7875,N_10764);
nor U13175 (N_13175,N_8105,N_9261);
and U13176 (N_13176,N_10787,N_10324);
or U13177 (N_13177,N_10670,N_8676);
or U13178 (N_13178,N_10428,N_6903);
or U13179 (N_13179,N_9774,N_8055);
and U13180 (N_13180,N_7292,N_6338);
or U13181 (N_13181,N_6717,N_8563);
or U13182 (N_13182,N_8430,N_11690);
nor U13183 (N_13183,N_10398,N_8007);
nor U13184 (N_13184,N_9122,N_8106);
xnor U13185 (N_13185,N_8341,N_10164);
nor U13186 (N_13186,N_10978,N_10133);
and U13187 (N_13187,N_10505,N_10922);
nand U13188 (N_13188,N_6690,N_7506);
or U13189 (N_13189,N_6507,N_8461);
and U13190 (N_13190,N_8977,N_9085);
nand U13191 (N_13191,N_7178,N_7380);
xor U13192 (N_13192,N_11673,N_9792);
nand U13193 (N_13193,N_6687,N_7422);
nand U13194 (N_13194,N_6824,N_6498);
or U13195 (N_13195,N_7144,N_6382);
or U13196 (N_13196,N_7138,N_6864);
xor U13197 (N_13197,N_12147,N_10432);
or U13198 (N_13198,N_9041,N_11909);
xor U13199 (N_13199,N_10350,N_10355);
nand U13200 (N_13200,N_11509,N_9964);
nand U13201 (N_13201,N_7000,N_11127);
nor U13202 (N_13202,N_7374,N_7483);
nand U13203 (N_13203,N_12342,N_11495);
or U13204 (N_13204,N_8347,N_8253);
nor U13205 (N_13205,N_9286,N_10478);
and U13206 (N_13206,N_10773,N_10961);
or U13207 (N_13207,N_8873,N_12225);
nand U13208 (N_13208,N_9838,N_11991);
or U13209 (N_13209,N_9893,N_11732);
nor U13210 (N_13210,N_8625,N_11741);
nor U13211 (N_13211,N_10075,N_9748);
nor U13212 (N_13212,N_11546,N_7919);
nand U13213 (N_13213,N_6316,N_10039);
nand U13214 (N_13214,N_11392,N_6891);
and U13215 (N_13215,N_7235,N_11914);
xnor U13216 (N_13216,N_10928,N_6308);
nor U13217 (N_13217,N_7517,N_9486);
xnor U13218 (N_13218,N_10916,N_7800);
xnor U13219 (N_13219,N_8156,N_7275);
nor U13220 (N_13220,N_11990,N_6258);
and U13221 (N_13221,N_9533,N_7388);
and U13222 (N_13222,N_6782,N_7787);
and U13223 (N_13223,N_11562,N_7434);
xor U13224 (N_13224,N_7551,N_11985);
nand U13225 (N_13225,N_7165,N_6923);
xor U13226 (N_13226,N_7096,N_11697);
or U13227 (N_13227,N_8037,N_7982);
nor U13228 (N_13228,N_8445,N_9140);
xnor U13229 (N_13229,N_11666,N_7693);
and U13230 (N_13230,N_6324,N_6398);
or U13231 (N_13231,N_9545,N_12422);
nand U13232 (N_13232,N_8690,N_7034);
xnor U13233 (N_13233,N_10901,N_8632);
xor U13234 (N_13234,N_9739,N_8424);
nand U13235 (N_13235,N_7105,N_8286);
nand U13236 (N_13236,N_9549,N_10636);
nor U13237 (N_13237,N_7755,N_12455);
nor U13238 (N_13238,N_6549,N_11332);
xor U13239 (N_13239,N_9171,N_7894);
nor U13240 (N_13240,N_9358,N_8019);
or U13241 (N_13241,N_12310,N_12263);
xor U13242 (N_13242,N_11762,N_11062);
nor U13243 (N_13243,N_7582,N_7845);
xor U13244 (N_13244,N_8659,N_10554);
xor U13245 (N_13245,N_7478,N_9736);
and U13246 (N_13246,N_8724,N_6500);
xnor U13247 (N_13247,N_6848,N_7774);
nand U13248 (N_13248,N_8575,N_7504);
xnor U13249 (N_13249,N_9898,N_9903);
and U13250 (N_13250,N_11450,N_7413);
nor U13251 (N_13251,N_6289,N_8345);
xnor U13252 (N_13252,N_8809,N_7078);
nor U13253 (N_13253,N_12417,N_8386);
or U13254 (N_13254,N_12251,N_12239);
and U13255 (N_13255,N_11035,N_10423);
or U13256 (N_13256,N_6263,N_10040);
nand U13257 (N_13257,N_8672,N_7432);
nand U13258 (N_13258,N_12226,N_12311);
nand U13259 (N_13259,N_6461,N_8788);
and U13260 (N_13260,N_11565,N_8411);
nor U13261 (N_13261,N_6655,N_11874);
nand U13262 (N_13262,N_12288,N_7844);
nor U13263 (N_13263,N_7470,N_7532);
xnor U13264 (N_13264,N_12064,N_11242);
or U13265 (N_13265,N_11382,N_11328);
nand U13266 (N_13266,N_6359,N_8311);
nand U13267 (N_13267,N_7753,N_7654);
and U13268 (N_13268,N_10656,N_9279);
or U13269 (N_13269,N_10628,N_10993);
nand U13270 (N_13270,N_7126,N_8936);
and U13271 (N_13271,N_10484,N_11287);
and U13272 (N_13272,N_12252,N_9944);
or U13273 (N_13273,N_9541,N_10674);
nand U13274 (N_13274,N_8830,N_11645);
nor U13275 (N_13275,N_11293,N_6442);
and U13276 (N_13276,N_7643,N_6722);
and U13277 (N_13277,N_10650,N_7746);
nand U13278 (N_13278,N_10750,N_8301);
xor U13279 (N_13279,N_10102,N_6571);
and U13280 (N_13280,N_9293,N_11037);
or U13281 (N_13281,N_10384,N_8162);
or U13282 (N_13282,N_10561,N_9740);
nor U13283 (N_13283,N_8527,N_7103);
or U13284 (N_13284,N_11688,N_12375);
xnor U13285 (N_13285,N_8635,N_9344);
nor U13286 (N_13286,N_7120,N_11992);
nor U13287 (N_13287,N_12046,N_6913);
or U13288 (N_13288,N_10331,N_6802);
or U13289 (N_13289,N_8511,N_8126);
xor U13290 (N_13290,N_6582,N_6274);
and U13291 (N_13291,N_6264,N_10285);
nor U13292 (N_13292,N_7309,N_6818);
nor U13293 (N_13293,N_9958,N_7395);
and U13294 (N_13294,N_12401,N_7691);
nand U13295 (N_13295,N_11863,N_10029);
or U13296 (N_13296,N_7647,N_8944);
xnor U13297 (N_13297,N_7674,N_7669);
or U13298 (N_13298,N_12181,N_8951);
and U13299 (N_13299,N_11359,N_11169);
nand U13300 (N_13300,N_8066,N_7573);
nand U13301 (N_13301,N_9093,N_10668);
xnor U13302 (N_13302,N_8359,N_10196);
and U13303 (N_13303,N_11235,N_12072);
or U13304 (N_13304,N_7692,N_6736);
nor U13305 (N_13305,N_7224,N_10054);
nor U13306 (N_13306,N_8138,N_10207);
and U13307 (N_13307,N_7921,N_7116);
nor U13308 (N_13308,N_6688,N_10796);
or U13309 (N_13309,N_12205,N_7929);
or U13310 (N_13310,N_10392,N_7087);
xnor U13311 (N_13311,N_12065,N_7303);
xor U13312 (N_13312,N_9495,N_6265);
nand U13313 (N_13313,N_9626,N_7285);
nand U13314 (N_13314,N_11461,N_11521);
and U13315 (N_13315,N_9900,N_7828);
xnor U13316 (N_13316,N_6607,N_6739);
nor U13317 (N_13317,N_10419,N_7519);
nor U13318 (N_13318,N_6477,N_8666);
xor U13319 (N_13319,N_7400,N_7487);
and U13320 (N_13320,N_12331,N_12332);
xor U13321 (N_13321,N_7770,N_8079);
or U13322 (N_13322,N_6356,N_12223);
nor U13323 (N_13323,N_12129,N_8985);
or U13324 (N_13324,N_8297,N_11962);
nand U13325 (N_13325,N_9025,N_11251);
and U13326 (N_13326,N_11627,N_11304);
nand U13327 (N_13327,N_8159,N_10665);
xor U13328 (N_13328,N_10985,N_11432);
xor U13329 (N_13329,N_11397,N_6641);
nor U13330 (N_13330,N_12213,N_11469);
and U13331 (N_13331,N_9813,N_7397);
nor U13332 (N_13332,N_7897,N_11734);
xor U13333 (N_13333,N_12156,N_6262);
xor U13334 (N_13334,N_7714,N_12344);
nor U13335 (N_13335,N_9908,N_10161);
nor U13336 (N_13336,N_10032,N_7815);
nor U13337 (N_13337,N_10532,N_7414);
nor U13338 (N_13338,N_11891,N_11269);
nor U13339 (N_13339,N_11400,N_6490);
nor U13340 (N_13340,N_11771,N_7430);
xor U13341 (N_13341,N_11848,N_7139);
nor U13342 (N_13342,N_9212,N_12157);
or U13343 (N_13343,N_6711,N_10080);
xnor U13344 (N_13344,N_9116,N_12320);
xnor U13345 (N_13345,N_9579,N_10427);
or U13346 (N_13346,N_7734,N_11894);
and U13347 (N_13347,N_10137,N_9451);
and U13348 (N_13348,N_9786,N_9690);
and U13349 (N_13349,N_10710,N_8337);
nor U13350 (N_13350,N_6669,N_8765);
or U13351 (N_13351,N_11491,N_6796);
or U13352 (N_13352,N_11890,N_8591);
nand U13353 (N_13353,N_6914,N_8711);
xor U13354 (N_13354,N_10347,N_9105);
nand U13355 (N_13355,N_12073,N_10476);
xor U13356 (N_13356,N_10417,N_12114);
and U13357 (N_13357,N_11423,N_6391);
nand U13358 (N_13358,N_10328,N_9528);
nor U13359 (N_13359,N_8121,N_9901);
xnor U13360 (N_13360,N_12121,N_8831);
nor U13361 (N_13361,N_10383,N_10969);
nor U13362 (N_13362,N_9288,N_11548);
nand U13363 (N_13363,N_9848,N_7823);
xnor U13364 (N_13364,N_10446,N_6795);
xnor U13365 (N_13365,N_11208,N_12055);
xnor U13366 (N_13366,N_7198,N_11168);
and U13367 (N_13367,N_8539,N_8392);
or U13368 (N_13368,N_10791,N_10165);
nand U13369 (N_13369,N_9254,N_9013);
or U13370 (N_13370,N_6591,N_7182);
or U13371 (N_13371,N_8439,N_11715);
nand U13372 (N_13372,N_11773,N_9585);
and U13373 (N_13373,N_8729,N_8490);
nor U13374 (N_13374,N_7534,N_6474);
xnor U13375 (N_13375,N_11018,N_6680);
nor U13376 (N_13376,N_11444,N_9581);
and U13377 (N_13377,N_7838,N_11558);
xnor U13378 (N_13378,N_11215,N_12165);
or U13379 (N_13379,N_7531,N_10666);
nor U13380 (N_13380,N_9029,N_8657);
and U13381 (N_13381,N_8303,N_8200);
xor U13382 (N_13382,N_6401,N_7108);
or U13383 (N_13383,N_8482,N_8234);
or U13384 (N_13384,N_8456,N_11000);
xnor U13385 (N_13385,N_8026,N_8466);
or U13386 (N_13386,N_9864,N_7569);
nor U13387 (N_13387,N_7261,N_9602);
nand U13388 (N_13388,N_7173,N_8697);
or U13389 (N_13389,N_10031,N_11111);
nand U13390 (N_13390,N_8365,N_10673);
nor U13391 (N_13391,N_11084,N_8277);
nand U13392 (N_13392,N_7047,N_9012);
nor U13393 (N_13393,N_8294,N_8418);
and U13394 (N_13394,N_8001,N_7163);
nor U13395 (N_13395,N_7341,N_9173);
and U13396 (N_13396,N_7197,N_11981);
and U13397 (N_13397,N_7037,N_8460);
and U13398 (N_13398,N_12321,N_6326);
xor U13399 (N_13399,N_12126,N_10468);
or U13400 (N_13400,N_9092,N_7109);
nor U13401 (N_13401,N_11172,N_10356);
nand U13402 (N_13402,N_8420,N_12023);
nor U13403 (N_13403,N_8869,N_7935);
nand U13404 (N_13404,N_10956,N_8572);
nand U13405 (N_13405,N_10239,N_7137);
or U13406 (N_13406,N_9195,N_7865);
or U13407 (N_13407,N_8404,N_6456);
or U13408 (N_13408,N_6283,N_7070);
xor U13409 (N_13409,N_7438,N_10290);
nor U13410 (N_13410,N_11709,N_11820);
xor U13411 (N_13411,N_11102,N_7779);
nor U13412 (N_13412,N_11447,N_7320);
xor U13413 (N_13413,N_6444,N_8124);
nand U13414 (N_13414,N_8222,N_9484);
or U13415 (N_13415,N_7983,N_11404);
or U13416 (N_13416,N_7537,N_11298);
or U13417 (N_13417,N_11680,N_6311);
nor U13418 (N_13418,N_7680,N_9825);
or U13419 (N_13419,N_7295,N_10181);
xnor U13420 (N_13420,N_10792,N_11318);
xnor U13421 (N_13421,N_6411,N_11919);
xor U13422 (N_13422,N_10402,N_11315);
nand U13423 (N_13423,N_10970,N_6583);
xnor U13424 (N_13424,N_9476,N_10442);
and U13425 (N_13425,N_11362,N_11210);
nor U13426 (N_13426,N_9749,N_8940);
or U13427 (N_13427,N_9126,N_11668);
xor U13428 (N_13428,N_9474,N_6433);
and U13429 (N_13429,N_9053,N_10454);
or U13430 (N_13430,N_11256,N_9997);
xnor U13431 (N_13431,N_11695,N_8308);
or U13432 (N_13432,N_11342,N_7831);
and U13433 (N_13433,N_9336,N_7063);
nor U13434 (N_13434,N_8028,N_8733);
nor U13435 (N_13435,N_11993,N_6850);
xnor U13436 (N_13436,N_10841,N_11519);
nor U13437 (N_13437,N_8638,N_11512);
or U13438 (N_13438,N_12217,N_6729);
or U13439 (N_13439,N_9523,N_11311);
or U13440 (N_13440,N_9046,N_7476);
and U13441 (N_13441,N_8233,N_10785);
nor U13442 (N_13442,N_11604,N_6833);
or U13443 (N_13443,N_9208,N_12203);
and U13444 (N_13444,N_10150,N_10663);
and U13445 (N_13445,N_12295,N_6562);
or U13446 (N_13446,N_10644,N_7940);
xnor U13447 (N_13447,N_12407,N_9249);
xnor U13448 (N_13448,N_10198,N_10507);
nor U13449 (N_13449,N_11657,N_8888);
xnor U13450 (N_13450,N_11564,N_11737);
nor U13451 (N_13451,N_8413,N_7036);
or U13452 (N_13452,N_9743,N_8381);
nor U13453 (N_13453,N_6523,N_6602);
and U13454 (N_13454,N_10469,N_11727);
or U13455 (N_13455,N_7112,N_6645);
nand U13456 (N_13456,N_9297,N_8330);
xnor U13457 (N_13457,N_9716,N_8267);
or U13458 (N_13458,N_9186,N_12265);
and U13459 (N_13459,N_6988,N_10349);
and U13460 (N_13460,N_9234,N_12364);
or U13461 (N_13461,N_7619,N_11280);
xnor U13462 (N_13462,N_10775,N_7805);
nand U13463 (N_13463,N_12318,N_12054);
nor U13464 (N_13464,N_11559,N_7237);
and U13465 (N_13465,N_9449,N_11056);
nand U13466 (N_13466,N_10267,N_7231);
or U13467 (N_13467,N_8960,N_8203);
nor U13468 (N_13468,N_11054,N_8703);
or U13469 (N_13469,N_8146,N_10187);
and U13470 (N_13470,N_9970,N_7979);
xnor U13471 (N_13471,N_8652,N_6775);
nor U13472 (N_13472,N_11641,N_6724);
or U13473 (N_13473,N_8941,N_6288);
nand U13474 (N_13474,N_8040,N_10731);
nor U13475 (N_13475,N_12303,N_6306);
xor U13476 (N_13476,N_10657,N_6683);
nand U13477 (N_13477,N_6561,N_11661);
nor U13478 (N_13478,N_10806,N_8307);
nor U13479 (N_13479,N_9986,N_11857);
or U13480 (N_13480,N_10404,N_9164);
nor U13481 (N_13481,N_7577,N_11309);
and U13482 (N_13482,N_10512,N_7319);
or U13483 (N_13483,N_12272,N_7827);
and U13484 (N_13484,N_8120,N_10182);
nand U13485 (N_13485,N_7495,N_8186);
nand U13486 (N_13486,N_8032,N_6331);
and U13487 (N_13487,N_9150,N_6920);
xor U13488 (N_13488,N_12338,N_12429);
nor U13489 (N_13489,N_7681,N_9435);
and U13490 (N_13490,N_6300,N_8855);
or U13491 (N_13491,N_12075,N_11497);
nand U13492 (N_13492,N_9388,N_9291);
nand U13493 (N_13493,N_10138,N_6619);
or U13494 (N_13494,N_8843,N_11498);
nor U13495 (N_13495,N_10569,N_12307);
xor U13496 (N_13496,N_7712,N_12116);
nand U13497 (N_13497,N_10240,N_6575);
nor U13498 (N_13498,N_11802,N_9911);
nand U13499 (N_13499,N_9769,N_10369);
and U13500 (N_13500,N_7810,N_10752);
xor U13501 (N_13501,N_11166,N_9251);
xnor U13502 (N_13502,N_7791,N_7642);
and U13503 (N_13503,N_7686,N_12347);
xor U13504 (N_13504,N_7003,N_9470);
and U13505 (N_13505,N_12243,N_10921);
or U13506 (N_13506,N_11785,N_9331);
nand U13507 (N_13507,N_10794,N_6527);
and U13508 (N_13508,N_8091,N_9381);
or U13509 (N_13509,N_7989,N_6413);
nand U13510 (N_13510,N_11294,N_10555);
nand U13511 (N_13511,N_7342,N_9431);
or U13512 (N_13512,N_6715,N_6944);
nand U13513 (N_13513,N_9448,N_10531);
xnor U13514 (N_13514,N_11812,N_10407);
or U13515 (N_13515,N_7308,N_11947);
nor U13516 (N_13516,N_6421,N_12325);
or U13517 (N_13517,N_12405,N_6656);
nand U13518 (N_13518,N_11131,N_12427);
nor U13519 (N_13519,N_7713,N_8206);
and U13520 (N_13520,N_7082,N_8259);
xnor U13521 (N_13521,N_7064,N_10110);
or U13522 (N_13522,N_8895,N_10675);
nor U13523 (N_13523,N_8090,N_8238);
nor U13524 (N_13524,N_7061,N_7545);
xor U13525 (N_13525,N_7454,N_7332);
nand U13526 (N_13526,N_11349,N_11411);
xor U13527 (N_13527,N_6574,N_12040);
xor U13528 (N_13528,N_6370,N_11223);
nand U13529 (N_13529,N_8924,N_9401);
xor U13530 (N_13530,N_8785,N_6815);
xnor U13531 (N_13531,N_10414,N_9733);
xor U13532 (N_13532,N_10448,N_6941);
nor U13533 (N_13533,N_6295,N_9094);
or U13534 (N_13534,N_12220,N_10986);
or U13535 (N_13535,N_9197,N_8289);
nor U13536 (N_13536,N_11966,N_10714);
nand U13537 (N_13537,N_7223,N_8402);
nor U13538 (N_13538,N_6762,N_10647);
and U13539 (N_13539,N_7640,N_7985);
xor U13540 (N_13540,N_8629,N_7666);
and U13541 (N_13541,N_7312,N_7541);
nand U13542 (N_13542,N_9731,N_10258);
or U13543 (N_13543,N_11822,N_12366);
or U13544 (N_13544,N_12270,N_10660);
xnor U13545 (N_13545,N_6629,N_9747);
and U13546 (N_13546,N_11487,N_8900);
nand U13547 (N_13547,N_6790,N_10622);
nor U13548 (N_13548,N_6309,N_7981);
nand U13549 (N_13549,N_8483,N_11704);
nand U13550 (N_13550,N_7093,N_10201);
nor U13551 (N_13551,N_11122,N_8085);
nand U13552 (N_13552,N_12052,N_6888);
and U13553 (N_13553,N_11761,N_6726);
nand U13554 (N_13554,N_6803,N_7971);
and U13555 (N_13555,N_8582,N_11886);
nor U13556 (N_13556,N_12425,N_7778);
nor U13557 (N_13557,N_7092,N_7322);
and U13558 (N_13558,N_6588,N_9704);
xor U13559 (N_13559,N_11484,N_9594);
nand U13560 (N_13560,N_8088,N_9294);
nor U13561 (N_13561,N_7229,N_9521);
and U13562 (N_13562,N_6835,N_10338);
xnor U13563 (N_13563,N_11155,N_12169);
nand U13564 (N_13564,N_10684,N_8734);
or U13565 (N_13565,N_6792,N_10275);
or U13566 (N_13566,N_10538,N_7784);
or U13567 (N_13567,N_10094,N_10246);
xor U13568 (N_13568,N_11179,N_11970);
nand U13569 (N_13569,N_6476,N_10535);
xnor U13570 (N_13570,N_7263,N_10053);
nor U13571 (N_13571,N_9906,N_6560);
xnor U13572 (N_13572,N_9866,N_11592);
nor U13573 (N_13573,N_10988,N_7248);
or U13574 (N_13574,N_6831,N_11723);
or U13575 (N_13575,N_9463,N_9894);
nor U13576 (N_13576,N_6532,N_9429);
and U13577 (N_13577,N_8903,N_8619);
or U13578 (N_13578,N_9808,N_10194);
nor U13579 (N_13579,N_7236,N_11772);
xor U13580 (N_13580,N_6965,N_10519);
nor U13581 (N_13581,N_11698,N_7630);
nor U13582 (N_13582,N_10859,N_9591);
nand U13583 (N_13583,N_7780,N_9204);
nand U13584 (N_13584,N_12443,N_12016);
nand U13585 (N_13585,N_12447,N_6652);
nand U13586 (N_13586,N_10509,N_11356);
xor U13587 (N_13587,N_11029,N_7704);
or U13588 (N_13588,N_12025,N_9442);
nand U13589 (N_13589,N_8847,N_11847);
nor U13590 (N_13590,N_12304,N_11274);
nand U13591 (N_13591,N_7415,N_8458);
or U13592 (N_13592,N_11438,N_7594);
or U13593 (N_13593,N_11353,N_8662);
xnor U13594 (N_13594,N_7012,N_10942);
and U13595 (N_13595,N_11524,N_10955);
nor U13596 (N_13596,N_9957,N_8314);
nand U13597 (N_13597,N_9421,N_8015);
or U13598 (N_13598,N_8768,N_10596);
xor U13599 (N_13599,N_7752,N_6553);
nand U13600 (N_13600,N_6594,N_9271);
xnor U13601 (N_13601,N_6446,N_9405);
nor U13602 (N_13602,N_9016,N_11455);
xor U13603 (N_13603,N_12092,N_12224);
nor U13604 (N_13604,N_10135,N_8859);
nor U13605 (N_13605,N_7055,N_12329);
or U13606 (N_13606,N_8000,N_11624);
nor U13607 (N_13607,N_7765,N_8877);
nor U13608 (N_13608,N_11245,N_9833);
nor U13609 (N_13609,N_9618,N_9170);
or U13610 (N_13610,N_9865,N_10436);
nor U13611 (N_13611,N_12050,N_11928);
nand U13612 (N_13612,N_8675,N_9802);
and U13613 (N_13613,N_12102,N_8753);
nand U13614 (N_13614,N_12077,N_6352);
and U13615 (N_13615,N_6565,N_9955);
xnor U13616 (N_13616,N_6521,N_11319);
and U13617 (N_13617,N_7934,N_7957);
nand U13618 (N_13618,N_7335,N_12410);
or U13619 (N_13619,N_6468,N_6399);
and U13620 (N_13620,N_7603,N_10860);
nand U13621 (N_13621,N_7035,N_11096);
and U13622 (N_13622,N_9207,N_8199);
nor U13623 (N_13623,N_7471,N_6744);
nand U13624 (N_13624,N_7809,N_10643);
and U13625 (N_13625,N_7437,N_6981);
nor U13626 (N_13626,N_8818,N_9391);
xnor U13627 (N_13627,N_8462,N_10669);
xor U13628 (N_13628,N_6314,N_8634);
xnor U13629 (N_13629,N_11869,N_10652);
nand U13630 (N_13630,N_6315,N_9074);
and U13631 (N_13631,N_7738,N_6417);
and U13632 (N_13632,N_8904,N_6927);
nand U13633 (N_13633,N_7662,N_10250);
nor U13634 (N_13634,N_7467,N_12476);
nand U13635 (N_13635,N_12453,N_7956);
or U13636 (N_13636,N_12021,N_11911);
nand U13637 (N_13637,N_7575,N_9616);
and U13638 (N_13638,N_9067,N_11776);
or U13639 (N_13639,N_11925,N_7028);
xnor U13640 (N_13640,N_6992,N_7644);
nor U13641 (N_13641,N_8528,N_8030);
or U13642 (N_13642,N_10449,N_10754);
nand U13643 (N_13643,N_9573,N_8833);
nor U13644 (N_13644,N_8201,N_10606);
xor U13645 (N_13645,N_8934,N_7268);
and U13646 (N_13646,N_9120,N_10936);
nor U13647 (N_13647,N_11643,N_10862);
and U13648 (N_13648,N_10050,N_7554);
or U13649 (N_13649,N_6568,N_10097);
nand U13650 (N_13650,N_10541,N_10795);
xor U13651 (N_13651,N_7361,N_8499);
or U13652 (N_13652,N_10202,N_7607);
nand U13653 (N_13653,N_11745,N_11011);
xor U13654 (N_13654,N_8920,N_9020);
xnor U13655 (N_13655,N_8390,N_6318);
xor U13656 (N_13656,N_10216,N_6671);
xor U13657 (N_13657,N_10058,N_8795);
or U13658 (N_13658,N_10722,N_11931);
nor U13659 (N_13659,N_7338,N_7381);
nor U13660 (N_13660,N_7001,N_10703);
nor U13661 (N_13661,N_8964,N_9142);
nand U13662 (N_13662,N_12194,N_10655);
nor U13663 (N_13663,N_6333,N_12315);
xor U13664 (N_13664,N_9350,N_8098);
nand U13665 (N_13665,N_9760,N_6512);
or U13666 (N_13666,N_10570,N_9661);
xor U13667 (N_13667,N_9650,N_12485);
nand U13668 (N_13668,N_8429,N_7887);
nor U13669 (N_13669,N_8132,N_7645);
xnor U13670 (N_13670,N_8440,N_7220);
and U13671 (N_13671,N_8209,N_6467);
xnor U13672 (N_13672,N_9507,N_12299);
nor U13673 (N_13673,N_11774,N_11164);
or U13674 (N_13674,N_11344,N_7443);
nand U13675 (N_13675,N_9108,N_6869);
or U13676 (N_13676,N_8322,N_7822);
or U13677 (N_13677,N_9130,N_10008);
and U13678 (N_13678,N_7872,N_11803);
or U13679 (N_13679,N_9697,N_11364);
nand U13680 (N_13680,N_6939,N_11046);
nand U13681 (N_13681,N_7411,N_8696);
nor U13682 (N_13682,N_6900,N_10131);
nor U13683 (N_13683,N_7777,N_6861);
and U13684 (N_13684,N_9339,N_7978);
xnor U13685 (N_13685,N_11068,N_7368);
or U13686 (N_13686,N_9631,N_8041);
nand U13687 (N_13687,N_11211,N_10450);
nand U13688 (N_13688,N_12041,N_12030);
and U13689 (N_13689,N_9506,N_9402);
or U13690 (N_13690,N_9218,N_10807);
nor U13691 (N_13691,N_12345,N_10604);
or U13692 (N_13692,N_9651,N_10812);
nand U13693 (N_13693,N_10747,N_12269);
or U13694 (N_13694,N_11810,N_10871);
xor U13695 (N_13695,N_6341,N_11845);
nor U13696 (N_13696,N_8754,N_7162);
nor U13697 (N_13697,N_10116,N_12155);
nor U13698 (N_13698,N_8601,N_7939);
or U13699 (N_13699,N_7976,N_6837);
xnor U13700 (N_13700,N_10927,N_6612);
and U13701 (N_13701,N_11465,N_11545);
xnor U13702 (N_13702,N_9076,N_10838);
nand U13703 (N_13703,N_8646,N_8389);
or U13704 (N_13704,N_7334,N_9805);
xor U13705 (N_13705,N_10437,N_11638);
or U13706 (N_13706,N_10286,N_7316);
or U13707 (N_13707,N_7475,N_9707);
xnor U13708 (N_13708,N_8984,N_7751);
or U13709 (N_13709,N_6587,N_10667);
nor U13710 (N_13710,N_7889,N_9583);
nand U13711 (N_13711,N_11938,N_6980);
and U13712 (N_13712,N_11613,N_10374);
or U13713 (N_13713,N_7459,N_10168);
and U13714 (N_13714,N_9689,N_7896);
xor U13715 (N_13715,N_8921,N_8856);
nand U13716 (N_13716,N_8363,N_10963);
or U13717 (N_13717,N_8606,N_8416);
or U13718 (N_13718,N_9375,N_10226);
nor U13719 (N_13719,N_9862,N_10272);
and U13720 (N_13720,N_6440,N_7824);
and U13721 (N_13721,N_8614,N_8565);
xor U13722 (N_13722,N_8530,N_11767);
nand U13723 (N_13723,N_12024,N_12174);
nor U13724 (N_13724,N_11213,N_7111);
nor U13725 (N_13725,N_7633,N_8262);
or U13726 (N_13726,N_8749,N_6743);
and U13727 (N_13727,N_7745,N_10489);
and U13728 (N_13728,N_9073,N_7493);
or U13729 (N_13729,N_11079,N_7481);
xor U13730 (N_13730,N_9837,N_9227);
and U13731 (N_13731,N_8668,N_7883);
nand U13732 (N_13732,N_10086,N_7949);
xnor U13733 (N_13733,N_11502,N_7634);
or U13734 (N_13734,N_8780,N_7661);
nand U13735 (N_13735,N_8514,N_7129);
and U13736 (N_13736,N_9776,N_6286);
and U13737 (N_13737,N_7801,N_9772);
and U13738 (N_13738,N_11964,N_10915);
nor U13739 (N_13739,N_11187,N_6668);
or U13740 (N_13740,N_9936,N_6639);
and U13741 (N_13741,N_9097,N_9968);
or U13742 (N_13742,N_8239,N_8450);
nand U13743 (N_13743,N_8154,N_9855);
nor U13744 (N_13744,N_7050,N_8502);
or U13745 (N_13745,N_9498,N_10366);
xnor U13746 (N_13746,N_10851,N_8627);
and U13747 (N_13747,N_7854,N_6437);
xor U13748 (N_13748,N_6373,N_12397);
nand U13749 (N_13749,N_9315,N_10472);
or U13750 (N_13750,N_11367,N_8679);
or U13751 (N_13751,N_11065,N_6463);
nand U13752 (N_13752,N_10737,N_9974);
nand U13753 (N_13753,N_8945,N_11010);
or U13754 (N_13754,N_6458,N_9829);
or U13755 (N_13755,N_6544,N_10262);
and U13756 (N_13756,N_12128,N_8326);
or U13757 (N_13757,N_9782,N_10149);
and U13758 (N_13758,N_6872,N_12191);
and U13759 (N_13759,N_8174,N_9037);
xor U13760 (N_13760,N_7188,N_10439);
nor U13761 (N_13761,N_8752,N_6931);
nor U13762 (N_13762,N_6438,N_12398);
xor U13763 (N_13763,N_8536,N_11977);
or U13764 (N_13764,N_11625,N_6752);
or U13765 (N_13765,N_6647,N_9871);
nand U13766 (N_13766,N_7015,N_7404);
nor U13767 (N_13767,N_7728,N_6296);
xor U13768 (N_13768,N_11777,N_11057);
nand U13769 (N_13769,N_8078,N_11180);
and U13770 (N_13770,N_8986,N_10488);
xnor U13771 (N_13771,N_7641,N_7128);
xor U13772 (N_13772,N_6670,N_10438);
nand U13773 (N_13773,N_11656,N_9953);
nor U13774 (N_13774,N_10883,N_8916);
nor U13775 (N_13775,N_11407,N_7725);
xor U13776 (N_13776,N_10971,N_10463);
xnor U13777 (N_13777,N_9351,N_10199);
nand U13778 (N_13778,N_6329,N_7729);
or U13779 (N_13779,N_11406,N_11533);
xor U13780 (N_13780,N_9270,N_10270);
and U13781 (N_13781,N_11462,N_9089);
or U13782 (N_13782,N_9263,N_10085);
or U13783 (N_13783,N_6304,N_7570);
and U13784 (N_13784,N_9511,N_7304);
nor U13785 (N_13785,N_9853,N_12037);
nand U13786 (N_13786,N_10726,N_11137);
and U13787 (N_13787,N_10378,N_12341);
xnor U13788 (N_13788,N_7966,N_7005);
or U13789 (N_13789,N_9543,N_11132);
or U13790 (N_13790,N_7274,N_8879);
and U13791 (N_13791,N_8231,N_11752);
nor U13792 (N_13792,N_6945,N_7507);
nand U13793 (N_13793,N_8061,N_10623);
and U13794 (N_13794,N_8255,N_6898);
or U13795 (N_13795,N_7702,N_12164);
or U13796 (N_13796,N_8593,N_8798);
or U13797 (N_13797,N_8383,N_11381);
and U13798 (N_13798,N_11660,N_10291);
or U13799 (N_13799,N_6550,N_11135);
and U13800 (N_13800,N_10946,N_10043);
and U13801 (N_13801,N_11884,N_9008);
nor U13802 (N_13802,N_9231,N_8992);
nor U13803 (N_13803,N_11288,N_9475);
nand U13804 (N_13804,N_10834,N_6936);
or U13805 (N_13805,N_9253,N_7318);
nor U13806 (N_13806,N_6378,N_8188);
or U13807 (N_13807,N_7510,N_11665);
nor U13808 (N_13808,N_11504,N_10733);
xnor U13809 (N_13809,N_10302,N_9551);
xor U13810 (N_13810,N_8716,N_7016);
xnor U13811 (N_13811,N_8446,N_8633);
nor U13812 (N_13812,N_9842,N_6791);
xnor U13813 (N_13813,N_6737,N_7657);
nand U13814 (N_13814,N_10739,N_10715);
and U13815 (N_13815,N_8857,N_7337);
xnor U13816 (N_13816,N_11965,N_8442);
and U13817 (N_13817,N_6821,N_6817);
nor U13818 (N_13818,N_9235,N_6889);
nand U13819 (N_13819,N_10206,N_7053);
and U13820 (N_13820,N_10470,N_9010);
nor U13821 (N_13821,N_8360,N_6673);
nand U13822 (N_13822,N_9715,N_7202);
nand U13823 (N_13823,N_9245,N_12043);
nor U13824 (N_13824,N_10044,N_6483);
xor U13825 (N_13825,N_9513,N_12414);
nor U13826 (N_13826,N_7371,N_12267);
nand U13827 (N_13827,N_8756,N_10316);
nor U13828 (N_13828,N_7771,N_9466);
nor U13829 (N_13829,N_10510,N_12143);
or U13830 (N_13830,N_7892,N_8452);
nor U13831 (N_13831,N_11042,N_10020);
or U13832 (N_13832,N_7301,N_6650);
or U13833 (N_13833,N_9021,N_11048);
xnor U13834 (N_13834,N_7622,N_6518);
nand U13835 (N_13835,N_10778,N_9033);
and U13836 (N_13836,N_8145,N_12100);
nor U13837 (N_13837,N_9246,N_12207);
and U13838 (N_13838,N_9115,N_11125);
nor U13839 (N_13839,N_11618,N_7996);
or U13840 (N_13840,N_9051,N_11331);
nor U13841 (N_13841,N_7997,N_8983);
or U13842 (N_13842,N_8886,N_12449);
and U13843 (N_13843,N_8799,N_9801);
xnor U13844 (N_13844,N_11971,N_8005);
nand U13845 (N_13845,N_11750,N_11183);
nand U13846 (N_13846,N_12402,N_9083);
nand U13847 (N_13847,N_9175,N_10746);
xor U13848 (N_13848,N_9123,N_6589);
xnor U13849 (N_13849,N_11654,N_9840);
or U13850 (N_13850,N_12355,N_8131);
nand U13851 (N_13851,N_8479,N_10061);
nor U13852 (N_13852,N_10077,N_7631);
and U13853 (N_13853,N_6267,N_7998);
nor U13854 (N_13854,N_11038,N_7081);
nor U13855 (N_13855,N_10247,N_9887);
and U13856 (N_13856,N_11320,N_9532);
nor U13857 (N_13857,N_10677,N_7119);
and U13858 (N_13858,N_6902,N_12361);
nor U13859 (N_13859,N_12080,N_9727);
nand U13860 (N_13860,N_8884,N_11778);
or U13861 (N_13861,N_9761,N_7426);
or U13862 (N_13862,N_9582,N_11601);
nand U13863 (N_13863,N_7258,N_12206);
nand U13864 (N_13864,N_6345,N_7069);
nor U13865 (N_13865,N_11980,N_12483);
nand U13866 (N_13866,N_6392,N_11333);
or U13867 (N_13867,N_9179,N_11481);
nand U13868 (N_13868,N_8905,N_6368);
and U13869 (N_13869,N_9885,N_6257);
and U13870 (N_13870,N_12063,N_7124);
or U13871 (N_13871,N_7189,N_12381);
nand U13872 (N_13872,N_6432,N_7615);
and U13873 (N_13873,N_9542,N_11602);
xnor U13874 (N_13874,N_7735,N_10308);
and U13875 (N_13875,N_8669,N_6693);
nand U13876 (N_13876,N_11594,N_10431);
nand U13877 (N_13877,N_9880,N_6789);
xor U13878 (N_13878,N_9555,N_11436);
nor U13879 (N_13879,N_7238,N_7817);
or U13880 (N_13880,N_12264,N_9444);
nor U13881 (N_13881,N_11912,N_10046);
or U13882 (N_13882,N_8212,N_9989);
xnor U13883 (N_13883,N_8070,N_11017);
nand U13884 (N_13884,N_12380,N_6859);
nand U13885 (N_13885,N_9196,N_9443);
nand U13886 (N_13886,N_6843,N_7408);
or U13887 (N_13887,N_10894,N_6273);
or U13888 (N_13888,N_7497,N_8970);
and U13889 (N_13889,N_6994,N_12393);
and U13890 (N_13890,N_7191,N_9360);
or U13891 (N_13891,N_8215,N_12305);
and U13892 (N_13892,N_11536,N_12091);
or U13893 (N_13893,N_6719,N_10924);
xnor U13894 (N_13894,N_8832,N_6935);
xor U13895 (N_13895,N_10269,N_11116);
nor U13896 (N_13896,N_7568,N_7344);
or U13897 (N_13897,N_9467,N_11972);
nor U13898 (N_13898,N_11301,N_8094);
or U13899 (N_13899,N_8128,N_7629);
nand U13900 (N_13900,N_9587,N_9228);
or U13901 (N_13901,N_9128,N_8762);
or U13902 (N_13902,N_9505,N_8073);
nand U13903 (N_13903,N_7484,N_8721);
xnor U13904 (N_13904,N_6770,N_6880);
or U13905 (N_13905,N_10284,N_10057);
and U13906 (N_13906,N_7775,N_12255);
xor U13907 (N_13907,N_8751,N_10038);
and U13908 (N_13908,N_8700,N_8953);
nor U13909 (N_13909,N_10940,N_9224);
nand U13910 (N_13910,N_12186,N_11167);
and U13911 (N_13911,N_6481,N_7501);
xor U13912 (N_13912,N_6332,N_7110);
nand U13913 (N_13913,N_8616,N_10263);
nand U13914 (N_13914,N_7951,N_8681);
or U13915 (N_13915,N_7362,N_8701);
nand U13916 (N_13916,N_10629,N_11865);
xor U13917 (N_13917,N_12188,N_8236);
nand U13918 (N_13918,N_12487,N_11076);
nor U13919 (N_13919,N_11142,N_11800);
nor U13920 (N_13920,N_11119,N_11402);
nor U13921 (N_13921,N_6581,N_10740);
and U13922 (N_13922,N_11843,N_7600);
xnor U13923 (N_13923,N_11748,N_12468);
xor U13924 (N_13924,N_9450,N_8053);
nand U13925 (N_13925,N_12391,N_10848);
and U13926 (N_13926,N_7048,N_8196);
nor U13927 (N_13927,N_9154,N_12428);
or U13928 (N_13928,N_12053,N_10950);
nand U13929 (N_13929,N_7995,N_8706);
or U13930 (N_13930,N_6741,N_9001);
nor U13931 (N_13931,N_11378,N_8529);
xnor U13932 (N_13932,N_10014,N_12353);
xor U13933 (N_13933,N_6495,N_11103);
or U13934 (N_13934,N_10766,N_9147);
or U13935 (N_13935,N_8569,N_9611);
xnor U13936 (N_13936,N_9072,N_8295);
or U13937 (N_13937,N_9879,N_10327);
or U13938 (N_13938,N_9612,N_11694);
nor U13939 (N_13939,N_12177,N_9548);
and U13940 (N_13940,N_7595,N_6365);
or U13941 (N_13941,N_7468,N_7522);
and U13942 (N_13942,N_7673,N_9726);
nor U13943 (N_13943,N_11178,N_11413);
nor U13944 (N_13944,N_9639,N_9796);
or U13945 (N_13945,N_7668,N_8902);
and U13946 (N_13946,N_8836,N_11219);
nor U13947 (N_13947,N_7696,N_12271);
and U13948 (N_13948,N_7291,N_7874);
xnor U13949 (N_13949,N_11801,N_9751);
xnor U13950 (N_13950,N_9504,N_11372);
xor U13951 (N_13951,N_10653,N_10709);
nand U13952 (N_13952,N_6343,N_9544);
nand U13953 (N_13953,N_9413,N_8782);
and U13954 (N_13954,N_8827,N_9942);
xor U13955 (N_13955,N_8939,N_7589);
or U13956 (N_13956,N_8620,N_11421);
nand U13957 (N_13957,N_7651,N_11511);
xor U13958 (N_13958,N_8518,N_9610);
or U13959 (N_13959,N_7682,N_6721);
xnor U13960 (N_13960,N_10881,N_12463);
nand U13961 (N_13961,N_6846,N_6596);
or U13962 (N_13962,N_11326,N_8315);
nand U13963 (N_13963,N_11729,N_10162);
or U13964 (N_13964,N_9575,N_9606);
nor U13965 (N_13965,N_10232,N_7252);
nand U13966 (N_13966,N_12352,N_7918);
nand U13967 (N_13967,N_10101,N_12228);
or U13968 (N_13968,N_12357,N_7698);
xor U13969 (N_13969,N_7830,N_9566);
or U13970 (N_13970,N_7626,N_8374);
xnor U13971 (N_13971,N_10579,N_7899);
nor U13972 (N_13972,N_8216,N_9695);
xnor U13973 (N_13973,N_11300,N_10741);
or U13974 (N_13974,N_9320,N_9788);
nor U13975 (N_13975,N_10642,N_12013);
nand U13976 (N_13976,N_10808,N_11087);
nand U13977 (N_13977,N_11002,N_10878);
xor U13978 (N_13978,N_7298,N_11261);
nor U13979 (N_13979,N_9415,N_7490);
or U13980 (N_13980,N_6450,N_9121);
nand U13981 (N_13981,N_7293,N_8391);
nand U13982 (N_13982,N_10615,N_10393);
nand U13983 (N_13983,N_11577,N_7325);
and U13984 (N_13984,N_8346,N_9084);
xnor U13985 (N_13985,N_11839,N_11066);
or U13986 (N_13986,N_8786,N_6637);
nor U13987 (N_13987,N_8348,N_12279);
xor U13988 (N_13988,N_9859,N_11237);
nand U13989 (N_13989,N_11984,N_6764);
nand U13990 (N_13990,N_10143,N_7637);
nand U13991 (N_13991,N_7024,N_7251);
nor U13992 (N_13992,N_8927,N_6298);
or U13993 (N_13993,N_12289,N_11472);
or U13994 (N_13994,N_11217,N_8214);
nor U13995 (N_13995,N_10397,N_9118);
and U13996 (N_13996,N_11786,N_11415);
nand U13997 (N_13997,N_12103,N_8373);
or U13998 (N_13998,N_6706,N_9151);
xor U13999 (N_13999,N_10490,N_10426);
nand U14000 (N_14000,N_9807,N_12058);
nor U14001 (N_14001,N_10685,N_8545);
or U14002 (N_14002,N_6829,N_10771);
xnor U14003 (N_14003,N_6772,N_10964);
nand U14004 (N_14004,N_12498,N_9347);
or U14005 (N_14005,N_8533,N_8641);
or U14006 (N_14006,N_12248,N_12362);
nor U14007 (N_14007,N_11369,N_7948);
nand U14008 (N_14008,N_6702,N_8148);
or U14009 (N_14009,N_8660,N_7959);
and U14010 (N_14010,N_10738,N_10453);
xnor U14011 (N_14011,N_8705,N_10496);
xor U14012 (N_14012,N_12198,N_7222);
nor U14013 (N_14013,N_10835,N_8166);
and U14014 (N_14014,N_6877,N_7583);
nor U14015 (N_14015,N_9190,N_10707);
and U14016 (N_14016,N_10234,N_9799);
nor U14017 (N_14017,N_9437,N_11999);
or U14018 (N_14018,N_11989,N_9460);
nor U14019 (N_14019,N_7715,N_10736);
xor U14020 (N_14020,N_6779,N_12440);
or U14021 (N_14021,N_11837,N_6783);
nor U14022 (N_14022,N_11448,N_6982);
nor U14023 (N_14023,N_8774,N_12283);
nand U14024 (N_14024,N_8592,N_8137);
nor U14025 (N_14025,N_7485,N_6471);
and U14026 (N_14026,N_9501,N_8187);
nor U14027 (N_14027,N_10461,N_12094);
and U14028 (N_14028,N_11022,N_7796);
or U14029 (N_14029,N_11557,N_7833);
nor U14030 (N_14030,N_7333,N_7578);
nor U14031 (N_14031,N_11614,N_8747);
xor U14032 (N_14032,N_7974,N_12445);
nor U14033 (N_14033,N_10645,N_7786);
or U14034 (N_14034,N_8946,N_8957);
nor U14035 (N_14035,N_9127,N_11089);
or U14036 (N_14036,N_12020,N_8858);
nor U14037 (N_14037,N_6716,N_10481);
nor U14038 (N_14038,N_8312,N_7592);
nor U14039 (N_14039,N_6954,N_9489);
or U14040 (N_14040,N_7234,N_8181);
and U14041 (N_14041,N_9327,N_8971);
nor U14042 (N_14042,N_6367,N_8948);
or U14043 (N_14043,N_8486,N_7147);
nor U14044 (N_14044,N_8008,N_7164);
nand U14045 (N_14045,N_6535,N_7393);
nor U14046 (N_14046,N_8901,N_8003);
nand U14047 (N_14047,N_6813,N_8587);
nor U14048 (N_14048,N_6801,N_8791);
nand U14049 (N_14049,N_9622,N_12257);
nor U14050 (N_14050,N_10635,N_10769);
nand U14051 (N_14051,N_9390,N_10917);
or U14052 (N_14052,N_7847,N_11528);
nand U14053 (N_14053,N_10452,N_9162);
and U14054 (N_14054,N_6418,N_11859);
xnor U14055 (N_14055,N_12424,N_11192);
and U14056 (N_14056,N_12039,N_9503);
nand U14057 (N_14057,N_10091,N_10241);
nand U14058 (N_14058,N_8399,N_7559);
and U14059 (N_14059,N_9723,N_8178);
and U14060 (N_14060,N_6611,N_6800);
or U14061 (N_14061,N_12437,N_7623);
nor U14062 (N_14062,N_8376,N_10729);
or U14063 (N_14063,N_7157,N_7546);
nor U14064 (N_14064,N_9605,N_12334);
or U14065 (N_14065,N_8702,N_9184);
and U14066 (N_14066,N_11336,N_10382);
nand U14067 (N_14067,N_11818,N_6572);
and U14068 (N_14068,N_6361,N_6462);
or U14069 (N_14069,N_7135,N_9420);
and U14070 (N_14070,N_11182,N_8275);
xnor U14071 (N_14071,N_7811,N_11986);
nor U14072 (N_14072,N_9199,N_7359);
nand U14073 (N_14073,N_7027,N_12125);
or U14074 (N_14074,N_10762,N_6313);
nand U14075 (N_14075,N_10228,N_7879);
nor U14076 (N_14076,N_9969,N_7219);
nand U14077 (N_14077,N_11013,N_9386);
and U14078 (N_14078,N_9032,N_10931);
and U14079 (N_14079,N_9785,N_9789);
and U14080 (N_14080,N_11190,N_6279);
nand U14081 (N_14081,N_8658,N_6414);
nor U14082 (N_14082,N_8644,N_7410);
xor U14083 (N_14083,N_11325,N_8865);
and U14084 (N_14084,N_8725,N_11678);
nor U14085 (N_14085,N_11949,N_12088);
and U14086 (N_14086,N_7477,N_6759);
nor U14087 (N_14087,N_8272,N_8384);
or U14088 (N_14088,N_9048,N_12459);
and U14089 (N_14089,N_9396,N_11276);
and U14090 (N_14090,N_7246,N_12010);
nand U14091 (N_14091,N_7758,N_11834);
nand U14092 (N_14092,N_6966,N_7671);
and U14093 (N_14093,N_9925,N_8095);
nor U14094 (N_14094,N_6632,N_10134);
nand U14095 (N_14095,N_9385,N_11445);
and U14096 (N_14096,N_6351,N_10662);
xnor U14097 (N_14097,N_9049,N_10517);
or U14098 (N_14098,N_10529,N_9300);
nor U14099 (N_14099,N_6686,N_10600);
and U14100 (N_14100,N_11241,N_7557);
nor U14101 (N_14101,N_11889,N_10412);
xor U14102 (N_14102,N_10788,N_7498);
and U14103 (N_14103,N_10790,N_10520);
and U14104 (N_14104,N_6709,N_7384);
and U14105 (N_14105,N_9624,N_9273);
nor U14106 (N_14106,N_12454,N_6569);
nand U14107 (N_14107,N_9461,N_6890);
nor U14108 (N_14108,N_9156,N_6376);
xor U14109 (N_14109,N_7207,N_8400);
and U14110 (N_14110,N_11805,N_9215);
and U14111 (N_14111,N_10968,N_11844);
and U14112 (N_14112,N_9980,N_7205);
and U14113 (N_14113,N_11563,N_8127);
and U14114 (N_14114,N_7685,N_7862);
nor U14115 (N_14115,N_10475,N_6436);
nand U14116 (N_14116,N_8067,N_9642);
nand U14117 (N_14117,N_9034,N_10858);
or U14118 (N_14118,N_12201,N_10536);
xor U14119 (N_14119,N_6385,N_11878);
nor U14120 (N_14120,N_10096,N_11793);
xor U14121 (N_14121,N_7029,N_10683);
xnor U14122 (N_14122,N_7331,N_12351);
nand U14123 (N_14123,N_10957,N_9646);
nor U14124 (N_14124,N_11852,N_10591);
and U14125 (N_14125,N_8717,N_10176);
and U14126 (N_14126,N_10877,N_11892);
nor U14127 (N_14127,N_9508,N_9346);
and U14128 (N_14128,N_8741,N_6618);
nor U14129 (N_14129,N_6578,N_9369);
and U14130 (N_14130,N_11129,N_9878);
nor U14131 (N_14131,N_9167,N_11687);
xnor U14132 (N_14132,N_10183,N_9259);
nor U14133 (N_14133,N_7370,N_7044);
xor U14134 (N_14134,N_6677,N_9614);
nand U14135 (N_14135,N_9066,N_12339);
and U14136 (N_14136,N_10092,N_8519);
nor U14137 (N_14137,N_9493,N_10166);
xor U14138 (N_14138,N_10148,N_8292);
xnor U14139 (N_14139,N_6657,N_8968);
nor U14140 (N_14140,N_7366,N_11758);
and U14141 (N_14141,N_11003,N_10388);
and U14142 (N_14142,N_10523,N_8488);
nand U14143 (N_14143,N_10376,N_7409);
xnor U14144 (N_14144,N_9800,N_9111);
and U14145 (N_14145,N_11815,N_6321);
nor U14146 (N_14146,N_8080,N_11960);
nor U14147 (N_14147,N_6839,N_11476);
and U14148 (N_14148,N_6853,N_8603);
nor U14149 (N_14149,N_10990,N_11218);
or U14150 (N_14150,N_7591,N_9635);
nor U14151 (N_14151,N_12467,N_12276);
xor U14152 (N_14152,N_11953,N_9163);
and U14153 (N_14153,N_6290,N_9758);
nor U14154 (N_14154,N_11265,N_11278);
and U14155 (N_14155,N_10553,N_12373);
xnor U14156 (N_14156,N_6282,N_8890);
xor U14157 (N_14157,N_9260,N_9615);
nand U14158 (N_14158,N_11198,N_9882);
nand U14159 (N_14159,N_6580,N_6685);
nand U14160 (N_14160,N_8107,N_8447);
or U14161 (N_14161,N_8653,N_9721);
or U14162 (N_14162,N_10440,N_7588);
nand U14163 (N_14163,N_9318,N_6819);
nor U14164 (N_14164,N_12231,N_10912);
nor U14165 (N_14165,N_10572,N_12168);
and U14166 (N_14166,N_10159,N_10885);
nor U14167 (N_14167,N_10104,N_11724);
and U14168 (N_14168,N_9604,N_8866);
and U14169 (N_14169,N_7474,N_12495);
or U14170 (N_14170,N_9428,N_12400);
nand U14171 (N_14171,N_10303,N_6651);
or U14172 (N_14172,N_6718,N_12081);
and U14173 (N_14173,N_8506,N_8779);
xor U14174 (N_14174,N_7834,N_11942);
and U14175 (N_14175,N_7509,N_10659);
and U14176 (N_14176,N_8850,N_11580);
nand U14177 (N_14177,N_6698,N_10237);
nor U14178 (N_14178,N_10056,N_10214);
or U14179 (N_14179,N_7803,N_9317);
nand U14180 (N_14180,N_11033,N_11004);
nor U14181 (N_14181,N_8410,N_8993);
and U14182 (N_14182,N_11676,N_10287);
and U14183 (N_14183,N_11531,N_6514);
nor U14184 (N_14184,N_8281,N_12280);
nor U14185 (N_14185,N_12323,N_11153);
nor U14186 (N_14186,N_8661,N_8876);
nor U14187 (N_14187,N_12420,N_9187);
nand U14188 (N_14188,N_11321,N_12250);
nand U14189 (N_14189,N_8165,N_7159);
xor U14190 (N_14190,N_6664,N_11520);
nand U14191 (N_14191,N_11832,N_11615);
or U14192 (N_14192,N_8736,N_6364);
and U14193 (N_14193,N_9232,N_6788);
or U14194 (N_14194,N_11983,N_8151);
or U14195 (N_14195,N_9910,N_7655);
nand U14196 (N_14196,N_7695,N_10433);
nor U14197 (N_14197,N_6497,N_6388);
nor U14198 (N_14198,N_9954,N_8987);
and U14199 (N_14199,N_12171,N_6912);
xnor U14200 (N_14200,N_9502,N_8288);
nor U14201 (N_14201,N_7002,N_8258);
nor U14202 (N_14202,N_11691,N_11823);
nor U14203 (N_14203,N_10337,N_6557);
xnor U14204 (N_14204,N_8552,N_12117);
or U14205 (N_14205,N_6597,N_8630);
or U14206 (N_14206,N_8554,N_6363);
nand U14207 (N_14207,N_11224,N_7825);
nor U14208 (N_14208,N_10309,N_6897);
or U14209 (N_14209,N_7482,N_9890);
nand U14210 (N_14210,N_11939,N_11535);
xor U14211 (N_14211,N_11446,N_9941);
nand U14212 (N_14212,N_7169,N_7855);
or U14213 (N_14213,N_7289,N_9857);
nor U14214 (N_14214,N_6847,N_11014);
xor U14215 (N_14215,N_9079,N_8811);
xnor U14216 (N_14216,N_11623,N_6780);
and U14217 (N_14217,N_11121,N_7923);
nor U14218 (N_14218,N_9982,N_7011);
nor U14219 (N_14219,N_11644,N_11764);
nand U14220 (N_14220,N_9305,N_8058);
nand U14221 (N_14221,N_6270,N_9006);
and U14222 (N_14222,N_10556,N_6362);
xnor U14223 (N_14223,N_10527,N_12465);
nand U14224 (N_14224,N_10501,N_7267);
or U14225 (N_14225,N_9081,N_6620);
nor U14226 (N_14226,N_8291,N_7878);
or U14227 (N_14227,N_10502,N_10180);
nand U14228 (N_14228,N_9663,N_11940);
nor U14229 (N_14229,N_8543,N_9636);
xor U14230 (N_14230,N_9988,N_12253);
xnor U14231 (N_14231,N_7908,N_8248);
xor U14232 (N_14232,N_9806,N_7762);
nor U14233 (N_14233,N_8006,N_11679);
xor U14234 (N_14234,N_8394,N_10698);
xor U14235 (N_14235,N_9976,N_11050);
and U14236 (N_14236,N_11233,N_10844);
or U14237 (N_14237,N_7098,N_8929);
xnor U14238 (N_14238,N_10781,N_6319);
nor U14239 (N_14239,N_8296,N_11518);
or U14240 (N_14240,N_10067,N_7180);
xor U14241 (N_14241,N_9828,N_8860);
nand U14242 (N_14242,N_9418,N_11195);
nor U14243 (N_14243,N_11220,N_6600);
nor U14244 (N_14244,N_11232,N_9706);
or U14245 (N_14245,N_12337,N_8748);
or U14246 (N_14246,N_7808,N_9559);
nor U14247 (N_14247,N_7689,N_7085);
nand U14248 (N_14248,N_7428,N_8451);
nor U14249 (N_14249,N_11705,N_11059);
nor U14250 (N_14250,N_7590,N_9176);
or U14251 (N_14251,N_7099,N_9490);
nand U14252 (N_14252,N_6745,N_10932);
nor U14253 (N_14253,N_7278,N_10530);
nor U14254 (N_14254,N_9960,N_11766);
xor U14255 (N_14255,N_7511,N_9169);
xor U14256 (N_14256,N_7877,N_10682);
and U14257 (N_14257,N_9483,N_8923);
and U14258 (N_14258,N_6548,N_7621);
nand U14259 (N_14259,N_9939,N_8823);
or U14260 (N_14260,N_8327,N_6678);
xor U14261 (N_14261,N_10298,N_8532);
and U14262 (N_14262,N_6989,N_7794);
nor U14263 (N_14263,N_8464,N_12461);
and U14264 (N_14264,N_8803,N_7703);
or U14265 (N_14265,N_11606,N_12446);
and U14266 (N_14266,N_10873,N_9472);
xor U14267 (N_14267,N_8144,N_11253);
and U14268 (N_14268,N_7610,N_10464);
or U14269 (N_14269,N_12319,N_11414);
nor U14270 (N_14270,N_9720,N_11642);
and U14271 (N_14271,N_10065,N_6496);
nand U14272 (N_14272,N_8504,N_10420);
nor U14273 (N_14273,N_7211,N_10974);
xnor U14274 (N_14274,N_9404,N_9546);
nor U14275 (N_14275,N_7321,N_11685);
or U14276 (N_14276,N_8981,N_7524);
xnor U14277 (N_14277,N_8263,N_9497);
and U14278 (N_14278,N_6584,N_12481);
and U14279 (N_14279,N_6254,N_8583);
nand U14280 (N_14280,N_11650,N_8763);
nand U14281 (N_14281,N_6404,N_8191);
or U14282 (N_14282,N_9052,N_12078);
xnor U14283 (N_14283,N_11118,N_10037);
and U14284 (N_14284,N_10926,N_8874);
nor U14285 (N_14285,N_10371,N_7094);
and U14286 (N_14286,N_11061,N_6866);
xor U14287 (N_14287,N_7377,N_10479);
xnor U14288 (N_14288,N_7727,N_12452);
xnor U14289 (N_14289,N_12421,N_11917);
nand U14290 (N_14290,N_7170,N_10278);
and U14291 (N_14291,N_6684,N_10977);
or U14292 (N_14292,N_11539,N_9742);
nand U14293 (N_14293,N_9359,N_11067);
and U14294 (N_14294,N_10079,N_7871);
and U14295 (N_14295,N_8408,N_11662);
and U14296 (N_14296,N_6519,N_11930);
nor U14297 (N_14297,N_9783,N_11755);
nor U14298 (N_14298,N_8800,N_10112);
or U14299 (N_14299,N_9468,N_9436);
nor U14300 (N_14300,N_6494,N_6448);
nor U14301 (N_14301,N_8841,N_8677);
and U14302 (N_14302,N_11295,N_7271);
nor U14303 (N_14303,N_11156,N_6430);
nand U14304 (N_14304,N_11425,N_10132);
xor U14305 (N_14305,N_6863,N_7257);
and U14306 (N_14306,N_12178,N_9491);
and U14307 (N_14307,N_8155,N_8401);
xnor U14308 (N_14308,N_7915,N_9990);
nor U14309 (N_14309,N_6738,N_9637);
nor U14310 (N_14310,N_11619,N_7687);
nor U14311 (N_14311,N_8299,N_11730);
and U14312 (N_14312,N_9995,N_10471);
xnor U14313 (N_14313,N_12196,N_11870);
or U14314 (N_14314,N_8534,N_7856);
or U14315 (N_14315,N_6415,N_7814);
or U14316 (N_14316,N_7444,N_7071);
nand U14317 (N_14317,N_7017,N_9570);
and U14318 (N_14318,N_6653,N_10546);
or U14319 (N_14319,N_12448,N_8498);
nand U14320 (N_14320,N_8033,N_8197);
nor U14321 (N_14321,N_6475,N_8965);
and U14322 (N_14322,N_12163,N_6322);
nand U14323 (N_14323,N_12132,N_9793);
and U14324 (N_14324,N_12324,N_12281);
nand U14325 (N_14325,N_6525,N_8089);
or U14326 (N_14326,N_11696,N_10759);
xnor U14327 (N_14327,N_8431,N_6598);
or U14328 (N_14328,N_8520,N_10221);
and U14329 (N_14329,N_9895,N_10574);
xor U14330 (N_14330,N_10534,N_6635);
and U14331 (N_14331,N_11107,N_10514);
or U14332 (N_14332,N_12082,N_7530);
or U14333 (N_14333,N_9323,N_7382);
or U14334 (N_14334,N_8142,N_6710);
nor U14335 (N_14335,N_7697,N_12135);
or U14336 (N_14336,N_11250,N_8806);
or U14337 (N_14337,N_10059,N_11201);
or U14338 (N_14338,N_12474,N_8761);
nand U14339 (N_14339,N_11570,N_6586);
xor U14340 (N_14340,N_8372,N_8906);
and U14341 (N_14341,N_11824,N_6536);
nor U14342 (N_14342,N_7462,N_9827);
nand U14343 (N_14343,N_8801,N_10024);
or U14344 (N_14344,N_9031,N_7245);
and U14345 (N_14345,N_12134,N_9070);
nand U14346 (N_14346,N_9433,N_8489);
and U14347 (N_14347,N_12374,N_11584);
xnor U14348 (N_14348,N_8184,N_11838);
xor U14349 (N_14349,N_8507,N_12166);
nor U14350 (N_14350,N_6554,N_9334);
nor U14351 (N_14351,N_10105,N_7132);
or U14352 (N_14352,N_8854,N_11581);
or U14353 (N_14353,N_7502,N_8574);
nand U14354 (N_14354,N_12099,N_8707);
xor U14355 (N_14355,N_12245,N_9701);
xor U14356 (N_14356,N_11814,N_6466);
or U14357 (N_14357,N_12062,N_6676);
xnor U14358 (N_14358,N_6765,N_11385);
and U14359 (N_14359,N_6347,N_9826);
xor U14360 (N_14360,N_6730,N_8051);
nand U14361 (N_14361,N_11064,N_8825);
nand U14362 (N_14362,N_10693,N_7465);
xnor U14363 (N_14363,N_8093,N_8538);
and U14364 (N_14364,N_6701,N_12029);
or U14365 (N_14365,N_8417,N_6511);
and U14366 (N_14366,N_9057,N_6838);
nor U14367 (N_14367,N_10700,N_12434);
and U14368 (N_14368,N_10353,N_7442);
xor U14369 (N_14369,N_11568,N_10189);
xnor U14370 (N_14370,N_10345,N_6875);
nor U14371 (N_14371,N_6672,N_6646);
nor U14372 (N_14372,N_9027,N_9026);
and U14373 (N_14373,N_6867,N_11209);
nand U14374 (N_14374,N_9711,N_9242);
and U14375 (N_14375,N_9102,N_12308);
nand U14376 (N_14376,N_6592,N_10687);
or U14377 (N_14377,N_9447,N_8475);
nor U14378 (N_14378,N_8444,N_8194);
nand U14379 (N_14379,N_6751,N_12187);
and U14380 (N_14380,N_9676,N_11023);
or U14381 (N_14381,N_12083,N_6334);
xor U14382 (N_14382,N_8501,N_12382);
and U14383 (N_14383,N_8407,N_9932);
xor U14384 (N_14384,N_7130,N_12456);
nor U14385 (N_14385,N_10107,N_11388);
xor U14386 (N_14386,N_6268,N_7733);
nor U14387 (N_14387,N_10503,N_10152);
or U14388 (N_14388,N_10365,N_9430);
xnor U14389 (N_14389,N_6962,N_9926);
nand U14390 (N_14390,N_9481,N_10802);
and U14391 (N_14391,N_7286,N_7349);
and U14392 (N_14392,N_11763,N_11635);
xor U14393 (N_14393,N_12471,N_11510);
and U14394 (N_14394,N_9732,N_12074);
nor U14395 (N_14395,N_9407,N_8129);
or U14396 (N_14396,N_11477,N_11109);
and U14397 (N_14397,N_11873,N_6403);
nor U14398 (N_14398,N_6999,N_7282);
xnor U14399 (N_14399,N_12435,N_8268);
and U14400 (N_14400,N_6881,N_11725);
nor U14401 (N_14401,N_12173,N_9553);
or U14402 (N_14402,N_11184,N_8794);
or U14403 (N_14403,N_9979,N_12431);
nor U14404 (N_14404,N_9131,N_9846);
nor U14405 (N_14405,N_8357,N_12105);
nand U14406 (N_14406,N_7884,N_9180);
nor U14407 (N_14407,N_7150,N_9647);
nor U14408 (N_14408,N_7924,N_11647);
nor U14409 (N_14409,N_9355,N_10334);
xor U14410 (N_14410,N_11835,N_6666);
xnor U14411 (N_14411,N_6934,N_9816);
xor U14412 (N_14412,N_6545,N_9325);
xnor U14413 (N_14413,N_6734,N_8513);
or U14414 (N_14414,N_12036,N_11117);
or U14415 (N_14415,N_11277,N_10003);
xor U14416 (N_14416,N_10631,N_9923);
xor U14417 (N_14417,N_8230,N_10800);
nand U14418 (N_14418,N_10745,N_7960);
and U14419 (N_14419,N_8557,N_10911);
or U14420 (N_14420,N_12215,N_7171);
xnor U14421 (N_14421,N_8820,N_7385);
or U14422 (N_14422,N_10098,N_8048);
or U14423 (N_14423,N_9668,N_11954);
or U14424 (N_14424,N_8117,N_9096);
or U14425 (N_14425,N_10049,N_8891);
or U14426 (N_14426,N_10435,N_7806);
or U14427 (N_14427,N_9607,N_10965);
and U14428 (N_14428,N_9219,N_9144);
or U14429 (N_14429,N_11648,N_11508);
and U14430 (N_14430,N_6260,N_6277);
xnor U14431 (N_14431,N_8042,N_10991);
nand U14432 (N_14432,N_10627,N_9845);
or U14433 (N_14433,N_11101,N_8611);
nand U14434 (N_14434,N_9138,N_10319);
nor U14435 (N_14435,N_7255,N_10624);
nand U14436 (N_14436,N_11682,N_6826);
xor U14437 (N_14437,N_6760,N_9693);
nor U14438 (N_14438,N_9134,N_8692);
nand U14439 (N_14439,N_6768,N_6856);
nand U14440 (N_14440,N_6558,N_11866);
nor U14441 (N_14441,N_6447,N_7881);
or U14442 (N_14442,N_7230,N_11633);
nor U14443 (N_14443,N_10128,N_8320);
xnor U14444 (N_14444,N_12009,N_10130);
xnor U14445 (N_14445,N_11861,N_8911);
or U14446 (N_14446,N_7683,N_7711);
and U14447 (N_14447,N_10342,N_11238);
nand U14448 (N_14448,N_9741,N_11659);
or U14449 (N_14449,N_10939,N_8698);
xnor U14450 (N_14450,N_11943,N_8141);
xnor U14451 (N_14451,N_9124,N_10857);
nand U14452 (N_14452,N_6860,N_6665);
nor U14453 (N_14453,N_6692,N_9818);
xor U14454 (N_14454,N_9722,N_8018);
or U14455 (N_14455,N_11747,N_10723);
and U14456 (N_14456,N_7209,N_11683);
nor U14457 (N_14457,N_9303,N_11451);
nor U14458 (N_14458,N_7066,N_12145);
nand U14459 (N_14459,N_7606,N_6603);
or U14460 (N_14460,N_6756,N_9153);
xor U14461 (N_14461,N_8306,N_7101);
or U14462 (N_14462,N_6423,N_12087);
and U14463 (N_14463,N_7789,N_8576);
nor U14464 (N_14464,N_6886,N_11515);
and U14465 (N_14465,N_12499,N_9987);
nor U14466 (N_14466,N_7601,N_12296);
xnor U14467 (N_14467,N_10063,N_8715);
nor U14468 (N_14468,N_7938,N_6909);
nor U14469 (N_14469,N_8604,N_6280);
nor U14470 (N_14470,N_12466,N_8025);
nor U14471 (N_14471,N_6524,N_7242);
nand U14472 (N_14472,N_10001,N_10074);
nor U14473 (N_14473,N_10259,N_7140);
nand U14474 (N_14474,N_6940,N_6377);
nand U14475 (N_14475,N_9729,N_11836);
xor U14476 (N_14476,N_10387,N_10494);
nand U14477 (N_14477,N_8054,N_9896);
nor U14478 (N_14478,N_9977,N_11200);
nand U14479 (N_14479,N_7041,N_7538);
nand U14480 (N_14480,N_11742,N_8989);
xor U14481 (N_14481,N_10185,N_11409);
and U14482 (N_14482,N_6793,N_6310);
nor U14483 (N_14483,N_11357,N_10982);
nand U14484 (N_14484,N_10332,N_10310);
and U14485 (N_14485,N_6879,N_11384);
or U14486 (N_14486,N_8329,N_7464);
nand U14487 (N_14487,N_8835,N_11922);
nand U14488 (N_14488,N_12457,N_11148);
xnor U14489 (N_14489,N_9063,N_10293);
nor U14490 (N_14490,N_7580,N_6952);
and U14491 (N_14491,N_7688,N_8772);
xnor U14492 (N_14492,N_9943,N_12086);
nor U14493 (N_14493,N_11858,N_9734);
and U14494 (N_14494,N_8883,N_6633);
and U14495 (N_14495,N_10245,N_11442);
nand U14496 (N_14496,N_7276,N_8436);
nand U14497 (N_14497,N_9613,N_11671);
nor U14498 (N_14498,N_10562,N_9299);
nand U14499 (N_14499,N_9904,N_10352);
nor U14500 (N_14500,N_8730,N_6918);
or U14501 (N_14501,N_8568,N_10006);
nor U14502 (N_14502,N_10601,N_9376);
and U14503 (N_14503,N_8414,N_12193);
or U14504 (N_14504,N_11377,N_6350);
and U14505 (N_14505,N_8838,N_8139);
xnor U14506 (N_14506,N_11351,N_6767);
xnor U14507 (N_14507,N_8994,N_6478);
xnor U14508 (N_14508,N_7731,N_8453);
and U14509 (N_14509,N_7431,N_11449);
xor U14510 (N_14510,N_11621,N_12033);
or U14511 (N_14511,N_9298,N_10909);
xnor U14512 (N_14512,N_9571,N_12162);
and U14513 (N_14513,N_10034,N_6380);
and U14514 (N_14514,N_7265,N_9210);
or U14515 (N_14515,N_6799,N_8693);
and U14516 (N_14516,N_8709,N_7088);
nor U14517 (N_14517,N_12479,N_8044);
or U14518 (N_14518,N_7652,N_6278);
nand U14519 (N_14519,N_6797,N_8571);
or U14520 (N_14520,N_7928,N_10951);
xor U14521 (N_14521,N_10825,N_6434);
and U14522 (N_14522,N_9149,N_10500);
xnor U14523 (N_14523,N_10573,N_10849);
nand U14524 (N_14524,N_9047,N_10233);
xnor U14525 (N_14525,N_6493,N_7905);
xor U14526 (N_14526,N_7149,N_8828);
and U14527 (N_14527,N_8035,N_10473);
nand U14528 (N_14528,N_11516,N_10613);
and U14529 (N_14529,N_9705,N_12142);
and U14530 (N_14530,N_7861,N_12450);
nor U14531 (N_14531,N_6552,N_9645);
xnor U14532 (N_14532,N_7077,N_9709);
xnor U14533 (N_14533,N_10445,N_9752);
xor U14534 (N_14534,N_11813,N_10418);
and U14535 (N_14535,N_8581,N_8210);
xnor U14536 (N_14536,N_12051,N_8361);
or U14537 (N_14537,N_8776,N_11030);
nor U14538 (N_14538,N_8631,N_8433);
nor U14539 (N_14539,N_6699,N_7279);
xnor U14540 (N_14540,N_10948,N_10616);
nand U14541 (N_14541,N_8500,N_9763);
nand U14542 (N_14542,N_8147,N_9669);
xor U14543 (N_14543,N_10753,N_8049);
nor U14544 (N_14544,N_9540,N_10686);
xnor U14545 (N_14545,N_10218,N_6406);
and U14546 (N_14546,N_10605,N_11566);
nand U14547 (N_14547,N_6472,N_8686);
or U14548 (N_14548,N_12246,N_11401);
or U14549 (N_14549,N_7376,N_10595);
xnor U14550 (N_14550,N_10441,N_7916);
xor U14551 (N_14551,N_10093,N_10379);
nor U14552 (N_14552,N_7225,N_12007);
nand U14553 (N_14553,N_8412,N_9290);
nor U14554 (N_14554,N_10720,N_6624);
xor U14555 (N_14555,N_6921,N_8548);
or U14556 (N_14556,N_6482,N_7307);
xor U14557 (N_14557,N_6885,N_10151);
nor U14558 (N_14558,N_8999,N_7658);
xnor U14559 (N_14559,N_9819,N_10295);
xnor U14560 (N_14560,N_10777,N_7392);
or U14561 (N_14561,N_10013,N_12160);
nand U14562 (N_14562,N_11587,N_7804);
and U14563 (N_14563,N_8995,N_6649);
and U14564 (N_14564,N_9209,N_8101);
nand U14565 (N_14565,N_9514,N_6707);
and U14566 (N_14566,N_12262,N_7720);
xor U14567 (N_14567,N_7403,N_8813);
nand U14568 (N_14568,N_9458,N_9927);
nor U14569 (N_14569,N_8907,N_9039);
nand U14570 (N_14570,N_8241,N_11345);
nor U14571 (N_14571,N_6631,N_12278);
and U14572 (N_14572,N_11652,N_10724);
nor U14573 (N_14573,N_10984,N_10933);
and U14574 (N_14574,N_6452,N_12404);
xnor U14575 (N_14575,N_10893,N_10422);
or U14576 (N_14576,N_7419,N_7113);
nand U14577 (N_14577,N_11663,N_11811);
nand U14578 (N_14578,N_11379,N_7967);
xnor U14579 (N_14579,N_11081,N_7233);
or U14580 (N_14580,N_11934,N_8403);
and U14581 (N_14581,N_12275,N_12137);
nand U14582 (N_14582,N_6408,N_10888);
and U14583 (N_14583,N_9778,N_8586);
or U14584 (N_14584,N_7396,N_11105);
and U14585 (N_14585,N_9877,N_8931);
nor U14586 (N_14586,N_8596,N_10887);
nor U14587 (N_14587,N_9735,N_11082);
xnor U14588 (N_14588,N_12076,N_7439);
and U14589 (N_14589,N_11975,N_12441);
or U14590 (N_14590,N_7386,N_6983);
nor U14591 (N_14591,N_12096,N_7287);
or U14592 (N_14592,N_6613,N_7665);
nand U14593 (N_14593,N_8667,N_8471);
and U14594 (N_14594,N_12489,N_12284);
and U14595 (N_14595,N_8448,N_8928);
nand U14596 (N_14596,N_9352,N_11094);
nand U14597 (N_14597,N_10782,N_12412);
or U14598 (N_14598,N_10103,N_10465);
nand U14599 (N_14599,N_7461,N_11051);
xor U14600 (N_14600,N_11016,N_6328);
and U14601 (N_14601,N_11308,N_7931);
nor U14602 (N_14602,N_6825,N_7297);
nand U14603 (N_14603,N_9278,N_10323);
nand U14604 (N_14604,N_9071,N_7195);
or U14605 (N_14605,N_8457,N_10117);
or U14606 (N_14606,N_7721,N_11664);
nor U14607 (N_14607,N_11263,N_7596);
or U14608 (N_14608,N_8004,N_8787);
or U14609 (N_14609,N_8198,N_6275);
nor U14610 (N_14610,N_9307,N_9322);
nor U14611 (N_14611,N_9370,N_7512);
nor U14612 (N_14612,N_12212,N_10455);
nor U14613 (N_14613,N_9526,N_10866);
and U14614 (N_14614,N_11867,N_6293);
nand U14615 (N_14615,N_7239,N_6259);
nor U14616 (N_14616,N_11091,N_9471);
nand U14617 (N_14617,N_9672,N_9870);
or U14618 (N_14618,N_8260,N_6882);
or U14619 (N_14619,N_11006,N_8423);
xor U14620 (N_14620,N_6857,N_10973);
and U14621 (N_14621,N_8176,N_10577);
or U14622 (N_14622,N_7104,N_10830);
xor U14623 (N_14623,N_9338,N_11932);
xnor U14624 (N_14624,N_8540,N_9133);
and U14625 (N_14625,N_8350,N_10592);
and U14626 (N_14626,N_11674,N_11726);
nor U14627 (N_14627,N_11790,N_8556);
nor U14628 (N_14628,N_8228,N_12110);
nor U14629 (N_14629,N_10368,N_8219);
or U14630 (N_14630,N_6531,N_9962);
or U14631 (N_14631,N_7212,N_10007);
and U14632 (N_14632,N_6530,N_9059);
and U14633 (N_14633,N_6963,N_8637);
xnor U14634 (N_14634,N_6396,N_11176);
xor U14635 (N_14635,N_6732,N_7492);
xnor U14636 (N_14636,N_7489,N_9780);
xor U14637 (N_14637,N_9189,N_9480);
nand U14638 (N_14638,N_6372,N_9408);
nor U14639 (N_14639,N_10113,N_8512);
and U14640 (N_14640,N_12249,N_10962);
and U14641 (N_14641,N_10907,N_7204);
nand U14642 (N_14642,N_8887,N_11740);
nor U14643 (N_14643,N_9255,N_10041);
or U14644 (N_14644,N_7977,N_6339);
nor U14645 (N_14645,N_10760,N_12372);
xor U14646 (N_14646,N_9177,N_11247);
and U14647 (N_14647,N_11505,N_8947);
and U14648 (N_14648,N_7250,N_8566);
nor U14649 (N_14649,N_10000,N_9597);
or U14650 (N_14650,N_11264,N_9380);
and U14651 (N_14651,N_7526,N_7914);
nand U14652 (N_14652,N_7782,N_10805);
or U14653 (N_14653,N_10265,N_11249);
or U14654 (N_14654,N_7667,N_9454);
and U14655 (N_14655,N_10141,N_10583);
nor U14656 (N_14656,N_8517,N_8205);
nand U14657 (N_14657,N_11903,N_7636);
nand U14658 (N_14658,N_6464,N_9284);
and U14659 (N_14659,N_11019,N_9168);
nand U14660 (N_14660,N_11658,N_12167);
nor U14661 (N_14661,N_11124,N_10654);
nor U14662 (N_14662,N_8535,N_6266);
xnor U14663 (N_14663,N_8352,N_6786);
nand U14664 (N_14664,N_11738,N_10640);
and U14665 (N_14665,N_8612,N_10210);
or U14666 (N_14666,N_7650,N_8438);
nand U14667 (N_14667,N_11069,N_7123);
nor U14668 (N_14668,N_10908,N_7598);
nand U14669 (N_14669,N_8382,N_7950);
nor U14670 (N_14670,N_7174,N_8321);
and U14671 (N_14671,N_11416,N_8338);
and U14672 (N_14672,N_10947,N_9333);
nand U14673 (N_14673,N_7040,N_9106);
nand U14674 (N_14674,N_9295,N_9766);
xor U14675 (N_14675,N_10864,N_8577);
and U14676 (N_14676,N_10296,N_9306);
nor U14677 (N_14677,N_10052,N_11373);
nor U14678 (N_14678,N_9934,N_6608);
nor U14679 (N_14679,N_9967,N_10889);
and U14680 (N_14680,N_12022,N_8938);
xnor U14681 (N_14681,N_9090,N_8160);
and U14682 (N_14682,N_11426,N_9136);
or U14683 (N_14683,N_10618,N_6689);
nor U14684 (N_14684,N_7926,N_9835);
or U14685 (N_14685,N_7913,N_11343);
xor U14686 (N_14686,N_8602,N_6563);
and U14687 (N_14687,N_9847,N_10575);
nor U14688 (N_14688,N_11130,N_7427);
and U14689 (N_14689,N_9274,N_9349);
and U14690 (N_14690,N_8975,N_9373);
or U14691 (N_14691,N_9416,N_9520);
xor U14692 (N_14692,N_9947,N_8955);
and U14693 (N_14693,N_10030,N_10405);
nor U14694 (N_14694,N_11969,N_6694);
xnor U14695 (N_14695,N_10906,N_12247);
nand U14696 (N_14696,N_10847,N_7010);
and U14697 (N_14697,N_9075,N_12000);
xnor U14698 (N_14698,N_9994,N_8287);
or U14699 (N_14699,N_6287,N_8046);
nor U14700 (N_14700,N_10292,N_7616);
xor U14701 (N_14701,N_7625,N_8497);
and U14702 (N_14702,N_6946,N_11720);
nand U14703 (N_14703,N_8119,N_9759);
or U14704 (N_14704,N_9137,N_7447);
nand U14705 (N_14705,N_10069,N_8897);
nor U14706 (N_14706,N_10377,N_12426);
and U14707 (N_14707,N_10690,N_6412);
nand U14708 (N_14708,N_7574,N_6691);
nand U14709 (N_14709,N_10599,N_11454);
or U14710 (N_14710,N_11174,N_12458);
and U14711 (N_14711,N_7952,N_11399);
xor U14712 (N_14712,N_11634,N_8484);
nand U14713 (N_14713,N_7473,N_7521);
nand U14714 (N_14714,N_6747,N_9965);
and U14715 (N_14715,N_11273,N_11779);
or U14716 (N_14716,N_8767,N_7941);
xor U14717 (N_14717,N_6508,N_9040);
nor U14718 (N_14718,N_9757,N_12360);
xnor U14719 (N_14719,N_10274,N_7350);
and U14720 (N_14720,N_12150,N_8171);
and U14721 (N_14721,N_9488,N_12423);
or U14722 (N_14722,N_7146,N_12389);
nand U14723 (N_14723,N_12154,N_8789);
xnor U14724 (N_14724,N_11260,N_6905);
or U14725 (N_14725,N_9002,N_10749);
nor U14726 (N_14726,N_11063,N_10855);
xor U14727 (N_14727,N_9265,N_11501);
and U14728 (N_14728,N_7618,N_7608);
xor U14729 (N_14729,N_8963,N_10958);
nand U14730 (N_14730,N_7870,N_7792);
xnor U14731 (N_14731,N_6556,N_7405);
nor U14732 (N_14732,N_7412,N_9578);
and U14733 (N_14733,N_11337,N_9572);
or U14734 (N_14734,N_11703,N_11430);
and U14735 (N_14735,N_9211,N_8169);
nand U14736 (N_14736,N_11398,N_9886);
and U14737 (N_14737,N_10220,N_10648);
and U14738 (N_14738,N_10341,N_6627);
and U14739 (N_14739,N_7373,N_8474);
or U14740 (N_14740,N_11086,N_6733);
nor U14741 (N_14741,N_8476,N_8310);
nand U14742 (N_14742,N_8477,N_9417);
xor U14743 (N_14743,N_9191,N_7060);
or U14744 (N_14744,N_10312,N_8177);
or U14745 (N_14745,N_11248,N_7802);
and U14746 (N_14746,N_11628,N_11434);
and U14747 (N_14747,N_11915,N_9364);
nand U14748 (N_14748,N_9539,N_9756);
nor U14749 (N_14749,N_7701,N_8991);
nor U14750 (N_14750,N_11998,N_7273);
or U14751 (N_14751,N_11735,N_6883);
or U14752 (N_14752,N_8651,N_12349);
and U14753 (N_14753,N_11097,N_11285);
nor U14754 (N_14754,N_8708,N_6943);
or U14755 (N_14755,N_9770,N_8185);
or U14756 (N_14756,N_7586,N_11374);
and U14757 (N_14757,N_8344,N_7706);
nand U14758 (N_14758,N_9272,N_6252);
nor U14759 (N_14759,N_8510,N_10735);
nor U14760 (N_14760,N_10679,N_9998);
nand U14761 (N_14761,N_8342,N_11856);
nor U14762 (N_14762,N_8349,N_7441);
nand U14763 (N_14763,N_8111,N_8332);
or U14764 (N_14764,N_8227,N_9357);
xor U14765 (N_14765,N_8010,N_9285);
and U14766 (N_14766,N_12060,N_12234);
and U14767 (N_14767,N_7821,N_11982);
nor U14768 (N_14768,N_12313,N_12172);
xor U14769 (N_14769,N_11941,N_9632);
nor U14770 (N_14770,N_7699,N_9292);
and U14771 (N_14771,N_10460,N_9377);
nor U14772 (N_14772,N_9482,N_7440);
and U14773 (N_14773,N_7435,N_7192);
nand U14774 (N_14774,N_6662,N_8368);
and U14775 (N_14775,N_9363,N_12136);
nor U14776 (N_14776,N_10283,N_6749);
or U14777 (N_14777,N_6526,N_12199);
xnor U14778 (N_14778,N_12371,N_10593);
or U14779 (N_14779,N_9256,N_9287);
or U14780 (N_14780,N_8217,N_10566);
and U14781 (N_14781,N_10630,N_10716);
nand U14782 (N_14782,N_12291,N_11946);
nand U14783 (N_14783,N_8663,N_9874);
nor U14784 (N_14784,N_10403,N_7187);
xor U14785 (N_14785,N_11191,N_12098);
nor U14786 (N_14786,N_9125,N_6623);
and U14787 (N_14787,N_10354,N_11754);
nand U14788 (N_14788,N_7186,N_11163);
xor U14789 (N_14789,N_10421,N_11204);
xnor U14790 (N_14790,N_7604,N_11088);
or U14791 (N_14791,N_10153,N_6551);
xnor U14792 (N_14792,N_12208,N_8334);
nand U14793 (N_14793,N_9902,N_10814);
nor U14794 (N_14794,N_11480,N_10146);
and U14795 (N_14795,N_6294,N_11728);
nor U14796 (N_14796,N_7313,N_10271);
nor U14797 (N_14797,N_11850,N_10023);
or U14798 (N_14798,N_6723,N_11532);
nor U14799 (N_14799,N_8837,N_8257);
nand U14800 (N_14800,N_7930,N_6681);
and U14801 (N_14801,N_7115,N_9326);
or U14802 (N_14802,N_8494,N_9313);
or U14803 (N_14803,N_12044,N_9409);
nand U14804 (N_14804,N_11389,N_9512);
or U14805 (N_14805,N_12482,N_11787);
nor U14806 (N_14806,N_9403,N_11390);
nor U14807 (N_14807,N_8588,N_6919);
and U14808 (N_14808,N_10344,N_9692);
xnor U14809 (N_14809,N_12170,N_9374);
or U14810 (N_14810,N_12242,N_9398);
or U14811 (N_14811,N_9562,N_12486);
xor U14812 (N_14812,N_10918,N_11540);
and U14813 (N_14813,N_11437,N_11159);
xor U14814 (N_14814,N_12386,N_7888);
and U14815 (N_14815,N_6948,N_8324);
or U14816 (N_14816,N_10551,N_6754);
nand U14817 (N_14817,N_8405,N_9899);
or U14818 (N_14818,N_10632,N_7038);
or U14819 (N_14819,N_7663,N_7452);
or U14820 (N_14820,N_11282,N_10070);
nor U14821 (N_14821,N_8112,N_11422);
nand U14822 (N_14822,N_11948,N_8331);
nor U14823 (N_14823,N_9952,N_7456);
nor U14824 (N_14824,N_7329,N_10547);
xor U14825 (N_14825,N_8449,N_12240);
or U14826 (N_14826,N_8370,N_7117);
or U14827 (N_14827,N_8039,N_10567);
and U14828 (N_14828,N_10088,N_11297);
nand U14829 (N_14829,N_6926,N_8379);
and U14830 (N_14830,N_11573,N_11334);
nand U14831 (N_14831,N_9524,N_11196);
nand U14832 (N_14832,N_7083,N_9113);
and U14833 (N_14833,N_11312,N_10204);
nor U14834 (N_14834,N_9181,N_12035);
nand U14835 (N_14835,N_9600,N_9400);
xnor U14836 (N_14836,N_10466,N_10966);
and U14837 (N_14837,N_11588,N_7560);
nor U14838 (N_14838,N_9477,N_7177);
and U14839 (N_14839,N_10702,N_10542);
xor U14840 (N_14840,N_8826,N_7848);
xor U14841 (N_14841,N_9361,N_10195);
nor U14842 (N_14842,N_7525,N_11997);
nand U14843 (N_14843,N_7907,N_9861);
or U14844 (N_14844,N_8317,N_12286);
nand U14845 (N_14845,N_6814,N_11193);
nand U14846 (N_14846,N_8274,N_7609);
nand U14847 (N_14847,N_9921,N_11240);
nand U14848 (N_14848,N_11629,N_10672);
or U14849 (N_14849,N_11047,N_10457);
xnor U14850 (N_14850,N_6488,N_7911);
and U14851 (N_14851,N_11162,N_11879);
and U14852 (N_14852,N_10763,N_9054);
and U14853 (N_14853,N_7748,N_10524);
and U14854 (N_14854,N_8922,N_6758);
and U14855 (N_14855,N_10839,N_6547);
nor U14856 (N_14856,N_7080,N_9183);
or U14857 (N_14857,N_11816,N_10770);
nand U14858 (N_14858,N_9791,N_11902);
nor U14859 (N_14859,N_8441,N_10638);
and U14860 (N_14860,N_8881,N_8135);
xor U14861 (N_14861,N_6644,N_7945);
or U14862 (N_14862,N_10322,N_11710);
nand U14863 (N_14863,N_8797,N_10021);
nor U14864 (N_14864,N_12141,N_8819);
nand U14865 (N_14865,N_9500,N_9914);
and U14866 (N_14866,N_10706,N_9205);
and U14867 (N_14867,N_10658,N_6394);
and U14868 (N_14868,N_8839,N_7999);
nor U14869 (N_14869,N_9343,N_6979);
nand U14870 (N_14870,N_8745,N_7617);
and U14871 (N_14871,N_9198,N_7613);
and U14872 (N_14872,N_8065,N_10815);
nand U14873 (N_14873,N_7075,N_10584);
nor U14874 (N_14874,N_7763,N_9267);
nor U14875 (N_14875,N_6317,N_11031);
nor U14876 (N_14876,N_8426,N_8834);
nor U14877 (N_14877,N_12015,N_11005);
nor U14878 (N_14878,N_10897,N_8861);
and U14879 (N_14879,N_7424,N_11626);
xnor U14880 (N_14880,N_12219,N_7241);
nor U14881 (N_14881,N_9379,N_8087);
or U14882 (N_14882,N_8313,N_7564);
or U14883 (N_14883,N_12258,N_10372);
or U14884 (N_14884,N_9973,N_9280);
nand U14885 (N_14885,N_9755,N_7826);
nor U14886 (N_14886,N_9028,N_6360);
or U14887 (N_14887,N_8848,N_11591);
nand U14888 (N_14888,N_9340,N_10351);
and U14889 (N_14889,N_11781,N_7627);
and U14890 (N_14890,N_8062,N_11310);
xnor U14891 (N_14891,N_11514,N_8561);
or U14892 (N_14892,N_9875,N_7363);
nand U14893 (N_14893,N_10045,N_11216);
xor U14894 (N_14894,N_11239,N_9158);
or U14895 (N_14895,N_12185,N_7232);
nand U14896 (N_14896,N_11083,N_12419);
nor U14897 (N_14897,N_8013,N_8168);
xor U14898 (N_14898,N_10633,N_10191);
or U14899 (N_14899,N_9427,N_9055);
or U14900 (N_14900,N_9913,N_6868);
xor U14901 (N_14901,N_8115,N_7315);
nor U14902 (N_14902,N_12274,N_11757);
xnor U14903 (N_14903,N_8871,N_8910);
and U14904 (N_14904,N_9103,N_6327);
and U14905 (N_14905,N_7369,N_6757);
nand U14906 (N_14906,N_9316,N_9384);
and U14907 (N_14907,N_10856,N_9798);
and U14908 (N_14908,N_11885,N_7886);
and U14909 (N_14909,N_7051,N_11221);
and U14910 (N_14910,N_12244,N_9625);
and U14911 (N_14911,N_10251,N_11807);
nor U14912 (N_14912,N_11567,N_10282);
nand U14913 (N_14913,N_11307,N_7768);
or U14914 (N_14914,N_9230,N_11933);
or U14915 (N_14915,N_8549,N_9174);
xnor U14916 (N_14916,N_12333,N_6272);
nand U14917 (N_14917,N_12184,N_12232);
xnor U14918 (N_14918,N_8739,N_10386);
or U14919 (N_14919,N_12413,N_11871);
nor U14920 (N_14920,N_8912,N_9143);
xnor U14921 (N_14921,N_10222,N_10602);
xor U14922 (N_14922,N_11113,N_11368);
nand U14923 (N_14923,N_11467,N_9457);
xor U14924 (N_14924,N_7773,N_7518);
and U14925 (N_14925,N_11817,N_7785);
nand U14926 (N_14926,N_12290,N_11330);
nor U14927 (N_14927,N_9387,N_9412);
nor U14928 (N_14928,N_7084,N_7936);
or U14929 (N_14929,N_6577,N_6320);
nor U14930 (N_14930,N_10493,N_9966);
nand U14931 (N_14931,N_11689,N_11417);
or U14932 (N_14932,N_8719,N_7418);
xnor U14933 (N_14933,N_6284,N_7500);
and U14934 (N_14934,N_10768,N_12017);
xnor U14935 (N_14935,N_7740,N_10809);
or U14936 (N_14936,N_10868,N_10155);
and U14937 (N_14937,N_11906,N_9309);
nor U14938 (N_14938,N_12004,N_8547);
nor U14939 (N_14939,N_10444,N_12122);
nor U14940 (N_14940,N_6335,N_12490);
or U14941 (N_14941,N_11599,N_11412);
nand U14942 (N_14942,N_10340,N_9787);
xor U14943 (N_14943,N_7155,N_7488);
nand U14944 (N_14944,N_8211,N_10243);
and U14945 (N_14945,N_8914,N_11041);
or U14946 (N_14946,N_7543,N_8459);
xor U14947 (N_14947,N_9803,N_10068);
or U14948 (N_14948,N_8305,N_11589);
xnor U14949 (N_14949,N_9366,N_6957);
xor U14950 (N_14950,N_11479,N_6990);
nand U14951 (N_14951,N_8773,N_6431);
or U14952 (N_14952,N_7062,N_12392);
or U14953 (N_14953,N_12277,N_11736);
xor U14954 (N_14954,N_12211,N_6901);
xnor U14955 (N_14955,N_9534,N_9060);
or U14956 (N_14956,N_9948,N_9310);
or U14957 (N_14957,N_12151,N_8164);
nand U14958 (N_14958,N_11370,N_10845);
nand U14959 (N_14959,N_10743,N_12376);
nor U14960 (N_14960,N_7450,N_7018);
and U14961 (N_14961,N_10614,N_8072);
nor U14962 (N_14962,N_7964,N_10732);
nand U14963 (N_14963,N_11227,N_11722);
or U14964 (N_14964,N_11338,N_8750);
nand U14965 (N_14965,N_6451,N_11140);
and U14966 (N_14966,N_8687,N_10925);
nor U14967 (N_14967,N_10380,N_8579);
nand U14968 (N_14968,N_8908,N_7867);
or U14969 (N_14969,N_9525,N_10919);
nand U14970 (N_14970,N_7990,N_7253);
nand U14971 (N_14971,N_10972,N_10801);
nor U14972 (N_14972,N_9634,N_6794);
nor U14973 (N_14973,N_9529,N_11503);
or U14974 (N_14974,N_9738,N_7898);
and U14975 (N_14975,N_10751,N_11854);
and U14976 (N_14976,N_9844,N_10174);
nor U14977 (N_14977,N_11527,N_7820);
and U14978 (N_14978,N_9790,N_7009);
or U14979 (N_14979,N_8265,N_10252);
nand U14980 (N_14980,N_6397,N_9045);
nand U14981 (N_14981,N_8525,N_7423);
nand U14982 (N_14982,N_6894,N_6695);
nand U14983 (N_14983,N_8491,N_10937);
nand U14984 (N_14984,N_10765,N_7819);
xor U14985 (N_14985,N_11145,N_11494);
nor U14986 (N_14986,N_10335,N_6609);
nor U14987 (N_14987,N_7317,N_6840);
nor U14988 (N_14988,N_7086,N_6485);
xor U14989 (N_14989,N_10429,N_11541);
xnor U14990 (N_14990,N_12067,N_7364);
nand U14991 (N_14991,N_9220,N_11474);
xor U14992 (N_14992,N_7090,N_8232);
and U14993 (N_14993,N_11828,N_8495);
and U14994 (N_14994,N_9487,N_11150);
and U14995 (N_14995,N_6842,N_10728);
nor U14996 (N_14996,N_8764,N_8683);
nor U14997 (N_14997,N_10279,N_6809);
nor U14998 (N_14998,N_6969,N_11770);
nand U14999 (N_14999,N_10533,N_10820);
nand U15000 (N_15000,N_10348,N_7031);
nand U15001 (N_15001,N_8175,N_12011);
and U15002 (N_15002,N_6499,N_9515);
xor U15003 (N_15003,N_7624,N_11821);
or U15004 (N_15004,N_8435,N_8952);
xnor U15005 (N_15005,N_9975,N_11809);
or U15006 (N_15006,N_10260,N_12182);
xor U15007 (N_15007,N_7494,N_11188);
nand U15008 (N_15008,N_12478,N_7769);
nand U15009 (N_15009,N_6510,N_12442);
and U15010 (N_15010,N_7073,N_6871);
or U15011 (N_15011,N_11896,N_7764);
or U15012 (N_15012,N_8564,N_10173);
and U15013 (N_15013,N_9623,N_10987);
xnor U15014 (N_15014,N_11043,N_11716);
and U15015 (N_15015,N_10748,N_7154);
and U15016 (N_15016,N_12399,N_11978);
or U15017 (N_15017,N_11322,N_6424);
and U15018 (N_15018,N_11572,N_11335);
nor U15019 (N_15019,N_11895,N_8290);
nor U15020 (N_15020,N_10813,N_9362);
or U15021 (N_15021,N_9301,N_10090);
nor U15022 (N_15022,N_11189,N_7262);
xnor U15023 (N_15023,N_6823,N_9985);
nand U15024 (N_15024,N_7030,N_7876);
xor U15025 (N_15025,N_11393,N_6660);
nand U15026 (N_15026,N_7158,N_7008);
nand U15027 (N_15027,N_9406,N_12287);
and U15028 (N_15028,N_9797,N_9993);
or U15029 (N_15029,N_9392,N_7059);
or U15030 (N_15030,N_7797,N_11313);
or U15031 (N_15031,N_7466,N_9684);
nand U15032 (N_15032,N_9745,N_6520);
and U15033 (N_15033,N_9050,N_10920);
or U15034 (N_15034,N_8282,N_9462);
nand U15035 (N_15035,N_7813,N_8118);
or U15036 (N_15036,N_12496,N_10357);
xor U15037 (N_15037,N_8770,N_10084);
or U15038 (N_15038,N_9527,N_8978);
nand U15039 (N_15039,N_7181,N_10983);
or U15040 (N_15040,N_9992,N_7210);
or U15041 (N_15041,N_7756,N_10019);
and U15042 (N_15042,N_10325,N_11080);
or U15043 (N_15043,N_11340,N_10401);
or U15044 (N_15044,N_9332,N_9166);
or U15045 (N_15045,N_10249,N_6590);
xnor U15046 (N_15046,N_8740,N_8728);
xor U15047 (N_15047,N_8161,N_6616);
and U15048 (N_15048,N_9660,N_10895);
nand U15049 (N_15049,N_10389,N_9238);
and U15050 (N_15050,N_11775,N_8213);
and U15051 (N_15051,N_6778,N_6505);
or U15052 (N_15052,N_6509,N_6667);
or U15053 (N_15053,N_11583,N_12140);
nand U15054 (N_15054,N_7943,N_10511);
and U15055 (N_15055,N_10767,N_11229);
nand U15056 (N_15056,N_10362,N_8685);
nand U15057 (N_15057,N_9810,N_6955);
or U15058 (N_15058,N_6654,N_9640);
nand U15059 (N_15059,N_8225,N_7328);
nand U15060 (N_15060,N_8021,N_11525);
or U15061 (N_15061,N_8982,N_9250);
nand U15062 (N_15062,N_9139,N_11468);
nor U15063 (N_15063,N_8769,N_12028);
or U15064 (N_15064,N_6479,N_11194);
and U15065 (N_15065,N_6942,N_8059);
or U15066 (N_15066,N_11493,N_9192);
and U15067 (N_15067,N_12059,N_8189);
nor U15068 (N_15068,N_8778,N_9628);
or U15069 (N_15069,N_6269,N_9863);
and U15070 (N_15070,N_9099,N_6977);
or U15071 (N_15071,N_7323,N_7421);
nand U15072 (N_15072,N_6910,N_7020);
and U15073 (N_15073,N_9269,N_9399);
nand U15074 (N_15074,N_9999,N_7853);
nor U15075 (N_15075,N_11428,N_6491);
nor U15076 (N_15076,N_9609,N_10833);
nand U15077 (N_15077,N_11272,N_6390);
xor U15078 (N_15078,N_11126,N_6473);
nand U15079 (N_15079,N_6951,N_10400);
nor U15080 (N_15080,N_6827,N_6950);
and U15081 (N_15081,N_6576,N_11032);
xor U15082 (N_15082,N_6728,N_9659);
xnor U15083 (N_15083,N_10071,N_8732);
and U15084 (N_15084,N_9658,N_8270);
nor U15085 (N_15085,N_9981,N_6489);
or U15086 (N_15086,N_10142,N_6930);
xor U15087 (N_15087,N_10257,N_8870);
or U15088 (N_15088,N_8624,N_12190);
xor U15089 (N_15089,N_9552,N_6455);
xor U15090 (N_15090,N_7463,N_8664);
nand U15091 (N_15091,N_8060,N_10108);
nor U15092 (N_15092,N_10843,N_9593);
xnor U15093 (N_15093,N_8988,N_11799);
xor U15094 (N_15094,N_12306,N_6546);
and U15095 (N_15095,N_11846,N_11074);
xor U15096 (N_15096,N_8023,N_11391);
and U15097 (N_15097,N_12317,N_6626);
nor U15098 (N_15098,N_9700,N_7659);
and U15099 (N_15099,N_9239,N_7022);
and U15100 (N_15100,N_10757,N_10363);
xor U15101 (N_15101,N_10118,N_8110);
and U15102 (N_15102,N_9928,N_10144);
or U15103 (N_15103,N_10620,N_9565);
nor U15104 (N_15104,N_7675,N_8790);
and U15105 (N_15105,N_10959,N_11711);
nor U15106 (N_15106,N_8076,N_10560);
xor U15107 (N_15107,N_8793,N_11488);
nand U15108 (N_15108,N_7354,N_7638);
nor U15109 (N_15109,N_7046,N_12048);
nand U15110 (N_15110,N_8467,N_8304);
nand U15111 (N_15111,N_10456,N_8195);
nand U15112 (N_15112,N_10304,N_12363);
or U15113 (N_15113,N_10122,N_6503);
or U15114 (N_15114,N_10571,N_11670);
nand U15115 (N_15115,N_6976,N_9023);
xnor U15116 (N_15116,N_10816,N_8208);
xor U15117 (N_15117,N_10186,N_11853);
xor U15118 (N_15118,N_7910,N_10999);
and U15119 (N_15119,N_10485,N_10062);
xor U15120 (N_15120,N_10289,N_7095);
and U15121 (N_15121,N_12488,N_8868);
or U15122 (N_15122,N_9411,N_12192);
nand U15123 (N_15123,N_8617,N_6808);
nand U15124 (N_15124,N_6502,N_12014);
nor U15125 (N_15125,N_8470,N_7839);
xnor U15126 (N_15126,N_7406,N_8092);
nor U15127 (N_15127,N_7664,N_12034);
and U15128 (N_15128,N_6459,N_11463);
and U15129 (N_15129,N_11603,N_9950);
nand U15130 (N_15130,N_7772,N_8353);
nor U15131 (N_15131,N_11547,N_11045);
or U15132 (N_15132,N_10586,N_6617);
nand U15133 (N_15133,N_6506,N_9243);
nor U15134 (N_15134,N_11070,N_10582);
nor U15135 (N_15135,N_7700,N_11093);
or U15136 (N_15136,N_10447,N_12254);
xor U15137 (N_15137,N_7339,N_12026);
or U15138 (N_15138,N_11420,N_10913);
xor U15139 (N_15139,N_10705,N_8116);
nand U15140 (N_15140,N_6978,N_11782);
nor U15141 (N_15141,N_7389,N_9221);
and U15142 (N_15142,N_11405,N_11486);
and U15143 (N_15143,N_11226,N_11222);
xor U15144 (N_15144,N_9080,N_7145);
and U15145 (N_15145,N_9004,N_9456);
or U15146 (N_15146,N_10076,N_6769);
and U15147 (N_15147,N_9850,N_7533);
nand U15148 (N_15148,N_10545,N_8688);
nand U15149 (N_15149,N_8980,N_7383);
and U15150 (N_15150,N_10261,N_11383);
nor U15151 (N_15151,N_7953,N_10385);
or U15152 (N_15152,N_9345,N_10886);
or U15153 (N_15153,N_11361,N_12378);
or U15154 (N_15154,N_9424,N_6674);
nor U15155 (N_15155,N_9619,N_8084);
nor U15156 (N_15156,N_10903,N_7707);
nor U15157 (N_15157,N_7757,N_8541);
or U15158 (N_15158,N_12071,N_9312);
nor U15159 (N_15159,N_7033,N_10989);
nand U15160 (N_15160,N_10169,N_12379);
xnor U15161 (N_15161,N_9777,N_6887);
and U15162 (N_15162,N_11721,N_11075);
or U15163 (N_15163,N_9768,N_8285);
xnor U15164 (N_15164,N_7579,N_7561);
and U15165 (N_15165,N_8097,N_10425);
nand U15166 (N_15166,N_6630,N_11958);
xor U15167 (N_15167,N_7141,N_10581);
xor U15168 (N_15168,N_7175,N_12079);
nand U15169 (N_15169,N_8179,N_11881);
or U15170 (N_15170,N_9036,N_10588);
nand U15171 (N_15171,N_8050,N_7843);
nand U15172 (N_15172,N_11496,N_10018);
nand U15173 (N_15173,N_9662,N_12097);
xor U15174 (N_15174,N_8183,N_7902);
or U15175 (N_15175,N_8804,N_7901);
or U15176 (N_15176,N_8802,N_11590);
nand U15177 (N_15177,N_11134,N_12200);
xor U15178 (N_15178,N_11955,N_10905);
nand U15179 (N_15179,N_7014,N_9681);
xor U15180 (N_15180,N_6501,N_8247);
nand U15181 (N_15181,N_6640,N_7179);
or U15182 (N_15182,N_8276,N_9832);
xnor U15183 (N_15183,N_6917,N_12430);
and U15184 (N_15184,N_7550,N_11036);
nand U15185 (N_15185,N_7679,N_7965);
xor U15186 (N_15186,N_12350,N_11598);
and U15187 (N_15187,N_11483,N_11901);
nor U15188 (N_15188,N_11078,N_6929);
and U15189 (N_15189,N_12409,N_11783);
and U15190 (N_15190,N_11060,N_7605);
xor U15191 (N_15191,N_10498,N_12418);
or U15192 (N_15192,N_7716,N_9937);
nand U15193 (N_15193,N_8505,N_8937);
nor U15194 (N_15194,N_10256,N_8694);
or U15195 (N_15195,N_11630,N_7676);
and U15196 (N_15196,N_7677,N_8319);
nand U15197 (N_15197,N_10305,N_10784);
nor U15198 (N_15198,N_11039,N_10359);
xor U15199 (N_15199,N_10025,N_9812);
nor U15200 (N_15200,N_11924,N_8842);
nor U15201 (N_15201,N_8173,N_11864);
nand U15202 (N_15202,N_10129,N_8419);
nor U15203 (N_15203,N_11460,N_7216);
or U15204 (N_15204,N_12408,N_10550);
nor U15205 (N_15205,N_10114,N_12462);
nor U15206 (N_15206,N_10789,N_11951);
xnor U15207 (N_15207,N_6735,N_7021);
and U15208 (N_15208,N_8251,N_8063);
and U15209 (N_15209,N_8735,N_7143);
nor U15210 (N_15210,N_8193,N_7097);
nor U15211 (N_15211,N_11439,N_10208);
or U15212 (N_15212,N_7840,N_8560);
xor U15213 (N_15213,N_12109,N_9935);
or U15214 (N_15214,N_9069,N_7520);
or U15215 (N_15215,N_10610,N_9779);
and U15216 (N_15216,N_9022,N_10727);
and U15217 (N_15217,N_8759,N_7290);
and U15218 (N_15218,N_10504,N_11862);
nor U15219 (N_15219,N_7100,N_11151);
xnor U15220 (N_15220,N_9916,N_10276);
and U15221 (N_15221,N_11929,N_8665);
nor U15222 (N_15222,N_6515,N_11876);
or U15223 (N_15223,N_9393,N_7457);
nand U15224 (N_15224,N_7305,N_6585);
and U15225 (N_15225,N_10443,N_12301);
or U15226 (N_15226,N_6893,N_12120);
nor U15227 (N_15227,N_8335,N_6896);
and U15228 (N_15228,N_11052,N_8256);
or U15229 (N_15229,N_10154,N_7653);
nor U15230 (N_15230,N_11826,N_8956);
and U15231 (N_15231,N_10188,N_12237);
or U15232 (N_15232,N_10360,N_10552);
or U15233 (N_15233,N_7127,N_6469);
nor U15234 (N_15234,N_10224,N_8516);
and U15235 (N_15235,N_12312,N_7558);
and U15236 (N_15236,N_9056,N_11120);
nand U15237 (N_15237,N_8726,N_10297);
nand U15238 (N_15238,N_8167,N_6615);
nand U15239 (N_15239,N_10391,N_9194);
or U15240 (N_15240,N_10516,N_7690);
or U15241 (N_15241,N_11875,N_12480);
nand U15242 (N_15242,N_11099,N_11973);
nand U15243 (N_15243,N_8224,N_9919);
nor U15244 (N_15244,N_8020,N_8671);
nand U15245 (N_15245,N_7160,N_10646);
nor U15246 (N_15246,N_8333,N_11578);
nand U15247 (N_15247,N_9687,N_10704);
nand U15248 (N_15248,N_8898,N_8997);
and U15249 (N_15249,N_11988,N_6420);
or U15250 (N_15250,N_11916,N_7367);
and U15251 (N_15251,N_8371,N_11751);
nand U15252 (N_15252,N_6907,N_11974);
and U15253 (N_15253,N_10994,N_9321);
nor U15254 (N_15254,N_9465,N_12233);
and U15255 (N_15255,N_9519,N_10219);
nor U15256 (N_15256,N_6439,N_11027);
nor U15257 (N_15257,N_11471,N_9971);
and U15258 (N_15258,N_6323,N_9956);
or U15259 (N_15259,N_10590,N_6985);
xor U15260 (N_15260,N_10073,N_9441);
or U15261 (N_15261,N_8812,N_8153);
and U15262 (N_15262,N_10028,N_10235);
or U15263 (N_15263,N_7968,N_11611);
and U15264 (N_15264,N_7264,N_10139);
nor U15265 (N_15265,N_8872,N_7416);
nor U15266 (N_15266,N_11765,N_8996);
xor U15267 (N_15267,N_9873,N_9815);
or U15268 (N_15268,N_8544,N_12222);
and U15269 (N_15269,N_11976,N_7215);
and U15270 (N_15270,N_7549,N_8024);
and U15271 (N_15271,N_10876,N_11286);
xor U15272 (N_15272,N_11419,N_7750);
nor U15273 (N_15273,N_9098,N_8075);
and U15274 (N_15274,N_9892,N_9109);
nand U15275 (N_15275,N_11609,N_9296);
or U15276 (N_15276,N_11552,N_9262);
nand U15277 (N_15277,N_11104,N_11024);
and U15278 (N_15278,N_7718,N_8915);
or U15279 (N_15279,N_8109,N_11605);
or U15280 (N_15280,N_6991,N_11700);
and U15281 (N_15281,N_10089,N_10004);
and U15282 (N_15282,N_9077,N_7324);
nand U15283 (N_15283,N_11513,N_7091);
or U15284 (N_15284,N_10625,N_11143);
or U15285 (N_15285,N_8388,N_7984);
and U15286 (N_15286,N_9945,N_9673);
nor U15287 (N_15287,N_7345,N_7254);
nand U15288 (N_15288,N_9185,N_6899);
and U15289 (N_15289,N_11073,N_11314);
and U15290 (N_15290,N_8852,N_10980);
and U15291 (N_15291,N_8077,N_6604);
or U15292 (N_15292,N_12153,N_8894);
xnor U15293 (N_15293,N_8180,N_7880);
xnor U15294 (N_15294,N_11640,N_12158);
nor U15295 (N_15295,N_7429,N_7566);
nand U15296 (N_15296,N_12227,N_6529);
or U15297 (N_15297,N_8570,N_11808);
nor U15298 (N_15298,N_6696,N_8369);
and U15299 (N_15299,N_7479,N_11979);
and U15300 (N_15300,N_7563,N_8553);
and U15301 (N_15301,N_8875,N_8844);
nor U15302 (N_15302,N_8204,N_7052);
or U15303 (N_15303,N_12006,N_12159);
nor U15304 (N_15304,N_8150,N_8673);
or U15305 (N_15305,N_11575,N_6566);
xor U15306 (N_15306,N_6261,N_6449);
or U15307 (N_15307,N_7201,N_10346);
nand U15308 (N_15308,N_7581,N_8069);
xnor U15309 (N_15309,N_10136,N_7407);
or U15310 (N_15310,N_10396,N_6874);
and U15311 (N_15311,N_10048,N_11692);
and U15312 (N_15312,N_6968,N_6773);
nand U15313 (N_15313,N_10513,N_11435);
or U15314 (N_15314,N_10280,N_8713);
nor U15315 (N_15315,N_10853,N_9680);
and U15316 (N_15316,N_11098,N_10719);
or U15317 (N_15317,N_7760,N_8704);
nand U15318 (N_15318,N_9464,N_10408);
and U15319 (N_15319,N_8240,N_11355);
and U15320 (N_15320,N_10301,N_8607);
nor U15321 (N_15321,N_6798,N_7352);
or U15322 (N_15322,N_7973,N_12138);
and U15323 (N_15323,N_8011,N_10406);
xor U15324 (N_15324,N_7759,N_11108);
or U15325 (N_15325,N_9007,N_7043);
nor U15326 (N_15326,N_10870,N_7632);
and U15327 (N_15327,N_8979,N_8244);
or U15328 (N_15328,N_8925,N_9765);
xor U15329 (N_15329,N_6460,N_10217);
nor U15330 (N_15330,N_9794,N_6470);
nor U15331 (N_15331,N_9217,N_7614);
xor U15332 (N_15332,N_7992,N_6534);
nor U15333 (N_15333,N_11904,N_10066);
nand U15334 (N_15334,N_9656,N_12085);
or U15335 (N_15335,N_11040,N_11243);
or U15336 (N_15336,N_8481,N_9666);
and U15337 (N_15337,N_12093,N_10761);
nand U15338 (N_15338,N_12383,N_11443);
xor U15339 (N_15339,N_9924,N_11610);
or U15340 (N_15340,N_9522,N_7148);
or U15341 (N_15341,N_7326,N_10339);
and U15342 (N_15342,N_8727,N_6297);
nor U15343 (N_15343,N_10879,N_7045);
and U15344 (N_15344,N_8559,N_10364);
nand U15345 (N_15345,N_7988,N_10836);
nor U15346 (N_15346,N_6492,N_11231);
or U15347 (N_15347,N_9909,N_11517);
xor U15348 (N_15348,N_9897,N_8760);
and U15349 (N_15349,N_6465,N_10467);
xor U15350 (N_15350,N_9557,N_9843);
or U15351 (N_15351,N_7505,N_10882);
xor U15352 (N_15352,N_6700,N_12406);
and U15353 (N_15353,N_8362,N_9836);
and U15354 (N_15354,N_10082,N_9750);
and U15355 (N_15355,N_8777,N_7585);
nor U15356 (N_15356,N_10544,N_6416);
nand U15357 (N_15357,N_7975,N_9867);
or U15358 (N_15358,N_6330,N_8822);
or U15359 (N_15359,N_8339,N_11214);
and U15360 (N_15360,N_12216,N_8699);
and U15361 (N_15361,N_10434,N_12127);
nand U15362 (N_15362,N_7281,N_9330);
and U15363 (N_15363,N_8853,N_11371);
nand U15364 (N_15364,N_10495,N_7499);
nor U15365 (N_15365,N_9643,N_7513);
nor U15366 (N_15366,N_9496,N_9652);
nor U15367 (N_15367,N_8815,N_7226);
xor U15368 (N_15368,N_8567,N_10190);
nor U15369 (N_15369,N_10929,N_6354);
or U15370 (N_15370,N_6884,N_10273);
nand U15371 (N_15371,N_8573,N_7007);
nor U15372 (N_15372,N_10381,N_9831);
nand U15373 (N_15373,N_10863,N_11008);
xnor U15374 (N_15374,N_11152,N_8293);
or U15375 (N_15375,N_7067,N_8163);
xnor U15376 (N_15376,N_7628,N_11792);
xor U15377 (N_15377,N_9453,N_10772);
and U15378 (N_15378,N_8656,N_6559);
nor U15379 (N_15379,N_7793,N_7925);
or U15380 (N_15380,N_10026,N_7747);
or U15381 (N_15381,N_12003,N_11585);
or U15382 (N_15382,N_12415,N_7420);
and U15383 (N_15383,N_9058,N_8744);
or U15384 (N_15384,N_12131,N_6777);
nand U15385 (N_15385,N_11631,N_9665);
nor U15386 (N_15386,N_9912,N_9248);
nor U15387 (N_15387,N_8096,N_10343);
nand U15388 (N_15388,N_7584,N_8893);
nand U15389 (N_15389,N_11798,N_9685);
and U15390 (N_15390,N_9627,N_10209);
xor U15391 (N_15391,N_8152,N_6832);
xnor U15392 (N_15392,N_6705,N_8057);
xnor U15393 (N_15393,N_6342,N_9348);
nand U15394 (N_15394,N_6785,N_11586);
xnor U15395 (N_15395,N_6967,N_11620);
nor U15396 (N_15396,N_9550,N_7963);
xnor U15397 (N_15397,N_9978,N_11789);
nand U15398 (N_15398,N_11768,N_8998);
or U15399 (N_15399,N_11185,N_11386);
or U15400 (N_15400,N_6725,N_9419);
and U15401 (N_15401,N_8252,N_9851);
or U15402 (N_15402,N_10255,N_9724);
xnor U15403 (N_15403,N_7635,N_9930);
and U15404 (N_15404,N_10934,N_9599);
nand U15405 (N_15405,N_6811,N_7836);
or U15406 (N_15406,N_6622,N_9132);
and U15407 (N_15407,N_7266,N_8926);
xnor U15408 (N_15408,N_9342,N_8243);
and U15409 (N_15409,N_9492,N_11408);
nor U15410 (N_15410,N_9311,N_8792);
or U15411 (N_15411,N_10875,N_9688);
nor U15412 (N_15412,N_6675,N_11655);
and U15413 (N_15413,N_7736,N_8758);
xnor U15414 (N_15414,N_11363,N_9949);
nand U15415 (N_15415,N_6753,N_6542);
nand U15416 (N_15416,N_8455,N_7107);
or U15417 (N_15417,N_8218,N_10696);
and U15418 (N_15418,N_8829,N_8143);
xnor U15419 (N_15419,N_11883,N_6457);
nor U15420 (N_15420,N_10375,N_7571);
xnor U15421 (N_15421,N_7969,N_8246);
xor U15422 (N_15422,N_8045,N_10390);
nand U15423 (N_15423,N_8742,N_8880);
and U15424 (N_15424,N_10178,N_10212);
xor U15425 (N_15425,N_12293,N_8031);
nand U15426 (N_15426,N_9200,N_10200);
nor U15427 (N_15427,N_10192,N_11110);
xor U15428 (N_15428,N_12444,N_9746);
or U15429 (N_15429,N_9044,N_10884);
or U15430 (N_15430,N_10482,N_11967);
and U15431 (N_15431,N_6964,N_12302);
or U15432 (N_15432,N_6810,N_12494);
xnor U15433 (N_15433,N_10671,N_9371);
xor U15434 (N_15434,N_10022,N_6599);
nand U15435 (N_15435,N_8250,N_9917);
and U15436 (N_15436,N_11281,N_8885);
or U15437 (N_15437,N_7597,N_9091);
nand U15438 (N_15438,N_11555,N_8655);
nand U15439 (N_15439,N_7535,N_11470);
nor U15440 (N_15440,N_11923,N_11806);
xnor U15441 (N_15441,N_6407,N_12259);
and U15442 (N_15442,N_9946,N_11769);
xnor U15443 (N_15443,N_10831,N_11804);
and U15444 (N_15444,N_7849,N_12229);
xor U15445 (N_15445,N_12411,N_7206);
or U15446 (N_15446,N_12367,N_8136);
and U15447 (N_15447,N_9019,N_10651);
or U15448 (N_15448,N_6973,N_10170);
nand U15449 (N_15449,N_7539,N_9860);
and U15450 (N_15450,N_11292,N_8882);
or U15451 (N_15451,N_7857,N_6998);
and U15452 (N_15452,N_11701,N_10015);
nor U15453 (N_15453,N_6285,N_10060);
and U15454 (N_15454,N_11554,N_10578);
or U15455 (N_15455,N_7829,N_6805);
and U15456 (N_15456,N_10850,N_8594);
or U15457 (N_15457,N_6303,N_9649);
and U15458 (N_15458,N_9561,N_10140);
nor U15459 (N_15459,N_9161,N_7167);
xor U15460 (N_15460,N_6960,N_6366);
and U15461 (N_15461,N_11956,N_11161);
xor U15462 (N_15462,N_11612,N_12008);
nand U15463 (N_15463,N_7390,N_7217);
xor U15464 (N_15464,N_9696,N_10557);
nand U15465 (N_15465,N_6255,N_9129);
xor U15466 (N_15466,N_12491,N_8626);
nor U15467 (N_15467,N_11794,N_11199);
or U15468 (N_15468,N_7529,N_11936);
or U15469 (N_15469,N_7436,N_10462);
and U15470 (N_15470,N_9439,N_7378);
nor U15471 (N_15471,N_8002,N_8237);
and U15472 (N_15472,N_10010,N_7076);
or U15473 (N_15473,N_7208,N_7272);
nor U15474 (N_15474,N_7744,N_12001);
and U15475 (N_15475,N_12107,N_11459);
nand U15476 (N_15476,N_7749,N_7355);
or U15477 (N_15477,N_8623,N_10264);
xor U15478 (N_15478,N_11560,N_8950);
xnor U15479 (N_15479,N_11327,N_6820);
or U15480 (N_15480,N_7351,N_12101);
nor U15481 (N_15481,N_7058,N_12327);
and U15482 (N_15482,N_11473,N_8375);
or U15483 (N_15483,N_11115,N_9686);
xor U15484 (N_15484,N_9753,N_6395);
xor U15485 (N_15485,N_7387,N_11529);
or U15486 (N_15486,N_12369,N_10311);
nor U15487 (N_15487,N_10639,N_11275);
and U15488 (N_15488,N_10415,N_7218);
xor U15489 (N_15489,N_10837,N_8284);
and U15490 (N_15490,N_8917,N_10649);
and U15491 (N_15491,N_9335,N_7991);
or U15492 (N_15492,N_7572,N_10175);
nand U15493 (N_15493,N_7183,N_9675);
or U15494 (N_15494,N_6537,N_6384);
and U15495 (N_15495,N_6642,N_6543);
and U15496 (N_15496,N_9304,N_9383);
nand U15497 (N_15497,N_11482,N_10410);
nand U15498 (N_15498,N_11072,N_11649);
xnor U15499 (N_15499,N_8580,N_7776);
nor U15500 (N_15500,N_11677,N_6648);
or U15501 (N_15501,N_12057,N_8974);
nand U15502 (N_15502,N_10943,N_10713);
and U15503 (N_15503,N_8229,N_12294);
nand U15504 (N_15504,N_12387,N_10744);
or U15505 (N_15505,N_7152,N_9469);
nor U15506 (N_15506,N_10492,N_11597);
and U15507 (N_15507,N_6763,N_8628);
nand U15508 (N_15508,N_12473,N_11595);
or U15509 (N_15509,N_7987,N_9678);
nor U15510 (N_15510,N_11458,N_11380);
and U15511 (N_15511,N_8608,N_11796);
and U15512 (N_15512,N_11788,N_10904);
xnor U15513 (N_15513,N_7065,N_11257);
nor U15514 (N_15514,N_6605,N_11138);
nor U15515 (N_15515,N_10558,N_8990);
xor U15516 (N_15516,N_9881,N_7327);
or U15517 (N_15517,N_10967,N_6301);
nand U15518 (N_15518,N_6517,N_10394);
xnor U15519 (N_15519,N_10891,N_6643);
or U15520 (N_15520,N_10711,N_7284);
and U15521 (N_15521,N_11840,N_10480);
xor U15522 (N_15522,N_11569,N_9499);
or U15523 (N_15523,N_6312,N_6516);
nor U15524 (N_15524,N_9888,N_7469);
and U15525 (N_15525,N_11607,N_10158);
or U15526 (N_15526,N_11667,N_11833);
and U15527 (N_15527,N_10211,N_11316);
xor U15528 (N_15528,N_9088,N_8036);
and U15529 (N_15529,N_11699,N_7508);
nand U15530 (N_15530,N_7168,N_9580);
xor U15531 (N_15531,N_11608,N_8318);
nand U15532 (N_15532,N_6703,N_8029);
or U15533 (N_15533,N_8783,N_10160);
or U15534 (N_15534,N_9455,N_11058);
nor U15535 (N_15535,N_6712,N_11329);
xnor U15536 (N_15536,N_8808,N_8207);
and U15537 (N_15537,N_6949,N_9922);
nor U15538 (N_15538,N_7552,N_7399);
nor U15539 (N_15539,N_8396,N_11827);
nor U15540 (N_15540,N_11296,N_6854);
and U15541 (N_15541,N_12256,N_10051);
or U15542 (N_15542,N_11323,N_8746);
nor U15543 (N_15543,N_11920,N_9644);
xor U15544 (N_15544,N_7986,N_7737);
xor U15545 (N_15545,N_6344,N_12322);
and U15546 (N_15546,N_8584,N_7314);
nor U15547 (N_15547,N_11669,N_7942);
or U15548 (N_15548,N_12056,N_6748);
and U15549 (N_15549,N_12068,N_9277);
or U15550 (N_15550,N_9030,N_11290);
xnor U15551 (N_15551,N_10033,N_12358);
and U15552 (N_15552,N_7343,N_12436);
and U15553 (N_15553,N_6250,N_7004);
or U15554 (N_15554,N_9426,N_8969);
and U15555 (N_15555,N_9822,N_9064);
xor U15556 (N_15556,N_11702,N_10823);
and U15557 (N_15557,N_8108,N_12119);
nand U15558 (N_15558,N_11141,N_11944);
nand U15559 (N_15559,N_8589,N_10793);
xor U15560 (N_15560,N_11007,N_10193);
nor U15561 (N_15561,N_7754,N_11544);
or U15562 (N_15562,N_10231,N_10537);
nor U15563 (N_15563,N_8082,N_10786);
xnor U15564 (N_15564,N_9564,N_12464);
and U15565 (N_15565,N_11440,N_10954);
and U15566 (N_15566,N_8526,N_7799);
nand U15567 (N_15567,N_8192,N_8340);
and U15568 (N_15568,N_10458,N_6504);
nand U15569 (N_15569,N_8647,N_10236);
and U15570 (N_15570,N_7458,N_6325);
nand U15571 (N_15571,N_11622,N_6595);
nor U15572 (N_15572,N_9883,N_9536);
nand U15573 (N_15573,N_11987,N_12124);
or U15574 (N_15574,N_10111,N_11395);
or U15575 (N_15575,N_11646,N_11317);
nor U15576 (N_15576,N_9590,N_7106);
or U15577 (N_15577,N_8271,N_8738);
nor U15578 (N_15578,N_6522,N_12195);
nand U15579 (N_15579,N_7705,N_8973);
xnor U15580 (N_15580,N_11394,N_8967);
or U15581 (N_15581,N_12330,N_12300);
nand U15582 (N_15582,N_6487,N_6340);
xnor U15583 (N_15583,N_6533,N_7730);
nor U15584 (N_15584,N_8086,N_11542);
or U15585 (N_15585,N_10203,N_11830);
xnor U15586 (N_15586,N_11279,N_6601);
nor U15587 (N_15587,N_9933,N_12113);
and U15588 (N_15588,N_11718,N_9781);
and U15589 (N_15589,N_9485,N_8354);
xnor U15590 (N_15590,N_9410,N_8325);
xnor U15591 (N_15591,N_10819,N_6742);
or U15592 (N_15592,N_10225,N_9554);
nor U15593 (N_15593,N_8432,N_9135);
xnor U15594 (N_15594,N_7858,N_6513);
xor U15595 (N_15595,N_9078,N_11490);
nor U15596 (N_15596,N_10002,N_9329);
nand U15597 (N_15597,N_9434,N_11228);
or U15598 (N_15598,N_7890,N_7310);
nor U15599 (N_15599,N_12118,N_10564);
nor U15600 (N_15600,N_8202,N_7247);
and U15601 (N_15601,N_9494,N_10721);
nand U15602 (N_15602,N_7961,N_9432);
xnor U15603 (N_15603,N_10568,N_11961);
xnor U15604 (N_15604,N_10367,N_6870);
nand U15605 (N_15605,N_7646,N_7391);
nand U15606 (N_15606,N_7496,N_7372);
and U15607 (N_15607,N_6996,N_8473);
nor U15608 (N_15608,N_10126,N_7185);
and U15609 (N_15609,N_10826,N_8650);
nand U15610 (N_15610,N_7904,N_6426);
nor U15611 (N_15611,N_9996,N_11128);
xnor U15612 (N_15612,N_11466,N_9015);
or U15613 (N_15613,N_9764,N_10277);
nor U15614 (N_15614,N_10430,N_9931);
or U15615 (N_15615,N_8427,N_7783);
nor U15616 (N_15616,N_10072,N_11352);
nor U15617 (N_15617,N_7013,N_9268);
nand U15618 (N_15618,N_6435,N_10549);
xor U15619 (N_15619,N_11431,N_6906);
and U15620 (N_15620,N_11632,N_11719);
nand U15621 (N_15621,N_12027,N_6353);
and U15622 (N_15622,N_8503,N_9530);
or U15623 (N_15623,N_10609,N_7026);
nand U15624 (N_15624,N_9869,N_7166);
nand U15625 (N_15625,N_6916,N_12075);
xor U15626 (N_15626,N_6387,N_10863);
or U15627 (N_15627,N_11180,N_10624);
nand U15628 (N_15628,N_9069,N_6269);
or U15629 (N_15629,N_10856,N_12177);
xnor U15630 (N_15630,N_11522,N_8475);
nand U15631 (N_15631,N_11198,N_8189);
nor U15632 (N_15632,N_11458,N_8374);
and U15633 (N_15633,N_8406,N_11248);
xnor U15634 (N_15634,N_7138,N_7712);
xnor U15635 (N_15635,N_11311,N_6938);
xor U15636 (N_15636,N_7789,N_7938);
xnor U15637 (N_15637,N_10168,N_6625);
nor U15638 (N_15638,N_6911,N_11523);
and U15639 (N_15639,N_6819,N_10152);
or U15640 (N_15640,N_12194,N_6731);
nor U15641 (N_15641,N_8658,N_11032);
nand U15642 (N_15642,N_6561,N_8468);
xnor U15643 (N_15643,N_8861,N_12083);
or U15644 (N_15644,N_8428,N_12263);
and U15645 (N_15645,N_8280,N_8222);
nand U15646 (N_15646,N_7477,N_10137);
xnor U15647 (N_15647,N_10004,N_11677);
or U15648 (N_15648,N_8239,N_8706);
xor U15649 (N_15649,N_12263,N_9600);
nor U15650 (N_15650,N_9911,N_11913);
nand U15651 (N_15651,N_7873,N_10059);
nor U15652 (N_15652,N_11493,N_7488);
xor U15653 (N_15653,N_9093,N_9761);
xnor U15654 (N_15654,N_11171,N_11186);
nand U15655 (N_15655,N_11193,N_10570);
xnor U15656 (N_15656,N_6482,N_11910);
and U15657 (N_15657,N_11039,N_10251);
nand U15658 (N_15658,N_9780,N_6981);
nor U15659 (N_15659,N_12162,N_7466);
and U15660 (N_15660,N_12108,N_10071);
xor U15661 (N_15661,N_7872,N_11611);
nor U15662 (N_15662,N_6347,N_8811);
and U15663 (N_15663,N_6284,N_10719);
xnor U15664 (N_15664,N_9250,N_6656);
or U15665 (N_15665,N_11892,N_9000);
xor U15666 (N_15666,N_11244,N_7806);
nor U15667 (N_15667,N_11631,N_9340);
nand U15668 (N_15668,N_6317,N_9475);
and U15669 (N_15669,N_10100,N_6515);
and U15670 (N_15670,N_8360,N_9398);
nor U15671 (N_15671,N_7769,N_9801);
or U15672 (N_15672,N_7153,N_11123);
and U15673 (N_15673,N_10148,N_8841);
nand U15674 (N_15674,N_7341,N_6945);
or U15675 (N_15675,N_9055,N_11830);
nand U15676 (N_15676,N_8230,N_6625);
and U15677 (N_15677,N_10024,N_10741);
nor U15678 (N_15678,N_10078,N_8432);
nor U15679 (N_15679,N_11819,N_8729);
nand U15680 (N_15680,N_8281,N_10401);
nand U15681 (N_15681,N_9238,N_12049);
or U15682 (N_15682,N_8164,N_11151);
and U15683 (N_15683,N_11106,N_7672);
or U15684 (N_15684,N_11629,N_10832);
or U15685 (N_15685,N_8408,N_12163);
or U15686 (N_15686,N_6488,N_6647);
nor U15687 (N_15687,N_7078,N_10402);
or U15688 (N_15688,N_7700,N_11426);
or U15689 (N_15689,N_8746,N_11480);
nor U15690 (N_15690,N_6586,N_6967);
nor U15691 (N_15691,N_12271,N_9993);
nand U15692 (N_15692,N_6975,N_12191);
nor U15693 (N_15693,N_9252,N_9643);
or U15694 (N_15694,N_7410,N_9311);
xnor U15695 (N_15695,N_12197,N_7820);
nor U15696 (N_15696,N_7343,N_11123);
xnor U15697 (N_15697,N_7004,N_10181);
xnor U15698 (N_15698,N_7877,N_10182);
and U15699 (N_15699,N_8923,N_7388);
or U15700 (N_15700,N_9988,N_7213);
nand U15701 (N_15701,N_6815,N_9073);
nor U15702 (N_15702,N_7692,N_12340);
or U15703 (N_15703,N_9074,N_9386);
xnor U15704 (N_15704,N_6919,N_7835);
and U15705 (N_15705,N_7589,N_6866);
or U15706 (N_15706,N_11976,N_7974);
and U15707 (N_15707,N_7279,N_11051);
and U15708 (N_15708,N_8741,N_10610);
nand U15709 (N_15709,N_8662,N_10046);
and U15710 (N_15710,N_7270,N_7658);
or U15711 (N_15711,N_10360,N_12287);
xnor U15712 (N_15712,N_7046,N_9146);
nor U15713 (N_15713,N_8801,N_7485);
nand U15714 (N_15714,N_10680,N_11561);
nor U15715 (N_15715,N_11436,N_9606);
nor U15716 (N_15716,N_10236,N_7875);
or U15717 (N_15717,N_9033,N_10352);
or U15718 (N_15718,N_9275,N_11368);
and U15719 (N_15719,N_10460,N_11630);
nand U15720 (N_15720,N_9752,N_12422);
nor U15721 (N_15721,N_6582,N_11718);
or U15722 (N_15722,N_11890,N_10611);
nor U15723 (N_15723,N_6435,N_6845);
xor U15724 (N_15724,N_10471,N_9499);
nand U15725 (N_15725,N_8994,N_8687);
and U15726 (N_15726,N_10345,N_7202);
xnor U15727 (N_15727,N_12431,N_7878);
nand U15728 (N_15728,N_8015,N_12286);
xnor U15729 (N_15729,N_8994,N_12287);
or U15730 (N_15730,N_7749,N_7360);
or U15731 (N_15731,N_8301,N_9395);
and U15732 (N_15732,N_6365,N_9499);
and U15733 (N_15733,N_6620,N_11793);
xor U15734 (N_15734,N_11847,N_9047);
or U15735 (N_15735,N_9025,N_11402);
or U15736 (N_15736,N_7922,N_6359);
nor U15737 (N_15737,N_7900,N_8322);
nand U15738 (N_15738,N_8670,N_7059);
nand U15739 (N_15739,N_8618,N_9377);
and U15740 (N_15740,N_11726,N_9157);
and U15741 (N_15741,N_7052,N_8572);
nor U15742 (N_15742,N_6519,N_8080);
nor U15743 (N_15743,N_7911,N_8646);
nor U15744 (N_15744,N_7166,N_11232);
and U15745 (N_15745,N_9169,N_8875);
nand U15746 (N_15746,N_9229,N_11399);
nor U15747 (N_15747,N_10272,N_12076);
xor U15748 (N_15748,N_11948,N_10421);
nor U15749 (N_15749,N_11653,N_12198);
or U15750 (N_15750,N_10571,N_6959);
nor U15751 (N_15751,N_9845,N_11005);
nand U15752 (N_15752,N_9914,N_10075);
and U15753 (N_15753,N_12243,N_11969);
nor U15754 (N_15754,N_7992,N_8345);
and U15755 (N_15755,N_7144,N_10137);
nor U15756 (N_15756,N_8143,N_10912);
and U15757 (N_15757,N_11937,N_7893);
nand U15758 (N_15758,N_8967,N_7864);
and U15759 (N_15759,N_11028,N_6718);
or U15760 (N_15760,N_9938,N_10493);
nor U15761 (N_15761,N_10273,N_8045);
nor U15762 (N_15762,N_10479,N_7941);
nor U15763 (N_15763,N_9488,N_6900);
nor U15764 (N_15764,N_11861,N_7605);
nand U15765 (N_15765,N_10101,N_9778);
xnor U15766 (N_15766,N_8423,N_8888);
nor U15767 (N_15767,N_11391,N_8434);
nor U15768 (N_15768,N_7942,N_8774);
or U15769 (N_15769,N_11643,N_12268);
nor U15770 (N_15770,N_9422,N_6808);
nand U15771 (N_15771,N_11284,N_12389);
or U15772 (N_15772,N_11701,N_11572);
or U15773 (N_15773,N_8732,N_7894);
or U15774 (N_15774,N_9497,N_9005);
nor U15775 (N_15775,N_12116,N_7644);
nand U15776 (N_15776,N_9466,N_7764);
nor U15777 (N_15777,N_7923,N_11563);
or U15778 (N_15778,N_9902,N_7576);
and U15779 (N_15779,N_10586,N_10462);
xnor U15780 (N_15780,N_11585,N_9180);
xnor U15781 (N_15781,N_6818,N_10613);
or U15782 (N_15782,N_8388,N_11081);
nand U15783 (N_15783,N_8880,N_6628);
nor U15784 (N_15784,N_8359,N_9132);
and U15785 (N_15785,N_6537,N_6629);
nand U15786 (N_15786,N_12134,N_9673);
xnor U15787 (N_15787,N_6253,N_7354);
or U15788 (N_15788,N_6294,N_10941);
and U15789 (N_15789,N_7987,N_8222);
or U15790 (N_15790,N_6974,N_8457);
nand U15791 (N_15791,N_9624,N_10038);
nor U15792 (N_15792,N_7504,N_9721);
and U15793 (N_15793,N_6797,N_7302);
and U15794 (N_15794,N_7750,N_7241);
or U15795 (N_15795,N_6340,N_12078);
and U15796 (N_15796,N_12492,N_9412);
xnor U15797 (N_15797,N_8379,N_9884);
or U15798 (N_15798,N_6671,N_8121);
nor U15799 (N_15799,N_7860,N_8763);
nand U15800 (N_15800,N_12312,N_12473);
or U15801 (N_15801,N_12080,N_10130);
nand U15802 (N_15802,N_9856,N_8804);
nor U15803 (N_15803,N_10636,N_8717);
xor U15804 (N_15804,N_10998,N_7202);
nand U15805 (N_15805,N_6839,N_9541);
nand U15806 (N_15806,N_9380,N_9293);
xor U15807 (N_15807,N_7896,N_7646);
xor U15808 (N_15808,N_7929,N_10212);
nand U15809 (N_15809,N_8264,N_7065);
xnor U15810 (N_15810,N_7191,N_6480);
or U15811 (N_15811,N_7549,N_11712);
nand U15812 (N_15812,N_7159,N_8942);
nor U15813 (N_15813,N_11930,N_11482);
nand U15814 (N_15814,N_7332,N_10096);
and U15815 (N_15815,N_7495,N_9934);
xnor U15816 (N_15816,N_10262,N_11515);
and U15817 (N_15817,N_12158,N_11635);
nand U15818 (N_15818,N_7296,N_6627);
or U15819 (N_15819,N_8619,N_10692);
xor U15820 (N_15820,N_10590,N_11793);
or U15821 (N_15821,N_9058,N_12349);
nand U15822 (N_15822,N_12194,N_11771);
and U15823 (N_15823,N_12049,N_8709);
or U15824 (N_15824,N_8279,N_10407);
nand U15825 (N_15825,N_10103,N_7226);
and U15826 (N_15826,N_7811,N_6997);
nor U15827 (N_15827,N_12359,N_6979);
xnor U15828 (N_15828,N_10760,N_10327);
or U15829 (N_15829,N_9541,N_10204);
nand U15830 (N_15830,N_8531,N_7166);
nand U15831 (N_15831,N_7238,N_7507);
xnor U15832 (N_15832,N_10029,N_10350);
nand U15833 (N_15833,N_8272,N_11495);
nor U15834 (N_15834,N_8047,N_9811);
nor U15835 (N_15835,N_8470,N_8593);
and U15836 (N_15836,N_8567,N_11842);
nor U15837 (N_15837,N_9534,N_7676);
nor U15838 (N_15838,N_11630,N_8932);
nor U15839 (N_15839,N_10626,N_11295);
nand U15840 (N_15840,N_6511,N_7959);
and U15841 (N_15841,N_6927,N_11098);
and U15842 (N_15842,N_9764,N_9488);
or U15843 (N_15843,N_10166,N_11815);
and U15844 (N_15844,N_9231,N_11628);
and U15845 (N_15845,N_6319,N_11614);
xor U15846 (N_15846,N_6568,N_11272);
or U15847 (N_15847,N_10916,N_6995);
and U15848 (N_15848,N_12137,N_9083);
and U15849 (N_15849,N_9602,N_9911);
and U15850 (N_15850,N_6280,N_9709);
nor U15851 (N_15851,N_11888,N_11834);
nor U15852 (N_15852,N_8906,N_11533);
and U15853 (N_15853,N_12113,N_7973);
nor U15854 (N_15854,N_7054,N_10939);
and U15855 (N_15855,N_11388,N_6355);
and U15856 (N_15856,N_8574,N_7774);
nor U15857 (N_15857,N_10548,N_7054);
xnor U15858 (N_15858,N_8150,N_11033);
xor U15859 (N_15859,N_12401,N_11315);
or U15860 (N_15860,N_7774,N_10689);
nand U15861 (N_15861,N_8357,N_7194);
or U15862 (N_15862,N_9032,N_8713);
or U15863 (N_15863,N_7233,N_7354);
nand U15864 (N_15864,N_11457,N_7843);
nand U15865 (N_15865,N_6960,N_10224);
and U15866 (N_15866,N_6285,N_10612);
nand U15867 (N_15867,N_6285,N_12306);
nand U15868 (N_15868,N_8189,N_6980);
nor U15869 (N_15869,N_7733,N_8849);
nor U15870 (N_15870,N_10928,N_9084);
or U15871 (N_15871,N_9397,N_6512);
or U15872 (N_15872,N_8104,N_9623);
or U15873 (N_15873,N_11402,N_8643);
and U15874 (N_15874,N_10791,N_10940);
nor U15875 (N_15875,N_10399,N_11966);
nor U15876 (N_15876,N_8038,N_12344);
nor U15877 (N_15877,N_10163,N_9095);
xnor U15878 (N_15878,N_9913,N_7652);
or U15879 (N_15879,N_7692,N_8703);
xor U15880 (N_15880,N_6473,N_9292);
and U15881 (N_15881,N_11639,N_11566);
nor U15882 (N_15882,N_6598,N_8440);
xnor U15883 (N_15883,N_8972,N_6689);
or U15884 (N_15884,N_11463,N_11163);
and U15885 (N_15885,N_8394,N_10824);
and U15886 (N_15886,N_12018,N_11609);
or U15887 (N_15887,N_8082,N_7621);
xnor U15888 (N_15888,N_12068,N_12414);
or U15889 (N_15889,N_6478,N_6941);
and U15890 (N_15890,N_10874,N_10659);
nand U15891 (N_15891,N_10189,N_9382);
or U15892 (N_15892,N_12022,N_7078);
nand U15893 (N_15893,N_9005,N_7681);
xor U15894 (N_15894,N_11453,N_11708);
nand U15895 (N_15895,N_7982,N_8858);
nand U15896 (N_15896,N_6560,N_9099);
xnor U15897 (N_15897,N_7469,N_8244);
nor U15898 (N_15898,N_8959,N_9438);
nor U15899 (N_15899,N_7279,N_11483);
nand U15900 (N_15900,N_10374,N_7601);
xnor U15901 (N_15901,N_6650,N_12429);
xor U15902 (N_15902,N_11405,N_11411);
xor U15903 (N_15903,N_7812,N_7349);
nor U15904 (N_15904,N_11652,N_9672);
or U15905 (N_15905,N_7431,N_9991);
nor U15906 (N_15906,N_7376,N_11945);
xor U15907 (N_15907,N_7735,N_9097);
nand U15908 (N_15908,N_6917,N_10595);
nand U15909 (N_15909,N_8465,N_12097);
xor U15910 (N_15910,N_9456,N_7439);
nor U15911 (N_15911,N_7525,N_6886);
or U15912 (N_15912,N_10577,N_6562);
nand U15913 (N_15913,N_10123,N_8192);
nor U15914 (N_15914,N_11056,N_9652);
nor U15915 (N_15915,N_11858,N_8680);
nor U15916 (N_15916,N_10886,N_8999);
and U15917 (N_15917,N_9847,N_8311);
or U15918 (N_15918,N_8061,N_7374);
nand U15919 (N_15919,N_10795,N_7965);
nand U15920 (N_15920,N_10521,N_12291);
nor U15921 (N_15921,N_12353,N_11953);
nor U15922 (N_15922,N_8379,N_8682);
and U15923 (N_15923,N_12432,N_7447);
and U15924 (N_15924,N_10169,N_11679);
xor U15925 (N_15925,N_6312,N_11556);
or U15926 (N_15926,N_9219,N_9337);
or U15927 (N_15927,N_11579,N_8284);
nand U15928 (N_15928,N_8707,N_11622);
or U15929 (N_15929,N_9963,N_10609);
nand U15930 (N_15930,N_6322,N_9062);
nand U15931 (N_15931,N_10687,N_11746);
xor U15932 (N_15932,N_12166,N_10175);
nor U15933 (N_15933,N_11917,N_10394);
or U15934 (N_15934,N_6290,N_10729);
and U15935 (N_15935,N_12130,N_7693);
nand U15936 (N_15936,N_8747,N_10367);
or U15937 (N_15937,N_9328,N_9709);
nand U15938 (N_15938,N_12359,N_10224);
and U15939 (N_15939,N_8216,N_12311);
or U15940 (N_15940,N_7022,N_12098);
or U15941 (N_15941,N_10929,N_12240);
xnor U15942 (N_15942,N_7429,N_11133);
nor U15943 (N_15943,N_9849,N_7449);
and U15944 (N_15944,N_7215,N_10415);
xor U15945 (N_15945,N_6940,N_9783);
xor U15946 (N_15946,N_6463,N_6995);
and U15947 (N_15947,N_9654,N_9128);
and U15948 (N_15948,N_10723,N_9389);
nor U15949 (N_15949,N_11944,N_8361);
nor U15950 (N_15950,N_10634,N_11799);
nor U15951 (N_15951,N_8466,N_7664);
and U15952 (N_15952,N_7663,N_6449);
nor U15953 (N_15953,N_7134,N_7634);
xnor U15954 (N_15954,N_8725,N_12394);
or U15955 (N_15955,N_10218,N_11817);
nor U15956 (N_15956,N_10928,N_9143);
and U15957 (N_15957,N_7451,N_6639);
nand U15958 (N_15958,N_7848,N_11717);
or U15959 (N_15959,N_8865,N_8340);
nand U15960 (N_15960,N_9563,N_7217);
xor U15961 (N_15961,N_7654,N_7199);
xnor U15962 (N_15962,N_6311,N_9597);
xnor U15963 (N_15963,N_6423,N_8540);
xnor U15964 (N_15964,N_7561,N_9593);
nor U15965 (N_15965,N_9229,N_10379);
nand U15966 (N_15966,N_7100,N_7157);
and U15967 (N_15967,N_6808,N_7810);
nor U15968 (N_15968,N_11000,N_10976);
xnor U15969 (N_15969,N_11429,N_10572);
xnor U15970 (N_15970,N_7758,N_8154);
xnor U15971 (N_15971,N_9251,N_8576);
nor U15972 (N_15972,N_8888,N_7931);
and U15973 (N_15973,N_9231,N_6459);
xnor U15974 (N_15974,N_6305,N_11958);
nand U15975 (N_15975,N_9929,N_10288);
nand U15976 (N_15976,N_10174,N_12302);
xnor U15977 (N_15977,N_8945,N_9839);
xnor U15978 (N_15978,N_9372,N_9423);
xor U15979 (N_15979,N_11645,N_7961);
and U15980 (N_15980,N_8179,N_11710);
nand U15981 (N_15981,N_8580,N_11404);
xor U15982 (N_15982,N_9880,N_11365);
xnor U15983 (N_15983,N_8412,N_10012);
xor U15984 (N_15984,N_11483,N_6502);
nand U15985 (N_15985,N_10252,N_10619);
nor U15986 (N_15986,N_8844,N_8417);
nand U15987 (N_15987,N_8857,N_9496);
or U15988 (N_15988,N_6382,N_10197);
xnor U15989 (N_15989,N_7231,N_12489);
or U15990 (N_15990,N_10784,N_6303);
xnor U15991 (N_15991,N_11748,N_8962);
or U15992 (N_15992,N_10708,N_11474);
and U15993 (N_15993,N_8977,N_9033);
or U15994 (N_15994,N_7234,N_10806);
nand U15995 (N_15995,N_6532,N_9468);
and U15996 (N_15996,N_11100,N_10742);
or U15997 (N_15997,N_8337,N_8326);
nor U15998 (N_15998,N_11120,N_11224);
xnor U15999 (N_15999,N_8409,N_7319);
or U16000 (N_16000,N_10852,N_10985);
xor U16001 (N_16001,N_11988,N_8088);
nor U16002 (N_16002,N_10613,N_11246);
and U16003 (N_16003,N_10463,N_10549);
or U16004 (N_16004,N_10325,N_9012);
and U16005 (N_16005,N_11485,N_7103);
or U16006 (N_16006,N_8034,N_9821);
xnor U16007 (N_16007,N_8205,N_11987);
nand U16008 (N_16008,N_7822,N_9259);
and U16009 (N_16009,N_6463,N_11605);
or U16010 (N_16010,N_7328,N_12388);
nor U16011 (N_16011,N_12192,N_12207);
nand U16012 (N_16012,N_11374,N_8979);
nand U16013 (N_16013,N_9611,N_11718);
or U16014 (N_16014,N_6742,N_6813);
nand U16015 (N_16015,N_10642,N_6578);
and U16016 (N_16016,N_11349,N_11627);
nor U16017 (N_16017,N_9102,N_10457);
xor U16018 (N_16018,N_11808,N_7164);
nor U16019 (N_16019,N_12012,N_6421);
xor U16020 (N_16020,N_11478,N_11898);
nor U16021 (N_16021,N_7562,N_6565);
and U16022 (N_16022,N_9434,N_7592);
nand U16023 (N_16023,N_9748,N_11408);
nor U16024 (N_16024,N_7113,N_11788);
or U16025 (N_16025,N_8835,N_8191);
and U16026 (N_16026,N_8229,N_6543);
nor U16027 (N_16027,N_11420,N_8492);
and U16028 (N_16028,N_7300,N_11447);
nor U16029 (N_16029,N_7486,N_6606);
and U16030 (N_16030,N_11781,N_10684);
xor U16031 (N_16031,N_10968,N_8734);
and U16032 (N_16032,N_8142,N_11403);
and U16033 (N_16033,N_9587,N_9838);
and U16034 (N_16034,N_10163,N_11184);
nor U16035 (N_16035,N_8580,N_7304);
and U16036 (N_16036,N_9933,N_7663);
nor U16037 (N_16037,N_10276,N_11627);
and U16038 (N_16038,N_9654,N_7598);
and U16039 (N_16039,N_9766,N_8004);
nor U16040 (N_16040,N_8872,N_11426);
nand U16041 (N_16041,N_10998,N_6338);
and U16042 (N_16042,N_7750,N_10085);
or U16043 (N_16043,N_7500,N_8315);
xnor U16044 (N_16044,N_9487,N_8113);
nand U16045 (N_16045,N_6295,N_6753);
and U16046 (N_16046,N_7814,N_7702);
or U16047 (N_16047,N_9401,N_7187);
xor U16048 (N_16048,N_9324,N_8609);
nand U16049 (N_16049,N_7426,N_8802);
nand U16050 (N_16050,N_9177,N_6832);
nor U16051 (N_16051,N_7993,N_9648);
nor U16052 (N_16052,N_6534,N_7118);
xnor U16053 (N_16053,N_11004,N_8183);
xor U16054 (N_16054,N_9139,N_8532);
nor U16055 (N_16055,N_6648,N_7537);
nor U16056 (N_16056,N_11584,N_10569);
nor U16057 (N_16057,N_8706,N_7041);
and U16058 (N_16058,N_9531,N_9162);
nand U16059 (N_16059,N_9934,N_11930);
xor U16060 (N_16060,N_11768,N_6886);
xnor U16061 (N_16061,N_7703,N_8337);
nor U16062 (N_16062,N_6454,N_9959);
and U16063 (N_16063,N_6974,N_6602);
nor U16064 (N_16064,N_6593,N_6335);
xnor U16065 (N_16065,N_10898,N_12359);
nand U16066 (N_16066,N_8317,N_8082);
nand U16067 (N_16067,N_11787,N_8464);
nand U16068 (N_16068,N_11690,N_7227);
nor U16069 (N_16069,N_8468,N_9122);
xor U16070 (N_16070,N_10518,N_6313);
or U16071 (N_16071,N_8321,N_9495);
xor U16072 (N_16072,N_9891,N_11589);
and U16073 (N_16073,N_9498,N_11669);
and U16074 (N_16074,N_11444,N_9193);
xnor U16075 (N_16075,N_10099,N_10059);
nand U16076 (N_16076,N_6429,N_7225);
or U16077 (N_16077,N_12126,N_10988);
nand U16078 (N_16078,N_7582,N_9893);
nor U16079 (N_16079,N_9605,N_8829);
or U16080 (N_16080,N_9816,N_6805);
nor U16081 (N_16081,N_11746,N_10406);
or U16082 (N_16082,N_8972,N_8870);
xnor U16083 (N_16083,N_8116,N_7202);
nor U16084 (N_16084,N_9690,N_10477);
or U16085 (N_16085,N_12463,N_12249);
nand U16086 (N_16086,N_7091,N_10298);
nor U16087 (N_16087,N_11904,N_11616);
nor U16088 (N_16088,N_6466,N_6916);
or U16089 (N_16089,N_6788,N_6908);
nand U16090 (N_16090,N_10231,N_7713);
xnor U16091 (N_16091,N_12282,N_10665);
and U16092 (N_16092,N_10613,N_11585);
nand U16093 (N_16093,N_12349,N_6645);
xor U16094 (N_16094,N_9223,N_11394);
and U16095 (N_16095,N_12484,N_10911);
or U16096 (N_16096,N_12182,N_12319);
or U16097 (N_16097,N_6299,N_7880);
xnor U16098 (N_16098,N_7150,N_7128);
and U16099 (N_16099,N_11033,N_8535);
or U16100 (N_16100,N_12181,N_6448);
xor U16101 (N_16101,N_7884,N_6799);
nand U16102 (N_16102,N_6699,N_12062);
nor U16103 (N_16103,N_9670,N_7383);
xnor U16104 (N_16104,N_8441,N_7424);
nor U16105 (N_16105,N_6319,N_12456);
xnor U16106 (N_16106,N_11699,N_8372);
or U16107 (N_16107,N_7015,N_8315);
nand U16108 (N_16108,N_11919,N_6379);
or U16109 (N_16109,N_6891,N_7155);
and U16110 (N_16110,N_6817,N_8157);
xnor U16111 (N_16111,N_10351,N_8923);
nor U16112 (N_16112,N_10206,N_11695);
or U16113 (N_16113,N_11574,N_6604);
and U16114 (N_16114,N_12391,N_9109);
xor U16115 (N_16115,N_10435,N_9404);
nor U16116 (N_16116,N_12340,N_9091);
and U16117 (N_16117,N_7482,N_6755);
or U16118 (N_16118,N_7499,N_9099);
nand U16119 (N_16119,N_12367,N_10442);
or U16120 (N_16120,N_6501,N_11784);
or U16121 (N_16121,N_9522,N_7571);
xnor U16122 (N_16122,N_6356,N_10915);
xnor U16123 (N_16123,N_11359,N_7549);
nand U16124 (N_16124,N_6822,N_10861);
or U16125 (N_16125,N_11121,N_6819);
and U16126 (N_16126,N_8411,N_8849);
and U16127 (N_16127,N_11996,N_10769);
and U16128 (N_16128,N_9023,N_8598);
or U16129 (N_16129,N_9981,N_10313);
xnor U16130 (N_16130,N_11299,N_10955);
and U16131 (N_16131,N_8627,N_10153);
or U16132 (N_16132,N_10421,N_11650);
nand U16133 (N_16133,N_12224,N_7989);
and U16134 (N_16134,N_12435,N_8125);
or U16135 (N_16135,N_8093,N_8414);
xor U16136 (N_16136,N_11670,N_10668);
xor U16137 (N_16137,N_11279,N_8514);
xor U16138 (N_16138,N_8194,N_8680);
xor U16139 (N_16139,N_6964,N_11375);
nand U16140 (N_16140,N_12038,N_11829);
and U16141 (N_16141,N_8648,N_7416);
nand U16142 (N_16142,N_6829,N_9336);
or U16143 (N_16143,N_10777,N_8063);
nand U16144 (N_16144,N_7633,N_11740);
or U16145 (N_16145,N_7987,N_10834);
or U16146 (N_16146,N_7367,N_8324);
nor U16147 (N_16147,N_6517,N_9694);
xor U16148 (N_16148,N_11409,N_8035);
nand U16149 (N_16149,N_12073,N_9772);
nor U16150 (N_16150,N_8467,N_9802);
or U16151 (N_16151,N_9208,N_6911);
nor U16152 (N_16152,N_9950,N_9185);
nand U16153 (N_16153,N_8236,N_8049);
nand U16154 (N_16154,N_10787,N_8648);
nand U16155 (N_16155,N_11469,N_8995);
xor U16156 (N_16156,N_12190,N_7678);
xor U16157 (N_16157,N_6937,N_11677);
or U16158 (N_16158,N_7816,N_9521);
and U16159 (N_16159,N_9239,N_8025);
and U16160 (N_16160,N_7011,N_7475);
and U16161 (N_16161,N_6665,N_9477);
nand U16162 (N_16162,N_12346,N_11081);
xor U16163 (N_16163,N_8906,N_7817);
xnor U16164 (N_16164,N_7223,N_10355);
nor U16165 (N_16165,N_6703,N_9181);
and U16166 (N_16166,N_9802,N_9515);
or U16167 (N_16167,N_7031,N_12385);
nor U16168 (N_16168,N_8115,N_11777);
and U16169 (N_16169,N_11256,N_12219);
xor U16170 (N_16170,N_11761,N_8381);
xnor U16171 (N_16171,N_7763,N_10449);
nand U16172 (N_16172,N_12288,N_12346);
xnor U16173 (N_16173,N_8294,N_12123);
nor U16174 (N_16174,N_9543,N_9328);
nor U16175 (N_16175,N_8023,N_8537);
and U16176 (N_16176,N_9540,N_6870);
xnor U16177 (N_16177,N_12189,N_8113);
nor U16178 (N_16178,N_10714,N_7272);
or U16179 (N_16179,N_12368,N_10856);
nor U16180 (N_16180,N_9740,N_6861);
nor U16181 (N_16181,N_7573,N_7392);
nand U16182 (N_16182,N_7843,N_8270);
nor U16183 (N_16183,N_9022,N_7957);
or U16184 (N_16184,N_9090,N_6365);
xor U16185 (N_16185,N_10387,N_8427);
nand U16186 (N_16186,N_11630,N_9064);
or U16187 (N_16187,N_6687,N_12290);
or U16188 (N_16188,N_12286,N_9019);
nand U16189 (N_16189,N_11325,N_7447);
and U16190 (N_16190,N_11946,N_8416);
xnor U16191 (N_16191,N_12429,N_9183);
xnor U16192 (N_16192,N_11387,N_11497);
xor U16193 (N_16193,N_7835,N_8530);
or U16194 (N_16194,N_10453,N_10144);
or U16195 (N_16195,N_10518,N_6549);
xnor U16196 (N_16196,N_7614,N_8278);
and U16197 (N_16197,N_11147,N_10275);
and U16198 (N_16198,N_7281,N_9644);
xor U16199 (N_16199,N_9126,N_6712);
xor U16200 (N_16200,N_6758,N_8989);
and U16201 (N_16201,N_8119,N_9056);
nor U16202 (N_16202,N_12463,N_8041);
or U16203 (N_16203,N_11937,N_11368);
and U16204 (N_16204,N_8883,N_9343);
xnor U16205 (N_16205,N_6505,N_7656);
nor U16206 (N_16206,N_9422,N_6579);
nor U16207 (N_16207,N_7683,N_12040);
or U16208 (N_16208,N_10303,N_11434);
or U16209 (N_16209,N_8284,N_11181);
nor U16210 (N_16210,N_8831,N_7165);
xnor U16211 (N_16211,N_7677,N_9335);
nand U16212 (N_16212,N_7447,N_10313);
xnor U16213 (N_16213,N_6881,N_9223);
xor U16214 (N_16214,N_8644,N_8222);
xnor U16215 (N_16215,N_7509,N_7910);
nor U16216 (N_16216,N_12474,N_6622);
xor U16217 (N_16217,N_8127,N_8264);
nor U16218 (N_16218,N_8427,N_12492);
xor U16219 (N_16219,N_8229,N_9624);
xor U16220 (N_16220,N_8814,N_9808);
nand U16221 (N_16221,N_9107,N_11687);
nor U16222 (N_16222,N_10074,N_7441);
xnor U16223 (N_16223,N_8700,N_11599);
or U16224 (N_16224,N_11984,N_9505);
xor U16225 (N_16225,N_9965,N_10391);
or U16226 (N_16226,N_10720,N_7767);
nand U16227 (N_16227,N_12174,N_6673);
xnor U16228 (N_16228,N_8342,N_8339);
or U16229 (N_16229,N_7046,N_8325);
or U16230 (N_16230,N_6913,N_11734);
nand U16231 (N_16231,N_10201,N_6915);
nor U16232 (N_16232,N_9034,N_8069);
nand U16233 (N_16233,N_12051,N_11132);
xnor U16234 (N_16234,N_8849,N_11261);
nand U16235 (N_16235,N_11045,N_8737);
and U16236 (N_16236,N_11014,N_7816);
and U16237 (N_16237,N_7391,N_8392);
and U16238 (N_16238,N_10899,N_12444);
nor U16239 (N_16239,N_10668,N_7024);
nor U16240 (N_16240,N_8813,N_8886);
nand U16241 (N_16241,N_11632,N_10161);
and U16242 (N_16242,N_10605,N_7524);
xor U16243 (N_16243,N_10968,N_6823);
or U16244 (N_16244,N_8214,N_9171);
nand U16245 (N_16245,N_8132,N_8661);
nand U16246 (N_16246,N_11975,N_11678);
nand U16247 (N_16247,N_7822,N_12402);
xnor U16248 (N_16248,N_6385,N_8315);
xnor U16249 (N_16249,N_10452,N_6781);
and U16250 (N_16250,N_10605,N_8069);
nor U16251 (N_16251,N_10140,N_6328);
nand U16252 (N_16252,N_9241,N_8431);
or U16253 (N_16253,N_8072,N_11181);
nor U16254 (N_16254,N_9669,N_11913);
xnor U16255 (N_16255,N_8080,N_6830);
or U16256 (N_16256,N_6611,N_9447);
nor U16257 (N_16257,N_9160,N_12436);
nor U16258 (N_16258,N_12296,N_7574);
nand U16259 (N_16259,N_8812,N_11456);
xnor U16260 (N_16260,N_9751,N_9505);
nor U16261 (N_16261,N_12149,N_11677);
or U16262 (N_16262,N_10997,N_10043);
xnor U16263 (N_16263,N_9290,N_9020);
nand U16264 (N_16264,N_8148,N_9197);
and U16265 (N_16265,N_9760,N_8046);
and U16266 (N_16266,N_7420,N_10248);
and U16267 (N_16267,N_12072,N_10621);
xor U16268 (N_16268,N_10061,N_10492);
nand U16269 (N_16269,N_6955,N_10024);
and U16270 (N_16270,N_11192,N_11296);
or U16271 (N_16271,N_11591,N_8910);
xor U16272 (N_16272,N_12255,N_10377);
and U16273 (N_16273,N_7782,N_6356);
nor U16274 (N_16274,N_12473,N_10027);
or U16275 (N_16275,N_11173,N_6789);
nor U16276 (N_16276,N_11662,N_6749);
nor U16277 (N_16277,N_6841,N_7901);
and U16278 (N_16278,N_9346,N_8181);
nor U16279 (N_16279,N_9459,N_8992);
or U16280 (N_16280,N_7676,N_6572);
and U16281 (N_16281,N_11323,N_10534);
nand U16282 (N_16282,N_6609,N_12385);
nand U16283 (N_16283,N_9523,N_11007);
nand U16284 (N_16284,N_7510,N_7678);
nor U16285 (N_16285,N_10492,N_6492);
nand U16286 (N_16286,N_10601,N_8903);
and U16287 (N_16287,N_12277,N_10676);
xor U16288 (N_16288,N_10286,N_7867);
xnor U16289 (N_16289,N_11648,N_8948);
or U16290 (N_16290,N_8100,N_6953);
and U16291 (N_16291,N_9089,N_8217);
or U16292 (N_16292,N_10630,N_11063);
nor U16293 (N_16293,N_7676,N_7184);
xor U16294 (N_16294,N_7857,N_9395);
and U16295 (N_16295,N_10994,N_11097);
and U16296 (N_16296,N_9762,N_7888);
nor U16297 (N_16297,N_9560,N_7760);
or U16298 (N_16298,N_12187,N_7524);
xnor U16299 (N_16299,N_10141,N_12424);
and U16300 (N_16300,N_9192,N_11589);
xor U16301 (N_16301,N_10738,N_7089);
xnor U16302 (N_16302,N_6361,N_8082);
nor U16303 (N_16303,N_8956,N_7100);
nand U16304 (N_16304,N_10599,N_10071);
nand U16305 (N_16305,N_8738,N_9527);
and U16306 (N_16306,N_10448,N_9195);
nor U16307 (N_16307,N_10395,N_11817);
and U16308 (N_16308,N_11214,N_8701);
nand U16309 (N_16309,N_9014,N_7972);
nor U16310 (N_16310,N_11833,N_10429);
nor U16311 (N_16311,N_10846,N_7902);
nand U16312 (N_16312,N_8963,N_8833);
or U16313 (N_16313,N_8985,N_10267);
xor U16314 (N_16314,N_8764,N_10919);
xor U16315 (N_16315,N_11165,N_8261);
xor U16316 (N_16316,N_10978,N_11106);
nand U16317 (N_16317,N_10910,N_8139);
nor U16318 (N_16318,N_7547,N_8768);
nand U16319 (N_16319,N_12062,N_10476);
nor U16320 (N_16320,N_9423,N_6480);
xnor U16321 (N_16321,N_7893,N_10177);
nor U16322 (N_16322,N_8452,N_11694);
xor U16323 (N_16323,N_7333,N_8077);
or U16324 (N_16324,N_6430,N_8455);
nand U16325 (N_16325,N_9818,N_10109);
and U16326 (N_16326,N_10101,N_11763);
xor U16327 (N_16327,N_6730,N_11277);
nor U16328 (N_16328,N_12118,N_11859);
nand U16329 (N_16329,N_7194,N_11504);
or U16330 (N_16330,N_9353,N_10118);
and U16331 (N_16331,N_11564,N_6397);
xor U16332 (N_16332,N_6750,N_6945);
nor U16333 (N_16333,N_8086,N_6704);
xnor U16334 (N_16334,N_6876,N_12101);
xnor U16335 (N_16335,N_6644,N_9940);
or U16336 (N_16336,N_6756,N_8083);
or U16337 (N_16337,N_9489,N_12303);
nand U16338 (N_16338,N_8847,N_9531);
nor U16339 (N_16339,N_11806,N_8209);
or U16340 (N_16340,N_9056,N_10926);
nand U16341 (N_16341,N_11546,N_11085);
xor U16342 (N_16342,N_8198,N_7200);
or U16343 (N_16343,N_6258,N_12199);
and U16344 (N_16344,N_12495,N_8927);
nor U16345 (N_16345,N_9567,N_6727);
xnor U16346 (N_16346,N_9617,N_11369);
nand U16347 (N_16347,N_11362,N_10003);
xor U16348 (N_16348,N_11659,N_11864);
or U16349 (N_16349,N_11552,N_9158);
nand U16350 (N_16350,N_8314,N_8887);
nand U16351 (N_16351,N_7550,N_10798);
nor U16352 (N_16352,N_9206,N_11794);
nor U16353 (N_16353,N_7221,N_7449);
nand U16354 (N_16354,N_11650,N_11319);
and U16355 (N_16355,N_6673,N_11405);
nor U16356 (N_16356,N_12424,N_6502);
and U16357 (N_16357,N_7408,N_9324);
or U16358 (N_16358,N_8155,N_10036);
xor U16359 (N_16359,N_7173,N_12321);
xnor U16360 (N_16360,N_9207,N_8542);
xor U16361 (N_16361,N_9387,N_11123);
xor U16362 (N_16362,N_8351,N_12151);
and U16363 (N_16363,N_6705,N_8316);
nand U16364 (N_16364,N_7673,N_10969);
nor U16365 (N_16365,N_9008,N_8692);
nor U16366 (N_16366,N_10051,N_8093);
and U16367 (N_16367,N_9027,N_8304);
nand U16368 (N_16368,N_6941,N_8250);
and U16369 (N_16369,N_11587,N_9137);
or U16370 (N_16370,N_10490,N_7216);
and U16371 (N_16371,N_6490,N_10783);
nand U16372 (N_16372,N_10730,N_6524);
or U16373 (N_16373,N_7129,N_8605);
nor U16374 (N_16374,N_9511,N_7477);
xor U16375 (N_16375,N_12238,N_11770);
xor U16376 (N_16376,N_7078,N_10933);
nor U16377 (N_16377,N_7186,N_12312);
xnor U16378 (N_16378,N_11572,N_11135);
or U16379 (N_16379,N_10445,N_10246);
nand U16380 (N_16380,N_11231,N_10968);
nand U16381 (N_16381,N_8911,N_8936);
nand U16382 (N_16382,N_8742,N_7419);
xor U16383 (N_16383,N_8138,N_10592);
and U16384 (N_16384,N_7911,N_9750);
nor U16385 (N_16385,N_9730,N_7337);
nand U16386 (N_16386,N_12310,N_10246);
nand U16387 (N_16387,N_9910,N_10532);
or U16388 (N_16388,N_8542,N_9986);
or U16389 (N_16389,N_10931,N_12154);
xor U16390 (N_16390,N_10026,N_12039);
xnor U16391 (N_16391,N_12381,N_12376);
xnor U16392 (N_16392,N_7207,N_9916);
xor U16393 (N_16393,N_11874,N_7686);
nand U16394 (N_16394,N_9607,N_10131);
and U16395 (N_16395,N_11139,N_9282);
or U16396 (N_16396,N_9808,N_10853);
or U16397 (N_16397,N_11457,N_7720);
and U16398 (N_16398,N_8456,N_12310);
or U16399 (N_16399,N_9207,N_9365);
or U16400 (N_16400,N_6463,N_6883);
nor U16401 (N_16401,N_10850,N_9848);
nor U16402 (N_16402,N_10271,N_6896);
xor U16403 (N_16403,N_9530,N_6840);
or U16404 (N_16404,N_6397,N_6716);
xor U16405 (N_16405,N_9235,N_7002);
and U16406 (N_16406,N_10131,N_10353);
nand U16407 (N_16407,N_9953,N_11147);
nand U16408 (N_16408,N_10771,N_12163);
nand U16409 (N_16409,N_12343,N_12427);
and U16410 (N_16410,N_8919,N_9653);
xnor U16411 (N_16411,N_8053,N_8837);
nor U16412 (N_16412,N_8932,N_9674);
or U16413 (N_16413,N_6814,N_11379);
nand U16414 (N_16414,N_9941,N_8008);
xnor U16415 (N_16415,N_7580,N_11827);
and U16416 (N_16416,N_10584,N_6708);
nor U16417 (N_16417,N_9606,N_7602);
nor U16418 (N_16418,N_10019,N_10724);
or U16419 (N_16419,N_9237,N_7355);
xnor U16420 (N_16420,N_12225,N_7444);
or U16421 (N_16421,N_7675,N_7157);
nor U16422 (N_16422,N_9943,N_8688);
or U16423 (N_16423,N_9933,N_9371);
xor U16424 (N_16424,N_11848,N_6485);
nand U16425 (N_16425,N_7883,N_9171);
nor U16426 (N_16426,N_11999,N_7700);
or U16427 (N_16427,N_9254,N_7808);
nand U16428 (N_16428,N_7136,N_8462);
xor U16429 (N_16429,N_9240,N_9571);
xnor U16430 (N_16430,N_6946,N_9907);
or U16431 (N_16431,N_7593,N_7228);
or U16432 (N_16432,N_6660,N_10096);
or U16433 (N_16433,N_7402,N_8724);
nand U16434 (N_16434,N_8474,N_10716);
and U16435 (N_16435,N_11390,N_12038);
nor U16436 (N_16436,N_6319,N_8660);
nand U16437 (N_16437,N_6720,N_6280);
nor U16438 (N_16438,N_6255,N_10074);
and U16439 (N_16439,N_8796,N_12220);
xnor U16440 (N_16440,N_10353,N_6774);
nand U16441 (N_16441,N_6923,N_7181);
xor U16442 (N_16442,N_8913,N_11528);
xor U16443 (N_16443,N_7600,N_9732);
or U16444 (N_16444,N_10512,N_7346);
or U16445 (N_16445,N_12298,N_8431);
and U16446 (N_16446,N_10762,N_8949);
and U16447 (N_16447,N_7433,N_9465);
or U16448 (N_16448,N_8378,N_11012);
xnor U16449 (N_16449,N_9225,N_7607);
and U16450 (N_16450,N_8173,N_9062);
xor U16451 (N_16451,N_9495,N_10142);
nor U16452 (N_16452,N_7452,N_11810);
nand U16453 (N_16453,N_6411,N_6352);
nand U16454 (N_16454,N_11877,N_6457);
nand U16455 (N_16455,N_9467,N_11945);
or U16456 (N_16456,N_7169,N_8411);
nand U16457 (N_16457,N_10790,N_12384);
xnor U16458 (N_16458,N_12486,N_12137);
nor U16459 (N_16459,N_9201,N_6846);
nand U16460 (N_16460,N_6629,N_11190);
xnor U16461 (N_16461,N_11549,N_8621);
or U16462 (N_16462,N_8054,N_11504);
nand U16463 (N_16463,N_11534,N_9998);
nand U16464 (N_16464,N_9248,N_9101);
nor U16465 (N_16465,N_9564,N_10240);
xnor U16466 (N_16466,N_11302,N_11193);
nand U16467 (N_16467,N_12428,N_9163);
nand U16468 (N_16468,N_11647,N_10619);
xor U16469 (N_16469,N_12113,N_6919);
nor U16470 (N_16470,N_11472,N_8485);
xor U16471 (N_16471,N_8564,N_10551);
xnor U16472 (N_16472,N_6845,N_7639);
and U16473 (N_16473,N_8289,N_7883);
xnor U16474 (N_16474,N_9570,N_10052);
or U16475 (N_16475,N_11116,N_7756);
or U16476 (N_16476,N_9797,N_11985);
or U16477 (N_16477,N_10065,N_8431);
nor U16478 (N_16478,N_11427,N_8105);
nor U16479 (N_16479,N_10952,N_8261);
and U16480 (N_16480,N_9294,N_6865);
nand U16481 (N_16481,N_8180,N_7143);
nor U16482 (N_16482,N_8254,N_11881);
nor U16483 (N_16483,N_7174,N_8069);
nand U16484 (N_16484,N_11575,N_12293);
xnor U16485 (N_16485,N_9694,N_6556);
and U16486 (N_16486,N_6427,N_11635);
nor U16487 (N_16487,N_9341,N_8570);
and U16488 (N_16488,N_6920,N_7759);
xnor U16489 (N_16489,N_6690,N_9812);
or U16490 (N_16490,N_11909,N_6804);
nand U16491 (N_16491,N_6438,N_8755);
nor U16492 (N_16492,N_11767,N_9566);
or U16493 (N_16493,N_10343,N_6482);
and U16494 (N_16494,N_10457,N_7174);
nand U16495 (N_16495,N_6974,N_9873);
nand U16496 (N_16496,N_11191,N_12197);
nand U16497 (N_16497,N_9178,N_7191);
nor U16498 (N_16498,N_11137,N_9043);
nand U16499 (N_16499,N_7234,N_7134);
or U16500 (N_16500,N_6800,N_12369);
and U16501 (N_16501,N_6375,N_8212);
or U16502 (N_16502,N_10565,N_7190);
or U16503 (N_16503,N_8583,N_6758);
or U16504 (N_16504,N_9778,N_6616);
or U16505 (N_16505,N_9331,N_8088);
and U16506 (N_16506,N_10866,N_6845);
nor U16507 (N_16507,N_9273,N_12048);
nor U16508 (N_16508,N_6717,N_6718);
xnor U16509 (N_16509,N_9767,N_9841);
nor U16510 (N_16510,N_7492,N_7164);
xor U16511 (N_16511,N_7856,N_6777);
nand U16512 (N_16512,N_9862,N_9072);
xor U16513 (N_16513,N_10130,N_9610);
xor U16514 (N_16514,N_7838,N_12029);
or U16515 (N_16515,N_9758,N_8944);
nor U16516 (N_16516,N_9275,N_7326);
nor U16517 (N_16517,N_6461,N_10696);
nor U16518 (N_16518,N_6383,N_8322);
nor U16519 (N_16519,N_7248,N_10462);
or U16520 (N_16520,N_6630,N_10954);
or U16521 (N_16521,N_6684,N_9192);
nor U16522 (N_16522,N_6437,N_11797);
and U16523 (N_16523,N_8418,N_7810);
xor U16524 (N_16524,N_10180,N_11094);
nand U16525 (N_16525,N_11375,N_12483);
or U16526 (N_16526,N_11582,N_8244);
and U16527 (N_16527,N_11288,N_8589);
xnor U16528 (N_16528,N_8642,N_6811);
xor U16529 (N_16529,N_7411,N_8304);
and U16530 (N_16530,N_9635,N_8664);
nor U16531 (N_16531,N_12001,N_9051);
and U16532 (N_16532,N_11743,N_10435);
nor U16533 (N_16533,N_7115,N_6940);
and U16534 (N_16534,N_6941,N_6914);
and U16535 (N_16535,N_9744,N_10101);
nand U16536 (N_16536,N_12462,N_10185);
nand U16537 (N_16537,N_6835,N_11080);
nor U16538 (N_16538,N_10865,N_12150);
nor U16539 (N_16539,N_11908,N_6571);
nor U16540 (N_16540,N_11427,N_11248);
or U16541 (N_16541,N_8316,N_10543);
nand U16542 (N_16542,N_6683,N_6600);
or U16543 (N_16543,N_11086,N_7726);
or U16544 (N_16544,N_8958,N_6380);
and U16545 (N_16545,N_7704,N_9525);
nor U16546 (N_16546,N_8255,N_7172);
nand U16547 (N_16547,N_11970,N_11575);
nand U16548 (N_16548,N_9051,N_6721);
or U16549 (N_16549,N_6408,N_8673);
or U16550 (N_16550,N_7486,N_11313);
or U16551 (N_16551,N_11156,N_7301);
nand U16552 (N_16552,N_12189,N_8748);
xor U16553 (N_16553,N_9612,N_9257);
nand U16554 (N_16554,N_9614,N_9485);
nand U16555 (N_16555,N_9531,N_12334);
xnor U16556 (N_16556,N_10131,N_9091);
and U16557 (N_16557,N_7421,N_10068);
nand U16558 (N_16558,N_10610,N_7375);
or U16559 (N_16559,N_9877,N_8350);
nand U16560 (N_16560,N_9700,N_8065);
nor U16561 (N_16561,N_6953,N_11124);
nor U16562 (N_16562,N_10393,N_8952);
nor U16563 (N_16563,N_8155,N_10218);
nor U16564 (N_16564,N_10494,N_9401);
and U16565 (N_16565,N_11181,N_10838);
xor U16566 (N_16566,N_12443,N_11421);
and U16567 (N_16567,N_6947,N_8393);
xor U16568 (N_16568,N_8262,N_6604);
and U16569 (N_16569,N_7247,N_6310);
nand U16570 (N_16570,N_11638,N_9297);
or U16571 (N_16571,N_9002,N_9309);
and U16572 (N_16572,N_11678,N_11442);
nor U16573 (N_16573,N_6428,N_7804);
nand U16574 (N_16574,N_10595,N_10855);
nor U16575 (N_16575,N_10210,N_11824);
or U16576 (N_16576,N_7212,N_7296);
nand U16577 (N_16577,N_6958,N_9466);
nor U16578 (N_16578,N_12052,N_8378);
and U16579 (N_16579,N_10896,N_9464);
and U16580 (N_16580,N_6970,N_10039);
or U16581 (N_16581,N_6620,N_10424);
nor U16582 (N_16582,N_7134,N_8422);
xnor U16583 (N_16583,N_9603,N_6540);
and U16584 (N_16584,N_11420,N_10045);
xnor U16585 (N_16585,N_7546,N_7731);
nand U16586 (N_16586,N_11745,N_11041);
nand U16587 (N_16587,N_11749,N_9997);
nor U16588 (N_16588,N_6851,N_10192);
nor U16589 (N_16589,N_6424,N_10028);
and U16590 (N_16590,N_12050,N_7679);
nor U16591 (N_16591,N_10120,N_10967);
nor U16592 (N_16592,N_12181,N_7164);
xor U16593 (N_16593,N_9127,N_7243);
nor U16594 (N_16594,N_7569,N_11268);
nor U16595 (N_16595,N_7106,N_9034);
nor U16596 (N_16596,N_9856,N_9999);
xor U16597 (N_16597,N_9895,N_12477);
and U16598 (N_16598,N_12329,N_11631);
and U16599 (N_16599,N_7607,N_10990);
or U16600 (N_16600,N_9379,N_7896);
and U16601 (N_16601,N_12402,N_7858);
nor U16602 (N_16602,N_6740,N_8731);
or U16603 (N_16603,N_11106,N_11053);
and U16604 (N_16604,N_6416,N_9343);
nor U16605 (N_16605,N_11335,N_10353);
nor U16606 (N_16606,N_6516,N_11187);
nor U16607 (N_16607,N_10788,N_6696);
nor U16608 (N_16608,N_10622,N_6688);
xor U16609 (N_16609,N_9926,N_9664);
and U16610 (N_16610,N_11722,N_12052);
or U16611 (N_16611,N_11097,N_9779);
xnor U16612 (N_16612,N_9042,N_9332);
nor U16613 (N_16613,N_9433,N_11968);
xor U16614 (N_16614,N_8502,N_7145);
nor U16615 (N_16615,N_11285,N_8505);
nor U16616 (N_16616,N_8807,N_6679);
xor U16617 (N_16617,N_7616,N_9338);
or U16618 (N_16618,N_6841,N_10059);
nor U16619 (N_16619,N_8998,N_6517);
nand U16620 (N_16620,N_7793,N_6571);
or U16621 (N_16621,N_7963,N_9719);
nand U16622 (N_16622,N_8374,N_6847);
and U16623 (N_16623,N_10090,N_8408);
xor U16624 (N_16624,N_7566,N_11262);
nand U16625 (N_16625,N_9599,N_8889);
xnor U16626 (N_16626,N_6963,N_6593);
nor U16627 (N_16627,N_11754,N_7681);
nand U16628 (N_16628,N_9403,N_8623);
nand U16629 (N_16629,N_10051,N_6841);
nor U16630 (N_16630,N_10135,N_9206);
xnor U16631 (N_16631,N_12212,N_7921);
nor U16632 (N_16632,N_10027,N_7562);
xnor U16633 (N_16633,N_11877,N_7002);
xnor U16634 (N_16634,N_9441,N_10725);
nand U16635 (N_16635,N_10447,N_8919);
nor U16636 (N_16636,N_9702,N_7502);
nor U16637 (N_16637,N_9592,N_12026);
xor U16638 (N_16638,N_9320,N_12375);
xnor U16639 (N_16639,N_9282,N_8310);
and U16640 (N_16640,N_11679,N_8067);
or U16641 (N_16641,N_9316,N_10365);
xnor U16642 (N_16642,N_6618,N_8668);
and U16643 (N_16643,N_11956,N_7107);
nor U16644 (N_16644,N_6385,N_6636);
nor U16645 (N_16645,N_7689,N_8556);
and U16646 (N_16646,N_6676,N_9683);
xnor U16647 (N_16647,N_6589,N_7132);
and U16648 (N_16648,N_9736,N_9344);
nor U16649 (N_16649,N_8102,N_6660);
or U16650 (N_16650,N_6374,N_10000);
nor U16651 (N_16651,N_6752,N_7885);
or U16652 (N_16652,N_8046,N_6354);
and U16653 (N_16653,N_10206,N_12454);
or U16654 (N_16654,N_9989,N_6954);
nand U16655 (N_16655,N_6383,N_7675);
nand U16656 (N_16656,N_6916,N_6780);
xnor U16657 (N_16657,N_9790,N_7629);
nor U16658 (N_16658,N_7881,N_10272);
and U16659 (N_16659,N_9866,N_9470);
nor U16660 (N_16660,N_12345,N_6843);
and U16661 (N_16661,N_9519,N_9807);
nand U16662 (N_16662,N_11623,N_8450);
xnor U16663 (N_16663,N_6767,N_9428);
and U16664 (N_16664,N_7378,N_6416);
and U16665 (N_16665,N_12258,N_12077);
nor U16666 (N_16666,N_7760,N_8613);
nor U16667 (N_16667,N_11754,N_9929);
xnor U16668 (N_16668,N_7293,N_8361);
or U16669 (N_16669,N_7566,N_8865);
xor U16670 (N_16670,N_10052,N_7472);
nor U16671 (N_16671,N_6303,N_8568);
nor U16672 (N_16672,N_10109,N_7770);
nand U16673 (N_16673,N_8360,N_8289);
or U16674 (N_16674,N_9460,N_7125);
xor U16675 (N_16675,N_8461,N_7842);
and U16676 (N_16676,N_9458,N_8422);
or U16677 (N_16677,N_7588,N_8409);
nand U16678 (N_16678,N_11513,N_9180);
xor U16679 (N_16679,N_11495,N_11333);
and U16680 (N_16680,N_6393,N_9855);
and U16681 (N_16681,N_9468,N_12112);
and U16682 (N_16682,N_7083,N_11112);
and U16683 (N_16683,N_7911,N_7685);
or U16684 (N_16684,N_10444,N_7532);
nor U16685 (N_16685,N_12131,N_9826);
and U16686 (N_16686,N_9660,N_9749);
and U16687 (N_16687,N_9867,N_9476);
and U16688 (N_16688,N_10730,N_12196);
xor U16689 (N_16689,N_12250,N_7787);
nand U16690 (N_16690,N_10414,N_8592);
nand U16691 (N_16691,N_8606,N_6670);
and U16692 (N_16692,N_6877,N_7075);
nor U16693 (N_16693,N_8967,N_8470);
or U16694 (N_16694,N_6543,N_9813);
nor U16695 (N_16695,N_10087,N_8445);
nor U16696 (N_16696,N_10154,N_8389);
nand U16697 (N_16697,N_11999,N_10914);
nand U16698 (N_16698,N_6755,N_9281);
xor U16699 (N_16699,N_7766,N_6435);
nand U16700 (N_16700,N_6968,N_7645);
nand U16701 (N_16701,N_6303,N_10080);
or U16702 (N_16702,N_6650,N_7054);
or U16703 (N_16703,N_11112,N_8324);
and U16704 (N_16704,N_9287,N_9678);
nand U16705 (N_16705,N_8393,N_9478);
nor U16706 (N_16706,N_10665,N_9019);
or U16707 (N_16707,N_9321,N_9305);
or U16708 (N_16708,N_7298,N_9329);
or U16709 (N_16709,N_9653,N_12357);
xnor U16710 (N_16710,N_9432,N_6427);
and U16711 (N_16711,N_11041,N_6734);
xnor U16712 (N_16712,N_12228,N_9663);
xor U16713 (N_16713,N_9361,N_8339);
and U16714 (N_16714,N_9132,N_9845);
and U16715 (N_16715,N_8028,N_9041);
or U16716 (N_16716,N_9519,N_10128);
xor U16717 (N_16717,N_10235,N_8978);
xnor U16718 (N_16718,N_9348,N_12193);
nor U16719 (N_16719,N_6668,N_8656);
xnor U16720 (N_16720,N_9666,N_8578);
or U16721 (N_16721,N_12043,N_7529);
nand U16722 (N_16722,N_11406,N_11298);
or U16723 (N_16723,N_7606,N_12129);
and U16724 (N_16724,N_8451,N_9989);
and U16725 (N_16725,N_9732,N_8015);
nor U16726 (N_16726,N_8354,N_7361);
xnor U16727 (N_16727,N_10261,N_7828);
nand U16728 (N_16728,N_8942,N_8463);
xnor U16729 (N_16729,N_11135,N_10039);
and U16730 (N_16730,N_7335,N_10412);
nand U16731 (N_16731,N_9211,N_9192);
nand U16732 (N_16732,N_11006,N_10836);
xor U16733 (N_16733,N_11787,N_11768);
or U16734 (N_16734,N_8652,N_9014);
and U16735 (N_16735,N_11426,N_7476);
or U16736 (N_16736,N_7399,N_11442);
xor U16737 (N_16737,N_12416,N_9699);
nor U16738 (N_16738,N_7745,N_7515);
nand U16739 (N_16739,N_8312,N_11914);
and U16740 (N_16740,N_10155,N_7444);
and U16741 (N_16741,N_12277,N_8671);
or U16742 (N_16742,N_12304,N_12073);
or U16743 (N_16743,N_7884,N_7404);
nand U16744 (N_16744,N_11799,N_10245);
xnor U16745 (N_16745,N_12116,N_7723);
or U16746 (N_16746,N_11318,N_7412);
xnor U16747 (N_16747,N_8391,N_11957);
or U16748 (N_16748,N_8113,N_9484);
and U16749 (N_16749,N_10467,N_7797);
or U16750 (N_16750,N_7214,N_6972);
nand U16751 (N_16751,N_9689,N_6865);
nor U16752 (N_16752,N_11228,N_9605);
xor U16753 (N_16753,N_7221,N_11127);
and U16754 (N_16754,N_7514,N_12115);
and U16755 (N_16755,N_7444,N_7463);
nor U16756 (N_16756,N_8080,N_8648);
nand U16757 (N_16757,N_10741,N_11447);
nor U16758 (N_16758,N_10164,N_9625);
xor U16759 (N_16759,N_6278,N_9805);
or U16760 (N_16760,N_12439,N_9349);
xor U16761 (N_16761,N_8339,N_10789);
xnor U16762 (N_16762,N_11778,N_7444);
and U16763 (N_16763,N_10923,N_7428);
and U16764 (N_16764,N_6482,N_11117);
xnor U16765 (N_16765,N_6697,N_6337);
nand U16766 (N_16766,N_9245,N_6922);
or U16767 (N_16767,N_10276,N_7719);
or U16768 (N_16768,N_9291,N_10336);
xnor U16769 (N_16769,N_10163,N_9749);
xnor U16770 (N_16770,N_6492,N_11470);
nor U16771 (N_16771,N_9131,N_9180);
or U16772 (N_16772,N_9572,N_7193);
xnor U16773 (N_16773,N_9989,N_7583);
and U16774 (N_16774,N_8983,N_10824);
nand U16775 (N_16775,N_6686,N_6925);
and U16776 (N_16776,N_7053,N_10522);
nand U16777 (N_16777,N_6997,N_9227);
nor U16778 (N_16778,N_10788,N_7093);
or U16779 (N_16779,N_9333,N_11436);
nor U16780 (N_16780,N_6277,N_6738);
or U16781 (N_16781,N_10111,N_8443);
nor U16782 (N_16782,N_8599,N_8340);
and U16783 (N_16783,N_10482,N_9351);
or U16784 (N_16784,N_7301,N_11429);
nand U16785 (N_16785,N_9799,N_8866);
and U16786 (N_16786,N_8118,N_9512);
xor U16787 (N_16787,N_8564,N_6691);
nand U16788 (N_16788,N_6640,N_6984);
and U16789 (N_16789,N_7891,N_8800);
nand U16790 (N_16790,N_9224,N_12300);
nand U16791 (N_16791,N_9858,N_8283);
nor U16792 (N_16792,N_9871,N_6645);
or U16793 (N_16793,N_11242,N_11482);
nand U16794 (N_16794,N_8985,N_9218);
and U16795 (N_16795,N_8614,N_12025);
and U16796 (N_16796,N_8483,N_9106);
and U16797 (N_16797,N_12261,N_8411);
nor U16798 (N_16798,N_11073,N_9087);
and U16799 (N_16799,N_9018,N_8194);
or U16800 (N_16800,N_10458,N_6668);
and U16801 (N_16801,N_9436,N_8027);
xnor U16802 (N_16802,N_11490,N_12108);
xor U16803 (N_16803,N_6747,N_7388);
or U16804 (N_16804,N_6769,N_10373);
nand U16805 (N_16805,N_11094,N_11403);
nor U16806 (N_16806,N_10109,N_8787);
xnor U16807 (N_16807,N_10747,N_7564);
and U16808 (N_16808,N_8797,N_7994);
nand U16809 (N_16809,N_11708,N_7592);
nor U16810 (N_16810,N_11179,N_6252);
nand U16811 (N_16811,N_9427,N_11397);
nor U16812 (N_16812,N_9122,N_9180);
nor U16813 (N_16813,N_10317,N_6377);
nor U16814 (N_16814,N_7415,N_10977);
nor U16815 (N_16815,N_10501,N_11047);
xor U16816 (N_16816,N_7164,N_7374);
or U16817 (N_16817,N_9556,N_8988);
and U16818 (N_16818,N_8901,N_10782);
and U16819 (N_16819,N_8943,N_9782);
and U16820 (N_16820,N_12480,N_10292);
and U16821 (N_16821,N_11839,N_9579);
nor U16822 (N_16822,N_8264,N_11363);
xor U16823 (N_16823,N_10168,N_11843);
xor U16824 (N_16824,N_7782,N_12330);
nand U16825 (N_16825,N_6455,N_6374);
or U16826 (N_16826,N_8829,N_8242);
xnor U16827 (N_16827,N_8422,N_10937);
and U16828 (N_16828,N_6937,N_6508);
xor U16829 (N_16829,N_6956,N_6269);
nor U16830 (N_16830,N_12176,N_10874);
nor U16831 (N_16831,N_6265,N_9407);
and U16832 (N_16832,N_8859,N_6633);
xor U16833 (N_16833,N_10725,N_6895);
nor U16834 (N_16834,N_11250,N_9702);
nand U16835 (N_16835,N_9774,N_11630);
nor U16836 (N_16836,N_11707,N_8026);
xor U16837 (N_16837,N_10606,N_6537);
xnor U16838 (N_16838,N_11960,N_12185);
xor U16839 (N_16839,N_9085,N_10990);
and U16840 (N_16840,N_11480,N_9778);
nor U16841 (N_16841,N_11885,N_12144);
and U16842 (N_16842,N_8228,N_7464);
and U16843 (N_16843,N_9767,N_10495);
and U16844 (N_16844,N_10707,N_12175);
nand U16845 (N_16845,N_10025,N_11396);
nor U16846 (N_16846,N_10730,N_8735);
nor U16847 (N_16847,N_8840,N_12133);
xnor U16848 (N_16848,N_11972,N_6283);
nor U16849 (N_16849,N_8079,N_7124);
xor U16850 (N_16850,N_11875,N_6555);
nand U16851 (N_16851,N_12018,N_8057);
and U16852 (N_16852,N_7948,N_6313);
xnor U16853 (N_16853,N_6274,N_6529);
nand U16854 (N_16854,N_11719,N_10423);
and U16855 (N_16855,N_9336,N_6352);
or U16856 (N_16856,N_8232,N_7083);
xor U16857 (N_16857,N_10798,N_7802);
or U16858 (N_16858,N_8054,N_10517);
or U16859 (N_16859,N_10284,N_11132);
xnor U16860 (N_16860,N_10986,N_10949);
or U16861 (N_16861,N_10633,N_9905);
and U16862 (N_16862,N_7542,N_7956);
nand U16863 (N_16863,N_7557,N_11873);
nor U16864 (N_16864,N_11013,N_7333);
xnor U16865 (N_16865,N_8850,N_8957);
nand U16866 (N_16866,N_12137,N_10301);
and U16867 (N_16867,N_8654,N_8843);
nand U16868 (N_16868,N_7520,N_11105);
or U16869 (N_16869,N_9074,N_8254);
xnor U16870 (N_16870,N_7691,N_11146);
nor U16871 (N_16871,N_8117,N_7757);
and U16872 (N_16872,N_8466,N_9022);
nor U16873 (N_16873,N_10659,N_6403);
nand U16874 (N_16874,N_7216,N_11310);
xnor U16875 (N_16875,N_11767,N_7898);
nor U16876 (N_16876,N_6517,N_9136);
nor U16877 (N_16877,N_9666,N_8101);
nand U16878 (N_16878,N_9348,N_7592);
and U16879 (N_16879,N_6759,N_9882);
xnor U16880 (N_16880,N_11119,N_7746);
nor U16881 (N_16881,N_8195,N_11663);
nand U16882 (N_16882,N_7134,N_12233);
nor U16883 (N_16883,N_7016,N_9806);
or U16884 (N_16884,N_8321,N_9852);
nand U16885 (N_16885,N_11938,N_10847);
nor U16886 (N_16886,N_8914,N_12125);
nor U16887 (N_16887,N_6603,N_12156);
nor U16888 (N_16888,N_9047,N_6685);
xor U16889 (N_16889,N_6472,N_7361);
xnor U16890 (N_16890,N_10167,N_11843);
nand U16891 (N_16891,N_7717,N_8770);
or U16892 (N_16892,N_9584,N_11091);
xnor U16893 (N_16893,N_9712,N_8587);
xnor U16894 (N_16894,N_7781,N_7733);
nand U16895 (N_16895,N_9522,N_7685);
nor U16896 (N_16896,N_8680,N_7394);
or U16897 (N_16897,N_10212,N_9323);
xnor U16898 (N_16898,N_9927,N_6901);
and U16899 (N_16899,N_6693,N_6945);
and U16900 (N_16900,N_6623,N_11476);
or U16901 (N_16901,N_10385,N_9022);
nor U16902 (N_16902,N_10066,N_7653);
xor U16903 (N_16903,N_7802,N_10310);
or U16904 (N_16904,N_9103,N_9262);
nor U16905 (N_16905,N_10752,N_7147);
nor U16906 (N_16906,N_7564,N_11366);
or U16907 (N_16907,N_7886,N_8692);
and U16908 (N_16908,N_9549,N_8829);
xor U16909 (N_16909,N_7570,N_9375);
or U16910 (N_16910,N_8403,N_8273);
nor U16911 (N_16911,N_12470,N_9590);
nor U16912 (N_16912,N_6931,N_12114);
xor U16913 (N_16913,N_7386,N_6783);
nand U16914 (N_16914,N_11906,N_9397);
nor U16915 (N_16915,N_8933,N_11186);
nand U16916 (N_16916,N_12088,N_7487);
nor U16917 (N_16917,N_7483,N_11886);
nand U16918 (N_16918,N_10618,N_11647);
and U16919 (N_16919,N_6829,N_11209);
nor U16920 (N_16920,N_8186,N_9074);
nor U16921 (N_16921,N_9514,N_11027);
nor U16922 (N_16922,N_11941,N_10971);
nor U16923 (N_16923,N_9452,N_10968);
nand U16924 (N_16924,N_6811,N_6960);
nor U16925 (N_16925,N_12108,N_9861);
nor U16926 (N_16926,N_7825,N_7710);
or U16927 (N_16927,N_11621,N_8314);
nor U16928 (N_16928,N_9588,N_12240);
and U16929 (N_16929,N_12088,N_8917);
xnor U16930 (N_16930,N_11424,N_12013);
and U16931 (N_16931,N_8177,N_11113);
and U16932 (N_16932,N_7035,N_8077);
nand U16933 (N_16933,N_10095,N_10313);
and U16934 (N_16934,N_11185,N_10338);
nor U16935 (N_16935,N_11412,N_10734);
xor U16936 (N_16936,N_11862,N_7476);
or U16937 (N_16937,N_8922,N_11818);
and U16938 (N_16938,N_6717,N_11681);
nand U16939 (N_16939,N_7843,N_9669);
xor U16940 (N_16940,N_10258,N_9039);
xnor U16941 (N_16941,N_7577,N_7873);
and U16942 (N_16942,N_10588,N_8464);
nor U16943 (N_16943,N_10203,N_11116);
nor U16944 (N_16944,N_7737,N_12400);
nor U16945 (N_16945,N_7345,N_10554);
nor U16946 (N_16946,N_11447,N_6628);
nand U16947 (N_16947,N_7139,N_7004);
or U16948 (N_16948,N_11380,N_7788);
and U16949 (N_16949,N_7231,N_11560);
nand U16950 (N_16950,N_10706,N_7497);
xor U16951 (N_16951,N_9947,N_6839);
or U16952 (N_16952,N_11431,N_10014);
or U16953 (N_16953,N_9105,N_9148);
or U16954 (N_16954,N_7948,N_8982);
xnor U16955 (N_16955,N_11474,N_6259);
nor U16956 (N_16956,N_8420,N_8177);
xnor U16957 (N_16957,N_7967,N_10701);
xor U16958 (N_16958,N_7082,N_10868);
and U16959 (N_16959,N_7567,N_9121);
or U16960 (N_16960,N_9655,N_10497);
nand U16961 (N_16961,N_10029,N_12094);
nand U16962 (N_16962,N_7384,N_11570);
and U16963 (N_16963,N_9777,N_7316);
or U16964 (N_16964,N_11446,N_6579);
or U16965 (N_16965,N_6641,N_12488);
xor U16966 (N_16966,N_11812,N_8086);
nand U16967 (N_16967,N_9263,N_8310);
xnor U16968 (N_16968,N_7409,N_10963);
xor U16969 (N_16969,N_9635,N_7633);
or U16970 (N_16970,N_7989,N_10459);
and U16971 (N_16971,N_11269,N_11832);
and U16972 (N_16972,N_9296,N_10872);
nor U16973 (N_16973,N_9179,N_10899);
xnor U16974 (N_16974,N_7740,N_10808);
nor U16975 (N_16975,N_7300,N_10754);
nor U16976 (N_16976,N_10999,N_11846);
or U16977 (N_16977,N_8486,N_11380);
and U16978 (N_16978,N_11393,N_11001);
xnor U16979 (N_16979,N_10557,N_7586);
nand U16980 (N_16980,N_12111,N_10229);
nor U16981 (N_16981,N_11963,N_10717);
or U16982 (N_16982,N_7762,N_11403);
or U16983 (N_16983,N_7318,N_10242);
or U16984 (N_16984,N_7284,N_6326);
nor U16985 (N_16985,N_12221,N_7829);
xnor U16986 (N_16986,N_7149,N_8978);
and U16987 (N_16987,N_6414,N_10361);
nand U16988 (N_16988,N_8409,N_7148);
nand U16989 (N_16989,N_7852,N_8670);
xor U16990 (N_16990,N_8667,N_11132);
and U16991 (N_16991,N_8580,N_7152);
and U16992 (N_16992,N_8711,N_9529);
nand U16993 (N_16993,N_8411,N_9680);
xor U16994 (N_16994,N_11827,N_12422);
or U16995 (N_16995,N_6638,N_6803);
and U16996 (N_16996,N_8670,N_7425);
or U16997 (N_16997,N_7547,N_7985);
nor U16998 (N_16998,N_10315,N_7658);
nand U16999 (N_16999,N_11883,N_7050);
or U17000 (N_17000,N_8278,N_8785);
nand U17001 (N_17001,N_11690,N_9381);
nand U17002 (N_17002,N_6989,N_10933);
nor U17003 (N_17003,N_9846,N_7158);
and U17004 (N_17004,N_7449,N_9008);
xor U17005 (N_17005,N_10431,N_10469);
and U17006 (N_17006,N_10711,N_10125);
and U17007 (N_17007,N_6812,N_10073);
nand U17008 (N_17008,N_12103,N_10135);
xor U17009 (N_17009,N_12443,N_11849);
and U17010 (N_17010,N_7046,N_10428);
nand U17011 (N_17011,N_8160,N_11180);
or U17012 (N_17012,N_11983,N_9097);
nor U17013 (N_17013,N_9198,N_7528);
and U17014 (N_17014,N_10771,N_12417);
xor U17015 (N_17015,N_9192,N_12315);
and U17016 (N_17016,N_9717,N_6933);
nor U17017 (N_17017,N_6364,N_7424);
nand U17018 (N_17018,N_11638,N_11169);
xor U17019 (N_17019,N_7161,N_7018);
xor U17020 (N_17020,N_8974,N_9672);
and U17021 (N_17021,N_9238,N_11238);
and U17022 (N_17022,N_12092,N_10667);
nor U17023 (N_17023,N_8556,N_8810);
xor U17024 (N_17024,N_7983,N_11943);
nand U17025 (N_17025,N_10003,N_10672);
nor U17026 (N_17026,N_9477,N_9463);
and U17027 (N_17027,N_7450,N_9032);
and U17028 (N_17028,N_11711,N_11660);
nor U17029 (N_17029,N_8427,N_11538);
nor U17030 (N_17030,N_8929,N_9046);
nand U17031 (N_17031,N_7496,N_9133);
nand U17032 (N_17032,N_9501,N_12001);
xnor U17033 (N_17033,N_6387,N_10810);
and U17034 (N_17034,N_6615,N_11027);
nor U17035 (N_17035,N_7064,N_11179);
xor U17036 (N_17036,N_7280,N_6757);
and U17037 (N_17037,N_7828,N_8603);
or U17038 (N_17038,N_12434,N_9210);
or U17039 (N_17039,N_10550,N_10305);
or U17040 (N_17040,N_11933,N_7824);
xnor U17041 (N_17041,N_11988,N_6755);
xor U17042 (N_17042,N_9502,N_11681);
or U17043 (N_17043,N_8805,N_7712);
xnor U17044 (N_17044,N_6356,N_10643);
xnor U17045 (N_17045,N_12183,N_10220);
and U17046 (N_17046,N_10925,N_9208);
or U17047 (N_17047,N_7744,N_9574);
nor U17048 (N_17048,N_8000,N_6309);
and U17049 (N_17049,N_7506,N_8368);
and U17050 (N_17050,N_11715,N_8224);
or U17051 (N_17051,N_10199,N_8132);
and U17052 (N_17052,N_7878,N_10949);
and U17053 (N_17053,N_6961,N_8438);
or U17054 (N_17054,N_8838,N_7658);
or U17055 (N_17055,N_7360,N_8144);
and U17056 (N_17056,N_11666,N_11561);
nand U17057 (N_17057,N_10466,N_11401);
nor U17058 (N_17058,N_6769,N_11557);
xnor U17059 (N_17059,N_8218,N_6879);
xor U17060 (N_17060,N_11502,N_10123);
and U17061 (N_17061,N_7652,N_11283);
and U17062 (N_17062,N_9301,N_9950);
xor U17063 (N_17063,N_6908,N_6493);
nor U17064 (N_17064,N_10031,N_9857);
xor U17065 (N_17065,N_11034,N_11196);
nand U17066 (N_17066,N_11190,N_6865);
and U17067 (N_17067,N_11417,N_9877);
nor U17068 (N_17068,N_6929,N_9819);
or U17069 (N_17069,N_9969,N_8968);
nor U17070 (N_17070,N_10214,N_10925);
nor U17071 (N_17071,N_8467,N_11878);
nand U17072 (N_17072,N_12459,N_9763);
or U17073 (N_17073,N_7579,N_8856);
and U17074 (N_17074,N_10062,N_6828);
nor U17075 (N_17075,N_6621,N_7499);
nand U17076 (N_17076,N_11191,N_8936);
nand U17077 (N_17077,N_6596,N_7117);
or U17078 (N_17078,N_8886,N_8549);
nand U17079 (N_17079,N_7704,N_6581);
nor U17080 (N_17080,N_6922,N_6812);
xor U17081 (N_17081,N_11758,N_6659);
or U17082 (N_17082,N_9979,N_10331);
or U17083 (N_17083,N_12394,N_8453);
xor U17084 (N_17084,N_11792,N_7280);
or U17085 (N_17085,N_6734,N_9925);
nand U17086 (N_17086,N_11970,N_7727);
xnor U17087 (N_17087,N_8378,N_10941);
and U17088 (N_17088,N_11461,N_11873);
nor U17089 (N_17089,N_10588,N_7060);
xnor U17090 (N_17090,N_10331,N_6870);
or U17091 (N_17091,N_8767,N_10568);
and U17092 (N_17092,N_10930,N_10450);
nand U17093 (N_17093,N_11904,N_8903);
nor U17094 (N_17094,N_8282,N_8645);
or U17095 (N_17095,N_7269,N_11639);
nand U17096 (N_17096,N_9007,N_10960);
xnor U17097 (N_17097,N_6392,N_11614);
xnor U17098 (N_17098,N_10108,N_11464);
or U17099 (N_17099,N_9154,N_11540);
and U17100 (N_17100,N_7282,N_9021);
nor U17101 (N_17101,N_8101,N_6621);
nor U17102 (N_17102,N_9126,N_8425);
and U17103 (N_17103,N_8201,N_11549);
or U17104 (N_17104,N_7415,N_9325);
nor U17105 (N_17105,N_11969,N_11332);
or U17106 (N_17106,N_8885,N_6668);
or U17107 (N_17107,N_9738,N_6807);
or U17108 (N_17108,N_7063,N_6493);
and U17109 (N_17109,N_11009,N_6647);
and U17110 (N_17110,N_7866,N_10634);
and U17111 (N_17111,N_8179,N_8241);
xor U17112 (N_17112,N_10041,N_8094);
and U17113 (N_17113,N_8935,N_7333);
nor U17114 (N_17114,N_6430,N_10288);
xor U17115 (N_17115,N_10171,N_8590);
xnor U17116 (N_17116,N_6925,N_11000);
nor U17117 (N_17117,N_6591,N_12420);
and U17118 (N_17118,N_9891,N_7241);
nand U17119 (N_17119,N_11003,N_6317);
nor U17120 (N_17120,N_7345,N_8631);
nand U17121 (N_17121,N_9471,N_9014);
and U17122 (N_17122,N_8189,N_6437);
and U17123 (N_17123,N_9347,N_11539);
xor U17124 (N_17124,N_9472,N_7526);
nand U17125 (N_17125,N_7298,N_11382);
xor U17126 (N_17126,N_9333,N_9793);
xnor U17127 (N_17127,N_7942,N_8733);
nand U17128 (N_17128,N_7453,N_10043);
nand U17129 (N_17129,N_11961,N_8172);
xnor U17130 (N_17130,N_8260,N_8917);
and U17131 (N_17131,N_7442,N_6616);
xnor U17132 (N_17132,N_8499,N_7680);
or U17133 (N_17133,N_8723,N_10921);
and U17134 (N_17134,N_12167,N_11159);
nand U17135 (N_17135,N_10708,N_7934);
and U17136 (N_17136,N_6481,N_8132);
or U17137 (N_17137,N_10516,N_7300);
nand U17138 (N_17138,N_7765,N_6656);
and U17139 (N_17139,N_10658,N_10434);
and U17140 (N_17140,N_11606,N_9439);
nor U17141 (N_17141,N_7343,N_12070);
nand U17142 (N_17142,N_10130,N_11464);
nor U17143 (N_17143,N_7723,N_9007);
and U17144 (N_17144,N_7053,N_9728);
nand U17145 (N_17145,N_12147,N_8556);
xnor U17146 (N_17146,N_9289,N_6991);
and U17147 (N_17147,N_7109,N_7499);
nand U17148 (N_17148,N_11897,N_7830);
xnor U17149 (N_17149,N_8127,N_12052);
or U17150 (N_17150,N_8112,N_10923);
nor U17151 (N_17151,N_8162,N_9364);
nor U17152 (N_17152,N_7961,N_10147);
nand U17153 (N_17153,N_9824,N_8751);
or U17154 (N_17154,N_7403,N_8726);
xor U17155 (N_17155,N_9894,N_10017);
xnor U17156 (N_17156,N_7161,N_9448);
nand U17157 (N_17157,N_6808,N_11174);
and U17158 (N_17158,N_12077,N_8003);
nand U17159 (N_17159,N_8523,N_8353);
and U17160 (N_17160,N_10111,N_6544);
or U17161 (N_17161,N_9035,N_7862);
xnor U17162 (N_17162,N_6250,N_10664);
nand U17163 (N_17163,N_7532,N_8111);
nand U17164 (N_17164,N_11007,N_9940);
or U17165 (N_17165,N_7575,N_11586);
nand U17166 (N_17166,N_10051,N_12166);
and U17167 (N_17167,N_9816,N_10019);
nor U17168 (N_17168,N_11885,N_11031);
xor U17169 (N_17169,N_7481,N_10833);
and U17170 (N_17170,N_11931,N_8063);
nor U17171 (N_17171,N_8877,N_9212);
xor U17172 (N_17172,N_8730,N_9363);
nand U17173 (N_17173,N_9112,N_9917);
xor U17174 (N_17174,N_9284,N_7620);
xnor U17175 (N_17175,N_9882,N_12118);
nand U17176 (N_17176,N_12081,N_7694);
and U17177 (N_17177,N_7417,N_6481);
or U17178 (N_17178,N_7082,N_7256);
nand U17179 (N_17179,N_12073,N_6352);
xnor U17180 (N_17180,N_9694,N_7170);
and U17181 (N_17181,N_10888,N_10410);
xnor U17182 (N_17182,N_7887,N_10254);
xnor U17183 (N_17183,N_11197,N_8822);
and U17184 (N_17184,N_8246,N_10460);
xnor U17185 (N_17185,N_8086,N_11273);
and U17186 (N_17186,N_7194,N_6833);
nand U17187 (N_17187,N_12160,N_12218);
or U17188 (N_17188,N_8479,N_8929);
nand U17189 (N_17189,N_9790,N_7443);
nor U17190 (N_17190,N_8547,N_9407);
xnor U17191 (N_17191,N_9286,N_6811);
xnor U17192 (N_17192,N_6898,N_10381);
xor U17193 (N_17193,N_7264,N_6784);
nor U17194 (N_17194,N_9829,N_9946);
xnor U17195 (N_17195,N_9082,N_6495);
and U17196 (N_17196,N_7735,N_8187);
nand U17197 (N_17197,N_7211,N_6274);
nor U17198 (N_17198,N_7452,N_12454);
xnor U17199 (N_17199,N_9828,N_12262);
nor U17200 (N_17200,N_10310,N_7381);
or U17201 (N_17201,N_9573,N_11678);
or U17202 (N_17202,N_9695,N_6437);
nor U17203 (N_17203,N_8746,N_9000);
and U17204 (N_17204,N_7404,N_11407);
nand U17205 (N_17205,N_9272,N_11379);
xnor U17206 (N_17206,N_11857,N_8739);
nand U17207 (N_17207,N_10289,N_7785);
nand U17208 (N_17208,N_10464,N_8400);
nor U17209 (N_17209,N_9225,N_8152);
or U17210 (N_17210,N_8721,N_7767);
nor U17211 (N_17211,N_6520,N_7501);
nand U17212 (N_17212,N_6805,N_7625);
nor U17213 (N_17213,N_7194,N_7377);
and U17214 (N_17214,N_7635,N_9078);
nand U17215 (N_17215,N_9557,N_10165);
and U17216 (N_17216,N_8549,N_11443);
or U17217 (N_17217,N_7580,N_10251);
nor U17218 (N_17218,N_6348,N_8491);
xor U17219 (N_17219,N_6731,N_8532);
xnor U17220 (N_17220,N_8773,N_11417);
or U17221 (N_17221,N_6426,N_10957);
and U17222 (N_17222,N_9713,N_8312);
or U17223 (N_17223,N_9149,N_10431);
xnor U17224 (N_17224,N_8392,N_10709);
nand U17225 (N_17225,N_8573,N_7833);
nor U17226 (N_17226,N_11286,N_11545);
xnor U17227 (N_17227,N_12194,N_9785);
and U17228 (N_17228,N_10040,N_11535);
or U17229 (N_17229,N_9857,N_7602);
xnor U17230 (N_17230,N_12298,N_8592);
nand U17231 (N_17231,N_10872,N_10134);
and U17232 (N_17232,N_10060,N_11670);
and U17233 (N_17233,N_9156,N_9380);
nor U17234 (N_17234,N_10608,N_10270);
xor U17235 (N_17235,N_7731,N_10498);
nor U17236 (N_17236,N_11883,N_8295);
and U17237 (N_17237,N_7613,N_11589);
nor U17238 (N_17238,N_11185,N_10914);
nor U17239 (N_17239,N_6482,N_6469);
or U17240 (N_17240,N_9944,N_8659);
or U17241 (N_17241,N_9927,N_12210);
xnor U17242 (N_17242,N_9571,N_11812);
and U17243 (N_17243,N_6299,N_9249);
xnor U17244 (N_17244,N_10697,N_9111);
or U17245 (N_17245,N_7335,N_6663);
xnor U17246 (N_17246,N_12283,N_8780);
or U17247 (N_17247,N_7076,N_10274);
nor U17248 (N_17248,N_8027,N_9177);
and U17249 (N_17249,N_8388,N_7796);
nor U17250 (N_17250,N_7209,N_9914);
nor U17251 (N_17251,N_6270,N_9917);
or U17252 (N_17252,N_10800,N_6341);
nand U17253 (N_17253,N_7112,N_8865);
xnor U17254 (N_17254,N_11081,N_11346);
xnor U17255 (N_17255,N_10120,N_11543);
nand U17256 (N_17256,N_11980,N_6438);
nor U17257 (N_17257,N_8056,N_8947);
and U17258 (N_17258,N_8941,N_12316);
nor U17259 (N_17259,N_9350,N_12465);
xor U17260 (N_17260,N_12480,N_10890);
and U17261 (N_17261,N_11048,N_11301);
nor U17262 (N_17262,N_9155,N_8935);
nor U17263 (N_17263,N_11339,N_6479);
nor U17264 (N_17264,N_10589,N_9145);
nand U17265 (N_17265,N_7746,N_10752);
or U17266 (N_17266,N_11793,N_8658);
or U17267 (N_17267,N_7364,N_8716);
xnor U17268 (N_17268,N_11068,N_11115);
xor U17269 (N_17269,N_8856,N_7609);
nor U17270 (N_17270,N_11513,N_11641);
nand U17271 (N_17271,N_9447,N_11130);
nand U17272 (N_17272,N_11157,N_7930);
xnor U17273 (N_17273,N_7576,N_10934);
or U17274 (N_17274,N_12428,N_11415);
xor U17275 (N_17275,N_8085,N_8380);
nor U17276 (N_17276,N_9672,N_11350);
and U17277 (N_17277,N_12488,N_11240);
and U17278 (N_17278,N_10571,N_7407);
and U17279 (N_17279,N_9940,N_7391);
xnor U17280 (N_17280,N_12138,N_11237);
xnor U17281 (N_17281,N_7172,N_11784);
or U17282 (N_17282,N_7640,N_7730);
xnor U17283 (N_17283,N_11295,N_8684);
nand U17284 (N_17284,N_7458,N_9733);
nor U17285 (N_17285,N_7446,N_8818);
nor U17286 (N_17286,N_10905,N_12444);
xor U17287 (N_17287,N_6938,N_7029);
xor U17288 (N_17288,N_11922,N_11604);
nand U17289 (N_17289,N_8136,N_10091);
nand U17290 (N_17290,N_10415,N_12368);
nor U17291 (N_17291,N_10305,N_10192);
and U17292 (N_17292,N_11345,N_10960);
or U17293 (N_17293,N_8924,N_9161);
xor U17294 (N_17294,N_7451,N_8728);
xor U17295 (N_17295,N_11740,N_11014);
nor U17296 (N_17296,N_10143,N_8768);
nand U17297 (N_17297,N_11729,N_11845);
nand U17298 (N_17298,N_9672,N_12414);
or U17299 (N_17299,N_8498,N_11519);
xnor U17300 (N_17300,N_8176,N_9056);
nor U17301 (N_17301,N_11850,N_6858);
or U17302 (N_17302,N_12316,N_10088);
nor U17303 (N_17303,N_6398,N_11622);
or U17304 (N_17304,N_7689,N_7375);
xnor U17305 (N_17305,N_12370,N_6583);
nor U17306 (N_17306,N_6626,N_12219);
nand U17307 (N_17307,N_6324,N_10152);
or U17308 (N_17308,N_8622,N_11926);
nand U17309 (N_17309,N_7885,N_7101);
and U17310 (N_17310,N_9742,N_10670);
or U17311 (N_17311,N_11787,N_10861);
or U17312 (N_17312,N_11690,N_9774);
xnor U17313 (N_17313,N_9294,N_10923);
xnor U17314 (N_17314,N_11523,N_11642);
xor U17315 (N_17315,N_8730,N_9425);
or U17316 (N_17316,N_9695,N_10997);
or U17317 (N_17317,N_7249,N_9089);
nor U17318 (N_17318,N_8346,N_6639);
xor U17319 (N_17319,N_8120,N_11175);
nand U17320 (N_17320,N_9434,N_7868);
or U17321 (N_17321,N_9984,N_6575);
nand U17322 (N_17322,N_7598,N_7769);
nand U17323 (N_17323,N_9284,N_11958);
or U17324 (N_17324,N_12477,N_8542);
xor U17325 (N_17325,N_7447,N_8456);
nor U17326 (N_17326,N_8355,N_8309);
and U17327 (N_17327,N_6557,N_7216);
or U17328 (N_17328,N_9733,N_9671);
xor U17329 (N_17329,N_7023,N_7416);
xnor U17330 (N_17330,N_7500,N_12373);
and U17331 (N_17331,N_9860,N_8175);
nand U17332 (N_17332,N_10059,N_10306);
and U17333 (N_17333,N_8593,N_10780);
or U17334 (N_17334,N_8880,N_10204);
nand U17335 (N_17335,N_7662,N_12035);
nand U17336 (N_17336,N_10288,N_8577);
and U17337 (N_17337,N_8259,N_12232);
nand U17338 (N_17338,N_11792,N_10066);
and U17339 (N_17339,N_9123,N_10108);
or U17340 (N_17340,N_10979,N_9921);
xnor U17341 (N_17341,N_11333,N_8725);
nor U17342 (N_17342,N_6549,N_12338);
nand U17343 (N_17343,N_12151,N_10538);
xnor U17344 (N_17344,N_9664,N_8783);
nand U17345 (N_17345,N_10818,N_7839);
nor U17346 (N_17346,N_11682,N_10908);
or U17347 (N_17347,N_10658,N_6411);
nor U17348 (N_17348,N_9401,N_9231);
nand U17349 (N_17349,N_12158,N_10520);
xnor U17350 (N_17350,N_10679,N_10781);
nand U17351 (N_17351,N_10594,N_9885);
nor U17352 (N_17352,N_7874,N_6514);
nand U17353 (N_17353,N_8283,N_10479);
nand U17354 (N_17354,N_8359,N_7386);
nor U17355 (N_17355,N_6356,N_7435);
nand U17356 (N_17356,N_12180,N_9883);
nand U17357 (N_17357,N_6392,N_10683);
or U17358 (N_17358,N_8295,N_6268);
nor U17359 (N_17359,N_6626,N_10222);
or U17360 (N_17360,N_8630,N_9919);
nor U17361 (N_17361,N_7239,N_12033);
nand U17362 (N_17362,N_9993,N_9983);
or U17363 (N_17363,N_11284,N_7683);
nor U17364 (N_17364,N_10025,N_11710);
and U17365 (N_17365,N_12430,N_6333);
or U17366 (N_17366,N_12247,N_7865);
xnor U17367 (N_17367,N_9797,N_10381);
and U17368 (N_17368,N_9352,N_11276);
xor U17369 (N_17369,N_9700,N_12441);
or U17370 (N_17370,N_10044,N_8704);
nand U17371 (N_17371,N_6302,N_11635);
nand U17372 (N_17372,N_12290,N_11642);
and U17373 (N_17373,N_8163,N_11141);
nand U17374 (N_17374,N_11254,N_8351);
nand U17375 (N_17375,N_8017,N_8961);
or U17376 (N_17376,N_9662,N_7764);
or U17377 (N_17377,N_11258,N_10389);
xnor U17378 (N_17378,N_6414,N_11755);
nor U17379 (N_17379,N_12058,N_8480);
nand U17380 (N_17380,N_6841,N_9751);
xnor U17381 (N_17381,N_9838,N_8864);
or U17382 (N_17382,N_10879,N_9649);
and U17383 (N_17383,N_10310,N_7235);
nand U17384 (N_17384,N_8822,N_12289);
xnor U17385 (N_17385,N_6310,N_11677);
or U17386 (N_17386,N_10141,N_8124);
and U17387 (N_17387,N_10949,N_6996);
and U17388 (N_17388,N_11420,N_7890);
or U17389 (N_17389,N_7561,N_9272);
and U17390 (N_17390,N_11601,N_6465);
xnor U17391 (N_17391,N_11516,N_8772);
xor U17392 (N_17392,N_6873,N_10335);
or U17393 (N_17393,N_9502,N_10507);
or U17394 (N_17394,N_8168,N_9598);
and U17395 (N_17395,N_9478,N_11913);
or U17396 (N_17396,N_11992,N_9254);
nor U17397 (N_17397,N_11209,N_11172);
xor U17398 (N_17398,N_7368,N_6940);
and U17399 (N_17399,N_7812,N_9177);
xnor U17400 (N_17400,N_11219,N_6804);
nor U17401 (N_17401,N_9476,N_6452);
and U17402 (N_17402,N_8034,N_6817);
nand U17403 (N_17403,N_7022,N_8797);
or U17404 (N_17404,N_11491,N_9618);
xnor U17405 (N_17405,N_9030,N_7337);
and U17406 (N_17406,N_8512,N_6684);
or U17407 (N_17407,N_7967,N_6950);
nor U17408 (N_17408,N_10808,N_7760);
nand U17409 (N_17409,N_6653,N_7689);
xor U17410 (N_17410,N_8305,N_8220);
and U17411 (N_17411,N_10861,N_10659);
or U17412 (N_17412,N_10726,N_9733);
or U17413 (N_17413,N_9629,N_6723);
nor U17414 (N_17414,N_9118,N_8073);
nand U17415 (N_17415,N_10396,N_6701);
nand U17416 (N_17416,N_11921,N_10087);
xor U17417 (N_17417,N_8451,N_11600);
nor U17418 (N_17418,N_11562,N_7811);
nand U17419 (N_17419,N_6996,N_7765);
or U17420 (N_17420,N_11599,N_11645);
or U17421 (N_17421,N_7055,N_12142);
and U17422 (N_17422,N_11962,N_8109);
nand U17423 (N_17423,N_10686,N_10308);
nand U17424 (N_17424,N_11194,N_9438);
nor U17425 (N_17425,N_6535,N_12268);
and U17426 (N_17426,N_8571,N_12224);
xnor U17427 (N_17427,N_8154,N_8226);
nand U17428 (N_17428,N_7525,N_9035);
and U17429 (N_17429,N_10636,N_9901);
or U17430 (N_17430,N_8184,N_11861);
nor U17431 (N_17431,N_9215,N_9554);
nor U17432 (N_17432,N_7436,N_12497);
or U17433 (N_17433,N_11029,N_8070);
and U17434 (N_17434,N_12043,N_12449);
or U17435 (N_17435,N_10090,N_10477);
or U17436 (N_17436,N_10797,N_10996);
nand U17437 (N_17437,N_8113,N_10579);
xor U17438 (N_17438,N_12335,N_7244);
xor U17439 (N_17439,N_6516,N_10629);
nor U17440 (N_17440,N_7155,N_8045);
nor U17441 (N_17441,N_7697,N_9800);
or U17442 (N_17442,N_10090,N_6646);
or U17443 (N_17443,N_10816,N_7851);
and U17444 (N_17444,N_10852,N_7173);
or U17445 (N_17445,N_11550,N_12328);
nand U17446 (N_17446,N_11508,N_10779);
and U17447 (N_17447,N_12333,N_8758);
or U17448 (N_17448,N_8331,N_12114);
or U17449 (N_17449,N_9008,N_9480);
and U17450 (N_17450,N_11380,N_9595);
xor U17451 (N_17451,N_9904,N_7837);
or U17452 (N_17452,N_7384,N_9425);
nor U17453 (N_17453,N_9452,N_11636);
xor U17454 (N_17454,N_11416,N_6299);
nand U17455 (N_17455,N_7170,N_7238);
and U17456 (N_17456,N_9096,N_6349);
or U17457 (N_17457,N_10468,N_6797);
and U17458 (N_17458,N_6421,N_7677);
nor U17459 (N_17459,N_11208,N_6400);
nor U17460 (N_17460,N_7798,N_10832);
nand U17461 (N_17461,N_9794,N_8914);
nor U17462 (N_17462,N_7224,N_11807);
xnor U17463 (N_17463,N_7537,N_11913);
or U17464 (N_17464,N_7432,N_7737);
xor U17465 (N_17465,N_8405,N_6864);
nor U17466 (N_17466,N_10538,N_10823);
or U17467 (N_17467,N_7814,N_10464);
or U17468 (N_17468,N_6417,N_7678);
and U17469 (N_17469,N_8031,N_7355);
nand U17470 (N_17470,N_11283,N_12196);
xor U17471 (N_17471,N_10688,N_11574);
nand U17472 (N_17472,N_11648,N_8756);
nor U17473 (N_17473,N_6661,N_8758);
nand U17474 (N_17474,N_11452,N_8520);
xnor U17475 (N_17475,N_9785,N_10297);
nand U17476 (N_17476,N_6637,N_7179);
and U17477 (N_17477,N_7065,N_10963);
or U17478 (N_17478,N_11529,N_12333);
nor U17479 (N_17479,N_10088,N_8521);
nor U17480 (N_17480,N_8925,N_9169);
and U17481 (N_17481,N_7922,N_11686);
xor U17482 (N_17482,N_6332,N_8911);
xnor U17483 (N_17483,N_11194,N_9639);
nand U17484 (N_17484,N_12373,N_7303);
and U17485 (N_17485,N_11395,N_6506);
and U17486 (N_17486,N_7614,N_12041);
nor U17487 (N_17487,N_8218,N_8772);
nor U17488 (N_17488,N_9071,N_8396);
nand U17489 (N_17489,N_9445,N_11884);
xnor U17490 (N_17490,N_8495,N_8652);
and U17491 (N_17491,N_11452,N_7264);
and U17492 (N_17492,N_10283,N_8940);
nor U17493 (N_17493,N_11978,N_8520);
and U17494 (N_17494,N_9458,N_10210);
xor U17495 (N_17495,N_9974,N_8945);
nor U17496 (N_17496,N_11216,N_9360);
xor U17497 (N_17497,N_9185,N_7279);
nand U17498 (N_17498,N_11839,N_7071);
nor U17499 (N_17499,N_7638,N_11307);
nand U17500 (N_17500,N_12211,N_8323);
or U17501 (N_17501,N_7992,N_10076);
nor U17502 (N_17502,N_9041,N_11318);
nor U17503 (N_17503,N_11305,N_7575);
and U17504 (N_17504,N_9760,N_11847);
nand U17505 (N_17505,N_7951,N_9580);
xnor U17506 (N_17506,N_6374,N_10518);
nor U17507 (N_17507,N_8354,N_9936);
or U17508 (N_17508,N_7140,N_9052);
nand U17509 (N_17509,N_10173,N_8346);
nor U17510 (N_17510,N_8900,N_10328);
or U17511 (N_17511,N_12462,N_8891);
xor U17512 (N_17512,N_8985,N_12162);
nand U17513 (N_17513,N_8022,N_7988);
and U17514 (N_17514,N_8981,N_8663);
or U17515 (N_17515,N_9949,N_10807);
nor U17516 (N_17516,N_8016,N_12487);
and U17517 (N_17517,N_8156,N_11820);
and U17518 (N_17518,N_7010,N_9433);
xnor U17519 (N_17519,N_8110,N_7520);
and U17520 (N_17520,N_12086,N_9712);
or U17521 (N_17521,N_11244,N_12085);
and U17522 (N_17522,N_10409,N_8584);
xor U17523 (N_17523,N_6928,N_6333);
nand U17524 (N_17524,N_11414,N_10375);
xnor U17525 (N_17525,N_7225,N_6605);
and U17526 (N_17526,N_11270,N_8471);
or U17527 (N_17527,N_11849,N_7872);
nor U17528 (N_17528,N_9277,N_6817);
nand U17529 (N_17529,N_6865,N_7004);
nor U17530 (N_17530,N_6853,N_7192);
nor U17531 (N_17531,N_7752,N_9481);
xor U17532 (N_17532,N_7111,N_11936);
and U17533 (N_17533,N_8503,N_7735);
and U17534 (N_17534,N_9188,N_10555);
and U17535 (N_17535,N_7702,N_10513);
or U17536 (N_17536,N_11402,N_8427);
or U17537 (N_17537,N_8080,N_8364);
nand U17538 (N_17538,N_11074,N_10526);
and U17539 (N_17539,N_6535,N_11291);
nand U17540 (N_17540,N_9414,N_12218);
nor U17541 (N_17541,N_6262,N_12139);
nor U17542 (N_17542,N_11322,N_6959);
xor U17543 (N_17543,N_6731,N_7741);
nand U17544 (N_17544,N_10483,N_8972);
or U17545 (N_17545,N_10910,N_11244);
and U17546 (N_17546,N_11921,N_9973);
nor U17547 (N_17547,N_11315,N_8454);
nand U17548 (N_17548,N_10111,N_10037);
or U17549 (N_17549,N_8605,N_9263);
xor U17550 (N_17550,N_6445,N_11266);
and U17551 (N_17551,N_11449,N_11621);
xor U17552 (N_17552,N_7401,N_7398);
or U17553 (N_17553,N_11412,N_11901);
nand U17554 (N_17554,N_7769,N_8220);
or U17555 (N_17555,N_6271,N_6428);
or U17556 (N_17556,N_9983,N_6465);
xnor U17557 (N_17557,N_9351,N_7237);
and U17558 (N_17558,N_8946,N_8782);
nand U17559 (N_17559,N_9542,N_6833);
nor U17560 (N_17560,N_9775,N_11214);
nand U17561 (N_17561,N_9245,N_11574);
and U17562 (N_17562,N_8146,N_11323);
or U17563 (N_17563,N_7817,N_6535);
nor U17564 (N_17564,N_11981,N_12019);
and U17565 (N_17565,N_7755,N_6614);
or U17566 (N_17566,N_11530,N_10596);
xnor U17567 (N_17567,N_9883,N_7813);
xor U17568 (N_17568,N_11946,N_9311);
xnor U17569 (N_17569,N_12426,N_6844);
and U17570 (N_17570,N_9751,N_7695);
xor U17571 (N_17571,N_11291,N_7426);
nand U17572 (N_17572,N_9286,N_9925);
nand U17573 (N_17573,N_10962,N_8889);
xnor U17574 (N_17574,N_7459,N_7843);
and U17575 (N_17575,N_11348,N_8131);
and U17576 (N_17576,N_8690,N_7185);
nand U17577 (N_17577,N_7496,N_9964);
nand U17578 (N_17578,N_11096,N_9304);
xor U17579 (N_17579,N_8082,N_7795);
nand U17580 (N_17580,N_10475,N_6594);
and U17581 (N_17581,N_11850,N_7967);
or U17582 (N_17582,N_11086,N_6621);
nor U17583 (N_17583,N_6291,N_12114);
nand U17584 (N_17584,N_8681,N_8956);
and U17585 (N_17585,N_11495,N_11233);
nand U17586 (N_17586,N_12214,N_9950);
nand U17587 (N_17587,N_12382,N_8390);
and U17588 (N_17588,N_11265,N_7732);
xnor U17589 (N_17589,N_11156,N_8817);
xnor U17590 (N_17590,N_11651,N_7750);
or U17591 (N_17591,N_8637,N_10616);
nand U17592 (N_17592,N_7829,N_8623);
nor U17593 (N_17593,N_7784,N_11600);
nor U17594 (N_17594,N_7084,N_10671);
or U17595 (N_17595,N_10040,N_7239);
nor U17596 (N_17596,N_11373,N_8994);
nor U17597 (N_17597,N_10680,N_11906);
xnor U17598 (N_17598,N_9418,N_9860);
nor U17599 (N_17599,N_10764,N_8148);
xor U17600 (N_17600,N_9715,N_6565);
or U17601 (N_17601,N_11181,N_11490);
nor U17602 (N_17602,N_10895,N_7495);
and U17603 (N_17603,N_9941,N_9794);
nand U17604 (N_17604,N_12475,N_8780);
xnor U17605 (N_17605,N_12447,N_12398);
xnor U17606 (N_17606,N_10992,N_9066);
nand U17607 (N_17607,N_10121,N_10703);
nor U17608 (N_17608,N_12499,N_10261);
nor U17609 (N_17609,N_8787,N_12453);
and U17610 (N_17610,N_6880,N_9916);
or U17611 (N_17611,N_11785,N_11174);
nand U17612 (N_17612,N_10622,N_12217);
nor U17613 (N_17613,N_11991,N_7939);
and U17614 (N_17614,N_12117,N_9905);
nor U17615 (N_17615,N_9043,N_8102);
nand U17616 (N_17616,N_10980,N_11030);
xnor U17617 (N_17617,N_11635,N_10982);
and U17618 (N_17618,N_6307,N_8738);
xnor U17619 (N_17619,N_10783,N_8612);
xnor U17620 (N_17620,N_6279,N_9380);
nand U17621 (N_17621,N_12287,N_10961);
or U17622 (N_17622,N_6997,N_11953);
or U17623 (N_17623,N_8707,N_9524);
and U17624 (N_17624,N_11776,N_8345);
nor U17625 (N_17625,N_8716,N_10270);
nor U17626 (N_17626,N_9188,N_7358);
xnor U17627 (N_17627,N_11612,N_6710);
and U17628 (N_17628,N_10019,N_7560);
xor U17629 (N_17629,N_7098,N_10241);
nor U17630 (N_17630,N_7487,N_10082);
and U17631 (N_17631,N_6379,N_8700);
nand U17632 (N_17632,N_8071,N_7422);
xnor U17633 (N_17633,N_11705,N_11787);
nand U17634 (N_17634,N_8469,N_11788);
or U17635 (N_17635,N_11515,N_9578);
or U17636 (N_17636,N_10122,N_8286);
nor U17637 (N_17637,N_6624,N_6299);
nor U17638 (N_17638,N_10700,N_8805);
or U17639 (N_17639,N_6728,N_10665);
nand U17640 (N_17640,N_9468,N_10708);
or U17641 (N_17641,N_8225,N_6959);
or U17642 (N_17642,N_10562,N_10055);
xor U17643 (N_17643,N_11732,N_12090);
and U17644 (N_17644,N_11662,N_7929);
nor U17645 (N_17645,N_10857,N_10086);
nand U17646 (N_17646,N_7529,N_12031);
xor U17647 (N_17647,N_6731,N_11787);
or U17648 (N_17648,N_10204,N_9439);
or U17649 (N_17649,N_7519,N_11449);
nor U17650 (N_17650,N_9610,N_10692);
xnor U17651 (N_17651,N_11560,N_11242);
and U17652 (N_17652,N_6672,N_9900);
nand U17653 (N_17653,N_9411,N_8269);
nand U17654 (N_17654,N_11123,N_10818);
xnor U17655 (N_17655,N_6873,N_11322);
xnor U17656 (N_17656,N_8740,N_8304);
or U17657 (N_17657,N_7187,N_11385);
or U17658 (N_17658,N_6896,N_11154);
nand U17659 (N_17659,N_6881,N_9766);
and U17660 (N_17660,N_7759,N_9112);
nor U17661 (N_17661,N_7753,N_11244);
and U17662 (N_17662,N_6869,N_11555);
nor U17663 (N_17663,N_10858,N_11660);
and U17664 (N_17664,N_6505,N_6528);
or U17665 (N_17665,N_11376,N_10486);
nand U17666 (N_17666,N_7086,N_10320);
xor U17667 (N_17667,N_6508,N_7201);
nand U17668 (N_17668,N_10379,N_10725);
or U17669 (N_17669,N_11005,N_10637);
or U17670 (N_17670,N_10577,N_11536);
and U17671 (N_17671,N_12103,N_7107);
xnor U17672 (N_17672,N_8154,N_10878);
nor U17673 (N_17673,N_9791,N_9451);
nand U17674 (N_17674,N_9127,N_10560);
or U17675 (N_17675,N_10430,N_6467);
xnor U17676 (N_17676,N_11123,N_12268);
xnor U17677 (N_17677,N_11591,N_6834);
xor U17678 (N_17678,N_10337,N_8617);
xnor U17679 (N_17679,N_8026,N_6557);
xor U17680 (N_17680,N_11374,N_10416);
xnor U17681 (N_17681,N_7613,N_6416);
or U17682 (N_17682,N_11265,N_12030);
and U17683 (N_17683,N_8052,N_7846);
nor U17684 (N_17684,N_12313,N_8233);
or U17685 (N_17685,N_8817,N_9878);
xnor U17686 (N_17686,N_10633,N_9140);
nand U17687 (N_17687,N_7104,N_7808);
nor U17688 (N_17688,N_7772,N_10214);
nand U17689 (N_17689,N_7199,N_11735);
nand U17690 (N_17690,N_8532,N_10561);
nor U17691 (N_17691,N_7894,N_7489);
nand U17692 (N_17692,N_9503,N_12316);
nor U17693 (N_17693,N_7480,N_11775);
nor U17694 (N_17694,N_11593,N_6849);
or U17695 (N_17695,N_6477,N_11414);
or U17696 (N_17696,N_6892,N_7349);
or U17697 (N_17697,N_7809,N_11289);
and U17698 (N_17698,N_10795,N_7201);
xnor U17699 (N_17699,N_9200,N_9863);
nor U17700 (N_17700,N_8865,N_9093);
or U17701 (N_17701,N_6289,N_11426);
or U17702 (N_17702,N_9221,N_6452);
nand U17703 (N_17703,N_9703,N_9312);
xor U17704 (N_17704,N_9150,N_7344);
or U17705 (N_17705,N_7922,N_7766);
nand U17706 (N_17706,N_7829,N_6855);
nand U17707 (N_17707,N_6693,N_8585);
nand U17708 (N_17708,N_8565,N_7922);
and U17709 (N_17709,N_12320,N_10457);
xor U17710 (N_17710,N_11469,N_8657);
nand U17711 (N_17711,N_11283,N_8596);
nor U17712 (N_17712,N_8867,N_10949);
and U17713 (N_17713,N_12012,N_6324);
and U17714 (N_17714,N_7934,N_10217);
nand U17715 (N_17715,N_11000,N_8245);
and U17716 (N_17716,N_12390,N_7910);
and U17717 (N_17717,N_9011,N_6618);
and U17718 (N_17718,N_8249,N_7483);
xor U17719 (N_17719,N_9921,N_8480);
nor U17720 (N_17720,N_7382,N_8800);
and U17721 (N_17721,N_11797,N_7971);
and U17722 (N_17722,N_6636,N_12196);
xnor U17723 (N_17723,N_9959,N_11909);
and U17724 (N_17724,N_8596,N_8835);
xnor U17725 (N_17725,N_6621,N_12186);
and U17726 (N_17726,N_7027,N_9167);
nand U17727 (N_17727,N_12387,N_11398);
or U17728 (N_17728,N_7512,N_7496);
xnor U17729 (N_17729,N_9755,N_11606);
and U17730 (N_17730,N_10800,N_12432);
xnor U17731 (N_17731,N_11296,N_7115);
nor U17732 (N_17732,N_7766,N_11820);
or U17733 (N_17733,N_6858,N_7605);
nor U17734 (N_17734,N_7577,N_8342);
nor U17735 (N_17735,N_7772,N_9369);
and U17736 (N_17736,N_12426,N_11838);
or U17737 (N_17737,N_10951,N_9906);
and U17738 (N_17738,N_11859,N_7781);
or U17739 (N_17739,N_12217,N_6426);
or U17740 (N_17740,N_11496,N_8001);
and U17741 (N_17741,N_6843,N_8402);
xor U17742 (N_17742,N_11128,N_6810);
nor U17743 (N_17743,N_12176,N_9629);
xnor U17744 (N_17744,N_8339,N_9963);
nor U17745 (N_17745,N_9976,N_9356);
nor U17746 (N_17746,N_6509,N_6320);
xor U17747 (N_17747,N_11198,N_7332);
and U17748 (N_17748,N_8172,N_6306);
or U17749 (N_17749,N_12297,N_7949);
and U17750 (N_17750,N_12158,N_7926);
nor U17751 (N_17751,N_11028,N_9136);
xor U17752 (N_17752,N_6817,N_11060);
xor U17753 (N_17753,N_7446,N_11123);
nand U17754 (N_17754,N_10725,N_6869);
nor U17755 (N_17755,N_10096,N_11757);
xor U17756 (N_17756,N_6417,N_8235);
nand U17757 (N_17757,N_10576,N_10836);
nand U17758 (N_17758,N_6529,N_10946);
or U17759 (N_17759,N_12287,N_11353);
nor U17760 (N_17760,N_7062,N_6596);
and U17761 (N_17761,N_11325,N_7997);
xor U17762 (N_17762,N_10593,N_11667);
xor U17763 (N_17763,N_10385,N_7377);
nand U17764 (N_17764,N_10564,N_7133);
and U17765 (N_17765,N_7152,N_11179);
and U17766 (N_17766,N_7545,N_7363);
nor U17767 (N_17767,N_6630,N_8727);
and U17768 (N_17768,N_12015,N_8628);
and U17769 (N_17769,N_9223,N_12343);
nor U17770 (N_17770,N_7752,N_9272);
nand U17771 (N_17771,N_8287,N_10729);
or U17772 (N_17772,N_11504,N_8619);
nor U17773 (N_17773,N_11513,N_6810);
nand U17774 (N_17774,N_9965,N_11316);
and U17775 (N_17775,N_11149,N_7779);
or U17776 (N_17776,N_10907,N_10456);
nor U17777 (N_17777,N_8491,N_12384);
nand U17778 (N_17778,N_8652,N_7032);
or U17779 (N_17779,N_11189,N_6551);
nand U17780 (N_17780,N_8172,N_7470);
or U17781 (N_17781,N_9116,N_11713);
and U17782 (N_17782,N_7385,N_8091);
nor U17783 (N_17783,N_8011,N_8831);
nand U17784 (N_17784,N_8422,N_8697);
xnor U17785 (N_17785,N_11956,N_11088);
and U17786 (N_17786,N_11552,N_11593);
nor U17787 (N_17787,N_9908,N_7603);
xnor U17788 (N_17788,N_10195,N_10390);
and U17789 (N_17789,N_10931,N_12033);
and U17790 (N_17790,N_7648,N_11564);
nor U17791 (N_17791,N_8319,N_9121);
nor U17792 (N_17792,N_10484,N_10864);
and U17793 (N_17793,N_11063,N_9772);
xor U17794 (N_17794,N_8780,N_7368);
nor U17795 (N_17795,N_9358,N_11325);
xor U17796 (N_17796,N_11623,N_12149);
xnor U17797 (N_17797,N_11564,N_10843);
xor U17798 (N_17798,N_11375,N_12145);
and U17799 (N_17799,N_11405,N_11831);
xor U17800 (N_17800,N_7390,N_8471);
xnor U17801 (N_17801,N_8125,N_10745);
nor U17802 (N_17802,N_8480,N_9854);
nor U17803 (N_17803,N_11070,N_8896);
nor U17804 (N_17804,N_9367,N_12310);
or U17805 (N_17805,N_8774,N_11487);
nor U17806 (N_17806,N_12127,N_11903);
and U17807 (N_17807,N_10103,N_9509);
and U17808 (N_17808,N_8040,N_8778);
xor U17809 (N_17809,N_8714,N_9027);
or U17810 (N_17810,N_7089,N_8037);
or U17811 (N_17811,N_6312,N_7620);
xor U17812 (N_17812,N_7116,N_7928);
nor U17813 (N_17813,N_7844,N_10635);
nand U17814 (N_17814,N_9251,N_6805);
xnor U17815 (N_17815,N_7048,N_9946);
nor U17816 (N_17816,N_8514,N_6712);
or U17817 (N_17817,N_8816,N_6631);
or U17818 (N_17818,N_10435,N_8479);
xnor U17819 (N_17819,N_11713,N_10941);
xor U17820 (N_17820,N_9254,N_9520);
nand U17821 (N_17821,N_8000,N_7061);
or U17822 (N_17822,N_10983,N_12352);
nand U17823 (N_17823,N_8287,N_12382);
nand U17824 (N_17824,N_10506,N_6604);
xor U17825 (N_17825,N_7641,N_8554);
xnor U17826 (N_17826,N_7816,N_11947);
xnor U17827 (N_17827,N_6411,N_6722);
xnor U17828 (N_17828,N_11784,N_6419);
or U17829 (N_17829,N_10611,N_11333);
nand U17830 (N_17830,N_11332,N_11636);
and U17831 (N_17831,N_7309,N_9995);
or U17832 (N_17832,N_7563,N_10226);
or U17833 (N_17833,N_6568,N_7365);
nor U17834 (N_17834,N_8249,N_7564);
and U17835 (N_17835,N_11632,N_8827);
nor U17836 (N_17836,N_9196,N_7778);
nand U17837 (N_17837,N_6583,N_6793);
or U17838 (N_17838,N_6801,N_8145);
nor U17839 (N_17839,N_9021,N_12012);
xor U17840 (N_17840,N_11087,N_7051);
xnor U17841 (N_17841,N_11150,N_6622);
nand U17842 (N_17842,N_11917,N_6494);
nand U17843 (N_17843,N_11990,N_12265);
nand U17844 (N_17844,N_8560,N_10233);
or U17845 (N_17845,N_9972,N_12167);
or U17846 (N_17846,N_6273,N_9328);
nand U17847 (N_17847,N_6825,N_11704);
xor U17848 (N_17848,N_11213,N_9933);
nor U17849 (N_17849,N_7002,N_8714);
nor U17850 (N_17850,N_6742,N_6559);
nor U17851 (N_17851,N_10164,N_11018);
and U17852 (N_17852,N_6267,N_7747);
and U17853 (N_17853,N_7723,N_11042);
and U17854 (N_17854,N_8289,N_6777);
or U17855 (N_17855,N_11393,N_10012);
and U17856 (N_17856,N_11728,N_10758);
and U17857 (N_17857,N_12058,N_8012);
or U17858 (N_17858,N_12460,N_6676);
nor U17859 (N_17859,N_11139,N_12067);
xor U17860 (N_17860,N_9968,N_7301);
xor U17861 (N_17861,N_6677,N_9822);
or U17862 (N_17862,N_10524,N_7706);
nand U17863 (N_17863,N_11107,N_6418);
nand U17864 (N_17864,N_6992,N_11621);
nor U17865 (N_17865,N_8597,N_10051);
nor U17866 (N_17866,N_9939,N_7745);
or U17867 (N_17867,N_7857,N_12272);
nor U17868 (N_17868,N_10462,N_11853);
nand U17869 (N_17869,N_12460,N_7054);
xnor U17870 (N_17870,N_8335,N_8179);
xor U17871 (N_17871,N_10747,N_6384);
xor U17872 (N_17872,N_8103,N_9798);
nand U17873 (N_17873,N_9298,N_11236);
or U17874 (N_17874,N_8083,N_8745);
nand U17875 (N_17875,N_10394,N_9598);
nor U17876 (N_17876,N_7618,N_9848);
nor U17877 (N_17877,N_8949,N_8039);
nand U17878 (N_17878,N_11956,N_8230);
xor U17879 (N_17879,N_7542,N_9253);
and U17880 (N_17880,N_8850,N_7303);
or U17881 (N_17881,N_9825,N_7300);
xor U17882 (N_17882,N_7682,N_11667);
nand U17883 (N_17883,N_10976,N_7154);
xnor U17884 (N_17884,N_11520,N_8490);
nor U17885 (N_17885,N_11405,N_7640);
and U17886 (N_17886,N_12371,N_12114);
and U17887 (N_17887,N_9178,N_6607);
or U17888 (N_17888,N_7120,N_9979);
nand U17889 (N_17889,N_7946,N_11058);
nand U17890 (N_17890,N_7849,N_8506);
xnor U17891 (N_17891,N_10981,N_9669);
or U17892 (N_17892,N_10630,N_7866);
nand U17893 (N_17893,N_8587,N_11033);
or U17894 (N_17894,N_7891,N_8492);
or U17895 (N_17895,N_7265,N_11059);
nand U17896 (N_17896,N_10360,N_9201);
nor U17897 (N_17897,N_9670,N_6420);
nor U17898 (N_17898,N_11458,N_10035);
and U17899 (N_17899,N_7457,N_10572);
nand U17900 (N_17900,N_8192,N_10483);
or U17901 (N_17901,N_10177,N_12199);
nor U17902 (N_17902,N_8802,N_9406);
nand U17903 (N_17903,N_7299,N_9926);
and U17904 (N_17904,N_12171,N_8476);
nand U17905 (N_17905,N_9732,N_10311);
nor U17906 (N_17906,N_9612,N_10528);
xnor U17907 (N_17907,N_6934,N_8038);
nor U17908 (N_17908,N_10937,N_11930);
xor U17909 (N_17909,N_7289,N_10261);
nor U17910 (N_17910,N_11202,N_9130);
nor U17911 (N_17911,N_8856,N_11268);
or U17912 (N_17912,N_9823,N_7071);
xnor U17913 (N_17913,N_10570,N_11834);
xor U17914 (N_17914,N_12072,N_11945);
xnor U17915 (N_17915,N_6728,N_8536);
nand U17916 (N_17916,N_10880,N_10948);
nand U17917 (N_17917,N_9510,N_9119);
or U17918 (N_17918,N_11055,N_8857);
and U17919 (N_17919,N_11603,N_9252);
and U17920 (N_17920,N_8918,N_7242);
or U17921 (N_17921,N_12436,N_7729);
and U17922 (N_17922,N_7713,N_6791);
nor U17923 (N_17923,N_11435,N_12076);
and U17924 (N_17924,N_9847,N_12370);
xor U17925 (N_17925,N_6410,N_7396);
xor U17926 (N_17926,N_11528,N_8929);
or U17927 (N_17927,N_10793,N_9659);
nor U17928 (N_17928,N_11980,N_6944);
nand U17929 (N_17929,N_11069,N_8379);
or U17930 (N_17930,N_12311,N_11868);
or U17931 (N_17931,N_9109,N_12152);
nand U17932 (N_17932,N_11229,N_10413);
or U17933 (N_17933,N_7762,N_9213);
xor U17934 (N_17934,N_11781,N_7873);
nand U17935 (N_17935,N_6994,N_10903);
and U17936 (N_17936,N_10209,N_7640);
or U17937 (N_17937,N_9769,N_12191);
and U17938 (N_17938,N_6352,N_9509);
xor U17939 (N_17939,N_6254,N_7619);
or U17940 (N_17940,N_9987,N_12054);
and U17941 (N_17941,N_10698,N_9052);
or U17942 (N_17942,N_11299,N_8495);
nor U17943 (N_17943,N_9673,N_9901);
nand U17944 (N_17944,N_11672,N_9848);
or U17945 (N_17945,N_6344,N_9329);
nor U17946 (N_17946,N_6594,N_8574);
or U17947 (N_17947,N_10598,N_7031);
or U17948 (N_17948,N_12435,N_10482);
nor U17949 (N_17949,N_8161,N_9493);
and U17950 (N_17950,N_7561,N_12236);
or U17951 (N_17951,N_7923,N_6978);
or U17952 (N_17952,N_11028,N_7204);
or U17953 (N_17953,N_12356,N_11019);
and U17954 (N_17954,N_12065,N_6282);
nor U17955 (N_17955,N_9327,N_11118);
and U17956 (N_17956,N_8526,N_10241);
nor U17957 (N_17957,N_9634,N_8965);
or U17958 (N_17958,N_11453,N_7786);
xnor U17959 (N_17959,N_11229,N_7381);
nor U17960 (N_17960,N_8951,N_7967);
or U17961 (N_17961,N_11169,N_9080);
nand U17962 (N_17962,N_6341,N_8345);
xor U17963 (N_17963,N_11185,N_9902);
or U17964 (N_17964,N_7396,N_7351);
nor U17965 (N_17965,N_7657,N_6917);
nand U17966 (N_17966,N_8141,N_11406);
nand U17967 (N_17967,N_8502,N_11410);
and U17968 (N_17968,N_9665,N_8328);
or U17969 (N_17969,N_11967,N_11805);
and U17970 (N_17970,N_6311,N_8293);
xnor U17971 (N_17971,N_8925,N_10215);
xor U17972 (N_17972,N_9425,N_8722);
xor U17973 (N_17973,N_11094,N_9463);
nor U17974 (N_17974,N_9026,N_7293);
nor U17975 (N_17975,N_11443,N_6836);
and U17976 (N_17976,N_11622,N_10793);
nor U17977 (N_17977,N_8065,N_11665);
nor U17978 (N_17978,N_11222,N_11473);
and U17979 (N_17979,N_8483,N_7666);
or U17980 (N_17980,N_11959,N_10830);
xor U17981 (N_17981,N_12370,N_9782);
nor U17982 (N_17982,N_10812,N_7701);
and U17983 (N_17983,N_10392,N_6901);
and U17984 (N_17984,N_11467,N_9340);
xor U17985 (N_17985,N_10011,N_9118);
nor U17986 (N_17986,N_8767,N_10452);
nand U17987 (N_17987,N_9025,N_6946);
and U17988 (N_17988,N_6786,N_8414);
nor U17989 (N_17989,N_10670,N_10112);
or U17990 (N_17990,N_6670,N_9852);
or U17991 (N_17991,N_9513,N_11254);
xor U17992 (N_17992,N_7382,N_8721);
nor U17993 (N_17993,N_6269,N_6704);
nor U17994 (N_17994,N_8411,N_11405);
nor U17995 (N_17995,N_10071,N_8928);
nor U17996 (N_17996,N_7962,N_7043);
nand U17997 (N_17997,N_7745,N_10711);
or U17998 (N_17998,N_6661,N_9262);
and U17999 (N_17999,N_11705,N_7372);
or U18000 (N_18000,N_7402,N_8706);
or U18001 (N_18001,N_10934,N_10801);
nand U18002 (N_18002,N_10411,N_7456);
nand U18003 (N_18003,N_11026,N_12301);
or U18004 (N_18004,N_9319,N_8301);
and U18005 (N_18005,N_8106,N_8183);
xnor U18006 (N_18006,N_9922,N_8824);
and U18007 (N_18007,N_11319,N_7534);
and U18008 (N_18008,N_11390,N_10231);
xnor U18009 (N_18009,N_11725,N_11019);
and U18010 (N_18010,N_8665,N_9479);
nor U18011 (N_18011,N_7144,N_7519);
and U18012 (N_18012,N_12083,N_9570);
xnor U18013 (N_18013,N_6682,N_9723);
nor U18014 (N_18014,N_7002,N_8101);
and U18015 (N_18015,N_11222,N_7347);
nand U18016 (N_18016,N_11547,N_8434);
xor U18017 (N_18017,N_9926,N_7995);
xor U18018 (N_18018,N_7042,N_6914);
nor U18019 (N_18019,N_6409,N_10339);
nand U18020 (N_18020,N_6295,N_8682);
nor U18021 (N_18021,N_7185,N_10393);
xor U18022 (N_18022,N_11842,N_8191);
nand U18023 (N_18023,N_10517,N_11269);
nand U18024 (N_18024,N_9714,N_9141);
and U18025 (N_18025,N_7779,N_8272);
nor U18026 (N_18026,N_12378,N_7398);
xnor U18027 (N_18027,N_10363,N_8416);
xor U18028 (N_18028,N_10904,N_11834);
or U18029 (N_18029,N_7723,N_10860);
nand U18030 (N_18030,N_11144,N_7763);
and U18031 (N_18031,N_7515,N_10339);
or U18032 (N_18032,N_8431,N_10716);
xor U18033 (N_18033,N_12493,N_11648);
nand U18034 (N_18034,N_10170,N_9312);
and U18035 (N_18035,N_9383,N_9525);
and U18036 (N_18036,N_12110,N_10740);
and U18037 (N_18037,N_6706,N_8058);
nor U18038 (N_18038,N_11090,N_12091);
nor U18039 (N_18039,N_11386,N_11952);
and U18040 (N_18040,N_10093,N_10328);
nand U18041 (N_18041,N_11131,N_11281);
nor U18042 (N_18042,N_9575,N_6778);
and U18043 (N_18043,N_8561,N_11562);
and U18044 (N_18044,N_12041,N_9045);
nor U18045 (N_18045,N_10999,N_11573);
or U18046 (N_18046,N_7117,N_10308);
nand U18047 (N_18047,N_6436,N_6458);
or U18048 (N_18048,N_8520,N_7810);
and U18049 (N_18049,N_8085,N_7494);
nand U18050 (N_18050,N_8420,N_9355);
nand U18051 (N_18051,N_6591,N_9250);
nor U18052 (N_18052,N_9123,N_9274);
and U18053 (N_18053,N_7259,N_6885);
nor U18054 (N_18054,N_10794,N_8976);
xor U18055 (N_18055,N_6308,N_9433);
or U18056 (N_18056,N_7386,N_11859);
and U18057 (N_18057,N_12240,N_7625);
nor U18058 (N_18058,N_6579,N_10606);
nor U18059 (N_18059,N_9372,N_10746);
and U18060 (N_18060,N_7027,N_11783);
and U18061 (N_18061,N_10739,N_7062);
nor U18062 (N_18062,N_7996,N_9395);
nor U18063 (N_18063,N_7797,N_8910);
and U18064 (N_18064,N_11258,N_11181);
or U18065 (N_18065,N_6671,N_7830);
and U18066 (N_18066,N_7696,N_12120);
xnor U18067 (N_18067,N_9560,N_8585);
or U18068 (N_18068,N_11699,N_9539);
nand U18069 (N_18069,N_7931,N_11888);
nand U18070 (N_18070,N_6449,N_7634);
and U18071 (N_18071,N_8698,N_11613);
and U18072 (N_18072,N_12189,N_7479);
nor U18073 (N_18073,N_6369,N_7099);
nor U18074 (N_18074,N_9600,N_11819);
nand U18075 (N_18075,N_8606,N_9865);
nand U18076 (N_18076,N_10803,N_11860);
or U18077 (N_18077,N_11474,N_10383);
nor U18078 (N_18078,N_11993,N_11106);
nand U18079 (N_18079,N_9605,N_10298);
and U18080 (N_18080,N_9200,N_12208);
xnor U18081 (N_18081,N_11684,N_9214);
xor U18082 (N_18082,N_11428,N_7149);
xnor U18083 (N_18083,N_7114,N_9585);
xor U18084 (N_18084,N_11157,N_7744);
xor U18085 (N_18085,N_9861,N_10655);
xnor U18086 (N_18086,N_8093,N_9102);
nor U18087 (N_18087,N_11397,N_12118);
nand U18088 (N_18088,N_8053,N_9919);
or U18089 (N_18089,N_12411,N_7236);
nor U18090 (N_18090,N_11010,N_9004);
or U18091 (N_18091,N_10738,N_7188);
xnor U18092 (N_18092,N_11261,N_9241);
nand U18093 (N_18093,N_11024,N_7062);
and U18094 (N_18094,N_8761,N_7874);
and U18095 (N_18095,N_10082,N_10778);
and U18096 (N_18096,N_8947,N_11254);
xnor U18097 (N_18097,N_12204,N_10829);
nand U18098 (N_18098,N_11418,N_10970);
nand U18099 (N_18099,N_7274,N_9429);
nand U18100 (N_18100,N_8284,N_8256);
and U18101 (N_18101,N_8042,N_10477);
xor U18102 (N_18102,N_11404,N_8082);
xnor U18103 (N_18103,N_10494,N_10458);
nand U18104 (N_18104,N_8443,N_6953);
and U18105 (N_18105,N_7152,N_10999);
or U18106 (N_18106,N_7088,N_11138);
nor U18107 (N_18107,N_11487,N_10886);
nand U18108 (N_18108,N_7266,N_6510);
and U18109 (N_18109,N_9641,N_6588);
or U18110 (N_18110,N_10387,N_9002);
and U18111 (N_18111,N_6482,N_7146);
and U18112 (N_18112,N_7356,N_12038);
and U18113 (N_18113,N_9469,N_10036);
and U18114 (N_18114,N_7085,N_7599);
nand U18115 (N_18115,N_9639,N_8629);
nand U18116 (N_18116,N_11920,N_9293);
xnor U18117 (N_18117,N_9426,N_7246);
and U18118 (N_18118,N_6265,N_7924);
xnor U18119 (N_18119,N_6291,N_11342);
or U18120 (N_18120,N_9478,N_10503);
or U18121 (N_18121,N_11258,N_11349);
nor U18122 (N_18122,N_7634,N_10480);
and U18123 (N_18123,N_11058,N_7174);
xor U18124 (N_18124,N_6331,N_11920);
xnor U18125 (N_18125,N_11461,N_10907);
xnor U18126 (N_18126,N_7804,N_12257);
or U18127 (N_18127,N_7795,N_10350);
or U18128 (N_18128,N_8050,N_9567);
nand U18129 (N_18129,N_12183,N_7166);
nor U18130 (N_18130,N_8686,N_7181);
xor U18131 (N_18131,N_8963,N_10363);
nand U18132 (N_18132,N_6979,N_11235);
nand U18133 (N_18133,N_10695,N_11730);
or U18134 (N_18134,N_6804,N_9084);
nor U18135 (N_18135,N_8624,N_11610);
xor U18136 (N_18136,N_8975,N_8045);
and U18137 (N_18137,N_8685,N_11710);
xor U18138 (N_18138,N_6873,N_12140);
or U18139 (N_18139,N_6258,N_10473);
nand U18140 (N_18140,N_11146,N_11773);
and U18141 (N_18141,N_8943,N_11829);
nor U18142 (N_18142,N_9450,N_7479);
and U18143 (N_18143,N_8118,N_12495);
xnor U18144 (N_18144,N_7245,N_7967);
nand U18145 (N_18145,N_11621,N_7237);
xor U18146 (N_18146,N_6517,N_6562);
and U18147 (N_18147,N_9446,N_11243);
xor U18148 (N_18148,N_9775,N_8841);
and U18149 (N_18149,N_10279,N_12399);
nand U18150 (N_18150,N_9009,N_7624);
nor U18151 (N_18151,N_8317,N_7680);
nand U18152 (N_18152,N_6798,N_10985);
or U18153 (N_18153,N_10667,N_9443);
and U18154 (N_18154,N_10175,N_6631);
nand U18155 (N_18155,N_10456,N_10553);
xor U18156 (N_18156,N_8024,N_9507);
nand U18157 (N_18157,N_11182,N_8621);
xnor U18158 (N_18158,N_12031,N_7849);
and U18159 (N_18159,N_9505,N_10494);
xor U18160 (N_18160,N_8410,N_6598);
nand U18161 (N_18161,N_9566,N_11573);
nor U18162 (N_18162,N_8789,N_11578);
xor U18163 (N_18163,N_9461,N_11141);
nor U18164 (N_18164,N_9558,N_12262);
nand U18165 (N_18165,N_10659,N_11153);
or U18166 (N_18166,N_12429,N_9192);
nor U18167 (N_18167,N_8495,N_10691);
nand U18168 (N_18168,N_6266,N_11074);
nor U18169 (N_18169,N_7806,N_9720);
nand U18170 (N_18170,N_11682,N_9635);
xnor U18171 (N_18171,N_12224,N_12142);
nand U18172 (N_18172,N_10410,N_8189);
and U18173 (N_18173,N_6612,N_12074);
or U18174 (N_18174,N_11798,N_7160);
nor U18175 (N_18175,N_11891,N_6666);
and U18176 (N_18176,N_8194,N_12136);
or U18177 (N_18177,N_9576,N_8121);
nor U18178 (N_18178,N_6284,N_11748);
xor U18179 (N_18179,N_7505,N_9454);
or U18180 (N_18180,N_11514,N_7515);
nor U18181 (N_18181,N_8770,N_11099);
and U18182 (N_18182,N_10743,N_9861);
nor U18183 (N_18183,N_11548,N_10563);
or U18184 (N_18184,N_7142,N_9952);
and U18185 (N_18185,N_7233,N_10819);
and U18186 (N_18186,N_8534,N_7731);
nor U18187 (N_18187,N_12432,N_10595);
and U18188 (N_18188,N_6878,N_8785);
or U18189 (N_18189,N_6460,N_7907);
or U18190 (N_18190,N_9118,N_6768);
nor U18191 (N_18191,N_12248,N_7338);
nor U18192 (N_18192,N_11607,N_9685);
xor U18193 (N_18193,N_12267,N_6394);
and U18194 (N_18194,N_8334,N_7902);
or U18195 (N_18195,N_9819,N_11541);
xnor U18196 (N_18196,N_9171,N_10737);
xnor U18197 (N_18197,N_7121,N_7816);
and U18198 (N_18198,N_7471,N_12446);
or U18199 (N_18199,N_8194,N_6588);
or U18200 (N_18200,N_8820,N_11727);
nand U18201 (N_18201,N_8282,N_9309);
xor U18202 (N_18202,N_12405,N_8372);
and U18203 (N_18203,N_8076,N_11837);
and U18204 (N_18204,N_11839,N_8693);
xor U18205 (N_18205,N_7077,N_7301);
nand U18206 (N_18206,N_10330,N_10718);
or U18207 (N_18207,N_9986,N_11331);
nor U18208 (N_18208,N_12096,N_11478);
nand U18209 (N_18209,N_8080,N_10692);
nor U18210 (N_18210,N_6556,N_10263);
or U18211 (N_18211,N_7711,N_11075);
and U18212 (N_18212,N_9485,N_10020);
xor U18213 (N_18213,N_7433,N_8540);
nor U18214 (N_18214,N_12043,N_12035);
and U18215 (N_18215,N_9238,N_8514);
and U18216 (N_18216,N_8836,N_10738);
or U18217 (N_18217,N_7455,N_9071);
and U18218 (N_18218,N_8875,N_9827);
and U18219 (N_18219,N_10455,N_6275);
nor U18220 (N_18220,N_8788,N_11999);
and U18221 (N_18221,N_10334,N_12112);
and U18222 (N_18222,N_9217,N_8205);
and U18223 (N_18223,N_7023,N_12227);
nand U18224 (N_18224,N_7803,N_8984);
and U18225 (N_18225,N_11309,N_11629);
xor U18226 (N_18226,N_8562,N_9505);
nand U18227 (N_18227,N_6530,N_8399);
or U18228 (N_18228,N_10492,N_7061);
or U18229 (N_18229,N_7962,N_11977);
nor U18230 (N_18230,N_6443,N_10932);
or U18231 (N_18231,N_8158,N_7604);
or U18232 (N_18232,N_7892,N_9988);
nor U18233 (N_18233,N_10690,N_11343);
nor U18234 (N_18234,N_11270,N_11006);
or U18235 (N_18235,N_11258,N_11774);
and U18236 (N_18236,N_8403,N_9684);
or U18237 (N_18237,N_7141,N_12376);
and U18238 (N_18238,N_8284,N_12370);
nor U18239 (N_18239,N_8336,N_8004);
nand U18240 (N_18240,N_10372,N_12413);
nand U18241 (N_18241,N_7144,N_8027);
nand U18242 (N_18242,N_11679,N_8524);
and U18243 (N_18243,N_8363,N_7584);
nor U18244 (N_18244,N_6712,N_9286);
or U18245 (N_18245,N_12309,N_8105);
and U18246 (N_18246,N_12247,N_7001);
and U18247 (N_18247,N_7920,N_10775);
nand U18248 (N_18248,N_12380,N_6644);
or U18249 (N_18249,N_8601,N_10473);
nand U18250 (N_18250,N_6691,N_11015);
xnor U18251 (N_18251,N_10411,N_11391);
nor U18252 (N_18252,N_6749,N_7026);
and U18253 (N_18253,N_11483,N_9896);
and U18254 (N_18254,N_11895,N_10687);
nand U18255 (N_18255,N_8565,N_6437);
xor U18256 (N_18256,N_7572,N_7392);
nand U18257 (N_18257,N_10822,N_8134);
nand U18258 (N_18258,N_11479,N_11487);
xor U18259 (N_18259,N_6712,N_8697);
or U18260 (N_18260,N_10302,N_11841);
and U18261 (N_18261,N_10983,N_9432);
and U18262 (N_18262,N_6747,N_8144);
nor U18263 (N_18263,N_8146,N_12307);
and U18264 (N_18264,N_8132,N_10103);
or U18265 (N_18265,N_7446,N_7659);
xnor U18266 (N_18266,N_6425,N_7464);
and U18267 (N_18267,N_8184,N_10245);
or U18268 (N_18268,N_7337,N_10716);
nor U18269 (N_18269,N_11526,N_7648);
nand U18270 (N_18270,N_12142,N_7836);
or U18271 (N_18271,N_8057,N_9092);
nand U18272 (N_18272,N_7496,N_9253);
nand U18273 (N_18273,N_10425,N_12019);
or U18274 (N_18274,N_9109,N_9629);
nand U18275 (N_18275,N_8197,N_12429);
or U18276 (N_18276,N_10562,N_10191);
or U18277 (N_18277,N_8034,N_9415);
or U18278 (N_18278,N_6418,N_8068);
nor U18279 (N_18279,N_8328,N_8941);
and U18280 (N_18280,N_7469,N_7560);
xnor U18281 (N_18281,N_6835,N_9647);
nand U18282 (N_18282,N_9933,N_10662);
nand U18283 (N_18283,N_12216,N_7966);
or U18284 (N_18284,N_6942,N_10955);
or U18285 (N_18285,N_10803,N_8322);
nand U18286 (N_18286,N_10383,N_10393);
and U18287 (N_18287,N_6280,N_6633);
nor U18288 (N_18288,N_8176,N_7765);
and U18289 (N_18289,N_8287,N_12076);
xor U18290 (N_18290,N_10644,N_8205);
nor U18291 (N_18291,N_9307,N_7395);
nor U18292 (N_18292,N_12486,N_11978);
nor U18293 (N_18293,N_10892,N_12246);
nand U18294 (N_18294,N_11099,N_9413);
xnor U18295 (N_18295,N_7386,N_7481);
or U18296 (N_18296,N_11926,N_10326);
and U18297 (N_18297,N_8024,N_9890);
and U18298 (N_18298,N_8173,N_7118);
and U18299 (N_18299,N_11373,N_6839);
and U18300 (N_18300,N_9616,N_12142);
or U18301 (N_18301,N_6544,N_11856);
nand U18302 (N_18302,N_12018,N_10219);
nor U18303 (N_18303,N_10986,N_6833);
nand U18304 (N_18304,N_11411,N_9217);
or U18305 (N_18305,N_7886,N_10261);
or U18306 (N_18306,N_12382,N_9043);
nor U18307 (N_18307,N_12060,N_10228);
or U18308 (N_18308,N_8346,N_8193);
and U18309 (N_18309,N_6403,N_7611);
or U18310 (N_18310,N_6975,N_7143);
xor U18311 (N_18311,N_11600,N_11855);
xnor U18312 (N_18312,N_8624,N_10937);
xnor U18313 (N_18313,N_11377,N_12168);
or U18314 (N_18314,N_9009,N_9440);
and U18315 (N_18315,N_9623,N_7370);
xor U18316 (N_18316,N_10717,N_11004);
xor U18317 (N_18317,N_8377,N_6884);
nor U18318 (N_18318,N_6281,N_8028);
nand U18319 (N_18319,N_11806,N_7543);
xor U18320 (N_18320,N_8512,N_11226);
and U18321 (N_18321,N_9810,N_9874);
nor U18322 (N_18322,N_8019,N_8632);
nor U18323 (N_18323,N_7203,N_8314);
and U18324 (N_18324,N_10511,N_11653);
nand U18325 (N_18325,N_10021,N_8571);
and U18326 (N_18326,N_11920,N_6291);
and U18327 (N_18327,N_8197,N_6986);
nor U18328 (N_18328,N_9963,N_9038);
or U18329 (N_18329,N_8508,N_7119);
nand U18330 (N_18330,N_11394,N_9371);
xnor U18331 (N_18331,N_10028,N_12421);
xor U18332 (N_18332,N_12396,N_10279);
xnor U18333 (N_18333,N_7082,N_8811);
xnor U18334 (N_18334,N_11147,N_7982);
nor U18335 (N_18335,N_8800,N_7998);
and U18336 (N_18336,N_12489,N_11641);
nand U18337 (N_18337,N_8315,N_11110);
and U18338 (N_18338,N_10489,N_7518);
nand U18339 (N_18339,N_9907,N_8469);
and U18340 (N_18340,N_10684,N_11720);
xor U18341 (N_18341,N_9158,N_7545);
xor U18342 (N_18342,N_9862,N_8366);
or U18343 (N_18343,N_7333,N_11632);
or U18344 (N_18344,N_12044,N_10178);
and U18345 (N_18345,N_11997,N_7749);
and U18346 (N_18346,N_12476,N_6876);
xor U18347 (N_18347,N_6371,N_8673);
nand U18348 (N_18348,N_11656,N_9913);
nand U18349 (N_18349,N_7002,N_11617);
nand U18350 (N_18350,N_11187,N_6802);
or U18351 (N_18351,N_7115,N_9407);
and U18352 (N_18352,N_7122,N_9095);
nor U18353 (N_18353,N_10653,N_6595);
and U18354 (N_18354,N_10193,N_10036);
and U18355 (N_18355,N_10182,N_6499);
and U18356 (N_18356,N_8851,N_12139);
nand U18357 (N_18357,N_10224,N_6923);
xnor U18358 (N_18358,N_10370,N_6841);
or U18359 (N_18359,N_10438,N_11050);
nand U18360 (N_18360,N_12301,N_12425);
and U18361 (N_18361,N_7016,N_7431);
xor U18362 (N_18362,N_9123,N_8266);
nor U18363 (N_18363,N_9261,N_7870);
or U18364 (N_18364,N_10085,N_8451);
nand U18365 (N_18365,N_6292,N_10860);
nand U18366 (N_18366,N_7663,N_7778);
nor U18367 (N_18367,N_6479,N_8720);
and U18368 (N_18368,N_6998,N_9096);
and U18369 (N_18369,N_10215,N_9192);
and U18370 (N_18370,N_9184,N_7680);
and U18371 (N_18371,N_6917,N_7257);
xnor U18372 (N_18372,N_10541,N_10609);
and U18373 (N_18373,N_11828,N_7336);
or U18374 (N_18374,N_11093,N_9378);
nand U18375 (N_18375,N_8471,N_10070);
nor U18376 (N_18376,N_8824,N_7930);
and U18377 (N_18377,N_6302,N_7423);
nand U18378 (N_18378,N_7654,N_10036);
nand U18379 (N_18379,N_11943,N_8642);
nand U18380 (N_18380,N_9390,N_12327);
and U18381 (N_18381,N_11662,N_10812);
or U18382 (N_18382,N_7074,N_9909);
xnor U18383 (N_18383,N_9357,N_9624);
and U18384 (N_18384,N_9440,N_7204);
and U18385 (N_18385,N_11536,N_8125);
nor U18386 (N_18386,N_10491,N_11726);
and U18387 (N_18387,N_8553,N_7390);
nor U18388 (N_18388,N_11534,N_9386);
nor U18389 (N_18389,N_7479,N_11358);
nand U18390 (N_18390,N_7652,N_11758);
xor U18391 (N_18391,N_7906,N_12064);
nor U18392 (N_18392,N_10591,N_8631);
nor U18393 (N_18393,N_11197,N_9275);
nor U18394 (N_18394,N_10563,N_11998);
and U18395 (N_18395,N_9560,N_11538);
or U18396 (N_18396,N_8768,N_9402);
or U18397 (N_18397,N_12483,N_9197);
xnor U18398 (N_18398,N_8587,N_11643);
xor U18399 (N_18399,N_9587,N_6887);
nand U18400 (N_18400,N_9102,N_11612);
nor U18401 (N_18401,N_6998,N_10960);
nor U18402 (N_18402,N_9649,N_9924);
nand U18403 (N_18403,N_6453,N_10715);
xor U18404 (N_18404,N_12446,N_10128);
nor U18405 (N_18405,N_9180,N_7833);
or U18406 (N_18406,N_12108,N_9610);
or U18407 (N_18407,N_7504,N_7206);
and U18408 (N_18408,N_6652,N_7266);
nor U18409 (N_18409,N_7045,N_9520);
nand U18410 (N_18410,N_10477,N_10092);
nor U18411 (N_18411,N_8983,N_11873);
nor U18412 (N_18412,N_11008,N_8468);
and U18413 (N_18413,N_10680,N_6698);
xnor U18414 (N_18414,N_7407,N_10328);
nand U18415 (N_18415,N_11033,N_9832);
nor U18416 (N_18416,N_7541,N_9929);
nor U18417 (N_18417,N_7427,N_8043);
nand U18418 (N_18418,N_11987,N_11888);
nand U18419 (N_18419,N_9595,N_8785);
and U18420 (N_18420,N_10734,N_9082);
xnor U18421 (N_18421,N_11917,N_11617);
and U18422 (N_18422,N_9675,N_10121);
and U18423 (N_18423,N_10826,N_7709);
nor U18424 (N_18424,N_9586,N_12115);
or U18425 (N_18425,N_9527,N_9378);
and U18426 (N_18426,N_7419,N_11761);
or U18427 (N_18427,N_12071,N_12232);
xor U18428 (N_18428,N_8743,N_11003);
nor U18429 (N_18429,N_10489,N_11989);
and U18430 (N_18430,N_11402,N_10033);
xnor U18431 (N_18431,N_8466,N_11519);
or U18432 (N_18432,N_8804,N_7971);
nor U18433 (N_18433,N_7906,N_7091);
xor U18434 (N_18434,N_6669,N_12223);
nor U18435 (N_18435,N_8123,N_9778);
and U18436 (N_18436,N_6438,N_11960);
nor U18437 (N_18437,N_11585,N_7972);
nor U18438 (N_18438,N_10637,N_6460);
and U18439 (N_18439,N_6645,N_6984);
nand U18440 (N_18440,N_6996,N_12212);
xor U18441 (N_18441,N_7495,N_8143);
xnor U18442 (N_18442,N_10422,N_11113);
or U18443 (N_18443,N_11584,N_8980);
nor U18444 (N_18444,N_9485,N_10084);
xor U18445 (N_18445,N_11216,N_11005);
and U18446 (N_18446,N_11341,N_6501);
nand U18447 (N_18447,N_8602,N_8274);
and U18448 (N_18448,N_11987,N_12232);
xor U18449 (N_18449,N_11885,N_11064);
or U18450 (N_18450,N_9936,N_9184);
nor U18451 (N_18451,N_11175,N_9163);
nand U18452 (N_18452,N_11093,N_8770);
xor U18453 (N_18453,N_7395,N_10863);
and U18454 (N_18454,N_7687,N_7908);
nor U18455 (N_18455,N_11249,N_8068);
nand U18456 (N_18456,N_6425,N_7310);
nand U18457 (N_18457,N_6260,N_6335);
nor U18458 (N_18458,N_10419,N_7011);
nand U18459 (N_18459,N_11813,N_10644);
nor U18460 (N_18460,N_7639,N_9631);
and U18461 (N_18461,N_8944,N_6650);
nand U18462 (N_18462,N_7377,N_6535);
or U18463 (N_18463,N_11374,N_11583);
xnor U18464 (N_18464,N_10262,N_9706);
or U18465 (N_18465,N_9741,N_9734);
and U18466 (N_18466,N_7357,N_6466);
xor U18467 (N_18467,N_9436,N_6924);
nor U18468 (N_18468,N_10907,N_8047);
and U18469 (N_18469,N_6904,N_6427);
xor U18470 (N_18470,N_10367,N_9164);
nand U18471 (N_18471,N_6315,N_9922);
xor U18472 (N_18472,N_7619,N_8354);
or U18473 (N_18473,N_12207,N_6934);
xnor U18474 (N_18474,N_8297,N_8439);
or U18475 (N_18475,N_9304,N_8312);
nor U18476 (N_18476,N_8247,N_9656);
xor U18477 (N_18477,N_10400,N_11767);
xnor U18478 (N_18478,N_7288,N_11419);
xnor U18479 (N_18479,N_9324,N_6833);
and U18480 (N_18480,N_9800,N_7660);
nand U18481 (N_18481,N_6408,N_6744);
xor U18482 (N_18482,N_11796,N_10001);
xor U18483 (N_18483,N_12177,N_12446);
and U18484 (N_18484,N_6724,N_9734);
nor U18485 (N_18485,N_8372,N_9551);
nand U18486 (N_18486,N_11703,N_6581);
and U18487 (N_18487,N_11582,N_10678);
nor U18488 (N_18488,N_8003,N_9802);
nand U18489 (N_18489,N_10250,N_6927);
or U18490 (N_18490,N_6628,N_9599);
and U18491 (N_18491,N_6352,N_9923);
and U18492 (N_18492,N_8399,N_6332);
xnor U18493 (N_18493,N_9703,N_9366);
nand U18494 (N_18494,N_6945,N_10688);
nor U18495 (N_18495,N_11693,N_6376);
nand U18496 (N_18496,N_9551,N_6690);
nand U18497 (N_18497,N_9800,N_11247);
nand U18498 (N_18498,N_8087,N_8380);
and U18499 (N_18499,N_11914,N_12306);
xor U18500 (N_18500,N_11395,N_7838);
nand U18501 (N_18501,N_10899,N_10264);
xor U18502 (N_18502,N_10844,N_12200);
nand U18503 (N_18503,N_8346,N_6647);
nor U18504 (N_18504,N_10240,N_6631);
or U18505 (N_18505,N_11374,N_9644);
nand U18506 (N_18506,N_11364,N_11957);
and U18507 (N_18507,N_6789,N_7600);
and U18508 (N_18508,N_6331,N_9220);
xor U18509 (N_18509,N_8205,N_9840);
and U18510 (N_18510,N_8422,N_11979);
or U18511 (N_18511,N_7959,N_10523);
and U18512 (N_18512,N_7221,N_9360);
nand U18513 (N_18513,N_11237,N_9904);
nand U18514 (N_18514,N_11811,N_9319);
nand U18515 (N_18515,N_8745,N_6605);
or U18516 (N_18516,N_10321,N_12390);
xor U18517 (N_18517,N_11442,N_11956);
xor U18518 (N_18518,N_9905,N_7223);
and U18519 (N_18519,N_12222,N_9365);
nand U18520 (N_18520,N_8428,N_8855);
xnor U18521 (N_18521,N_6497,N_10192);
xnor U18522 (N_18522,N_7336,N_7395);
or U18523 (N_18523,N_7260,N_11577);
xnor U18524 (N_18524,N_10322,N_6786);
and U18525 (N_18525,N_11549,N_10867);
or U18526 (N_18526,N_8011,N_10426);
nand U18527 (N_18527,N_10262,N_7974);
or U18528 (N_18528,N_7653,N_10165);
nor U18529 (N_18529,N_9373,N_9742);
xor U18530 (N_18530,N_9532,N_9933);
or U18531 (N_18531,N_9395,N_9017);
xor U18532 (N_18532,N_12127,N_11318);
or U18533 (N_18533,N_9601,N_8278);
nor U18534 (N_18534,N_11010,N_8944);
nor U18535 (N_18535,N_11385,N_6586);
and U18536 (N_18536,N_6883,N_8323);
xor U18537 (N_18537,N_9244,N_11914);
nand U18538 (N_18538,N_6946,N_7323);
xor U18539 (N_18539,N_7127,N_11513);
xnor U18540 (N_18540,N_7247,N_9358);
or U18541 (N_18541,N_8776,N_10012);
xor U18542 (N_18542,N_8663,N_10238);
nor U18543 (N_18543,N_8377,N_11394);
or U18544 (N_18544,N_9466,N_10467);
nand U18545 (N_18545,N_10168,N_10310);
and U18546 (N_18546,N_10659,N_9541);
or U18547 (N_18547,N_11221,N_10191);
nor U18548 (N_18548,N_8808,N_6336);
nor U18549 (N_18549,N_11697,N_7361);
nor U18550 (N_18550,N_11355,N_8525);
nand U18551 (N_18551,N_11321,N_6633);
nand U18552 (N_18552,N_11336,N_6689);
xor U18553 (N_18553,N_10712,N_10657);
and U18554 (N_18554,N_7917,N_10156);
xor U18555 (N_18555,N_9802,N_7525);
or U18556 (N_18556,N_11536,N_7091);
xor U18557 (N_18557,N_7563,N_6809);
xor U18558 (N_18558,N_8274,N_10781);
nand U18559 (N_18559,N_11314,N_7035);
and U18560 (N_18560,N_6812,N_11610);
or U18561 (N_18561,N_7035,N_8768);
nor U18562 (N_18562,N_8731,N_6725);
nor U18563 (N_18563,N_7751,N_9949);
and U18564 (N_18564,N_10345,N_8700);
or U18565 (N_18565,N_6465,N_10472);
nand U18566 (N_18566,N_7387,N_10804);
nand U18567 (N_18567,N_7389,N_7288);
nand U18568 (N_18568,N_7704,N_6549);
xor U18569 (N_18569,N_8189,N_7863);
and U18570 (N_18570,N_10265,N_6376);
xor U18571 (N_18571,N_6957,N_6525);
nor U18572 (N_18572,N_11320,N_11620);
and U18573 (N_18573,N_9906,N_6864);
nor U18574 (N_18574,N_10696,N_12028);
xor U18575 (N_18575,N_7483,N_9129);
and U18576 (N_18576,N_9216,N_9565);
and U18577 (N_18577,N_11491,N_7318);
xnor U18578 (N_18578,N_7972,N_10454);
and U18579 (N_18579,N_6256,N_6634);
xnor U18580 (N_18580,N_9477,N_11643);
xor U18581 (N_18581,N_6516,N_11322);
nand U18582 (N_18582,N_12352,N_8105);
nand U18583 (N_18583,N_11806,N_11278);
nor U18584 (N_18584,N_11747,N_12003);
xnor U18585 (N_18585,N_8891,N_7931);
and U18586 (N_18586,N_8873,N_10661);
nor U18587 (N_18587,N_12004,N_7378);
or U18588 (N_18588,N_10232,N_11580);
nand U18589 (N_18589,N_12397,N_11756);
xor U18590 (N_18590,N_6714,N_10797);
and U18591 (N_18591,N_6351,N_8766);
nor U18592 (N_18592,N_11874,N_12488);
or U18593 (N_18593,N_10647,N_7140);
and U18594 (N_18594,N_11907,N_10684);
nand U18595 (N_18595,N_9223,N_10391);
or U18596 (N_18596,N_6829,N_12120);
nor U18597 (N_18597,N_8245,N_11703);
and U18598 (N_18598,N_11214,N_6972);
and U18599 (N_18599,N_9240,N_7289);
and U18600 (N_18600,N_11966,N_8028);
or U18601 (N_18601,N_8752,N_10635);
xor U18602 (N_18602,N_12428,N_6419);
and U18603 (N_18603,N_10679,N_8810);
or U18604 (N_18604,N_7231,N_10818);
nand U18605 (N_18605,N_8109,N_12005);
xnor U18606 (N_18606,N_11855,N_6715);
nor U18607 (N_18607,N_12152,N_9376);
nand U18608 (N_18608,N_9677,N_9381);
or U18609 (N_18609,N_10283,N_11379);
nand U18610 (N_18610,N_12477,N_10990);
nor U18611 (N_18611,N_8373,N_8161);
or U18612 (N_18612,N_10510,N_9335);
nand U18613 (N_18613,N_8761,N_9051);
or U18614 (N_18614,N_11143,N_7876);
nand U18615 (N_18615,N_11055,N_12041);
or U18616 (N_18616,N_12197,N_9450);
or U18617 (N_18617,N_10422,N_6628);
and U18618 (N_18618,N_12314,N_7356);
nor U18619 (N_18619,N_11006,N_12110);
xor U18620 (N_18620,N_9399,N_12015);
xnor U18621 (N_18621,N_9281,N_9030);
nor U18622 (N_18622,N_11453,N_7123);
or U18623 (N_18623,N_11777,N_6314);
nor U18624 (N_18624,N_6466,N_6925);
nand U18625 (N_18625,N_6279,N_7619);
nand U18626 (N_18626,N_9934,N_11592);
and U18627 (N_18627,N_7040,N_12389);
xnor U18628 (N_18628,N_6821,N_6362);
nor U18629 (N_18629,N_10471,N_11000);
or U18630 (N_18630,N_7689,N_10127);
or U18631 (N_18631,N_7625,N_11477);
nor U18632 (N_18632,N_7581,N_7210);
xnor U18633 (N_18633,N_9871,N_12076);
xnor U18634 (N_18634,N_10836,N_9494);
nand U18635 (N_18635,N_6414,N_11494);
or U18636 (N_18636,N_6846,N_11420);
or U18637 (N_18637,N_10884,N_12317);
or U18638 (N_18638,N_9496,N_10882);
or U18639 (N_18639,N_7535,N_6509);
nand U18640 (N_18640,N_9118,N_7100);
nand U18641 (N_18641,N_10652,N_10024);
and U18642 (N_18642,N_8103,N_9963);
nand U18643 (N_18643,N_12462,N_7144);
nand U18644 (N_18644,N_12121,N_6489);
or U18645 (N_18645,N_6658,N_7045);
or U18646 (N_18646,N_8997,N_10766);
nand U18647 (N_18647,N_7167,N_9669);
xnor U18648 (N_18648,N_7086,N_7652);
nor U18649 (N_18649,N_9891,N_8058);
or U18650 (N_18650,N_12122,N_11353);
or U18651 (N_18651,N_6762,N_9234);
xnor U18652 (N_18652,N_9474,N_8254);
nand U18653 (N_18653,N_10347,N_6839);
nor U18654 (N_18654,N_10248,N_8497);
or U18655 (N_18655,N_12341,N_6439);
and U18656 (N_18656,N_10018,N_10967);
and U18657 (N_18657,N_11175,N_10599);
or U18658 (N_18658,N_11838,N_8209);
or U18659 (N_18659,N_11892,N_6857);
xor U18660 (N_18660,N_8635,N_12291);
nor U18661 (N_18661,N_11358,N_12337);
or U18662 (N_18662,N_11961,N_9864);
nand U18663 (N_18663,N_6944,N_8453);
xor U18664 (N_18664,N_10933,N_6661);
nor U18665 (N_18665,N_9597,N_10608);
nand U18666 (N_18666,N_11885,N_6813);
or U18667 (N_18667,N_11191,N_8989);
and U18668 (N_18668,N_10694,N_11489);
or U18669 (N_18669,N_9043,N_10503);
nor U18670 (N_18670,N_9973,N_10507);
nand U18671 (N_18671,N_8817,N_8618);
and U18672 (N_18672,N_8579,N_8332);
or U18673 (N_18673,N_7046,N_8840);
xnor U18674 (N_18674,N_11246,N_7464);
and U18675 (N_18675,N_11816,N_6890);
nand U18676 (N_18676,N_9323,N_8206);
nand U18677 (N_18677,N_7887,N_7776);
nand U18678 (N_18678,N_8477,N_8037);
and U18679 (N_18679,N_11552,N_11013);
xor U18680 (N_18680,N_9349,N_9981);
xor U18681 (N_18681,N_8196,N_8871);
and U18682 (N_18682,N_8177,N_6591);
xor U18683 (N_18683,N_11617,N_7345);
nor U18684 (N_18684,N_10220,N_8031);
nor U18685 (N_18685,N_7095,N_7595);
or U18686 (N_18686,N_12108,N_11215);
nor U18687 (N_18687,N_12485,N_10084);
and U18688 (N_18688,N_10290,N_9141);
or U18689 (N_18689,N_8535,N_10772);
and U18690 (N_18690,N_10922,N_9856);
xor U18691 (N_18691,N_6846,N_7604);
nor U18692 (N_18692,N_6586,N_6805);
xnor U18693 (N_18693,N_11795,N_11679);
and U18694 (N_18694,N_9121,N_6288);
nand U18695 (N_18695,N_9251,N_9018);
or U18696 (N_18696,N_7547,N_9129);
or U18697 (N_18697,N_11714,N_8068);
and U18698 (N_18698,N_11448,N_6634);
or U18699 (N_18699,N_9802,N_7300);
nand U18700 (N_18700,N_7592,N_9449);
nor U18701 (N_18701,N_11600,N_7167);
xor U18702 (N_18702,N_10304,N_9686);
and U18703 (N_18703,N_8121,N_6251);
or U18704 (N_18704,N_6450,N_12232);
nand U18705 (N_18705,N_7556,N_12333);
xor U18706 (N_18706,N_7937,N_6709);
nand U18707 (N_18707,N_11855,N_9291);
xor U18708 (N_18708,N_8400,N_10447);
and U18709 (N_18709,N_9139,N_8408);
nand U18710 (N_18710,N_8602,N_6904);
and U18711 (N_18711,N_6950,N_11945);
xnor U18712 (N_18712,N_7980,N_12038);
nand U18713 (N_18713,N_7496,N_11584);
xor U18714 (N_18714,N_7824,N_10908);
nand U18715 (N_18715,N_8694,N_7212);
xor U18716 (N_18716,N_10541,N_6417);
and U18717 (N_18717,N_8068,N_7982);
xnor U18718 (N_18718,N_10976,N_7923);
or U18719 (N_18719,N_12187,N_10665);
nor U18720 (N_18720,N_9658,N_10365);
nor U18721 (N_18721,N_6636,N_11281);
nor U18722 (N_18722,N_10553,N_7012);
nand U18723 (N_18723,N_11014,N_12254);
nor U18724 (N_18724,N_11121,N_10968);
nand U18725 (N_18725,N_10373,N_6793);
or U18726 (N_18726,N_7960,N_10882);
nor U18727 (N_18727,N_8806,N_7892);
xor U18728 (N_18728,N_6743,N_8586);
and U18729 (N_18729,N_11335,N_11458);
xnor U18730 (N_18730,N_6427,N_6491);
or U18731 (N_18731,N_11720,N_6433);
nand U18732 (N_18732,N_9780,N_10184);
xor U18733 (N_18733,N_9046,N_12284);
or U18734 (N_18734,N_8614,N_12138);
and U18735 (N_18735,N_11141,N_9113);
and U18736 (N_18736,N_7546,N_10814);
nand U18737 (N_18737,N_11438,N_12273);
xnor U18738 (N_18738,N_9446,N_6926);
nor U18739 (N_18739,N_12106,N_11707);
or U18740 (N_18740,N_6421,N_6736);
nor U18741 (N_18741,N_8410,N_12260);
xor U18742 (N_18742,N_11268,N_12445);
xor U18743 (N_18743,N_9837,N_10890);
nor U18744 (N_18744,N_6940,N_7784);
or U18745 (N_18745,N_10190,N_12072);
nand U18746 (N_18746,N_11660,N_9139);
nand U18747 (N_18747,N_8229,N_7403);
or U18748 (N_18748,N_11179,N_9653);
or U18749 (N_18749,N_9167,N_12013);
or U18750 (N_18750,N_14362,N_12526);
and U18751 (N_18751,N_14751,N_17386);
or U18752 (N_18752,N_17606,N_14237);
nor U18753 (N_18753,N_16868,N_18426);
or U18754 (N_18754,N_14700,N_13306);
or U18755 (N_18755,N_15359,N_13100);
and U18756 (N_18756,N_16448,N_16812);
and U18757 (N_18757,N_17112,N_12887);
xor U18758 (N_18758,N_16871,N_15811);
and U18759 (N_18759,N_14696,N_18502);
or U18760 (N_18760,N_16381,N_16627);
nor U18761 (N_18761,N_16637,N_14518);
or U18762 (N_18762,N_13071,N_13632);
nand U18763 (N_18763,N_14243,N_15458);
nor U18764 (N_18764,N_18718,N_15639);
and U18765 (N_18765,N_14428,N_16929);
nand U18766 (N_18766,N_16853,N_17149);
and U18767 (N_18767,N_16006,N_14635);
and U18768 (N_18768,N_13359,N_16992);
nand U18769 (N_18769,N_17559,N_14994);
nor U18770 (N_18770,N_17587,N_17888);
nand U18771 (N_18771,N_18419,N_16898);
nand U18772 (N_18772,N_16553,N_12723);
nor U18773 (N_18773,N_14594,N_18545);
or U18774 (N_18774,N_14065,N_13085);
or U18775 (N_18775,N_17098,N_12966);
nor U18776 (N_18776,N_16796,N_18164);
xnor U18777 (N_18777,N_14936,N_17398);
xnor U18778 (N_18778,N_14271,N_14888);
and U18779 (N_18779,N_13491,N_18346);
and U18780 (N_18780,N_12873,N_18146);
or U18781 (N_18781,N_13504,N_13444);
and U18782 (N_18782,N_14231,N_13410);
nand U18783 (N_18783,N_16009,N_15554);
and U18784 (N_18784,N_15970,N_12758);
nor U18785 (N_18785,N_16767,N_14443);
nor U18786 (N_18786,N_15613,N_18012);
nand U18787 (N_18787,N_18403,N_16007);
or U18788 (N_18788,N_14970,N_13351);
nand U18789 (N_18789,N_14665,N_17582);
and U18790 (N_18790,N_18723,N_17927);
or U18791 (N_18791,N_12619,N_17315);
nand U18792 (N_18792,N_14124,N_18647);
nor U18793 (N_18793,N_15306,N_17567);
or U18794 (N_18794,N_15745,N_16499);
nand U18795 (N_18795,N_15752,N_18032);
nand U18796 (N_18796,N_17783,N_15495);
nand U18797 (N_18797,N_18575,N_15247);
or U18798 (N_18798,N_15427,N_12883);
nand U18799 (N_18799,N_13517,N_14430);
or U18800 (N_18800,N_14293,N_14456);
or U18801 (N_18801,N_13304,N_15885);
nor U18802 (N_18802,N_15942,N_16192);
nor U18803 (N_18803,N_18680,N_15606);
or U18804 (N_18804,N_15575,N_12964);
or U18805 (N_18805,N_17084,N_13553);
nor U18806 (N_18806,N_18183,N_17866);
xnor U18807 (N_18807,N_16800,N_14611);
and U18808 (N_18808,N_16822,N_13542);
nor U18809 (N_18809,N_13857,N_13484);
xor U18810 (N_18810,N_14176,N_13299);
and U18811 (N_18811,N_18058,N_17823);
nand U18812 (N_18812,N_14402,N_12598);
nor U18813 (N_18813,N_15157,N_18186);
or U18814 (N_18814,N_18100,N_12869);
xor U18815 (N_18815,N_12886,N_17312);
and U18816 (N_18816,N_16799,N_13640);
xnor U18817 (N_18817,N_12673,N_15461);
and U18818 (N_18818,N_15532,N_18658);
nor U18819 (N_18819,N_16075,N_16453);
nand U18820 (N_18820,N_17057,N_15605);
or U18821 (N_18821,N_15374,N_16820);
nand U18822 (N_18822,N_13250,N_15007);
nor U18823 (N_18823,N_17397,N_15878);
nand U18824 (N_18824,N_12581,N_16556);
nand U18825 (N_18825,N_15103,N_16559);
xor U18826 (N_18826,N_14960,N_16769);
nand U18827 (N_18827,N_16420,N_13683);
and U18828 (N_18828,N_18141,N_18537);
and U18829 (N_18829,N_16116,N_15210);
and U18830 (N_18830,N_17467,N_13841);
xor U18831 (N_18831,N_18224,N_17183);
nor U18832 (N_18832,N_15073,N_17611);
xor U18833 (N_18833,N_14731,N_14777);
nor U18834 (N_18834,N_13199,N_18685);
nor U18835 (N_18835,N_17486,N_16078);
and U18836 (N_18836,N_13988,N_14395);
and U18837 (N_18837,N_16176,N_15229);
or U18838 (N_18838,N_18061,N_16137);
and U18839 (N_18839,N_12753,N_16304);
xor U18840 (N_18840,N_17735,N_15350);
and U18841 (N_18841,N_17694,N_16832);
nand U18842 (N_18842,N_17409,N_16488);
xor U18843 (N_18843,N_16412,N_13004);
and U18844 (N_18844,N_13602,N_17920);
and U18845 (N_18845,N_15760,N_16484);
or U18846 (N_18846,N_16353,N_15650);
nor U18847 (N_18847,N_18678,N_18454);
or U18848 (N_18848,N_13577,N_17181);
and U18849 (N_18849,N_17480,N_13617);
nor U18850 (N_18850,N_16002,N_18399);
nor U18851 (N_18851,N_16883,N_15573);
xnor U18852 (N_18852,N_16524,N_15330);
or U18853 (N_18853,N_17333,N_14501);
xor U18854 (N_18854,N_16170,N_18359);
and U18855 (N_18855,N_16459,N_15382);
nand U18856 (N_18856,N_15317,N_14873);
or U18857 (N_18857,N_13293,N_18579);
and U18858 (N_18858,N_17995,N_17302);
or U18859 (N_18859,N_18083,N_13619);
or U18860 (N_18860,N_12669,N_14965);
nor U18861 (N_18861,N_12617,N_14471);
or U18862 (N_18862,N_17919,N_17516);
xor U18863 (N_18863,N_18079,N_16561);
and U18864 (N_18864,N_16461,N_16259);
xnor U18865 (N_18865,N_16810,N_13018);
or U18866 (N_18866,N_13819,N_18089);
or U18867 (N_18867,N_13978,N_16286);
nand U18868 (N_18868,N_18425,N_12672);
xnor U18869 (N_18869,N_13702,N_17107);
nor U18870 (N_18870,N_17330,N_13360);
nand U18871 (N_18871,N_16254,N_13618);
nand U18872 (N_18872,N_16631,N_18651);
nor U18873 (N_18873,N_18595,N_18740);
and U18874 (N_18874,N_16411,N_18090);
nor U18875 (N_18875,N_14669,N_16380);
nand U18876 (N_18876,N_13987,N_12709);
nand U18877 (N_18877,N_12501,N_16384);
nand U18878 (N_18878,N_15067,N_18182);
nand U18879 (N_18879,N_18603,N_14596);
nor U18880 (N_18880,N_16342,N_16869);
nand U18881 (N_18881,N_14793,N_14730);
or U18882 (N_18882,N_14376,N_17325);
nor U18883 (N_18883,N_13685,N_14300);
nor U18884 (N_18884,N_12659,N_16118);
xnor U18885 (N_18885,N_16602,N_12848);
nor U18886 (N_18886,N_13662,N_16709);
nor U18887 (N_18887,N_15984,N_13035);
nor U18888 (N_18888,N_12818,N_15328);
nor U18889 (N_18889,N_14804,N_14502);
and U18890 (N_18890,N_14150,N_17817);
nand U18891 (N_18891,N_17187,N_18179);
xor U18892 (N_18892,N_14286,N_13172);
nand U18893 (N_18893,N_17004,N_17189);
or U18894 (N_18894,N_14759,N_18366);
xor U18895 (N_18895,N_12916,N_17431);
and U18896 (N_18896,N_15720,N_15355);
nand U18897 (N_18897,N_14931,N_18457);
nor U18898 (N_18898,N_13733,N_17420);
nand U18899 (N_18899,N_17136,N_12509);
nand U18900 (N_18900,N_17083,N_14976);
xnor U18901 (N_18901,N_13198,N_14012);
xor U18902 (N_18902,N_13358,N_12529);
nand U18903 (N_18903,N_13333,N_12732);
nand U18904 (N_18904,N_14290,N_14741);
nand U18905 (N_18905,N_13060,N_13160);
xnor U18906 (N_18906,N_14424,N_16968);
nor U18907 (N_18907,N_15657,N_14263);
xor U18908 (N_18908,N_16379,N_14439);
nand U18909 (N_18909,N_16344,N_17827);
nor U18910 (N_18910,N_13276,N_16861);
nor U18911 (N_18911,N_17212,N_17160);
nand U18912 (N_18912,N_17166,N_13411);
nor U18913 (N_18913,N_16201,N_17127);
nor U18914 (N_18914,N_15365,N_15938);
or U18915 (N_18915,N_13891,N_15814);
nand U18916 (N_18916,N_14188,N_17544);
nor U18917 (N_18917,N_17028,N_17380);
and U18918 (N_18918,N_14824,N_15510);
nor U18919 (N_18919,N_13243,N_14305);
or U18920 (N_18920,N_18267,N_17791);
and U18921 (N_18921,N_18035,N_13835);
nand U18922 (N_18922,N_15663,N_16945);
xnor U18923 (N_18923,N_15221,N_18644);
nor U18924 (N_18924,N_17433,N_14229);
or U18925 (N_18925,N_18463,N_14423);
xor U18926 (N_18926,N_13000,N_15478);
or U18927 (N_18927,N_16248,N_13213);
xnor U18928 (N_18928,N_18563,N_17840);
nor U18929 (N_18929,N_12637,N_13500);
and U18930 (N_18930,N_16733,N_17048);
or U18931 (N_18931,N_12780,N_16977);
and U18932 (N_18932,N_16786,N_15957);
nor U18933 (N_18933,N_14584,N_17293);
nor U18934 (N_18934,N_14863,N_13335);
or U18935 (N_18935,N_14767,N_15160);
and U18936 (N_18936,N_17077,N_16635);
or U18937 (N_18937,N_17358,N_14809);
xor U18938 (N_18938,N_12696,N_15578);
or U18939 (N_18939,N_15834,N_15245);
and U18940 (N_18940,N_14509,N_14327);
nand U18941 (N_18941,N_16910,N_17422);
and U18942 (N_18942,N_14394,N_16538);
or U18943 (N_18943,N_17319,N_15806);
and U18944 (N_18944,N_17764,N_17718);
and U18945 (N_18945,N_13057,N_13945);
nor U18946 (N_18946,N_15545,N_16785);
nor U18947 (N_18947,N_17507,N_14850);
or U18948 (N_18948,N_13415,N_13046);
xor U18949 (N_18949,N_17378,N_16697);
nand U18950 (N_18950,N_12969,N_13793);
nand U18951 (N_18951,N_15493,N_13759);
and U18952 (N_18952,N_13762,N_18652);
nor U18953 (N_18953,N_15552,N_15920);
nor U18954 (N_18954,N_13191,N_13708);
nand U18955 (N_18955,N_13093,N_12502);
nor U18956 (N_18956,N_16748,N_16143);
or U18957 (N_18957,N_15633,N_17739);
and U18958 (N_18958,N_13461,N_18532);
and U18959 (N_18959,N_13775,N_17591);
xnor U18960 (N_18960,N_18187,N_14486);
nor U18961 (N_18961,N_13322,N_16497);
nor U18962 (N_18962,N_17273,N_15271);
or U18963 (N_18963,N_14952,N_12958);
or U18964 (N_18964,N_12524,N_16416);
and U18965 (N_18965,N_15025,N_15909);
xnor U18966 (N_18966,N_14590,N_13173);
and U18967 (N_18967,N_14384,N_17931);
nand U18968 (N_18968,N_13760,N_17584);
xor U18969 (N_18969,N_17229,N_16566);
and U18970 (N_18970,N_17942,N_15836);
nor U18971 (N_18971,N_13494,N_12639);
xnor U18972 (N_18972,N_17894,N_13611);
xnor U18973 (N_18973,N_16189,N_17184);
and U18974 (N_18974,N_13952,N_15860);
xnor U18975 (N_18975,N_15127,N_17432);
nor U18976 (N_18976,N_17052,N_14740);
xnor U18977 (N_18977,N_15068,N_15793);
xor U18978 (N_18978,N_14993,N_17944);
nor U18979 (N_18979,N_14179,N_12892);
nand U18980 (N_18980,N_12870,N_17326);
or U18981 (N_18981,N_17613,N_12534);
and U18982 (N_18982,N_15170,N_13590);
nor U18983 (N_18983,N_17768,N_14745);
or U18984 (N_18984,N_13209,N_17279);
nor U18985 (N_18985,N_17088,N_13256);
xnor U18986 (N_18986,N_18594,N_18275);
nor U18987 (N_18987,N_16105,N_16323);
and U18988 (N_18988,N_14997,N_14680);
and U18989 (N_18989,N_13859,N_14151);
xor U18990 (N_18990,N_17993,N_12629);
and U18991 (N_18991,N_16519,N_16866);
or U18992 (N_18992,N_12535,N_18263);
or U18993 (N_18993,N_14504,N_15916);
nand U18994 (N_18994,N_16848,N_15612);
or U18995 (N_18995,N_15230,N_16843);
and U18996 (N_18996,N_14879,N_16354);
nor U18997 (N_18997,N_15096,N_17214);
nand U18998 (N_18998,N_17970,N_15727);
nand U18999 (N_18999,N_15396,N_16090);
nor U19000 (N_19000,N_17691,N_15693);
or U19001 (N_19001,N_14815,N_14910);
and U19002 (N_19002,N_13439,N_15313);
xnor U19003 (N_19003,N_15826,N_15665);
nand U19004 (N_19004,N_12574,N_14415);
or U19005 (N_19005,N_14120,N_17956);
nand U19006 (N_19006,N_16443,N_14215);
xor U19007 (N_19007,N_14771,N_13750);
nor U19008 (N_19008,N_17301,N_17294);
nor U19009 (N_19009,N_15481,N_15700);
xor U19010 (N_19010,N_12541,N_13200);
or U19011 (N_19011,N_16134,N_15407);
and U19012 (N_19012,N_14410,N_16725);
xor U19013 (N_19013,N_14147,N_18496);
nand U19014 (N_19014,N_17755,N_17177);
xnor U19015 (N_19015,N_12936,N_13377);
nor U19016 (N_19016,N_18735,N_16204);
nand U19017 (N_19017,N_15069,N_15879);
nand U19018 (N_19018,N_12606,N_15258);
and U19019 (N_19019,N_13378,N_13706);
and U19020 (N_19020,N_14014,N_14512);
nor U19021 (N_19021,N_12905,N_13932);
xor U19022 (N_19022,N_18121,N_16974);
nor U19023 (N_19023,N_12897,N_17001);
nor U19024 (N_19024,N_15858,N_13551);
and U19025 (N_19025,N_15873,N_16964);
nor U19026 (N_19026,N_13823,N_18060);
nand U19027 (N_19027,N_15415,N_14346);
or U19028 (N_19028,N_17759,N_15467);
or U19029 (N_19029,N_16067,N_15505);
nand U19030 (N_19030,N_13274,N_15712);
nor U19031 (N_19031,N_14081,N_15882);
nor U19032 (N_19032,N_15747,N_16915);
and U19033 (N_19033,N_15804,N_13671);
nand U19034 (N_19034,N_16984,N_14906);
nand U19035 (N_19035,N_17494,N_15586);
nand U19036 (N_19036,N_18296,N_13156);
xnor U19037 (N_19037,N_16364,N_15234);
nor U19038 (N_19038,N_17223,N_15810);
nand U19039 (N_19039,N_16880,N_14102);
or U19040 (N_19040,N_14732,N_18327);
or U19041 (N_19041,N_13755,N_13223);
xor U19042 (N_19042,N_15244,N_12851);
xor U19043 (N_19043,N_16195,N_14046);
or U19044 (N_19044,N_13300,N_17983);
nand U19045 (N_19045,N_17437,N_18382);
xor U19046 (N_19046,N_17161,N_14608);
or U19047 (N_19047,N_17634,N_13538);
nand U19048 (N_19048,N_18731,N_17858);
or U19049 (N_19049,N_16670,N_14725);
xnor U19050 (N_19050,N_17720,N_16892);
and U19051 (N_19051,N_14870,N_14989);
nand U19052 (N_19052,N_17206,N_14978);
nand U19053 (N_19053,N_15162,N_17207);
or U19054 (N_19054,N_16493,N_14605);
and U19055 (N_19055,N_17816,N_14691);
nand U19056 (N_19056,N_14945,N_18042);
nor U19057 (N_19057,N_17317,N_17309);
nand U19058 (N_19058,N_13935,N_15490);
nand U19059 (N_19059,N_16473,N_14564);
nand U19060 (N_19060,N_14198,N_15807);
nor U19061 (N_19061,N_16302,N_13397);
and U19062 (N_19062,N_14056,N_17771);
nor U19063 (N_19063,N_15156,N_13711);
or U19064 (N_19064,N_17953,N_17255);
nand U19065 (N_19065,N_18004,N_17965);
nand U19066 (N_19066,N_13134,N_18041);
xor U19067 (N_19067,N_12847,N_17449);
and U19068 (N_19068,N_16082,N_17376);
nand U19069 (N_19069,N_12993,N_17389);
or U19070 (N_19070,N_12917,N_13024);
or U19071 (N_19071,N_14472,N_16893);
nor U19072 (N_19072,N_15917,N_18223);
nor U19073 (N_19073,N_14905,N_15119);
or U19074 (N_19074,N_16703,N_14947);
or U19075 (N_19075,N_18162,N_13443);
nand U19076 (N_19076,N_15038,N_15640);
nor U19077 (N_19077,N_15297,N_15023);
nand U19078 (N_19078,N_14649,N_13744);
xnor U19079 (N_19079,N_14230,N_17893);
or U19080 (N_19080,N_13574,N_15565);
xnor U19081 (N_19081,N_16084,N_17979);
nand U19082 (N_19082,N_12836,N_13818);
or U19083 (N_19083,N_18320,N_18139);
xor U19084 (N_19084,N_14967,N_15015);
nand U19085 (N_19085,N_15719,N_13796);
nand U19086 (N_19086,N_17321,N_18153);
xor U19087 (N_19087,N_12650,N_18117);
and U19088 (N_19088,N_15780,N_14752);
or U19089 (N_19089,N_13531,N_18295);
nor U19090 (N_19090,N_12794,N_13851);
xnor U19091 (N_19091,N_18548,N_15178);
nor U19092 (N_19092,N_16212,N_18197);
or U19093 (N_19093,N_13727,N_14126);
nand U19094 (N_19094,N_15818,N_17228);
nand U19095 (N_19095,N_17781,N_17425);
xor U19096 (N_19096,N_15908,N_13006);
nor U19097 (N_19097,N_15227,N_16230);
xnor U19098 (N_19098,N_15881,N_12862);
and U19099 (N_19099,N_14505,N_18298);
xor U19100 (N_19100,N_16356,N_16550);
and U19101 (N_19101,N_16200,N_13799);
nand U19102 (N_19102,N_13012,N_18504);
nor U19103 (N_19103,N_18167,N_13382);
xor U19104 (N_19104,N_17493,N_17335);
xnor U19105 (N_19105,N_15153,N_16015);
nand U19106 (N_19106,N_18726,N_18498);
or U19107 (N_19107,N_17991,N_14182);
xnor U19108 (N_19108,N_16875,N_18112);
nand U19109 (N_19109,N_13037,N_15838);
nor U19110 (N_19110,N_14999,N_13502);
or U19111 (N_19111,N_12583,N_14336);
or U19112 (N_19112,N_13597,N_18259);
xnor U19113 (N_19113,N_14158,N_17093);
and U19114 (N_19114,N_13120,N_15185);
xnor U19115 (N_19115,N_15829,N_14962);
and U19116 (N_19116,N_16594,N_12708);
or U19117 (N_19117,N_17589,N_12804);
nand U19118 (N_19118,N_13428,N_17683);
and U19119 (N_19119,N_13635,N_17950);
xor U19120 (N_19120,N_14218,N_14648);
xor U19121 (N_19121,N_16355,N_12587);
nand U19122 (N_19122,N_15683,N_18151);
nand U19123 (N_19123,N_13258,N_18069);
nor U19124 (N_19124,N_18171,N_15571);
and U19125 (N_19125,N_17887,N_12654);
or U19126 (N_19126,N_12904,N_13656);
nand U19127 (N_19127,N_16606,N_15848);
nand U19128 (N_19128,N_17086,N_14080);
nand U19129 (N_19129,N_15530,N_17285);
xor U19130 (N_19130,N_14184,N_12711);
nand U19131 (N_19131,N_17071,N_15401);
or U19132 (N_19132,N_16878,N_14917);
nor U19133 (N_19133,N_18174,N_12578);
or U19134 (N_19134,N_14074,N_16266);
or U19135 (N_19135,N_16440,N_14820);
or U19136 (N_19136,N_15610,N_15566);
xor U19137 (N_19137,N_15537,N_15161);
nand U19138 (N_19138,N_13314,N_18655);
xnor U19139 (N_19139,N_14044,N_17913);
and U19140 (N_19140,N_17536,N_12954);
xor U19141 (N_19141,N_17122,N_15627);
nand U19142 (N_19142,N_17205,N_12945);
nor U19143 (N_19143,N_16245,N_18690);
nand U19144 (N_19144,N_15304,N_13810);
xor U19145 (N_19145,N_18656,N_16405);
and U19146 (N_19146,N_13456,N_15997);
xnor U19147 (N_19147,N_13608,N_14569);
nand U19148 (N_19148,N_18220,N_14324);
nor U19149 (N_19149,N_17337,N_17802);
xnor U19150 (N_19150,N_18052,N_18622);
and U19151 (N_19151,N_13453,N_18148);
xor U19152 (N_19152,N_17353,N_15800);
nor U19153 (N_19153,N_17468,N_15539);
or U19154 (N_19154,N_15784,N_18404);
and U19155 (N_19155,N_18443,N_17186);
xnor U19156 (N_19156,N_16620,N_12593);
xnor U19157 (N_19157,N_14373,N_14790);
or U19158 (N_19158,N_14347,N_16887);
nand U19159 (N_19159,N_15116,N_18304);
or U19160 (N_19160,N_18456,N_13565);
and U19161 (N_19161,N_17361,N_18672);
xnor U19162 (N_19162,N_13704,N_14795);
or U19163 (N_19163,N_14713,N_15705);
xnor U19164 (N_19164,N_18620,N_16494);
nor U19165 (N_19165,N_13427,N_17241);
xnor U19166 (N_19166,N_18216,N_14447);
xor U19167 (N_19167,N_14921,N_15907);
nor U19168 (N_19168,N_18440,N_18458);
xnor U19169 (N_19169,N_18011,N_14534);
nor U19170 (N_19170,N_18172,N_16619);
xnor U19171 (N_19171,N_12622,N_16242);
nand U19172 (N_19172,N_16746,N_14316);
nand U19173 (N_19173,N_16735,N_17407);
and U19174 (N_19174,N_16456,N_18500);
xnor U19175 (N_19175,N_18073,N_13442);
nor U19176 (N_19176,N_13262,N_17966);
nor U19177 (N_19177,N_17436,N_13649);
nand U19178 (N_19178,N_14726,N_14566);
xnor U19179 (N_19179,N_17156,N_17147);
xnor U19180 (N_19180,N_17988,N_16166);
xnor U19181 (N_19181,N_18316,N_18325);
or U19182 (N_19182,N_17495,N_12590);
nor U19183 (N_19183,N_16431,N_17274);
nor U19184 (N_19184,N_15698,N_18480);
or U19185 (N_19185,N_18230,N_16393);
or U19186 (N_19186,N_13745,N_13748);
and U19187 (N_19187,N_16580,N_17286);
xor U19188 (N_19188,N_16528,N_18638);
and U19189 (N_19189,N_16607,N_13182);
xnor U19190 (N_19190,N_12559,N_15026);
and U19191 (N_19191,N_18293,N_18662);
or U19192 (N_19192,N_12986,N_13968);
nor U19193 (N_19193,N_16611,N_13970);
xor U19194 (N_19194,N_13568,N_16407);
and U19195 (N_19195,N_12591,N_13937);
nor U19196 (N_19196,N_18528,N_17660);
nor U19197 (N_19197,N_16958,N_16719);
xor U19198 (N_19198,N_15759,N_17344);
xnor U19199 (N_19199,N_13466,N_15975);
nand U19200 (N_19200,N_14701,N_15148);
and U19201 (N_19201,N_13127,N_14391);
nand U19202 (N_19202,N_15922,N_12850);
and U19203 (N_19203,N_15768,N_16682);
nor U19204 (N_19204,N_14496,N_13288);
nor U19205 (N_19205,N_12746,N_17461);
xnor U19206 (N_19206,N_15765,N_12728);
nand U19207 (N_19207,N_13921,N_16278);
or U19208 (N_19208,N_18503,N_18250);
nand U19209 (N_19209,N_17455,N_15830);
nand U19210 (N_19210,N_16979,N_14219);
nor U19211 (N_19211,N_17178,N_13152);
xnor U19212 (N_19212,N_15443,N_16401);
xor U19213 (N_19213,N_14356,N_16626);
or U19214 (N_19214,N_13680,N_13254);
nand U19215 (N_19215,N_16462,N_13639);
nand U19216 (N_19216,N_17388,N_15180);
nand U19217 (N_19217,N_15118,N_15164);
and U19218 (N_19218,N_17753,N_16274);
and U19219 (N_19219,N_18306,N_15043);
nor U19220 (N_19220,N_14500,N_16156);
and U19221 (N_19221,N_13731,N_15137);
and U19222 (N_19222,N_15716,N_13686);
or U19223 (N_19223,N_13946,N_17424);
nand U19224 (N_19224,N_14334,N_13666);
and U19225 (N_19225,N_16163,N_16667);
nand U19226 (N_19226,N_13789,N_17523);
nand U19227 (N_19227,N_15529,N_15238);
nor U19228 (N_19228,N_15187,N_18007);
and U19229 (N_19229,N_17264,N_17730);
or U19230 (N_19230,N_18077,N_17406);
and U19231 (N_19231,N_13079,N_17038);
nand U19232 (N_19232,N_17716,N_16737);
and U19233 (N_19233,N_14779,N_17999);
xnor U19234 (N_19234,N_15977,N_13944);
xnor U19235 (N_19235,N_18339,N_12665);
nor U19236 (N_19236,N_16403,N_12984);
and U19237 (N_19237,N_16229,N_16770);
xnor U19238 (N_19238,N_15788,N_15282);
nand U19239 (N_19239,N_17875,N_17261);
and U19240 (N_19240,N_13925,N_13080);
or U19241 (N_19241,N_16422,N_15513);
nand U19242 (N_19242,N_16310,N_13578);
nand U19243 (N_19243,N_16970,N_12894);
nor U19244 (N_19244,N_13971,N_14319);
nor U19245 (N_19245,N_13922,N_17778);
nor U19246 (N_19246,N_14148,N_14491);
or U19247 (N_19247,N_16782,N_17943);
nor U19248 (N_19248,N_13210,N_15528);
and U19249 (N_19249,N_14554,N_14156);
xnor U19250 (N_19250,N_16694,N_14762);
and U19251 (N_19251,N_12608,N_12519);
or U19252 (N_19252,N_15625,N_17396);
or U19253 (N_19253,N_13871,N_18297);
or U19254 (N_19254,N_16833,N_14221);
nor U19255 (N_19255,N_17322,N_18271);
nor U19256 (N_19256,N_15508,N_14133);
or U19257 (N_19257,N_17202,N_13168);
or U19258 (N_19258,N_14420,N_17041);
and U19259 (N_19259,N_18472,N_16701);
nand U19260 (N_19260,N_12652,N_17368);
or U19261 (N_19261,N_15732,N_16924);
nand U19262 (N_19262,N_13365,N_13188);
nor U19263 (N_19263,N_18542,N_13131);
nand U19264 (N_19264,N_16630,N_17900);
and U19265 (N_19265,N_13105,N_18257);
nand U19266 (N_19266,N_16299,N_16139);
nor U19267 (N_19267,N_12552,N_13918);
nor U19268 (N_19268,N_16724,N_18087);
or U19269 (N_19269,N_13959,N_13973);
nor U19270 (N_19270,N_17503,N_13251);
nor U19271 (N_19271,N_18336,N_12953);
nand U19272 (N_19272,N_12885,N_18364);
xnor U19273 (N_19273,N_15616,N_15817);
nor U19274 (N_19274,N_16076,N_14098);
or U19275 (N_19275,N_12983,N_12693);
or U19276 (N_19276,N_15548,N_16997);
or U19277 (N_19277,N_17000,N_15541);
nor U19278 (N_19278,N_14821,N_13985);
xor U19279 (N_19279,N_12730,N_13896);
nor U19280 (N_19280,N_12898,N_16375);
or U19281 (N_19281,N_17598,N_14988);
or U19282 (N_19282,N_13265,N_12760);
nor U19283 (N_19283,N_17377,N_12764);
xor U19284 (N_19284,N_12537,N_13836);
or U19285 (N_19285,N_16926,N_18437);
nand U19286 (N_19286,N_13317,N_18194);
xnor U19287 (N_19287,N_16710,N_18442);
and U19288 (N_19288,N_14058,N_18191);
or U19289 (N_19289,N_16882,N_12955);
or U19290 (N_19290,N_13070,N_18717);
nor U19291 (N_19291,N_17075,N_14154);
nor U19292 (N_19292,N_17841,N_14352);
nor U19293 (N_19293,N_17834,N_12856);
xnor U19294 (N_19294,N_18260,N_15470);
and U19295 (N_19295,N_14618,N_14753);
or U19296 (N_19296,N_17500,N_15494);
nand U19297 (N_19297,N_13626,N_18155);
nand U19298 (N_19298,N_17370,N_16944);
xnor U19299 (N_19299,N_15239,N_17331);
nand U19300 (N_19300,N_13515,N_15516);
nand U19301 (N_19301,N_14742,N_16496);
nor U19302 (N_19302,N_16243,N_16234);
and U19303 (N_19303,N_16565,N_15121);
xnor U19304 (N_19304,N_15389,N_12701);
xnor U19305 (N_19305,N_13364,N_15562);
nor U19306 (N_19306,N_15789,N_13872);
nand U19307 (N_19307,N_13147,N_18160);
nor U19308 (N_19308,N_14455,N_16368);
xnor U19309 (N_19309,N_18138,N_17579);
xnor U19310 (N_19310,N_12846,N_13117);
and U19311 (N_19311,N_14202,N_12807);
nand U19312 (N_19312,N_13047,N_13718);
nand U19313 (N_19313,N_12757,N_13730);
and U19314 (N_19314,N_14028,N_13029);
nor U19315 (N_19315,N_15843,N_15163);
or U19316 (N_19316,N_16938,N_13497);
nand U19317 (N_19317,N_15033,N_18064);
nor U19318 (N_19318,N_18596,N_13566);
nor U19319 (N_19319,N_17272,N_14388);
and U19320 (N_19320,N_13434,N_17070);
or U19321 (N_19321,N_14766,N_12819);
or U19322 (N_19322,N_13446,N_16805);
and U19323 (N_19323,N_12779,N_13190);
nor U19324 (N_19324,N_16196,N_15405);
xnor U19325 (N_19325,N_17566,N_17971);
nor U19326 (N_19326,N_13109,N_13884);
or U19327 (N_19327,N_15778,N_14240);
nand U19328 (N_19328,N_12994,N_13753);
xnor U19329 (N_19329,N_17746,N_17176);
xnor U19330 (N_19330,N_17085,N_15379);
and U19331 (N_19331,N_17479,N_15384);
and U19332 (N_19332,N_14170,N_15790);
or U19333 (N_19333,N_15837,N_17080);
or U19334 (N_19334,N_16228,N_13203);
or U19335 (N_19335,N_18521,N_16126);
or U19336 (N_19336,N_14658,N_16257);
or U19337 (N_19337,N_16723,N_17124);
nor U19338 (N_19338,N_17360,N_18084);
and U19339 (N_19339,N_12632,N_18415);
and U19340 (N_19340,N_13158,N_15966);
nor U19341 (N_19341,N_17509,N_12828);
or U19342 (N_19342,N_16054,N_13346);
and U19343 (N_19343,N_13996,N_18559);
nand U19344 (N_19344,N_14859,N_14654);
xor U19345 (N_19345,N_14880,N_15031);
nor U19346 (N_19346,N_16794,N_12747);
or U19347 (N_19347,N_15597,N_13725);
nand U19348 (N_19348,N_18623,N_14515);
xor U19349 (N_19349,N_17076,N_16969);
nor U19350 (N_19350,N_15272,N_13699);
and U19351 (N_19351,N_17058,N_16335);
or U19352 (N_19352,N_16083,N_18677);
xor U19353 (N_19353,N_15808,N_18650);
nor U19354 (N_19354,N_13086,N_13010);
and U19355 (N_19355,N_18489,N_18471);
nand U19356 (N_19356,N_13962,N_13722);
nand U19357 (N_19357,N_16652,N_16842);
or U19358 (N_19358,N_12651,N_13324);
and U19359 (N_19359,N_15213,N_15483);
nor U19360 (N_19360,N_18562,N_17247);
nand U19361 (N_19361,N_16577,N_13802);
xor U19362 (N_19362,N_15130,N_16809);
xor U19363 (N_19363,N_14091,N_16290);
and U19364 (N_19364,N_13624,N_12662);
xor U19365 (N_19365,N_12726,N_12790);
and U19366 (N_19366,N_16544,N_13513);
nor U19367 (N_19367,N_17933,N_12996);
nor U19368 (N_19368,N_13011,N_14693);
or U19369 (N_19369,N_16526,N_13239);
nor U19370 (N_19370,N_13936,N_14551);
or U19371 (N_19371,N_16154,N_17854);
nor U19372 (N_19372,N_15413,N_12724);
nor U19373 (N_19373,N_14422,N_15449);
and U19374 (N_19374,N_13230,N_16867);
or U19375 (N_19375,N_16656,N_13202);
or U19376 (N_19376,N_16736,N_17239);
xor U19377 (N_19377,N_18450,N_13772);
xnor U19378 (N_19378,N_14320,N_18255);
xnor U19379 (N_19379,N_17546,N_15165);
and U19380 (N_19380,N_14435,N_18491);
and U19381 (N_19381,N_13557,N_17514);
and U19382 (N_19382,N_16986,N_13143);
nor U19383 (N_19383,N_14475,N_17667);
nand U19384 (N_19384,N_18431,N_15482);
nand U19385 (N_19385,N_13267,N_13929);
xnor U19386 (N_19386,N_15702,N_18536);
nand U19387 (N_19387,N_12564,N_15391);
nand U19388 (N_19388,N_16390,N_14827);
xnor U19389 (N_19389,N_16436,N_15502);
nor U19390 (N_19390,N_18147,N_18002);
nand U19391 (N_19391,N_12549,N_17855);
or U19392 (N_19392,N_18406,N_14234);
xnor U19393 (N_19393,N_17459,N_18633);
nor U19394 (N_19394,N_13788,N_13228);
or U19395 (N_19395,N_14239,N_17157);
nor U19396 (N_19396,N_14171,N_17554);
xor U19397 (N_19397,N_15051,N_15674);
nor U19398 (N_19398,N_17822,N_17300);
and U19399 (N_19399,N_13616,N_14946);
nand U19400 (N_19400,N_13316,N_13690);
or U19401 (N_19401,N_13902,N_14294);
nand U19402 (N_19402,N_14338,N_18465);
xor U19403 (N_19403,N_15506,N_14285);
nor U19404 (N_19404,N_13545,N_17782);
or U19405 (N_19405,N_13653,N_14313);
nand U19406 (N_19406,N_15746,N_17193);
nand U19407 (N_19407,N_12933,N_14652);
and U19408 (N_19408,N_16674,N_15637);
nand U19409 (N_19409,N_15691,N_14159);
nand U19410 (N_19410,N_18253,N_16233);
or U19411 (N_19411,N_13009,N_15911);
and U19412 (N_19412,N_16600,N_15821);
or U19413 (N_19413,N_14205,N_16018);
and U19414 (N_19414,N_14481,N_13271);
or U19415 (N_19415,N_17678,N_13111);
xor U19416 (N_19416,N_18369,N_16669);
nand U19417 (N_19417,N_16857,N_17113);
nand U19418 (N_19418,N_13790,N_16877);
xnor U19419 (N_19419,N_13646,N_15351);
nor U19420 (N_19420,N_16114,N_15446);
or U19421 (N_19421,N_16865,N_18645);
nor U19422 (N_19422,N_16758,N_14671);
or U19423 (N_19423,N_17670,N_18175);
nand U19424 (N_19424,N_15722,N_17704);
xnor U19425 (N_19425,N_16072,N_15319);
nor U19426 (N_19426,N_13781,N_13061);
and U19427 (N_19427,N_15845,N_18639);
nor U19428 (N_19428,N_16688,N_16732);
xor U19429 (N_19429,N_13376,N_14132);
xor U19430 (N_19430,N_15684,N_15827);
nand U19431 (N_19431,N_13026,N_16942);
nand U19432 (N_19432,N_18374,N_15697);
and U19433 (N_19433,N_14049,N_13493);
xnor U19434 (N_19434,N_14358,N_18088);
and U19435 (N_19435,N_13148,N_15376);
nand U19436 (N_19436,N_12921,N_17941);
or U19437 (N_19437,N_14023,N_13524);
nor U19438 (N_19438,N_17074,N_15454);
or U19439 (N_19439,N_16558,N_18475);
and U19440 (N_19440,N_18238,N_13102);
and U19441 (N_19441,N_17045,N_12791);
and U19442 (N_19442,N_16772,N_17641);
nand U19443 (N_19443,N_13924,N_17952);
xnor U19444 (N_19444,N_17128,N_12614);
or U19445 (N_19445,N_18428,N_13598);
nor U19446 (N_19446,N_15061,N_17772);
nor U19447 (N_19447,N_14122,N_17698);
nand U19448 (N_19448,N_17539,N_13264);
nand U19449 (N_19449,N_16917,N_16152);
or U19450 (N_19450,N_18629,N_18280);
xor U19451 (N_19451,N_12861,N_17387);
xnor U19452 (N_19452,N_18357,N_13888);
xnor U19453 (N_19453,N_16681,N_16432);
nor U19454 (N_19454,N_14849,N_14961);
xnor U19455 (N_19455,N_14575,N_18149);
or U19456 (N_19456,N_13657,N_14991);
nor U19457 (N_19457,N_17818,N_13139);
nand U19458 (N_19458,N_17666,N_17911);
and U19459 (N_19459,N_17848,N_12748);
and U19460 (N_19460,N_16906,N_16708);
nand U19461 (N_19461,N_16959,N_14511);
or U19462 (N_19462,N_18006,N_16447);
nand U19463 (N_19463,N_15081,N_15986);
nand U19464 (N_19464,N_15890,N_18483);
xnor U19465 (N_19465,N_14623,N_17297);
and U19466 (N_19466,N_13087,N_18109);
or U19467 (N_19467,N_13450,N_18683);
and U19468 (N_19468,N_16704,N_14974);
nand U19469 (N_19469,N_17190,N_15093);
and U19470 (N_19470,N_17251,N_18133);
or U19471 (N_19471,N_12742,N_16616);
xnor U19472 (N_19472,N_18127,N_12799);
xor U19473 (N_19473,N_18691,N_13157);
nand U19474 (N_19474,N_15874,N_16209);
and U19475 (N_19475,N_15544,N_15583);
nor U19476 (N_19476,N_12781,N_16645);
nand U19477 (N_19477,N_14530,N_16471);
and U19478 (N_19478,N_18412,N_13467);
or U19479 (N_19479,N_16279,N_13125);
or U19480 (N_19480,N_15062,N_15932);
or U19481 (N_19481,N_13997,N_16252);
xnor U19482 (N_19482,N_16592,N_18305);
and U19483 (N_19483,N_18198,N_15559);
xnor U19484 (N_19484,N_12741,N_14163);
and U19485 (N_19485,N_17597,N_15123);
and U19486 (N_19486,N_12880,N_16470);
or U19487 (N_19487,N_14943,N_14872);
or U19488 (N_19488,N_16322,N_14470);
and U19489 (N_19489,N_18618,N_17624);
nand U19490 (N_19490,N_12520,N_18136);
xnor U19491 (N_19491,N_16428,N_15521);
nand U19492 (N_19492,N_16025,N_17868);
nand U19493 (N_19493,N_12692,N_16276);
nand U19494 (N_19494,N_15671,N_14525);
or U19495 (N_19495,N_14137,N_14944);
nor U19496 (N_19496,N_15886,N_15322);
or U19497 (N_19497,N_17814,N_16024);
xor U19498 (N_19498,N_16711,N_13715);
or U19499 (N_19499,N_15862,N_13739);
xnor U19500 (N_19500,N_12666,N_17140);
or U19501 (N_19501,N_14659,N_17013);
nor U19502 (N_19502,N_16280,N_18324);
and U19503 (N_19503,N_14959,N_13128);
xnor U19504 (N_19504,N_15375,N_16112);
nand U19505 (N_19505,N_13423,N_15243);
xor U19506 (N_19506,N_16159,N_13692);
or U19507 (N_19507,N_17690,N_17474);
and U19508 (N_19508,N_18326,N_18675);
nor U19509 (N_19509,N_16133,N_17935);
or U19510 (N_19510,N_16510,N_14340);
xor U19511 (N_19511,N_13926,N_15488);
nand U19512 (N_19512,N_12661,N_17023);
nand U19513 (N_19513,N_17901,N_17498);
nand U19514 (N_19514,N_14622,N_13647);
and U19515 (N_19515,N_13689,N_15371);
and U19516 (N_19516,N_14709,N_18592);
xor U19517 (N_19517,N_17363,N_13171);
xnor U19518 (N_19518,N_16657,N_12809);
or U19519 (N_19519,N_15204,N_16117);
nand U19520 (N_19520,N_13854,N_15588);
nor U19521 (N_19521,N_12876,N_12865);
nand U19522 (N_19522,N_15019,N_17864);
nand U19523 (N_19523,N_12875,N_14628);
and U19524 (N_19524,N_18301,N_13027);
xor U19525 (N_19525,N_17385,N_18173);
nor U19526 (N_19526,N_13280,N_15809);
nor U19527 (N_19527,N_13613,N_15568);
or U19528 (N_19528,N_18342,N_15531);
nand U19529 (N_19529,N_18640,N_13661);
or U19530 (N_19530,N_18283,N_16433);
nor U19531 (N_19531,N_13868,N_15342);
nand U19532 (N_19532,N_18696,N_16622);
nand U19533 (N_19533,N_14343,N_17853);
and U19534 (N_19534,N_13636,N_17676);
nand U19535 (N_19535,N_17578,N_13831);
xnor U19536 (N_19536,N_15592,N_18544);
nor U19537 (N_19537,N_18125,N_15618);
nand U19538 (N_19538,N_15520,N_14626);
or U19539 (N_19539,N_16542,N_14029);
xor U19540 (N_19540,N_17238,N_12788);
or U19541 (N_19541,N_16568,N_13233);
nand U19542 (N_19542,N_16040,N_17630);
nand U19543 (N_19543,N_17620,N_15992);
nand U19544 (N_19544,N_13528,N_18232);
nand U19545 (N_19545,N_17472,N_12530);
nand U19546 (N_19546,N_16983,N_16503);
nor U19547 (N_19547,N_16226,N_13792);
xnor U19548 (N_19548,N_16593,N_16444);
and U19549 (N_19549,N_14418,N_15285);
xor U19550 (N_19550,N_17365,N_16506);
nand U19551 (N_19551,N_18429,N_12570);
nand U19552 (N_19552,N_14514,N_16260);
nor U19553 (N_19553,N_15289,N_16068);
or U19554 (N_19554,N_18720,N_12547);
and U19555 (N_19555,N_15242,N_12700);
or U19556 (N_19556,N_14412,N_12838);
nor U19557 (N_19557,N_17576,N_12678);
nand U19558 (N_19558,N_18269,N_13435);
and U19559 (N_19559,N_14103,N_17773);
nand U19560 (N_19560,N_16849,N_15197);
nor U19561 (N_19561,N_15102,N_16659);
and U19562 (N_19562,N_12990,N_17525);
nand U19563 (N_19563,N_17230,N_14729);
xor U19564 (N_19564,N_17586,N_16264);
and U19565 (N_19565,N_13303,N_13540);
xnor U19566 (N_19566,N_12702,N_12769);
xnor U19567 (N_19567,N_16467,N_16549);
nor U19568 (N_19568,N_16445,N_13558);
nor U19569 (N_19569,N_15416,N_16615);
and U19570 (N_19570,N_14941,N_16164);
and U19571 (N_19571,N_18178,N_16173);
nand U19572 (N_19572,N_14309,N_14109);
xnor U19573 (N_19573,N_14189,N_14704);
xnor U19574 (N_19574,N_15024,N_17123);
nor U19575 (N_19575,N_17401,N_18461);
xnor U19576 (N_19576,N_14055,N_12874);
or U19577 (N_19577,N_14938,N_14459);
nand U19578 (N_19578,N_17529,N_17465);
nor U19579 (N_19579,N_13007,N_18660);
xnor U19580 (N_19580,N_17454,N_18334);
xor U19581 (N_19581,N_15591,N_18722);
nand U19582 (N_19582,N_13241,N_12716);
and U19583 (N_19583,N_13572,N_18361);
nand U19584 (N_19584,N_18054,N_18704);
and U19585 (N_19585,N_12911,N_17442);
xnor U19586 (N_19586,N_13478,N_14818);
or U19587 (N_19587,N_15464,N_14082);
xnor U19588 (N_19588,N_14744,N_14247);
or U19589 (N_19589,N_13437,N_16175);
and U19590 (N_19590,N_14601,N_15664);
xnor U19591 (N_19591,N_17572,N_18016);
or U19592 (N_19592,N_16668,N_12569);
nor U19593 (N_19593,N_17350,N_17762);
nor U19594 (N_19594,N_17460,N_16891);
and U19595 (N_19595,N_14421,N_14254);
xor U19596 (N_19596,N_15624,N_14964);
and U19597 (N_19597,N_15939,N_17664);
xnor U19598 (N_19598,N_18614,N_17340);
and U19599 (N_19599,N_12960,N_14369);
and U19600 (N_19600,N_14364,N_18287);
xnor U19601 (N_19601,N_16454,N_15561);
xor U19602 (N_19602,N_17895,N_14835);
xor U19603 (N_19603,N_13424,N_18527);
nand U19604 (N_19604,N_12531,N_12785);
xor U19605 (N_19605,N_16518,N_15005);
nor U19606 (N_19606,N_15218,N_18270);
or U19607 (N_19607,N_18434,N_15200);
xor U19608 (N_19608,N_18284,N_15621);
nand U19609 (N_19609,N_15028,N_16003);
or U19610 (N_19610,N_18075,N_14077);
xnor U19611 (N_19611,N_18315,N_15018);
nand U19612 (N_19612,N_14030,N_18131);
and U19613 (N_19613,N_18405,N_14383);
nor U19614 (N_19614,N_18018,N_14079);
xnor U19615 (N_19615,N_16598,N_16590);
and U19616 (N_19616,N_14377,N_17240);
xor U19617 (N_19617,N_14024,N_12841);
nand U19618 (N_19618,N_16564,N_17876);
nor U19619 (N_19619,N_16802,N_14956);
nand U19620 (N_19620,N_12896,N_14105);
xnor U19621 (N_19621,N_16579,N_13452);
and U19622 (N_19622,N_13212,N_16847);
and U19623 (N_19623,N_13507,N_17131);
or U19624 (N_19624,N_16340,N_14825);
nand U19625 (N_19625,N_14754,N_13820);
nand U19626 (N_19626,N_15824,N_15582);
nor U19627 (N_19627,N_16153,N_17051);
or U19628 (N_19628,N_12857,N_15349);
or U19629 (N_19629,N_15472,N_18034);
or U19630 (N_19630,N_18081,N_15252);
nor U19631 (N_19631,N_14676,N_13362);
xor U19632 (N_19632,N_18144,N_17192);
xnor U19633 (N_19633,N_18323,N_17362);
nor U19634 (N_19634,N_15232,N_13063);
nor U19635 (N_19635,N_17133,N_16008);
and U19636 (N_19636,N_18535,N_14368);
and U19637 (N_19637,N_15010,N_13938);
and U19638 (N_19638,N_15795,N_14661);
and U19639 (N_19639,N_16972,N_14266);
nand U19640 (N_19640,N_14557,N_16655);
xor U19641 (N_19641,N_16081,N_13058);
nand U19642 (N_19642,N_14076,N_18391);
nand U19643 (N_19643,N_17877,N_16178);
xor U19644 (N_19644,N_15710,N_14817);
and U19645 (N_19645,N_14773,N_15758);
or U19646 (N_19646,N_18583,N_13843);
and U19647 (N_19647,N_16570,N_14411);
and U19648 (N_19648,N_16171,N_16745);
xnor U19649 (N_19649,N_16005,N_16596);
nand U19650 (N_19650,N_16167,N_18045);
or U19651 (N_19651,N_13078,N_14647);
and U19652 (N_19652,N_14942,N_13244);
and U19653 (N_19653,N_12599,N_17992);
xor U19654 (N_19654,N_14492,N_17163);
nand U19655 (N_19655,N_18715,N_17471);
or U19656 (N_19656,N_13536,N_16225);
nor U19657 (N_19657,N_15256,N_17339);
and U19658 (N_19658,N_14517,N_15122);
xnor U19659 (N_19659,N_12705,N_17798);
or U19660 (N_19660,N_12727,N_15052);
and U19661 (N_19661,N_18132,N_17725);
nand U19662 (N_19662,N_16962,N_15453);
and U19663 (N_19663,N_16206,N_18128);
nor U19664 (N_19664,N_15195,N_17795);
nor U19665 (N_19665,N_13537,N_13155);
nor U19666 (N_19666,N_17040,N_17921);
or U19667 (N_19667,N_13589,N_13290);
or U19668 (N_19668,N_14092,N_18467);
and U19669 (N_19669,N_17236,N_17603);
nand U19670 (N_19670,N_12931,N_13883);
or U19671 (N_19671,N_14168,N_13559);
nor U19672 (N_19672,N_13166,N_16115);
nand U19673 (N_19673,N_18062,N_15755);
and U19674 (N_19674,N_17266,N_16062);
or U19675 (N_19675,N_15673,N_13055);
nor U19676 (N_19676,N_15145,N_17513);
nor U19677 (N_19677,N_16034,N_16825);
nand U19678 (N_19678,N_14549,N_12968);
nor U19679 (N_19679,N_17135,N_13349);
or U19680 (N_19680,N_16272,N_13881);
xor U19681 (N_19681,N_15078,N_13614);
or U19682 (N_19682,N_13700,N_15176);
nand U19683 (N_19683,N_17926,N_15864);
or U19684 (N_19684,N_17705,N_14478);
or U19685 (N_19685,N_15231,N_13328);
or U19686 (N_19686,N_18446,N_15783);
nand U19687 (N_19687,N_15944,N_15614);
and U19688 (N_19688,N_14232,N_16932);
nor U19689 (N_19689,N_13550,N_14916);
nand U19690 (N_19690,N_15773,N_16976);
nor U19691 (N_19691,N_17033,N_18373);
and U19692 (N_19692,N_14538,N_14672);
and U19693 (N_19693,N_17423,N_16650);
nand U19694 (N_19694,N_14668,N_13431);
xnor U19695 (N_19695,N_16811,N_15973);
and U19696 (N_19696,N_17839,N_17172);
nand U19697 (N_19697,N_14683,N_14887);
nand U19698 (N_19698,N_16256,N_13176);
and U19699 (N_19699,N_15635,N_16722);
or U19700 (N_19700,N_12514,N_16691);
and U19701 (N_19701,N_14548,N_14940);
and U19702 (N_19702,N_18749,N_17021);
or U19703 (N_19703,N_16552,N_13232);
or U19704 (N_19704,N_15027,N_14201);
xor U19705 (N_19705,N_12656,N_13141);
or U19706 (N_19706,N_13853,N_17533);
nand U19707 (N_19707,N_18524,N_14495);
and U19708 (N_19708,N_17874,N_15412);
or U19709 (N_19709,N_15226,N_18393);
or U19710 (N_19710,N_13681,N_15948);
xnor U19711 (N_19711,N_13767,N_18385);
xnor U19712 (N_19712,N_18518,N_14165);
or U19713 (N_19713,N_13668,N_18222);
and U19714 (N_19714,N_16306,N_12913);
xor U19715 (N_19715,N_17006,N_13146);
nand U19716 (N_19716,N_16477,N_18181);
nand U19717 (N_19717,N_16628,N_12867);
or U19718 (N_19718,N_16031,N_16729);
or U19719 (N_19719,N_15208,N_14950);
xnor U19720 (N_19720,N_17091,N_13094);
or U19721 (N_19721,N_14246,N_14020);
nor U19722 (N_19722,N_17542,N_16037);
xnor U19723 (N_19723,N_16581,N_15277);
nand U19724 (N_19724,N_14087,N_13791);
and U19725 (N_19725,N_16930,N_13837);
nand U19726 (N_19726,N_15474,N_15718);
and U19727 (N_19727,N_14900,N_14217);
nor U19728 (N_19728,N_18436,N_15799);
nor U19729 (N_19729,N_13754,N_13575);
nand U19730 (N_19730,N_15951,N_12554);
xor U19731 (N_19731,N_17652,N_15515);
xor U19732 (N_19732,N_14440,N_17687);
nor U19733 (N_19733,N_16684,N_13828);
or U19734 (N_19734,N_13413,N_16223);
and U19735 (N_19735,N_14749,N_14193);
nor U19736 (N_19736,N_18097,N_15311);
nor U19737 (N_19737,N_13165,N_17167);
nand U19738 (N_19738,N_17457,N_18056);
and U19739 (N_19739,N_16933,N_13153);
nor U19740 (N_19740,N_14797,N_18492);
and U19741 (N_19741,N_18363,N_18598);
nor U19742 (N_19742,N_16660,N_16013);
or U19743 (N_19743,N_15189,N_15517);
and U19744 (N_19744,N_13778,N_16754);
nor U19745 (N_19745,N_14721,N_16466);
and U19746 (N_19746,N_14090,N_16610);
or U19747 (N_19747,N_14288,N_18383);
nand U19748 (N_19748,N_14607,N_18274);
and U19749 (N_19749,N_13088,N_16515);
and U19750 (N_19750,N_14844,N_13370);
nor U19751 (N_19751,N_17987,N_18309);
nand U19752 (N_19752,N_15815,N_13389);
nor U19753 (N_19753,N_13980,N_17967);
xnor U19754 (N_19754,N_17150,N_16241);
and U19755 (N_19755,N_14645,N_16476);
nand U19756 (N_19756,N_15411,N_13170);
nand U19757 (N_19757,N_14996,N_13969);
nand U19758 (N_19758,N_16289,N_14528);
xnor U19759 (N_19759,N_14277,N_18474);
and U19760 (N_19760,N_14047,N_18362);
and U19761 (N_19761,N_15601,N_16988);
nand U19762 (N_19762,N_17308,N_17903);
and U19763 (N_19763,N_14909,N_13623);
nand U19764 (N_19764,N_18302,N_13752);
nor U19765 (N_19765,N_15166,N_13900);
xnor U19766 (N_19766,N_15223,N_15262);
and U19767 (N_19767,N_16774,N_17470);
xor U19768 (N_19768,N_13840,N_17569);
nor U19769 (N_19769,N_17015,N_18648);
xor U19770 (N_19770,N_13808,N_12893);
xnor U19771 (N_19771,N_12973,N_17102);
and U19772 (N_19772,N_13083,N_15356);
nand U19773 (N_19773,N_13554,N_13509);
and U19774 (N_19774,N_14180,N_13032);
and U19775 (N_19775,N_12849,N_15402);
or U19776 (N_19776,N_16705,N_14705);
and U19777 (N_19777,N_15168,N_18372);
or U19778 (N_19778,N_15340,N_13641);
nand U19779 (N_19779,N_16756,N_18030);
and U19780 (N_19780,N_14466,N_13374);
xor U19781 (N_19781,N_17708,N_14167);
and U19782 (N_19782,N_13811,N_13110);
or U19783 (N_19783,N_15631,N_16591);
or U19784 (N_19784,N_12550,N_15847);
nor U19785 (N_19785,N_15950,N_17025);
nor U19786 (N_19786,N_13547,N_15055);
xnor U19787 (N_19787,N_12538,N_13091);
and U19788 (N_19788,N_17126,N_18356);
and U19789 (N_19789,N_14746,N_14350);
or U19790 (N_19790,N_17957,N_18022);
and U19791 (N_19791,N_16485,N_15308);
nand U19792 (N_19792,N_13842,N_15960);
or U19793 (N_19793,N_13807,N_18628);
xnor U19794 (N_19794,N_17043,N_18396);
or U19795 (N_19795,N_17914,N_13295);
or U19796 (N_19796,N_15626,N_18605);
or U19797 (N_19797,N_14441,N_14322);
and U19798 (N_19798,N_17056,N_13448);
and U19799 (N_19799,N_16817,N_16852);
xnor U19800 (N_19800,N_17675,N_12948);
or U19801 (N_19801,N_17748,N_17744);
nor U19802 (N_19802,N_15699,N_13876);
and U19803 (N_19803,N_18102,N_18729);
or U19804 (N_19804,N_14527,N_16334);
or U19805 (N_19805,N_17618,N_13679);
or U19806 (N_19806,N_16349,N_12579);
nor U19807 (N_19807,N_15089,N_14241);
or U19808 (N_19808,N_14489,N_18247);
xor U19809 (N_19809,N_15507,N_14862);
and U19810 (N_19810,N_15546,N_15012);
and U19811 (N_19811,N_14064,N_17348);
nor U19812 (N_19812,N_15021,N_13081);
xnor U19813 (N_19813,N_13445,N_14016);
or U19814 (N_19814,N_14005,N_15632);
nand U19815 (N_19815,N_14560,N_18510);
or U19816 (N_19816,N_14655,N_16181);
nor U19817 (N_19817,N_16120,N_15871);
nor U19818 (N_19818,N_17359,N_14131);
or U19819 (N_19819,N_16791,N_17270);
and U19820 (N_19820,N_14537,N_12940);
or U19821 (N_19821,N_17132,N_16298);
nand U19822 (N_19822,N_12787,N_15057);
nor U19823 (N_19823,N_16707,N_13040);
or U19824 (N_19824,N_15949,N_18576);
or U19825 (N_19825,N_12947,N_16395);
nand U19826 (N_19826,N_16410,N_16151);
or U19827 (N_19827,N_16658,N_15958);
or U19828 (N_19828,N_17574,N_14053);
and U19829 (N_19829,N_16949,N_14051);
nand U19830 (N_19830,N_18567,N_13357);
nand U19831 (N_19831,N_13135,N_14497);
or U19832 (N_19832,N_14291,N_16673);
or U19833 (N_19833,N_14484,N_16102);
nor U19834 (N_19834,N_16788,N_13927);
nor U19835 (N_19835,N_12920,N_17299);
and U19836 (N_19836,N_16092,N_17200);
xnor U19837 (N_19837,N_16080,N_17211);
xor U19838 (N_19838,N_14589,N_15260);
or U19839 (N_19839,N_15542,N_14015);
nand U19840 (N_19840,N_12972,N_16987);
or U19841 (N_19841,N_13292,N_17760);
nand U19842 (N_19842,N_13181,N_16011);
or U19843 (N_19843,N_13028,N_18409);
nor U19844 (N_19844,N_15857,N_14567);
and U19845 (N_19845,N_16713,N_15403);
and U19846 (N_19846,N_16902,N_14595);
or U19847 (N_19847,N_14116,N_14448);
or U19848 (N_19848,N_16547,N_18669);
nor U19849 (N_19849,N_14287,N_18612);
and U19850 (N_19850,N_14245,N_16661);
or U19851 (N_19851,N_17408,N_13815);
xor U19852 (N_19852,N_14404,N_13688);
nand U19853 (N_19853,N_16831,N_14043);
nand U19854 (N_19854,N_16042,N_16185);
and U19855 (N_19855,N_18670,N_14339);
nand U19856 (N_19856,N_13312,N_16071);
or U19857 (N_19857,N_17908,N_15060);
and U19858 (N_19858,N_16672,N_13579);
or U19859 (N_19859,N_14389,N_15257);
or U19860 (N_19860,N_15112,N_17049);
nand U19861 (N_19861,N_16781,N_12909);
or U19862 (N_19862,N_18743,N_12814);
nand U19863 (N_19863,N_18604,N_18332);
nor U19864 (N_19864,N_15854,N_14363);
nand U19865 (N_19865,N_17626,N_16376);
xnor U19866 (N_19866,N_16387,N_13407);
xor U19867 (N_19867,N_12551,N_15343);
or U19868 (N_19868,N_13107,N_12597);
and U19869 (N_19869,N_15316,N_15792);
or U19870 (N_19870,N_16023,N_17924);
and U19871 (N_19871,N_16856,N_16419);
xnor U19872 (N_19872,N_12937,N_18520);
nand U19873 (N_19873,N_18340,N_15876);
or U19874 (N_19874,N_16750,N_17009);
xnor U19875 (N_19875,N_17413,N_17096);
xnor U19876 (N_19876,N_14401,N_15281);
nand U19877 (N_19877,N_17622,N_12633);
nor U19878 (N_19878,N_17754,N_16183);
and U19879 (N_19879,N_13327,N_15071);
nand U19880 (N_19880,N_16741,N_13804);
nand U19881 (N_19881,N_15609,N_18184);
nand U19882 (N_19882,N_15259,N_18118);
nand U19883 (N_19883,N_15076,N_15392);
nand U19884 (N_19884,N_16583,N_14235);
or U19885 (N_19885,N_16180,N_16557);
and U19886 (N_19886,N_15841,N_12516);
nand U19887 (N_19887,N_17958,N_14883);
nand U19888 (N_19888,N_18486,N_13399);
or U19889 (N_19889,N_18748,N_15422);
xor U19890 (N_19890,N_12603,N_18188);
and U19891 (N_19891,N_17394,N_16103);
nor U19892 (N_19892,N_17047,N_16425);
or U19893 (N_19893,N_13743,N_17305);
nand U19894 (N_19894,N_14796,N_15394);
nor U19895 (N_19895,N_13227,N_14298);
nor U19896 (N_19896,N_13898,N_17700);
or U19897 (N_19897,N_14477,N_15687);
xnor U19898 (N_19898,N_17969,N_18543);
nand U19899 (N_19899,N_15743,N_16437);
nor U19900 (N_19900,N_13468,N_12504);
or U19901 (N_19901,N_14317,N_16505);
nand U19902 (N_19902,N_14572,N_15828);
nand U19903 (N_19903,N_15756,N_16780);
nand U19904 (N_19904,N_14980,N_16325);
and U19905 (N_19905,N_15329,N_14462);
xor U19906 (N_19906,N_17886,N_14860);
xnor U19907 (N_19907,N_18558,N_18037);
xor U19908 (N_19908,N_12670,N_17029);
nor U19909 (N_19909,N_12607,N_17234);
nor U19910 (N_19910,N_13961,N_15968);
and U19911 (N_19911,N_15704,N_17757);
xor U19912 (N_19912,N_14857,N_14543);
nor U19913 (N_19913,N_14187,N_14405);
xnor U19914 (N_19914,N_12630,N_17328);
xnor U19915 (N_19915,N_16693,N_17399);
or U19916 (N_19916,N_14072,N_16345);
and U19917 (N_19917,N_15046,N_18701);
or U19918 (N_19918,N_17605,N_17354);
and U19919 (N_19919,N_17796,N_18351);
and U19920 (N_19920,N_17296,N_18086);
xnor U19921 (N_19921,N_16359,N_12576);
xor U19922 (N_19922,N_14021,N_15518);
xor U19923 (N_19923,N_16751,N_13163);
xor U19924 (N_19924,N_18355,N_13154);
and U19925 (N_19925,N_15525,N_14975);
and U19926 (N_19926,N_12930,N_13667);
or U19927 (N_19927,N_16666,N_15646);
xnor U19928 (N_19928,N_16639,N_16636);
nor U19929 (N_19929,N_18606,N_16815);
or U19930 (N_19930,N_18268,N_16283);
or U19931 (N_19931,N_17304,N_16752);
or U19932 (N_19932,N_18262,N_16055);
nor U19933 (N_19933,N_12773,N_15105);
and U19934 (N_19934,N_14650,N_17050);
and U19935 (N_19935,N_13795,N_15129);
nand U19936 (N_19936,N_15059,N_17182);
nand U19937 (N_19937,N_12513,N_17439);
nand U19938 (N_19938,N_14772,N_13321);
or U19939 (N_19939,N_16653,N_15273);
or U19940 (N_19940,N_13043,N_13381);
and U19941 (N_19941,N_14328,N_13992);
nor U19942 (N_19942,N_13609,N_12868);
or U19943 (N_19943,N_16955,N_14679);
nand U19944 (N_19944,N_15630,N_14130);
and U19945 (N_19945,N_16429,N_13041);
xnor U19946 (N_19946,N_15672,N_14711);
nand U19947 (N_19947,N_17208,N_14283);
xor U19948 (N_19948,N_14600,N_17235);
xor U19949 (N_19949,N_14017,N_17168);
nor U19950 (N_19950,N_12721,N_14819);
or U19951 (N_19951,N_14110,N_13797);
nand U19952 (N_19952,N_18470,N_14104);
xnor U19953 (N_19953,N_15307,N_12686);
nand U19954 (N_19954,N_18435,N_18487);
and U19955 (N_19955,N_15652,N_15173);
nor U19956 (N_19956,N_18095,N_17067);
nor U19957 (N_19957,N_13905,N_16187);
and U19958 (N_19958,N_17724,N_17518);
nor U19959 (N_19959,N_16586,N_18365);
nor U19960 (N_19960,N_17130,N_14449);
or U19961 (N_19961,N_16569,N_17022);
or U19962 (N_19962,N_13218,N_13889);
xnor U19963 (N_19963,N_12511,N_18013);
nand U19964 (N_19964,N_18335,N_16996);
and U19965 (N_19965,N_17481,N_17114);
nand U19966 (N_19966,N_18286,N_16830);
xnor U19967 (N_19967,N_18292,N_14261);
xor U19968 (N_19968,N_14009,N_17008);
and U19969 (N_19969,N_18453,N_16920);
or U19970 (N_19970,N_15774,N_18331);
and U19971 (N_19971,N_18272,N_15079);
nor U19972 (N_19972,N_14547,N_14252);
nand U19973 (N_19973,N_18432,N_16251);
nor U19974 (N_19974,N_13369,N_17039);
or U19975 (N_19975,N_12729,N_18210);
or U19976 (N_19976,N_12932,N_14256);
nor U19977 (N_19977,N_13238,N_13348);
or U19978 (N_19978,N_18494,N_17402);
xor U19979 (N_19979,N_16246,N_18741);
nand U19980 (N_19980,N_17723,N_13516);
nand U19981 (N_19981,N_13475,N_16472);
and U19982 (N_19982,N_14429,N_16801);
or U19983 (N_19983,N_13149,N_17948);
and U19984 (N_19984,N_13367,N_15397);
or U19985 (N_19985,N_15101,N_14160);
or U19986 (N_19986,N_13019,N_12507);
or U19987 (N_19987,N_14036,N_15651);
nand U19988 (N_19988,N_15685,N_17785);
nor U19989 (N_19989,N_17608,N_13684);
and U19990 (N_19990,N_12763,N_13999);
nand U19991 (N_19991,N_13334,N_13361);
or U19992 (N_19992,N_13870,N_12895);
xor U19993 (N_19993,N_13001,N_14136);
or U19994 (N_19994,N_16740,N_14054);
nor U19995 (N_19995,N_15209,N_17477);
xor U19996 (N_19996,N_17685,N_17517);
and U19997 (N_19997,N_16642,N_14380);
xor U19998 (N_19998,N_17929,N_18103);
or U19999 (N_19999,N_15499,N_13383);
xor U20000 (N_20000,N_15246,N_16876);
nor U20001 (N_20001,N_14177,N_15947);
nor U20002 (N_20002,N_17668,N_16625);
or U20003 (N_20003,N_13849,N_12649);
and U20004 (N_20004,N_17445,N_13224);
nor U20005 (N_20005,N_14444,N_14270);
xnor U20006 (N_20006,N_18019,N_14255);
xnor U20007 (N_20007,N_12528,N_18390);
and U20008 (N_20008,N_12558,N_18225);
and U20009 (N_20009,N_18039,N_15867);
nand U20010 (N_20010,N_16285,N_14536);
or U20011 (N_20011,N_16783,N_14718);
or U20012 (N_20012,N_15092,N_13279);
nand U20013 (N_20013,N_15390,N_13728);
and U20014 (N_20014,N_16382,N_18414);
xnor U20015 (N_20015,N_13185,N_14453);
and U20016 (N_20016,N_15976,N_13386);
xnor U20017 (N_20017,N_12655,N_14535);
nand U20018 (N_20018,N_14897,N_16396);
xnor U20019 (N_20019,N_12503,N_13941);
nor U20020 (N_20020,N_17146,N_15985);
nand U20021 (N_20021,N_15215,N_16963);
and U20022 (N_20022,N_13607,N_12770);
or U20023 (N_20023,N_16036,N_18036);
nand U20024 (N_20024,N_18193,N_17216);
or U20025 (N_20025,N_13875,N_16316);
xor U20026 (N_20026,N_13645,N_13133);
nor U20027 (N_20027,N_15159,N_17665);
and U20028 (N_20028,N_13270,N_13939);
nor U20029 (N_20029,N_15438,N_18533);
nand U20030 (N_20030,N_13180,N_17100);
or U20031 (N_20031,N_18422,N_14640);
or U20032 (N_20032,N_13738,N_16790);
and U20033 (N_20033,N_17592,N_15193);
nand U20034 (N_20034,N_15206,N_16687);
nor U20035 (N_20035,N_18338,N_14452);
or U20036 (N_20036,N_12688,N_17663);
nand U20037 (N_20037,N_13343,N_13017);
xnor U20038 (N_20038,N_12995,N_13771);
or U20039 (N_20039,N_16046,N_14928);
and U20040 (N_20040,N_16208,N_13530);
and U20041 (N_20041,N_13585,N_15280);
or U20042 (N_20042,N_17164,N_15188);
or U20043 (N_20043,N_16258,N_15352);
and U20044 (N_20044,N_17415,N_18318);
xnor U20045 (N_20045,N_13197,N_16268);
nor U20046 (N_20046,N_16975,N_14096);
xor U20047 (N_20047,N_14152,N_15054);
or U20048 (N_20048,N_17515,N_14413);
and U20049 (N_20049,N_13783,N_12938);
or U20050 (N_20050,N_12974,N_18313);
nand U20051 (N_20051,N_18240,N_17092);
nand U20052 (N_20052,N_12914,N_14598);
xnor U20053 (N_20053,N_16839,N_18345);
xnor U20054 (N_20054,N_16864,N_12647);
or U20055 (N_20055,N_14986,N_17262);
nand U20056 (N_20056,N_14289,N_17438);
xor U20057 (N_20057,N_13525,N_17375);
nor U20058 (N_20058,N_14519,N_13920);
nand U20059 (N_20059,N_14078,N_14568);
xor U20060 (N_20060,N_17871,N_14406);
and U20061 (N_20061,N_17907,N_13724);
nand U20062 (N_20062,N_18632,N_18619);
and U20063 (N_20063,N_18724,N_14335);
nor U20064 (N_20064,N_14763,N_12925);
nor U20065 (N_20065,N_13915,N_14644);
xnor U20066 (N_20066,N_18072,N_17813);
nand U20067 (N_20067,N_16269,N_15574);
xor U20068 (N_20068,N_15590,N_16841);
and U20069 (N_20069,N_17657,N_16074);
and U20070 (N_20070,N_12620,N_17310);
nand U20071 (N_20071,N_14127,N_16523);
xor U20072 (N_20072,N_18096,N_13832);
nor U20073 (N_20073,N_17733,N_14396);
or U20074 (N_20074,N_16501,N_14142);
and U20075 (N_20075,N_12636,N_13874);
or U20076 (N_20076,N_17103,N_17244);
and U20077 (N_20077,N_12621,N_16138);
nand U20078 (N_20078,N_16392,N_17811);
and U20079 (N_20079,N_18430,N_16389);
or U20080 (N_20080,N_17327,N_17742);
nand U20081 (N_20081,N_15207,N_15387);
or U20082 (N_20082,N_17580,N_13958);
nand U20083 (N_20083,N_17600,N_16478);
nand U20084 (N_20084,N_17732,N_16474);
xor U20085 (N_20085,N_15302,N_14609);
xnor U20086 (N_20086,N_12798,N_18281);
or U20087 (N_20087,N_18337,N_12582);
xnor U20088 (N_20088,N_16177,N_16604);
nand U20089 (N_20089,N_13564,N_15364);
nand U20090 (N_20090,N_15996,N_18671);
or U20091 (N_20091,N_14191,N_12859);
xor U20092 (N_20092,N_15888,N_15856);
xnor U20093 (N_20093,N_17978,N_13201);
xnor U20094 (N_20094,N_15042,N_13211);
nand U20095 (N_20095,N_17564,N_16578);
and U20096 (N_20096,N_13481,N_14840);
nor U20097 (N_20097,N_16889,N_12961);
xor U20098 (N_20098,N_13219,N_12863);
nand U20099 (N_20099,N_16899,N_14574);
nor U20100 (N_20100,N_17242,N_17932);
nor U20101 (N_20101,N_17373,N_16124);
and U20102 (N_20102,N_17427,N_17219);
and U20103 (N_20103,N_17788,N_12989);
and U20104 (N_20104,N_14780,N_17826);
nand U20105 (N_20105,N_13005,N_16789);
nand U20106 (N_20106,N_17400,N_17728);
nand U20107 (N_20107,N_18288,N_18001);
nand U20108 (N_20108,N_14912,N_15455);
or U20109 (N_20109,N_17928,N_15757);
or U20110 (N_20110,N_16095,N_16026);
and U20111 (N_20111,N_15489,N_13418);
and U20112 (N_20112,N_15840,N_15099);
or U20113 (N_20113,N_13409,N_13555);
xor U20114 (N_20114,N_16629,N_16469);
or U20115 (N_20115,N_14689,N_18553);
nor U20116 (N_20116,N_13847,N_16541);
nor U20117 (N_20117,N_14990,N_13286);
and U20118 (N_20118,N_15999,N_16312);
nand U20119 (N_20119,N_13490,N_14814);
nand U20120 (N_20120,N_14264,N_17604);
or U20121 (N_20121,N_16191,N_15335);
and U20122 (N_20122,N_15324,N_14522);
nor U20123 (N_20123,N_16136,N_16300);
nand U20124 (N_20124,N_13059,N_12682);
nor U20125 (N_20125,N_14695,N_17288);
nand U20126 (N_20126,N_13282,N_12959);
nand U20127 (N_20127,N_13595,N_12680);
nand U20128 (N_20128,N_18245,N_12628);
nor U20129 (N_20129,N_14583,N_16357);
nand U20130 (N_20130,N_18161,N_15254);
nor U20131 (N_20131,N_17152,N_16217);
xnor U20132 (N_20132,N_14494,N_17780);
or U20133 (N_20133,N_16649,N_18507);
nor U20134 (N_20134,N_13305,N_15150);
nor U20135 (N_20135,N_15433,N_18209);
nand U20136 (N_20136,N_13610,N_16978);
and U20137 (N_20137,N_13189,N_17832);
nand U20138 (N_20138,N_18092,N_18423);
xnor U20139 (N_20139,N_15737,N_18570);
or U20140 (N_20140,N_18150,N_12671);
nor U20141 (N_20141,N_12952,N_13195);
and U20142 (N_20142,N_17158,N_16281);
or U20143 (N_20143,N_13582,N_14630);
nand U20144 (N_20144,N_13782,N_15941);
nand U20145 (N_20145,N_16214,N_12557);
nor U20146 (N_20146,N_13067,N_18738);
nor U20147 (N_20147,N_14450,N_17222);
or U20148 (N_20148,N_13082,N_15742);
xnor U20149 (N_20149,N_12712,N_14117);
nand U20150 (N_20150,N_14552,N_17448);
nor U20151 (N_20151,N_16821,N_15661);
nand U20152 (N_20152,N_17435,N_17594);
or U20153 (N_20153,N_18410,N_16665);
nor U20154 (N_20154,N_16640,N_13615);
xnor U20155 (N_20155,N_13735,N_17391);
or U20156 (N_20156,N_13580,N_15050);
nand U20157 (N_20157,N_17556,N_16648);
nand U20158 (N_20158,N_16388,N_17658);
nor U20159 (N_20159,N_13956,N_17224);
or U20160 (N_20160,N_15717,N_18114);
xnor U20161 (N_20161,N_13038,N_15522);
and U20162 (N_20162,N_18094,N_13904);
nand U20163 (N_20163,N_15002,N_13694);
xnor U20164 (N_20164,N_14972,N_18169);
xor U20165 (N_20165,N_16012,N_17843);
or U20166 (N_20166,N_17726,N_14660);
and U20167 (N_20167,N_18123,N_15135);
nand U20168 (N_20168,N_16207,N_17968);
or U20169 (N_20169,N_13665,N_12553);
nor U20170 (N_20170,N_15736,N_15598);
or U20171 (N_20171,N_16773,N_15139);
nor U20172 (N_20172,N_17672,N_15410);
nor U20173 (N_20173,N_17345,N_13372);
nor U20174 (N_20174,N_15690,N_14144);
xnor U20175 (N_20175,N_18266,N_15670);
xnor U20176 (N_20176,N_18587,N_16104);
nand U20177 (N_20177,N_13401,N_14145);
nor U20178 (N_20178,N_13183,N_16222);
and U20179 (N_20179,N_15431,N_17712);
nand U20180 (N_20180,N_13571,N_14210);
and U20181 (N_20181,N_16205,N_17625);
xor U20182 (N_20182,N_18066,N_17697);
nor U20183 (N_20183,N_13852,N_15931);
xnor U20184 (N_20184,N_13629,N_13196);
nor U20185 (N_20185,N_12813,N_16702);
xor U20186 (N_20186,N_17899,N_18126);
or U20187 (N_20187,N_18333,N_12796);
or U20188 (N_20188,N_15373,N_15569);
nand U20189 (N_20189,N_13860,N_14898);
nand U20190 (N_20190,N_15761,N_13013);
nand U20191 (N_20191,N_16981,N_16900);
or U20192 (N_20192,N_13106,N_12690);
nand U20193 (N_20193,N_15450,N_16308);
xnor U20194 (N_20194,N_16903,N_13089);
and U20195 (N_20195,N_15017,N_15603);
nand U20196 (N_20196,N_14211,N_13663);
xnor U20197 (N_20197,N_13245,N_12645);
nor U20198 (N_20198,N_13907,N_18590);
nor U20199 (N_20199,N_14768,N_14958);
nor U20200 (N_20200,N_15331,N_18519);
and U20201 (N_20201,N_15993,N_13380);
nand U20202 (N_20202,N_12985,N_15734);
and U20203 (N_20203,N_17476,N_17828);
nor U20204 (N_20204,N_18330,N_17194);
xor U20205 (N_20205,N_13561,N_15419);
xnor U20206 (N_20206,N_13975,N_13546);
and U20207 (N_20207,N_17430,N_18449);
xor U20208 (N_20208,N_16925,N_18158);
xor U20209 (N_20209,N_14738,N_16109);
and U20210 (N_20210,N_17007,N_17997);
or U20211 (N_20211,N_16948,N_13539);
or U20212 (N_20212,N_17917,N_17318);
nand U20213 (N_20213,N_14199,N_15080);
nor U20214 (N_20214,N_14451,N_12720);
or U20215 (N_20215,N_16950,N_14474);
and U20216 (N_20216,N_16676,N_15990);
and U20217 (N_20217,N_14438,N_16912);
xor U20218 (N_20218,N_16327,N_14066);
and U20219 (N_20219,N_14895,N_15934);
nor U20220 (N_20220,N_17469,N_17220);
nand U20221 (N_20221,N_12613,N_17475);
nor U20222 (N_20222,N_17371,N_12929);
xor U20223 (N_20223,N_15361,N_13675);
and U20224 (N_20224,N_14686,N_15903);
or U20225 (N_20225,N_12853,N_18481);
and U20226 (N_20226,N_18028,N_18249);
and U20227 (N_20227,N_13751,N_13455);
and U20228 (N_20228,N_12827,N_15620);
nand U20229 (N_20229,N_16936,N_13420);
or U20230 (N_20230,N_16162,N_17393);
xnor U20231 (N_20231,N_12759,N_13021);
xnor U20232 (N_20232,N_17951,N_15667);
nand U20233 (N_20233,N_16922,N_17010);
and U20234 (N_20234,N_16662,N_12663);
or U20235 (N_20235,N_13672,N_13391);
or U20236 (N_20236,N_18244,N_13862);
nor U20237 (N_20237,N_14468,N_13887);
or U20238 (N_20238,N_15292,N_17599);
nor U20239 (N_20239,N_14508,N_13039);
or U20240 (N_20240,N_15369,N_18478);
nor U20241 (N_20241,N_16511,N_16293);
xnor U20242 (N_20242,N_15097,N_12902);
or U20243 (N_20243,N_17484,N_18254);
xnor U20244 (N_20244,N_13673,N_13573);
nand U20245 (N_20245,N_14172,N_13301);
xnor U20246 (N_20246,N_15770,N_16567);
xor U20247 (N_20247,N_17632,N_14083);
and U20248 (N_20248,N_15553,N_14222);
nor U20249 (N_20249,N_12615,N_13698);
nor U20250 (N_20250,N_15926,N_16621);
or U20251 (N_20251,N_16351,N_12889);
nor U20252 (N_20252,N_14791,N_14337);
nor U20253 (N_20253,N_15263,N_18636);
nor U20254 (N_20254,N_17709,N_15869);
and U20255 (N_20255,N_14579,N_18371);
nand U20256 (N_20256,N_16816,N_14908);
nand U20257 (N_20257,N_17654,N_14615);
xnor U20258 (N_20258,N_15100,N_18264);
nor U20259 (N_20259,N_14510,N_14657);
or U20260 (N_20260,N_15607,N_16418);
or U20261 (N_20261,N_15558,N_15623);
and U20262 (N_20262,N_12975,N_15915);
nor U20263 (N_20263,N_16872,N_15668);
nor U20264 (N_20264,N_16110,N_17790);
or U20265 (N_20265,N_17441,N_17563);
nor U20266 (N_20266,N_14682,N_16512);
and U20267 (N_20267,N_14295,N_18051);
and U20268 (N_20268,N_18534,N_17059);
xnor U20269 (N_20269,N_15776,N_18663);
nor U20270 (N_20270,N_17713,N_15095);
nand U20271 (N_20271,N_17867,N_18688);
xor U20272 (N_20272,N_16671,N_15654);
nor U20273 (N_20273,N_14781,N_15167);
nand U20274 (N_20274,N_16211,N_16048);
nand U20275 (N_20275,N_16324,N_17738);
nand U20276 (N_20276,N_15998,N_13387);
nor U20277 (N_20277,N_17629,N_14308);
xor U20278 (N_20278,N_16956,N_15721);
nor U20279 (N_20279,N_14899,N_13308);
or U20280 (N_20280,N_14467,N_15849);
nand U20281 (N_20281,N_17649,N_17138);
nor U20282 (N_20282,N_12756,N_13495);
nor U20283 (N_20283,N_17511,N_16998);
nand U20284 (N_20284,N_12806,N_12694);
and U20285 (N_20285,N_18427,N_16692);
and U20286 (N_20286,N_13588,N_17017);
nand U20287 (N_20287,N_15250,N_13621);
nor U20288 (N_20288,N_15527,N_16757);
nor U20289 (N_20289,N_13042,N_13205);
xor U20290 (N_20290,N_17909,N_15766);
nor U20291 (N_20291,N_17198,N_18742);
and U20292 (N_20292,N_13296,N_15143);
xor U20293 (N_20293,N_15141,N_15036);
or U20294 (N_20294,N_18156,N_15805);
nor U20295 (N_20295,N_14431,N_15647);
and U20296 (N_20296,N_17639,N_17729);
or U20297 (N_20297,N_13469,N_16458);
and U20298 (N_20298,N_17258,N_18597);
and U20299 (N_20299,N_18242,N_13758);
nor U20300 (N_20300,N_18246,N_15072);
nand U20301 (N_20301,N_14027,N_17278);
or U20302 (N_20302,N_17779,N_15551);
nor U20303 (N_20303,N_12778,N_16641);
nor U20304 (N_20304,N_14487,N_16038);
or U20305 (N_20305,N_15020,N_14524);
and U20306 (N_20306,N_13054,N_17996);
or U20307 (N_20307,N_13281,N_12832);
nand U20308 (N_20308,N_16793,N_14544);
xor U20309 (N_20309,N_16755,N_17701);
or U20310 (N_20310,N_17109,N_17831);
or U20311 (N_20311,N_12750,N_17372);
or U20312 (N_20312,N_18666,N_16113);
and U20313 (N_20313,N_16438,N_13008);
or U20314 (N_20314,N_13664,N_18712);
nor U20315 (N_20315,N_15045,N_14488);
nand U20316 (N_20316,N_14146,N_17256);
and U20317 (N_20317,N_14129,N_14521);
and U20318 (N_20318,N_13865,N_14854);
xnor U20319 (N_20319,N_17246,N_15604);
xor U20320 (N_20320,N_14006,N_17280);
nor U20321 (N_20321,N_18581,N_16060);
and U20322 (N_20322,N_14813,N_13800);
xor U20323 (N_20323,N_13229,N_12928);
nor U20324 (N_20324,N_18441,N_18021);
xor U20325 (N_20325,N_14707,N_12685);
nor U20326 (N_20326,N_18166,N_15927);
nor U20327 (N_20327,N_12634,N_13338);
nand U20328 (N_20328,N_12882,N_18299);
nor U20329 (N_20329,N_18582,N_16762);
or U20330 (N_20330,N_12935,N_16533);
and U20331 (N_20331,N_18654,N_15138);
nand U20332 (N_20332,N_13030,N_16347);
nor U20333 (N_20333,N_18065,N_13737);
nor U20334 (N_20334,N_14890,N_12771);
and U20335 (N_20335,N_17277,N_17466);
and U20336 (N_20336,N_15447,N_16828);
and U20337 (N_20337,N_18705,N_16844);
nand U20338 (N_20338,N_18530,N_13520);
and U20339 (N_20339,N_17532,N_15434);
and U20340 (N_20340,N_16731,N_14829);
nor U20341 (N_20341,N_15181,N_16096);
nor U20342 (N_20342,N_14723,N_15729);
or U20343 (N_20343,N_14279,N_18499);
nor U20344 (N_20344,N_13044,N_18142);
nor U20345 (N_20345,N_18300,N_15363);
or U20346 (N_20346,N_14385,N_17940);
nor U20347 (N_20347,N_15564,N_14688);
nor U20348 (N_20348,N_13830,N_17283);
or U20349 (N_20349,N_17850,N_14828);
nand U20350 (N_20350,N_13289,N_15940);
nand U20351 (N_20351,N_14236,N_17974);
xnor U20352 (N_20352,N_13015,N_15037);
nand U20353 (N_20353,N_18444,N_13993);
nand U20354 (N_20354,N_17925,N_14075);
nand U20355 (N_20355,N_13677,N_13480);
nor U20356 (N_20356,N_16001,N_13257);
xnor U20357 (N_20357,N_16957,N_17973);
nand U20358 (N_20358,N_13628,N_13701);
nor U20359 (N_20359,N_13773,N_17263);
nor U20360 (N_20360,N_13709,N_14088);
nand U20361 (N_20361,N_13307,N_13942);
nand U20362 (N_20362,N_16548,N_17213);
or U20363 (N_20363,N_16155,N_16328);
and U20364 (N_20364,N_14968,N_15498);
or U20365 (N_20365,N_15921,N_14482);
nor U20366 (N_20366,N_14933,N_14262);
nand U20367 (N_20367,N_18026,N_13142);
or U20368 (N_20368,N_15584,N_14203);
nor U20369 (N_20369,N_18024,N_12660);
nand U20370 (N_20370,N_16326,N_16363);
nand U20371 (N_20371,N_16562,N_17311);
nand U20372 (N_20372,N_17568,N_16317);
nand U20373 (N_20373,N_16901,N_12768);
or U20374 (N_20374,N_14684,N_13458);
nor U20375 (N_20375,N_18258,N_14856);
or U20376 (N_20376,N_16603,N_15235);
or U20377 (N_20377,N_14250,N_15669);
xor U20378 (N_20378,N_16540,N_16486);
nand U20379 (N_20379,N_15500,N_14393);
or U20380 (N_20380,N_14260,N_14619);
nand U20381 (N_20381,N_18378,N_14275);
or U20382 (N_20382,N_16455,N_13651);
nand U20383 (N_20383,N_15887,N_18135);
xnor U20384 (N_20384,N_14874,N_15775);
nor U20385 (N_20385,N_17066,N_16232);
nor U20386 (N_20386,N_16854,N_15832);
nand U20387 (N_20387,N_18312,N_16337);
nand U20388 (N_20388,N_15440,N_16971);
and U20389 (N_20389,N_15914,N_17491);
xor U20390 (N_20390,N_15158,N_16427);
nor U20391 (N_20391,N_13062,N_16391);
xnor U20392 (N_20392,N_18227,N_16500);
nand U20393 (N_20393,N_15594,N_16698);
or U20394 (N_20394,N_14399,N_13398);
or U20395 (N_20395,N_13394,N_13355);
xnor U20396 (N_20396,N_14458,N_16203);
and U20397 (N_20397,N_14476,N_15473);
nand U20398 (N_20398,N_14581,N_17825);
and U20399 (N_20399,N_13886,N_18546);
nand U20400 (N_20400,N_15237,N_17188);
nor U20401 (N_20401,N_15877,N_18555);
or U20402 (N_20402,N_18215,N_14062);
nand U20403 (N_20403,N_15486,N_13248);
or U20404 (N_20404,N_18251,N_18667);
nor U20405 (N_20405,N_13487,N_14001);
nand U20406 (N_20406,N_16288,N_14627);
xnor U20407 (N_20407,N_14810,N_18734);
xnor U20408 (N_20408,N_13963,N_16332);
and U20409 (N_20409,N_17125,N_15030);
nor U20410 (N_20410,N_15741,N_18617);
and U20411 (N_20411,N_13855,N_18577);
or U20412 (N_20412,N_15386,N_13947);
nand U20413 (N_20413,N_14985,N_14018);
nor U20414 (N_20414,N_15171,N_16077);
nor U20415 (N_20415,N_17976,N_16881);
xnor U20416 (N_20416,N_14939,N_16879);
nor U20417 (N_20417,N_18413,N_15338);
xnor U20418 (N_20418,N_15381,N_15839);
nand U20419 (N_20419,N_17412,N_15900);
xor U20420 (N_20420,N_13812,N_17185);
xor U20421 (N_20421,N_17562,N_16361);
nand U20422 (N_20422,N_13691,N_15883);
or U20423 (N_20423,N_15655,N_13237);
nand U20424 (N_20424,N_15179,N_18556);
or U20425 (N_20425,N_18176,N_13518);
nor U20426 (N_20426,N_17681,N_17426);
xnor U20427 (N_20427,N_17803,N_12684);
or U20428 (N_20428,N_17930,N_16572);
and U20429 (N_20429,N_15320,N_15408);
or U20430 (N_20430,N_16218,N_15550);
xor U20431 (N_20431,N_12698,N_17661);
or U20432 (N_20432,N_13864,N_13719);
and U20433 (N_20433,N_12988,N_18014);
or U20434 (N_20434,N_17037,N_13798);
nand U20435 (N_20435,N_16481,N_12555);
nor U20436 (N_20436,N_16027,N_13222);
and U20437 (N_20437,N_14785,N_17447);
or U20438 (N_20438,N_16311,N_18497);
nor U20439 (N_20439,N_18241,N_16378);
nand U20440 (N_20440,N_14769,N_16341);
nand U20441 (N_20441,N_13856,N_16122);
or U20442 (N_20442,N_13255,N_18319);
or U20443 (N_20443,N_13092,N_16873);
nor U20444 (N_20444,N_15850,N_15284);
nor U20445 (N_20445,N_15261,N_17910);
xnor U20446 (N_20446,N_13508,N_16696);
and U20447 (N_20447,N_13150,N_17464);
xor U20448 (N_20448,N_13273,N_16994);
or U20449 (N_20449,N_15201,N_13104);
or U20450 (N_20450,N_17859,N_16028);
or U20451 (N_20451,N_15066,N_17153);
xor U20452 (N_20452,N_16726,N_13596);
nand U20453 (N_20453,N_16135,N_15400);
nor U20454 (N_20454,N_15248,N_17990);
xnor U20455 (N_20455,N_17994,N_15459);
nor U20456 (N_20456,N_13523,N_13648);
or U20457 (N_20457,N_13897,N_14498);
nor U20458 (N_20458,N_15198,N_18322);
nand U20459 (N_20459,N_14212,N_17923);
xnor U20460 (N_20460,N_13479,N_15274);
or U20461 (N_20461,N_17543,N_13655);
nand U20462 (N_20462,N_18200,N_15132);
or U20463 (N_20463,N_16943,N_13113);
xnor U20464 (N_20464,N_14011,N_13177);
nand U20465 (N_20465,N_18388,N_16193);
nor U20466 (N_20466,N_16336,N_16319);
xor U20467 (N_20467,N_13310,N_14436);
or U20468 (N_20468,N_14724,N_14783);
nor U20469 (N_20469,N_16020,N_16150);
nor U20470 (N_20470,N_14194,N_13225);
or U20471 (N_20471,N_16623,N_17320);
nand U20472 (N_20472,N_15040,N_18512);
nor U20473 (N_20473,N_14084,N_12991);
nor U20474 (N_20474,N_15980,N_13829);
or U20475 (N_20475,N_17510,N_17616);
nand U20476 (N_20476,N_17880,N_12793);
nand U20477 (N_20477,N_15763,N_16147);
nand U20478 (N_20478,N_17060,N_14060);
nand U20479 (N_20479,N_14175,N_17492);
or U20480 (N_20480,N_12811,N_16597);
nor U20481 (N_20481,N_13249,N_12653);
xor U20482 (N_20482,N_16907,N_14834);
xnor U20483 (N_20483,N_15196,N_15124);
nor U20484 (N_20484,N_14224,N_16522);
nand U20485 (N_20485,N_15172,N_15199);
nand U20486 (N_20486,N_16358,N_18591);
xor U20487 (N_20487,N_15982,N_16720);
and U20488 (N_20488,N_14360,N_15644);
xnor U20489 (N_20489,N_15360,N_15547);
nor U20490 (N_20490,N_14651,N_13412);
nand U20491 (N_20491,N_17036,N_13869);
and U20492 (N_20492,N_15088,N_12965);
xor U20493 (N_20493,N_15692,N_15724);
or U20494 (N_20494,N_17703,N_18070);
nand U20495 (N_20495,N_13488,N_14281);
nor U20496 (N_20496,N_17954,N_12508);
and U20497 (N_20497,N_17489,N_18137);
nor U20498 (N_20498,N_13138,N_15893);
xnor U20499 (N_20499,N_13352,N_15501);
or U20500 (N_20500,N_18697,N_13204);
nand U20501 (N_20501,N_13879,N_16632);
or U20502 (N_20502,N_12631,N_12915);
xor U20503 (N_20503,N_16239,N_14871);
and U20504 (N_20504,N_16399,N_16588);
nor U20505 (N_20505,N_16633,N_14604);
or U20506 (N_20506,N_18733,N_16574);
xor U20507 (N_20507,N_16333,N_15393);
nand U20508 (N_20508,N_16896,N_14318);
nor U20509 (N_20509,N_16792,N_16058);
xor U20510 (N_20510,N_14143,N_18580);
nor U20511 (N_20511,N_14268,N_14621);
nor U20512 (N_20512,N_14115,N_17545);
nand U20513 (N_20513,N_18695,N_17019);
nand U20514 (N_20514,N_14788,N_15372);
or U20515 (N_20515,N_13342,N_13473);
xor U20516 (N_20516,N_12812,N_13746);
xor U20517 (N_20517,N_18068,N_14775);
xnor U20518 (N_20518,N_15075,N_17892);
and U20519 (N_20519,N_14400,N_14063);
nand U20520 (N_20520,N_13814,N_14865);
and U20521 (N_20521,N_18170,N_17897);
or U20522 (N_20522,N_14437,N_14733);
xnor U20523 (N_20523,N_13095,N_18192);
xnor U20524 (N_20524,N_18261,N_17540);
nor U20525 (N_20525,N_14297,N_15713);
or U20526 (N_20526,N_16927,N_15919);
xnor U20527 (N_20527,N_15819,N_16699);
and U20528 (N_20528,N_15368,N_16999);
and U20529 (N_20529,N_16739,N_17512);
and U20530 (N_20530,N_17323,N_13914);
and U20531 (N_20531,N_14893,N_13178);
nand U20532 (N_20532,N_16129,N_12624);
nor U20533 (N_20533,N_15334,N_18031);
and U20534 (N_20534,N_17254,N_15074);
nor U20535 (N_20535,N_17711,N_16919);
xnor U20536 (N_20536,N_12713,N_15047);
nand U20537 (N_20537,N_14831,N_18516);
or U20538 (N_20538,N_14361,N_15063);
xnor U20539 (N_20539,N_12580,N_15039);
or U20540 (N_20540,N_12584,N_13631);
and U20541 (N_20541,N_13298,N_16141);
xor U20542 (N_20542,N_16991,N_16263);
nor U20543 (N_20543,N_18689,N_16855);
and U20544 (N_20544,N_13670,N_17062);
nand U20545 (N_20545,N_18165,N_18291);
or U20546 (N_20546,N_13115,N_18737);
nor U20547 (N_20547,N_12674,N_13642);
xnor U20548 (N_20548,N_18460,N_14556);
and U20549 (N_20549,N_18059,N_14685);
nand U20550 (N_20550,N_13972,N_16061);
and U20551 (N_20551,N_14904,N_12924);
and U20552 (N_20552,N_14331,N_13605);
nand U20553 (N_20553,N_18111,N_15269);
nand U20554 (N_20554,N_16862,N_14414);
and U20555 (N_20555,N_13432,N_14333);
or U20556 (N_20556,N_17636,N_16107);
or U20557 (N_20557,N_14013,N_14816);
nor U20558 (N_20558,N_16601,N_18226);
nor U20559 (N_20559,N_12521,N_13033);
nand U20560 (N_20560,N_17596,N_12852);
or U20561 (N_20561,N_17615,N_14381);
nand U20562 (N_20562,N_17977,N_16608);
or U20563 (N_20563,N_13794,N_18387);
or U20564 (N_20564,N_14670,N_18063);
and U20565 (N_20565,N_17003,N_16539);
xor U20566 (N_20566,N_14629,N_18699);
nand U20567 (N_20567,N_15318,N_16270);
nor U20568 (N_20568,N_17381,N_16277);
nand U20569 (N_20569,N_16535,N_17758);
nor U20570 (N_20570,N_16818,N_13846);
nor U20571 (N_20571,N_18029,N_17521);
xnor U20572 (N_20572,N_16451,N_15715);
or U20573 (N_20573,N_17595,N_17417);
or U20574 (N_20574,N_17747,N_15327);
xnor U20575 (N_20575,N_18328,N_14839);
and U20576 (N_20576,N_14843,N_17349);
nor U20577 (N_20577,N_17769,N_18282);
and U20578 (N_20578,N_13451,N_14267);
nand U20579 (N_20579,N_14957,N_13916);
or U20580 (N_20580,N_16795,N_14632);
or U20581 (N_20581,N_17638,N_16099);
xor U20582 (N_20582,N_13187,N_13341);
or U20583 (N_20583,N_13890,N_14765);
and U20584 (N_20584,N_16372,N_14539);
or U20585 (N_20585,N_14002,N_14089);
nand U20586 (N_20586,N_14269,N_14823);
xnor U20587 (N_20587,N_15904,N_18626);
or U20588 (N_20588,N_18451,N_15580);
nor U20589 (N_20589,N_13873,N_13402);
and U20590 (N_20590,N_14562,N_14107);
and U20591 (N_20591,N_13593,N_16771);
xor U20592 (N_20592,N_15300,N_15383);
and U20593 (N_20593,N_14954,N_17801);
or U20594 (N_20594,N_13576,N_17534);
xnor U20595 (N_20595,N_13928,N_16010);
or U20596 (N_20596,N_15205,N_12565);
or U20597 (N_20597,N_15321,N_13844);
and U20598 (N_20598,N_17884,N_14307);
nor U20599 (N_20599,N_16753,N_17237);
or U20600 (N_20600,N_15636,N_18438);
nand U20601 (N_20601,N_18145,N_14694);
nor U20602 (N_20602,N_16532,N_12888);
nand U20603 (N_20603,N_13336,N_17027);
nor U20604 (N_20604,N_17030,N_14546);
nor U20605 (N_20605,N_17830,N_18609);
nor U20606 (N_20606,N_18057,N_17395);
nand U20607 (N_20607,N_15509,N_12797);
nand U20608 (N_20608,N_17583,N_14379);
xnor U20609 (N_20609,N_13951,N_17602);
xor U20610 (N_20610,N_15347,N_13581);
nor U20611 (N_20611,N_15395,N_14480);
and U20612 (N_20612,N_13036,N_14052);
nor U20613 (N_20613,N_14786,N_12616);
nand U20614 (N_20614,N_18684,N_13747);
xnor U20615 (N_20615,N_14398,N_14923);
nand U20616 (N_20616,N_13982,N_16554);
or U20617 (N_20617,N_17351,N_15169);
and U20618 (N_20618,N_18747,N_16897);
nand U20619 (N_20619,N_18190,N_16808);
nor U20620 (N_20620,N_14249,N_14922);
or U20621 (N_20621,N_16367,N_15190);
or U20622 (N_20622,N_14010,N_12822);
and U20623 (N_20623,N_15337,N_13682);
nand U20624 (N_20624,N_17898,N_13404);
nor U20625 (N_20625,N_14983,N_12602);
xor U20626 (N_20626,N_14022,N_13320);
xnor U20627 (N_20627,N_14864,N_14646);
and U20628 (N_20628,N_12912,N_16634);
and U20629 (N_20629,N_17134,N_17233);
and U20630 (N_20630,N_14108,N_17810);
and U20631 (N_20631,N_14748,N_17557);
xor U20632 (N_20632,N_15797,N_17756);
and U20633 (N_20633,N_12719,N_15216);
or U20634 (N_20634,N_14792,N_15011);
nand U20635 (N_20635,N_14641,N_14067);
nor U20636 (N_20636,N_16184,N_13917);
or U20637 (N_20637,N_15107,N_13323);
nor U20638 (N_20638,N_17143,N_12891);
nor U20639 (N_20639,N_16905,N_14004);
xnor U20640 (N_20640,N_14757,N_14073);
and U20641 (N_20641,N_13470,N_15653);
nor U20642 (N_20642,N_15414,N_15666);
xor U20643 (N_20643,N_13315,N_14969);
nand U20644 (N_20644,N_17651,N_16309);
nand U20645 (N_20645,N_14427,N_12548);
and U20646 (N_20646,N_16160,N_13124);
and U20647 (N_20647,N_15035,N_16303);
nand U20648 (N_20648,N_14059,N_18107);
xnor U20649 (N_20649,N_17741,N_16123);
and U20650 (N_20650,N_16514,N_15460);
and U20651 (N_20651,N_16585,N_13408);
xor U20652 (N_20652,N_14155,N_13122);
xor U20653 (N_20653,N_16838,N_13839);
nor U20654 (N_20654,N_18668,N_18571);
or U20655 (N_20655,N_13031,N_12998);
and U20656 (N_20656,N_16718,N_13247);
xnor U20657 (N_20657,N_17946,N_15476);
and U20658 (N_20658,N_15628,N_13768);
and U20659 (N_20659,N_17196,N_15504);
nor U20660 (N_20660,N_16985,N_17121);
nor U20661 (N_20661,N_14114,N_15785);
xor U20662 (N_20662,N_13721,N_12714);
xnor U20663 (N_20663,N_15853,N_14678);
and U20664 (N_20664,N_16939,N_18455);
xor U20665 (N_20665,N_15549,N_17936);
nor U20666 (N_20666,N_13366,N_16837);
xor U20667 (N_20667,N_16190,N_16916);
or U20668 (N_20668,N_14366,N_12575);
and U20669 (N_20669,N_15846,N_14280);
and U20670 (N_20670,N_13612,N_15897);
xnor U20671 (N_20671,N_16172,N_15963);
nand U20672 (N_20672,N_16747,N_15065);
xor U20673 (N_20673,N_18098,N_15923);
nor U20674 (N_20674,N_16255,N_13630);
nor U20675 (N_20675,N_14716,N_17857);
nor U20676 (N_20676,N_18564,N_18352);
nand U20677 (N_20677,N_16125,N_15723);
xnor U20678 (N_20678,N_18468,N_13075);
nand U20679 (N_20679,N_15048,N_18294);
and U20680 (N_20680,N_13118,N_17151);
xnor U20681 (N_20681,N_12585,N_17259);
xor U20682 (N_20682,N_15214,N_13216);
nand U20683 (N_20683,N_13594,N_15314);
or U20684 (N_20684,N_15147,N_17418);
and U20685 (N_20685,N_17366,N_16016);
nor U20686 (N_20686,N_17820,N_18539);
nor U20687 (N_20687,N_16679,N_15634);
or U20688 (N_20688,N_15465,N_15649);
nor U20689 (N_20689,N_12803,N_12512);
nand U20690 (N_20690,N_12676,N_15777);
or U20691 (N_20691,N_15136,N_17696);
and U20692 (N_20692,N_14971,N_16787);
nor U20693 (N_20693,N_13527,N_14169);
and U20694 (N_20694,N_17550,N_17012);
nand U20695 (N_20695,N_15680,N_14042);
or U20696 (N_20696,N_15451,N_17204);
or U20697 (N_20697,N_15589,N_13934);
nand U20698 (N_20698,N_15336,N_17139);
nor U20699 (N_20699,N_12816,N_14326);
and U20700 (N_20700,N_15844,N_14248);
nor U20701 (N_20701,N_14507,N_15053);
nor U20702 (N_20702,N_13764,N_14304);
and U20703 (N_20703,N_16716,N_14889);
nor U20704 (N_20704,N_15418,N_14973);
nand U20705 (N_20705,N_13877,N_15910);
nand U20706 (N_20706,N_16318,N_14602);
or U20707 (N_20707,N_16531,N_12784);
xor U20708 (N_20708,N_14878,N_15964);
and U20709 (N_20709,N_13643,N_12946);
nand U20710 (N_20710,N_14612,N_15577);
nand U20711 (N_20711,N_15358,N_15782);
or U20712 (N_20712,N_17642,N_14755);
xnor U20713 (N_20713,N_16937,N_15441);
and U20714 (N_20714,N_17044,N_17384);
xnor U20715 (N_20715,N_16019,N_18213);
or U20716 (N_20716,N_13911,N_17199);
nor U20717 (N_20717,N_13186,N_18673);
xnor U20718 (N_20718,N_13392,N_16267);
xnor U20719 (N_20719,N_15094,N_14068);
and U20720 (N_20720,N_16426,N_18511);
xor U20721 (N_20721,N_16491,N_15279);
or U20722 (N_20722,N_14847,N_18732);
nand U20723 (N_20723,N_15991,N_12908);
nand U20724 (N_20724,N_18119,N_12638);
nand U20725 (N_20725,N_18707,N_15694);
nor U20726 (N_20726,N_18189,N_14891);
or U20727 (N_20727,N_15703,N_13130);
nand U20728 (N_20728,N_16495,N_13801);
xnor U20729 (N_20729,N_14926,N_17862);
xnor U20730 (N_20730,N_13240,N_18631);
xor U20731 (N_20731,N_15688,N_18085);
nand U20732 (N_20732,N_14220,N_14937);
nor U20733 (N_20733,N_17032,N_16029);
nand U20734 (N_20734,N_17289,N_17087);
xor U20735 (N_20735,N_14310,N_15290);
nor U20736 (N_20736,N_18017,N_15701);
or U20737 (N_20737,N_17155,N_14057);
nor U20738 (N_20738,N_14806,N_14805);
nand U20739 (N_20739,N_16295,N_16520);
nand U20740 (N_20740,N_18273,N_14445);
and U20741 (N_20741,N_13489,N_16573);
nor U20742 (N_20742,N_16409,N_15753);
nand U20743 (N_20743,N_16797,N_14832);
nor U20744 (N_20744,N_17734,N_17108);
nor U20745 (N_20745,N_18400,N_15463);
and U20746 (N_20746,N_18569,N_18708);
or U20747 (N_20747,N_16935,N_17538);
xor U20748 (N_20748,N_13606,N_13763);
nor U20749 (N_20749,N_13259,N_16434);
xnor U20750 (N_20750,N_14426,N_12560);
xnor U20751 (N_20751,N_12618,N_14276);
xor U20752 (N_20752,N_15855,N_18554);
or U20753 (N_20753,N_13756,N_12725);
nand U20754 (N_20754,N_17799,N_18349);
nand U20755 (N_20755,N_16439,N_13824);
xnor U20756 (N_20756,N_17064,N_15128);
nor U20757 (N_20757,N_15430,N_18473);
or U20758 (N_20758,N_14332,N_14121);
nor U20759 (N_20759,N_13821,N_14378);
and U20760 (N_20760,N_15905,N_14183);
or U20761 (N_20761,N_15600,N_13777);
nand U20762 (N_20762,N_13503,N_12525);
nand U20763 (N_20763,N_14708,N_16098);
nand U20764 (N_20764,N_13045,N_15016);
and U20765 (N_20765,N_14342,N_15906);
or U20766 (N_20766,N_14637,N_17905);
nor U20767 (N_20767,N_13784,N_16717);
and U20768 (N_20768,N_18418,N_18529);
nand U20769 (N_20769,N_16954,N_14735);
nand U20770 (N_20770,N_16457,N_13318);
and U20771 (N_20771,N_18698,N_15557);
and U20772 (N_20772,N_13097,N_17290);
nor U20773 (N_20773,N_15406,N_17411);
and U20774 (N_20774,N_13809,N_17644);
nor U20775 (N_20775,N_13779,N_17963);
or U20776 (N_20776,N_18154,N_12801);
nand U20777 (N_20777,N_15339,N_15835);
nor U20778 (N_20778,N_12878,N_15581);
or U20779 (N_20779,N_18140,N_18307);
and U20780 (N_20780,N_17267,N_14178);
or U20781 (N_20781,N_15398,N_15563);
xor U20782 (N_20782,N_17104,N_17714);
nor U20783 (N_20783,N_15678,N_17573);
and U20784 (N_20784,N_13583,N_17590);
nand U20785 (N_20785,N_15380,N_16990);
xnor U20786 (N_20786,N_16624,N_13311);
xnor U20787 (N_20787,N_15323,N_17159);
nand U20788 (N_20788,N_17896,N_17902);
xor U20789 (N_20789,N_13068,N_17869);
nor U20790 (N_20790,N_17053,N_14610);
xnor U20791 (N_20791,N_15264,N_18659);
and U20792 (N_20792,N_13669,N_12731);
or U20793 (N_20793,N_15728,N_12824);
xnor U20794 (N_20794,N_16402,N_14666);
nand U20795 (N_20795,N_14432,N_15378);
xor U20796 (N_20796,N_15587,N_16130);
or U20797 (N_20797,N_14173,N_16827);
or U20798 (N_20798,N_14099,N_18101);
nand U20799 (N_20799,N_15219,N_13552);
xor U20800 (N_20800,N_13396,N_13977);
nor U20801 (N_20801,N_16804,N_14881);
nand U20802 (N_20802,N_14085,N_18236);
or U20803 (N_20803,N_16220,N_17737);
or U20804 (N_20804,N_14918,N_14216);
nor U20805 (N_20805,N_14195,N_16492);
and U20806 (N_20806,N_13099,N_17845);
nor U20807 (N_20807,N_12604,N_13440);
nand U20808 (N_20808,N_12927,N_13217);
xnor U20809 (N_20809,N_15126,N_14161);
or U20810 (N_20810,N_16777,N_18703);
nand U20811 (N_20811,N_15648,N_18464);
nand U20812 (N_20812,N_16032,N_15969);
and U20813 (N_20813,N_13474,N_12830);
nand U20814 (N_20814,N_15708,N_18493);
and U20815 (N_20815,N_18395,N_12823);
nand U20816 (N_20816,N_18265,N_17721);
nand U20817 (N_20817,N_14206,N_18736);
or U20818 (N_20818,N_15543,N_17640);
or U20819 (N_20819,N_14593,N_13994);
and U20820 (N_20820,N_14981,N_18314);
and U20821 (N_20821,N_12963,N_14303);
nand U20822 (N_20822,N_15496,N_12600);
and U20823 (N_20823,N_18044,N_15859);
or U20824 (N_20824,N_12556,N_16813);
nor U20825 (N_20825,N_15602,N_16097);
nand U20826 (N_20826,N_15779,N_13272);
nand U20827 (N_20827,N_18015,N_18208);
xnor U20828 (N_20828,N_18417,N_18402);
xor U20829 (N_20829,N_16840,N_15924);
nand U20830 (N_20830,N_15823,N_13861);
nor U20831 (N_20831,N_13284,N_14597);
xnor U20832 (N_20832,N_17271,N_18204);
nor U20833 (N_20833,N_13953,N_18479);
or U20834 (N_20834,N_16966,N_18694);
or U20835 (N_20835,N_13654,N_18048);
and U20836 (N_20836,N_13592,N_12543);
nand U20837 (N_20837,N_16967,N_15417);
and U20838 (N_20838,N_18523,N_18152);
xor U20839 (N_20839,N_14930,N_18055);
nand U20840 (N_20840,N_15475,N_12510);
and U20841 (N_20841,N_14639,N_18515);
nor U20842 (N_20842,N_14097,N_14433);
nand U20843 (N_20843,N_17031,N_15870);
or U20844 (N_20844,N_12754,N_17482);
nor U20845 (N_20845,N_15385,N_13266);
and U20846 (N_20846,N_14911,N_14563);
nand U20847 (N_20847,N_14690,N_14951);
xor U20848 (N_20848,N_14998,N_15925);
or U20849 (N_20849,N_17306,N_17775);
nand U20850 (N_20850,N_18445,N_16014);
nor U20851 (N_20851,N_14613,N_15326);
and U20852 (N_20852,N_14807,N_16775);
nand U20853 (N_20853,N_15077,N_15344);
or U20854 (N_20854,N_14106,N_15186);
and U20855 (N_20855,N_18424,N_15049);
or U20856 (N_20856,N_17101,N_13806);
or U20857 (N_20857,N_12605,N_14019);
nand U20858 (N_20858,N_17549,N_14101);
and U20859 (N_20859,N_17334,N_18384);
and U20860 (N_20860,N_14559,N_18311);
and U20861 (N_20861,N_13309,N_15749);
and U20862 (N_20862,N_12934,N_17916);
nor U20863 (N_20863,N_14848,N_17693);
xnor U20864 (N_20864,N_16004,N_14826);
or U20865 (N_20865,N_18476,N_13441);
nor U20866 (N_20866,N_18078,N_17473);
or U20867 (N_20867,N_12772,N_14112);
nand U20868 (N_20868,N_13390,N_13833);
and U20869 (N_20869,N_17763,N_16888);
or U20870 (N_20870,N_15466,N_15457);
and U20871 (N_20871,N_13477,N_13813);
or U20872 (N_20872,N_16846,N_15113);
xor U20873 (N_20873,N_13287,N_17243);
and U20874 (N_20874,N_18578,N_14093);
nand U20875 (N_20875,N_15803,N_16571);
nand U20876 (N_20876,N_16730,N_14794);
nand U20877 (N_20877,N_14365,N_15388);
xor U20878 (N_20878,N_17527,N_14214);
nor U20879 (N_20879,N_16128,N_18108);
and U20880 (N_20880,N_12821,N_15642);
nand U20881 (N_20881,N_14446,N_18730);
and U20882 (N_20882,N_16073,N_15104);
or U20883 (N_20883,N_18348,N_14469);
and U20884 (N_20884,N_13419,N_15462);
nor U20885 (N_20885,N_13535,N_16371);
and U20886 (N_20886,N_16543,N_14697);
xnor U20887 (N_20887,N_18488,N_18495);
or U20888 (N_20888,N_15325,N_18104);
nor U20889 (N_20889,N_17504,N_15437);
nand U20890 (N_20890,N_17355,N_13025);
xor U20891 (N_20891,N_17118,N_14948);
nand U20892 (N_20892,N_18235,N_15967);
or U20893 (N_20893,N_18380,N_14330);
nand U20894 (N_20894,N_14094,N_17766);
xor U20895 (N_20895,N_13330,N_15480);
and U20896 (N_20896,N_14007,N_15346);
and U20897 (N_20897,N_16479,N_16236);
xnor U20898 (N_20898,N_14050,N_18180);
and U20899 (N_20899,N_15643,N_13129);
nor U20900 (N_20900,N_13242,N_17846);
nor U20901 (N_20901,N_18721,N_18630);
nor U20902 (N_20902,N_12884,N_13757);
nand U20903 (N_20903,N_15367,N_15439);
or U20904 (N_20904,N_13687,N_13268);
and U20905 (N_20905,N_18635,N_14265);
nor U20906 (N_20906,N_17765,N_13384);
or U20907 (N_20907,N_14540,N_16706);
nand U20908 (N_20908,N_12982,N_14302);
nor U20909 (N_20909,N_14282,N_13548);
and U20910 (N_20910,N_18634,N_17295);
xor U20911 (N_20911,N_17072,N_17488);
or U20912 (N_20912,N_17090,N_16406);
and U20913 (N_20913,N_17593,N_15833);
and U20914 (N_20914,N_16094,N_18185);
and U20915 (N_20915,N_14675,N_14204);
nand U20916 (N_20916,N_15294,N_14982);
nor U20917 (N_20917,N_17269,N_13697);
or U20918 (N_20918,N_18398,N_16338);
and U20919 (N_20919,N_16168,N_16000);
xor U20920 (N_20920,N_14578,N_18551);
xor U20921 (N_20921,N_15946,N_13741);
and U20922 (N_20922,N_14464,N_12586);
nor U20923 (N_20923,N_16287,N_18508);
and U20924 (N_20924,N_13834,N_13584);
or U20925 (N_20925,N_13729,N_14244);
nand U20926 (N_20926,N_14048,N_13600);
xnor U20927 (N_20927,N_14714,N_18202);
or U20928 (N_20928,N_17680,N_16210);
nand U20929 (N_20929,N_13169,N_16663);
and U20930 (N_20930,N_16182,N_16890);
or U20931 (N_20931,N_15534,N_18377);
xnor U20932 (N_20932,N_16525,N_14638);
and U20933 (N_20933,N_15769,N_13454);
xnor U20934 (N_20934,N_17530,N_16070);
nand U20935 (N_20935,N_13065,N_14208);
xnor U20936 (N_20936,N_16480,N_18329);
and U20937 (N_20937,N_12563,N_17631);
nand U20938 (N_20938,N_12707,N_17809);
and U20939 (N_20939,N_15681,N_16546);
xor U20940 (N_20940,N_15936,N_15852);
nor U20941 (N_20941,N_14866,N_15203);
nand U20942 (N_20942,N_13422,N_13825);
nand U20943 (N_20943,N_16765,N_16398);
nand U20944 (N_20944,N_15943,N_16951);
and U20945 (N_20945,N_16362,N_14526);
and U20946 (N_20946,N_15479,N_15032);
nand U20947 (N_20947,N_17784,N_12837);
xnor U20948 (N_20948,N_15918,N_13634);
and U20949 (N_20949,N_14698,N_18420);
or U20950 (N_20950,N_17111,N_18347);
xor U20951 (N_20951,N_14200,N_15341);
or U20952 (N_20952,N_14787,N_14739);
or U20953 (N_20953,N_16157,N_17298);
and U20954 (N_20954,N_13827,N_14273);
xor U20955 (N_20955,N_12815,N_13591);
and U20956 (N_20956,N_17761,N_15487);
nand U20957 (N_20957,N_15767,N_13126);
nand U20958 (N_20958,N_16235,N_12864);
xnor U20959 (N_20959,N_15913,N_18641);
or U20960 (N_20960,N_12745,N_13676);
xor U20961 (N_20961,N_15006,N_14416);
or U20962 (N_20962,N_17541,N_13414);
nor U20963 (N_20963,N_15357,N_13511);
nor U20964 (N_20964,N_17962,N_13919);
xor U20965 (N_20965,N_17253,N_13277);
or U20966 (N_20966,N_12577,N_15345);
or U20967 (N_20967,N_18462,N_12752);
or U20968 (N_20968,N_18020,N_12977);
and U20969 (N_20969,N_12765,N_17450);
and U20970 (N_20970,N_15117,N_14118);
xnor U20971 (N_20971,N_15677,N_15266);
xor U20972 (N_20972,N_16320,N_17531);
or U20973 (N_20973,N_18653,N_14296);
or U20974 (N_20974,N_17961,N_12523);
and U20975 (N_20975,N_14636,N_13637);
xor U20976 (N_20976,N_16035,N_16664);
or U20977 (N_20977,N_14190,N_16612);
xnor U20978 (N_20978,N_12691,N_16654);
xor U20979 (N_20979,N_13979,N_14934);
nand U20980 (N_20980,N_13587,N_16314);
and U20981 (N_20981,N_12518,N_12667);
nor U20982 (N_20982,N_13285,N_15933);
nand U20983 (N_20983,N_16712,N_17833);
nor U20984 (N_20984,N_15278,N_16021);
and U20985 (N_20985,N_15111,N_14392);
nand U20986 (N_20986,N_16904,N_16487);
xor U20987 (N_20987,N_16100,N_13447);
nand U20988 (N_20988,N_18093,N_18719);
or U20989 (N_20989,N_16940,N_15445);
or U20990 (N_20990,N_18228,N_15125);
and U20991 (N_20991,N_18674,N_14196);
and U20992 (N_20992,N_15267,N_16346);
or U20993 (N_20993,N_18381,N_12761);
nand U20994 (N_20994,N_15492,N_12718);
xor U20995 (N_20995,N_15875,N_16647);
or U20996 (N_20996,N_17346,N_14770);
nand U20997 (N_20997,N_14425,N_13121);
and U20998 (N_20998,N_17414,N_15884);
xnor U20999 (N_20999,N_14606,N_12743);
nand U21000 (N_21000,N_12820,N_14603);
or U21001 (N_21001,N_13601,N_15133);
or U21002 (N_21002,N_18159,N_14321);
or U21003 (N_21003,N_13534,N_17117);
and U21004 (N_21004,N_15409,N_13893);
xnor U21005 (N_21005,N_16050,N_14192);
nand U21006 (N_21006,N_13940,N_12767);
or U21007 (N_21007,N_17986,N_17073);
xnor U21008 (N_21008,N_17548,N_16348);
or U21009 (N_21009,N_17443,N_18122);
or U21010 (N_21010,N_12527,N_13541);
or U21011 (N_21011,N_12738,N_16845);
nor U21012 (N_21012,N_12943,N_15224);
xor U21013 (N_21013,N_17883,N_15812);
xnor U21014 (N_21014,N_12942,N_17020);
xnor U21015 (N_21015,N_17248,N_17870);
nand U21016 (N_21016,N_18550,N_16527);
or U21017 (N_21017,N_16121,N_15082);
xor U21018 (N_21018,N_16224,N_12979);
xnor U21019 (N_21019,N_13162,N_17736);
and U21020 (N_21020,N_15056,N_16250);
xnor U21021 (N_21021,N_13066,N_17947);
nand U21022 (N_21022,N_13429,N_16053);
or U21023 (N_21023,N_13765,N_15041);
nor U21024 (N_21024,N_16086,N_16908);
nand U21025 (N_21025,N_12596,N_13246);
xor U21026 (N_21026,N_14041,N_16294);
xnor U21027 (N_21027,N_16807,N_15435);
nor U21028 (N_21028,N_12522,N_16414);
nand U21029 (N_21029,N_15098,N_18231);
xnor U21030 (N_21030,N_13931,N_17844);
or U21031 (N_21031,N_18411,N_12643);
and U21032 (N_21032,N_13866,N_18025);
nand U21033 (N_21033,N_16408,N_12871);
nand U21034 (N_21034,N_14643,N_14141);
nor U21035 (N_21035,N_17575,N_14599);
nand U21036 (N_21036,N_18692,N_18129);
nor U21037 (N_21037,N_16360,N_14125);
xnor U21038 (N_21038,N_13848,N_12872);
nand U21039 (N_21039,N_15540,N_17499);
nor U21040 (N_21040,N_13114,N_13215);
xnor U21041 (N_21041,N_12997,N_12949);
or U21042 (N_21042,N_15953,N_17382);
nor U21043 (N_21043,N_15310,N_16534);
or U21044 (N_21044,N_15725,N_17805);
and U21045 (N_21045,N_18343,N_13449);
or U21046 (N_21046,N_15656,N_14355);
xnor U21047 (N_21047,N_16377,N_16197);
nor U21048 (N_21048,N_12567,N_17807);
and U21049 (N_21049,N_13863,N_14582);
xnor U21050 (N_21050,N_17332,N_13556);
or U21051 (N_21051,N_14550,N_15987);
nand U21052 (N_21052,N_14251,N_16051);
and U21053 (N_21053,N_17662,N_12950);
xnor U21054 (N_21054,N_13416,N_13137);
xnor U21055 (N_21055,N_15596,N_15802);
nand U21056 (N_21056,N_18624,N_13625);
or U21057 (N_21057,N_17865,N_17110);
and U21058 (N_21058,N_13406,N_13885);
or U21059 (N_21059,N_16836,N_18727);
and U21060 (N_21060,N_18509,N_14164);
xor U21061 (N_21061,N_17635,N_17836);
nor U21062 (N_21062,N_17148,N_14323);
or U21063 (N_21063,N_13913,N_15989);
and U21064 (N_21064,N_17565,N_12903);
or U21065 (N_21065,N_15348,N_14529);
nand U21066 (N_21066,N_16331,N_14325);
and U21067 (N_21067,N_16851,N_18505);
xor U21068 (N_21068,N_15801,N_14715);
nor U21069 (N_21069,N_13375,N_17165);
or U21070 (N_21070,N_14852,N_16960);
or U21071 (N_21071,N_12736,N_16131);
nor U21072 (N_21072,N_14345,N_15353);
nand U21073 (N_21073,N_17524,N_16759);
or U21074 (N_21074,N_17180,N_16941);
nand U21075 (N_21075,N_15192,N_17637);
and U21076 (N_21076,N_18585,N_16521);
xor U21077 (N_21077,N_16030,N_15309);
and U21078 (N_21078,N_13786,N_13073);
nand U21079 (N_21079,N_17249,N_14473);
nand U21080 (N_21080,N_16814,N_12546);
and U21081 (N_21081,N_16689,N_12687);
nand U21082 (N_21082,N_16760,N_17656);
nand U21083 (N_21083,N_14311,N_16069);
nand U21084 (N_21084,N_14375,N_18177);
xor U21085 (N_21085,N_16973,N_18321);
xnor U21086 (N_21086,N_13340,N_15675);
nor U21087 (N_21087,N_14919,N_13995);
nor U21088 (N_21088,N_13716,N_18049);
xor U21089 (N_21089,N_17872,N_12689);
nand U21090 (N_21090,N_17581,N_17699);
xor U21091 (N_21091,N_16146,N_13693);
and U21092 (N_21092,N_18397,N_18038);
nor U21093 (N_21093,N_12697,N_17727);
nor U21094 (N_21094,N_12571,N_12808);
nand U21095 (N_21095,N_13981,N_17175);
nand U21096 (N_21096,N_18661,N_16744);
nor U21097 (N_21097,N_14374,N_13050);
or U21098 (N_21098,N_13522,N_18700);
or U21099 (N_21099,N_13294,N_15739);
nand U21100 (N_21100,N_14284,N_17552);
xor U21101 (N_21101,N_12957,N_17042);
xnor U21102 (N_21102,N_14706,N_17367);
or U21103 (N_21103,N_18279,N_15436);
and U21104 (N_21104,N_13964,N_16576);
or U21105 (N_21105,N_17116,N_13867);
nor U21106 (N_21106,N_17452,N_14750);
nand U21107 (N_21107,N_18234,N_15287);
nand U21108 (N_21108,N_17141,N_14674);
nand U21109 (N_21109,N_17462,N_16989);
and U21110 (N_21110,N_13260,N_17404);
or U21111 (N_21111,N_13459,N_15174);
xor U21112 (N_21112,N_17232,N_15615);
or U21113 (N_21113,N_12944,N_16595);
nand U21114 (N_21114,N_16145,N_14656);
nor U21115 (N_21115,N_18517,N_16297);
nand U21116 (N_21116,N_12532,N_16301);
and U21117 (N_21117,N_17528,N_15109);
xor U21118 (N_21118,N_14836,N_18237);
and U21119 (N_21119,N_17751,N_17918);
nor U21120 (N_21120,N_16545,N_12517);
and U21121 (N_21121,N_15751,N_13353);
and U21122 (N_21122,N_18285,N_17343);
nor U21123 (N_21123,N_17428,N_18601);
nand U21124 (N_21124,N_18589,N_13749);
nor U21125 (N_21125,N_16132,N_15064);
nor U21126 (N_21126,N_12544,N_15106);
or U21127 (N_21127,N_14720,N_16045);
or U21128 (N_21128,N_17659,N_12722);
or U21129 (N_21129,N_16695,N_17054);
or U21130 (N_21130,N_16041,N_12679);
and U21131 (N_21131,N_15608,N_12592);
nor U21132 (N_21132,N_17684,N_13954);
or U21133 (N_21133,N_13769,N_12506);
xor U21134 (N_21134,N_16343,N_12855);
and U21135 (N_21135,N_18308,N_17677);
or U21136 (N_21136,N_18256,N_13923);
or U21137 (N_21137,N_15000,N_13253);
nand U21138 (N_21138,N_13976,N_17390);
or U21139 (N_21139,N_12664,N_13261);
nor U21140 (N_21140,N_14503,N_14634);
nor U21141 (N_21141,N_17171,N_17035);
or U21142 (N_21142,N_18401,N_18074);
and U21143 (N_21143,N_14454,N_16560);
nor U21144 (N_21144,N_15182,N_12939);
or U21145 (N_21145,N_15536,N_17998);
and U21146 (N_21146,N_14838,N_14371);
xor U21147 (N_21147,N_14894,N_18106);
nor U21148 (N_21148,N_15469,N_17835);
or U21149 (N_21149,N_15619,N_13562);
and U21150 (N_21150,N_14703,N_17889);
and U21151 (N_21151,N_13231,N_12626);
or U21152 (N_21152,N_18379,N_15787);
nor U21153 (N_21153,N_16148,N_18000);
nand U21154 (N_21154,N_14070,N_14357);
nor U21155 (N_21155,N_16273,N_16742);
nor U21156 (N_21156,N_16776,N_13184);
and U21157 (N_21157,N_15468,N_15567);
xnor U21158 (N_21158,N_15772,N_14591);
or U21159 (N_21159,N_18353,N_18233);
or U21160 (N_21160,N_18408,N_18613);
and U21161 (N_21161,N_15144,N_13740);
nor U21162 (N_21162,N_14758,N_12710);
or U21163 (N_21163,N_18522,N_14541);
nand U21164 (N_21164,N_12795,N_16509);
nand U21165 (N_21165,N_14925,N_12611);
nand U21166 (N_21166,N_15629,N_16063);
or U21167 (N_21167,N_14677,N_14228);
xor U21168 (N_21168,N_15298,N_14743);
and U21169 (N_21169,N_17034,N_17526);
nand U21170 (N_21170,N_16144,N_13785);
or U21171 (N_21171,N_15851,N_12648);
and U21172 (N_21172,N_15225,N_17707);
nand U21173 (N_21173,N_16468,N_16079);
and U21174 (N_21174,N_16142,N_13505);
nor U21175 (N_21175,N_15972,N_17695);
and U21176 (N_21176,N_13344,N_15428);
nand U21177 (N_21177,N_16430,N_14407);
xor U21178 (N_21178,N_18452,N_17612);
nand U21179 (N_21179,N_14782,N_16213);
nor U21180 (N_21180,N_12625,N_14692);
and U21181 (N_21181,N_16424,N_18706);
or U21182 (N_21182,N_13521,N_17621);
and U21183 (N_21183,N_16366,N_12980);
and U21184 (N_21184,N_12568,N_13909);
nand U21185 (N_21185,N_13471,N_16227);
nand U21186 (N_21186,N_18196,N_14038);
nand U21187 (N_21187,N_16921,N_15866);
nor U21188 (N_21188,N_13116,N_16165);
nor U21189 (N_21189,N_17314,N_18050);
and U21190 (N_21190,N_18643,N_18484);
or U21191 (N_21191,N_17329,N_16350);
xnor U21192 (N_21192,N_17740,N_14382);
nor U21193 (N_21193,N_17743,N_13476);
and U21194 (N_21194,N_17281,N_13838);
or U21195 (N_21195,N_15764,N_13373);
and U21196 (N_21196,N_13136,N_15491);
and U21197 (N_21197,N_17792,N_17535);
nor U21198 (N_21198,N_13436,N_16198);
xor U21199 (N_21199,N_18657,N_13822);
nand U21200 (N_21200,N_16980,N_13506);
nor U21201 (N_21201,N_12703,N_13560);
or U21202 (N_21202,N_15058,N_18637);
and U21203 (N_21203,N_13603,N_18214);
or U21204 (N_21204,N_14868,N_15891);
xnor U21205 (N_21205,N_17055,N_16374);
xnor U21206 (N_21206,N_14397,N_17313);
nand U21207 (N_21207,N_13016,N_15014);
nand U21208 (N_21208,N_13339,N_14915);
xor U21209 (N_21209,N_18076,N_14242);
nand U21210 (N_21210,N_15004,N_14181);
nor U21211 (N_21211,N_18248,N_18367);
nor U21212 (N_21212,N_14197,N_17610);
xor U21213 (N_21213,N_18709,N_14561);
nor U21214 (N_21214,N_15497,N_16928);
nor U21215 (N_21215,N_15617,N_18219);
nand U21216 (N_21216,N_18394,N_12926);
nand U21217 (N_21217,N_17646,N_17794);
nand U21218 (N_21218,N_15731,N_12901);
nor U21219 (N_21219,N_13983,N_18716);
nor U21220 (N_21220,N_16734,N_15952);
xor U21221 (N_21221,N_15312,N_16738);
xnor U21222 (N_21222,N_15689,N_17463);
nor U21223 (N_21223,N_12810,N_17142);
nand U21224 (N_21224,N_12843,N_12540);
xor U21225 (N_21225,N_18725,N_17303);
or U21226 (N_21226,N_16449,N_13514);
or U21227 (N_21227,N_17252,N_17674);
or U21228 (N_21228,N_15029,N_16835);
or U21229 (N_21229,N_16101,N_17873);
nand U21230 (N_21230,N_15523,N_18552);
or U21231 (N_21231,N_18317,N_16946);
nor U21232 (N_21232,N_15895,N_17560);
and U21233 (N_21233,N_12786,N_13263);
nand U21234 (N_21234,N_14553,N_17607);
xor U21235 (N_21235,N_14367,N_15120);
or U21236 (N_21236,N_13074,N_16161);
xor U21237 (N_21237,N_14687,N_16826);
and U21238 (N_21238,N_16065,N_12683);
and U21239 (N_21239,N_17369,N_13090);
and U21240 (N_21240,N_15825,N_12623);
nand U21241 (N_21241,N_17095,N_16064);
xnor U21242 (N_21242,N_17829,N_12545);
nand U21243 (N_21243,N_16275,N_13570);
nand U21244 (N_21244,N_15822,N_17815);
and U21245 (N_21245,N_16530,N_15217);
or U21246 (N_21246,N_14702,N_13901);
or U21247 (N_21247,N_18201,N_15423);
and U21248 (N_21248,N_17197,N_13048);
and U21249 (N_21249,N_12992,N_18501);
and U21250 (N_21250,N_17806,N_17555);
or U21251 (N_21251,N_13880,N_16965);
and U21252 (N_21252,N_17497,N_17485);
xnor U21253 (N_21253,N_14008,N_17842);
or U21254 (N_21254,N_14833,N_12505);
nor U21255 (N_21255,N_17955,N_15978);
or U21256 (N_21256,N_14882,N_15579);
and U21257 (N_21257,N_16858,N_14822);
and U21258 (N_21258,N_15399,N_16265);
nor U21259 (N_21259,N_17937,N_18621);
or U21260 (N_21260,N_13234,N_14722);
or U21261 (N_21261,N_16617,N_13742);
nor U21262 (N_21262,N_15270,N_14035);
xor U21263 (N_21263,N_14417,N_18469);
nor U21264 (N_21264,N_16244,N_15253);
xnor U21265 (N_21265,N_17434,N_17679);
nand U21266 (N_21266,N_18745,N_15184);
nor U21267 (N_21267,N_16330,N_18728);
and U21268 (N_21268,N_16106,N_14717);
nand U21269 (N_21269,N_17617,N_16582);
nor U21270 (N_21270,N_16909,N_14896);
or U21271 (N_21271,N_18627,N_14186);
xor U21272 (N_21272,N_13460,N_17819);
and U21273 (N_21273,N_14506,N_17553);
nor U21274 (N_21274,N_18466,N_13077);
or U21275 (N_21275,N_17609,N_12542);
nand U21276 (N_21276,N_16047,N_16140);
xor U21277 (N_21277,N_14003,N_14571);
xnor U21278 (N_21278,N_17458,N_15956);
xor U21279 (N_21279,N_18541,N_17231);
xnor U21280 (N_21280,N_12923,N_17980);
xor U21281 (N_21281,N_18557,N_18586);
and U21282 (N_21282,N_16108,N_17221);
nor U21283 (N_21283,N_15696,N_12774);
nor U21284 (N_21284,N_14927,N_14576);
nor U21285 (N_21285,N_15599,N_17614);
and U21286 (N_21286,N_17702,N_16563);
and U21287 (N_21287,N_17645,N_12681);
xnor U21288 (N_21288,N_18687,N_14617);
nor U21289 (N_21289,N_13022,N_13966);
and U21290 (N_21290,N_16365,N_13393);
xnor U21291 (N_21291,N_16686,N_15251);
nand U21292 (N_21292,N_13660,N_13319);
xor U21293 (N_21293,N_17451,N_14040);
xnor U21294 (N_21294,N_12751,N_17227);
nor U21295 (N_21295,N_16291,N_15301);
xor U21296 (N_21296,N_15622,N_16394);
nand U21297 (N_21297,N_16059,N_12829);
nor U21298 (N_21298,N_13569,N_17985);
nand U21299 (N_21299,N_13236,N_15868);
or U21300 (N_21300,N_12562,N_15995);
nor U21301 (N_21301,N_15425,N_17129);
or U21302 (N_21302,N_15538,N_13974);
nand U21303 (N_21303,N_13486,N_15929);
and U21304 (N_21304,N_15194,N_15863);
nor U21305 (N_21305,N_14033,N_15945);
or U21306 (N_21306,N_13161,N_16093);
xnor U21307 (N_21307,N_18433,N_13950);
xnor U21308 (N_21308,N_16763,N_17505);
nand U21309 (N_21309,N_14119,N_14315);
nor U21310 (N_21310,N_16819,N_16088);
or U21311 (N_21311,N_15212,N_17719);
and U21312 (N_21312,N_14681,N_13532);
nand U21313 (N_21313,N_16329,N_16536);
and U21314 (N_21314,N_13726,N_14861);
and U21315 (N_21315,N_15377,N_17777);
nor U21316 (N_21316,N_17520,N_15236);
and U21317 (N_21317,N_17094,N_14620);
and U21318 (N_21318,N_18584,N_18350);
and U21319 (N_21319,N_16961,N_13510);
xnor U21320 (N_21320,N_13703,N_14061);
nand U21321 (N_21321,N_13252,N_17601);
xor U21322 (N_21322,N_17356,N_16238);
and U21323 (N_21323,N_13912,N_14516);
or U21324 (N_21324,N_16315,N_16529);
or U21325 (N_21325,N_16870,N_18243);
or U21326 (N_21326,N_18120,N_14867);
nor U21327 (N_21327,N_17715,N_15485);
nor U21328 (N_21328,N_16613,N_14272);
xnor U21329 (N_21329,N_17861,N_18360);
nand U21330 (N_21330,N_14885,N_18538);
nor U21331 (N_21331,N_13892,N_14135);
nand U21332 (N_21332,N_12601,N_15008);
and U21333 (N_21333,N_13363,N_16537);
and U21334 (N_21334,N_17949,N_12755);
xnor U21335 (N_21335,N_17065,N_14811);
or U21336 (N_21336,N_13283,N_13221);
xor U21337 (N_21337,N_14719,N_13850);
nor U21338 (N_21338,N_12641,N_18526);
nor U21339 (N_21339,N_17570,N_12572);
xor U21340 (N_21340,N_13465,N_18206);
nor U21341 (N_21341,N_15988,N_18447);
and U21342 (N_21342,N_13734,N_16386);
xnor U21343 (N_21343,N_12744,N_16914);
nand U21344 (N_21344,N_14736,N_12879);
or U21345 (N_21345,N_16677,N_13492);
or U21346 (N_21346,N_15276,N_13770);
xor U21347 (N_21347,N_17653,N_17453);
nand U21348 (N_21348,N_17063,N_17226);
and U21349 (N_21349,N_14372,N_16952);
nor U21350 (N_21350,N_16417,N_14565);
nor U21351 (N_21351,N_15484,N_16085);
or U21352 (N_21352,N_13930,N_13034);
nand U21353 (N_21353,N_16352,N_15733);
and U21354 (N_21354,N_15524,N_12907);
nor U21355 (N_21355,N_18080,N_16609);
and U21356 (N_21356,N_13326,N_17245);
nor U21357 (N_21357,N_15456,N_16860);
or U21358 (N_21358,N_15971,N_18392);
nor U21359 (N_21359,N_12536,N_17024);
or U21360 (N_21360,N_14545,N_17209);
nor U21361 (N_21361,N_12644,N_13385);
xnor U21362 (N_21362,N_18047,N_14434);
or U21363 (N_21363,N_16039,N_14134);
or U21364 (N_21364,N_17786,N_14238);
and U21365 (N_21365,N_14633,N_14039);
nor U21366 (N_21366,N_13291,N_16413);
and U21367 (N_21367,N_17018,N_15514);
or U21368 (N_21368,N_16911,N_15798);
nor U21369 (N_21369,N_16199,N_17061);
xnor U21370 (N_21370,N_15593,N_16644);
or U21371 (N_21371,N_14157,N_14673);
nor U21372 (N_21372,N_13101,N_13732);
and U21373 (N_21373,N_17324,N_15641);
nand U21374 (N_21374,N_16296,N_15750);
nand U21375 (N_21375,N_13350,N_12834);
nor U21376 (N_21376,N_16834,N_14784);
xnor U21377 (N_21377,N_14354,N_14924);
nand U21378 (N_21378,N_18091,N_14460);
or U21379 (N_21379,N_13766,N_15726);
xnor U21380 (N_21380,N_15730,N_12866);
xor U21381 (N_21381,N_13761,N_12858);
or U21382 (N_21382,N_17577,N_13356);
xor U21383 (N_21383,N_13499,N_12970);
nand U21384 (N_21384,N_14587,N_15452);
nand U21385 (N_21385,N_17824,N_15424);
xnor U21386 (N_21386,N_18303,N_17648);
nor U21387 (N_21387,N_14153,N_18540);
and U21388 (N_21388,N_17522,N_13145);
xnor U21389 (N_21389,N_15146,N_15305);
or U21390 (N_21390,N_17099,N_18099);
nor U21391 (N_21391,N_12845,N_18514);
or U21392 (N_21392,N_13053,N_16043);
and U21393 (N_21393,N_13056,N_14370);
nor U21394 (N_21394,N_14162,N_16651);
nor U21395 (N_21395,N_12967,N_14359);
nand U21396 (N_21396,N_15954,N_15889);
or U21397 (N_21397,N_15155,N_12817);
and U21398 (N_21398,N_14140,N_15151);
or U21399 (N_21399,N_17912,N_14756);
and U21400 (N_21400,N_15134,N_13533);
nor U21401 (N_21401,N_14258,N_14841);
nand U21402 (N_21402,N_14226,N_15994);
and U21403 (N_21403,N_16450,N_16934);
or U21404 (N_21404,N_14490,N_16240);
nor U21405 (N_21405,N_18593,N_18130);
xnor U21406 (N_21406,N_17287,N_12762);
xor U21407 (N_21407,N_17561,N_13899);
or U21408 (N_21408,N_16158,N_12766);
or U21409 (N_21409,N_17650,N_15354);
nor U21410 (N_21410,N_15115,N_16017);
nand U21411 (N_21411,N_17643,N_16305);
nor U21412 (N_21412,N_13949,N_15202);
nor U21413 (N_21413,N_17938,N_13076);
or U21414 (N_21414,N_16253,N_13179);
or U21415 (N_21415,N_14953,N_18711);
nand U21416 (N_21416,N_17079,N_18143);
nand U21417 (N_21417,N_14348,N_17276);
and U21418 (N_21418,N_17145,N_17502);
xnor U21419 (N_21419,N_14776,N_13354);
nand U21420 (N_21420,N_17440,N_15426);
nand U21421 (N_21421,N_15471,N_18547);
nor U21422 (N_21422,N_16507,N_17225);
nor U21423 (N_21423,N_17669,N_13986);
or U21424 (N_21424,N_13903,N_15709);
nor U21425 (N_21425,N_14992,N_17421);
xor U21426 (N_21426,N_18681,N_16683);
and U21427 (N_21427,N_15519,N_17257);
or U21428 (N_21428,N_17975,N_14984);
or U21429 (N_21429,N_17906,N_16202);
nor U21430 (N_21430,N_14555,N_17268);
nand U21431 (N_21431,N_14846,N_14138);
nand U21432 (N_21432,N_12981,N_17547);
nand U21433 (N_21433,N_14577,N_15370);
or U21434 (N_21434,N_17416,N_16186);
and U21435 (N_21435,N_15022,N_13140);
and U21436 (N_21436,N_15013,N_14667);
and U21437 (N_21437,N_16778,N_17847);
or U21438 (N_21438,N_14025,N_16149);
and U21439 (N_21439,N_14801,N_16678);
or U21440 (N_21440,N_18207,N_16806);
xnor U21441 (N_21441,N_18168,N_14662);
or U21442 (N_21442,N_14278,N_17837);
xnor U21443 (N_21443,N_13933,N_13098);
nor U21444 (N_21444,N_17939,N_17752);
xor U21445 (N_21445,N_18649,N_13463);
nor U21446 (N_21446,N_16385,N_18710);
nor U21447 (N_21447,N_13194,N_14227);
nor U21448 (N_21448,N_15820,N_13347);
nor U21449 (N_21449,N_16373,N_13159);
xnor U21450 (N_21450,N_18713,N_16953);
nand U21451 (N_21451,N_15477,N_15291);
nor U21452 (N_21452,N_17686,N_17849);
nand U21453 (N_21453,N_15560,N_18009);
nand U21454 (N_21454,N_18625,N_16894);
nand U21455 (N_21455,N_16247,N_15762);
xor U21456 (N_21456,N_16803,N_16249);
xor U21457 (N_21457,N_18389,N_16918);
or U21458 (N_21458,N_15965,N_14139);
xnor U21459 (N_21459,N_12792,N_14111);
xor U21460 (N_21460,N_16779,N_16995);
nand U21461 (N_21461,N_18203,N_16089);
and U21462 (N_21462,N_17082,N_15288);
nand U21463 (N_21463,N_16931,N_13051);
nor U21464 (N_21464,N_13696,N_13175);
nand U21465 (N_21465,N_15177,N_15034);
xor U21466 (N_21466,N_17446,N_14799);
nand U21467 (N_21467,N_14903,N_16584);
xor U21468 (N_21468,N_14902,N_16169);
xor U21469 (N_21469,N_15735,N_18607);
nand U21470 (N_21470,N_14734,N_18375);
and U21471 (N_21471,N_14798,N_15249);
and U21472 (N_21472,N_15865,N_15711);
and U21473 (N_21473,N_16784,N_13529);
xnor U21474 (N_21474,N_16638,N_13164);
nand U21475 (N_21475,N_15961,N_16743);
or U21476 (N_21476,N_18386,N_14166);
or U21477 (N_21477,N_13388,N_13144);
or U21478 (N_21478,N_16489,N_13457);
or U21479 (N_21479,N_15816,N_12910);
nor U21480 (N_21480,N_17154,N_13002);
xnor U21481 (N_21481,N_15191,N_15296);
nor U21482 (N_21482,N_15070,N_16127);
nand U21483 (N_21483,N_14624,N_15892);
nand U21484 (N_21484,N_17770,N_15738);
or U21485 (N_21485,N_15044,N_14086);
and U21486 (N_21486,N_12668,N_15183);
or U21487 (N_21487,N_18439,N_18344);
nand U21488 (N_21488,N_14026,N_14123);
or U21489 (N_21489,N_12844,N_18027);
or U21490 (N_21490,N_15695,N_15090);
or U21491 (N_21491,N_17689,N_15293);
nand U21492 (N_21492,N_17558,N_12842);
nor U21493 (N_21493,N_14837,N_12500);
and U21494 (N_21494,N_15662,N_13955);
xnor U21495 (N_21495,N_17673,N_15740);
xor U21496 (N_21496,N_17749,N_15303);
nor U21497 (N_21497,N_16215,N_18746);
and U21498 (N_21498,N_12840,N_18221);
or U21499 (N_21499,N_12826,N_13604);
nand U21500 (N_21500,N_14875,N_15880);
nor U21501 (N_21501,N_17046,N_17487);
nor U21502 (N_21502,N_13003,N_14808);
nand U21503 (N_21503,N_12877,N_13991);
or U21504 (N_21504,N_15794,N_17089);
nor U21505 (N_21505,N_13780,N_13297);
and U21506 (N_21506,N_13774,N_18218);
nor U21507 (N_21507,N_16464,N_13627);
xnor U21508 (N_21508,N_15255,N_17352);
nor U21509 (N_21509,N_15404,N_16874);
nand U21510 (N_21510,N_15429,N_14977);
or U21511 (N_21511,N_17972,N_15240);
xor U21512 (N_21512,N_16680,N_14558);
or U21513 (N_21513,N_18459,N_12640);
nor U21514 (N_21514,N_13325,N_12999);
nor U21515 (N_21515,N_14100,N_14966);
nor U21516 (N_21516,N_18033,N_16690);
or U21517 (N_21517,N_15955,N_13207);
nand U21518 (N_21518,N_13805,N_16605);
nand U21519 (N_21519,N_13425,N_15009);
nand U21520 (N_21520,N_13108,N_14886);
and U21521 (N_21521,N_17750,N_14533);
nand U21522 (N_21522,N_14631,N_16516);
nand U21523 (N_21523,N_17808,N_15842);
nand U21524 (N_21524,N_15108,N_15533);
and U21525 (N_21525,N_12740,N_15366);
nor U21526 (N_21526,N_17002,N_15083);
and U21527 (N_21527,N_16369,N_16452);
and U21528 (N_21528,N_17250,N_18134);
xnor U21529 (N_21529,N_13302,N_12588);
nand U21530 (N_21530,N_13275,N_16766);
and U21531 (N_21531,N_12610,N_14032);
nor U21532 (N_21532,N_13403,N_13052);
nand U21533 (N_21533,N_15211,N_17537);
and U21534 (N_21534,N_18693,N_13132);
xnor U21535 (N_21535,N_13167,N_15444);
nor U21536 (N_21536,N_18341,N_13519);
nor U21537 (N_21537,N_14803,N_16798);
or U21538 (N_21538,N_14387,N_16400);
nand U21539 (N_21539,N_17852,N_12612);
or U21540 (N_21540,N_13395,N_18239);
nand U21541 (N_21541,N_14069,N_13206);
and U21542 (N_21542,N_15748,N_12699);
or U21543 (N_21543,N_18277,N_12561);
nor U21544 (N_21544,N_18212,N_14442);
or U21545 (N_21545,N_15110,N_15981);
xnor U21546 (N_21546,N_13713,N_12919);
xor U21547 (N_21547,N_14045,N_17722);
and U21548 (N_21548,N_15228,N_14573);
or U21549 (N_21549,N_13119,N_18023);
nand U21550 (N_21550,N_16423,N_13345);
xor U21551 (N_21551,N_12675,N_17585);
and U21552 (N_21552,N_15744,N_14542);
and U21553 (N_21553,N_16179,N_17068);
nor U21554 (N_21554,N_18310,N_17265);
or U21555 (N_21555,N_13313,N_14592);
nor U21556 (N_21556,N_13193,N_15333);
nand U21557 (N_21557,N_12776,N_14699);
xor U21558 (N_21558,N_12533,N_15898);
and U21559 (N_21559,N_17787,N_15432);
and U21560 (N_21560,N_13482,N_16715);
nand U21561 (N_21561,N_14760,N_12594);
xor U21562 (N_21562,N_14585,N_13485);
xnor U21563 (N_21563,N_17551,N_14306);
xor U21564 (N_21564,N_12906,N_13543);
or U21565 (N_21565,N_14386,N_18482);
or U21566 (N_21566,N_18676,N_13472);
nor U21567 (N_21567,N_14949,N_16044);
nor U21568 (N_21568,N_18714,N_17379);
and U21569 (N_21569,N_15570,N_12717);
nor U21570 (N_21570,N_17496,N_17878);
and U21571 (N_21571,N_12609,N_17623);
or U21572 (N_21572,N_13620,N_18370);
or U21573 (N_21573,N_17588,N_14764);
nor U21574 (N_21574,N_18358,N_13705);
or U21575 (N_21575,N_13151,N_16675);
nor U21576 (N_21576,N_12805,N_18105);
or U21577 (N_21577,N_14932,N_13990);
xnor U21578 (N_21578,N_13712,N_15638);
or U21579 (N_21579,N_16768,N_16886);
xor U21580 (N_21580,N_17215,N_13496);
nand U21581 (N_21581,N_16575,N_16188);
nand U21582 (N_21582,N_13483,N_16685);
nor U21583 (N_21583,N_13957,N_14463);
xor U21584 (N_21584,N_18010,N_14884);
and U21585 (N_21585,N_15084,N_17989);
or U21586 (N_21586,N_14580,N_14419);
nand U21587 (N_21587,N_17374,N_15085);
nor U21588 (N_21588,N_15707,N_17774);
xnor U21589 (N_21589,N_14149,N_16465);
nand U21590 (N_21590,N_15754,N_15658);
or U21591 (N_21591,N_15974,N_12825);
nor U21592 (N_21592,N_15979,N_18600);
nand U21593 (N_21593,N_12839,N_15595);
and U21594 (N_21594,N_17403,N_17429);
or U21595 (N_21595,N_16823,N_12737);
nand U21596 (N_21596,N_14037,N_16049);
and U21597 (N_21597,N_14727,N_12539);
xnor U21598 (N_21598,N_16091,N_18005);
nor U21599 (N_21599,N_15087,N_17201);
and U21600 (N_21600,N_14253,N_13948);
and U21601 (N_21601,N_14351,N_17005);
or U21602 (N_21602,N_17627,N_13096);
nor U21603 (N_21603,N_16421,N_15901);
nor U21604 (N_21604,N_15555,N_18067);
and U21605 (N_21605,N_14664,N_18252);
or U21606 (N_21606,N_15091,N_12941);
nand U21607 (N_21607,N_15512,N_13882);
nor U21608 (N_21608,N_16504,N_12802);
or U21609 (N_21609,N_17882,N_18163);
and U21610 (N_21610,N_14778,N_15299);
xnor U21611 (N_21611,N_16589,N_12739);
nor U21612 (N_21612,N_14344,N_16174);
nor U21613 (N_21613,N_15315,N_18113);
xor U21614 (N_21614,N_13720,N_15983);
nor U21615 (N_21615,N_15421,N_16643);
and U21616 (N_21616,N_12657,N_14842);
or U21617 (N_21617,N_14233,N_16216);
and U21618 (N_21618,N_18217,N_15912);
nor U21619 (N_21619,N_17170,N_13331);
nor U21620 (N_21620,N_12890,N_14301);
nand U21621 (N_21621,N_14520,N_13989);
and U21622 (N_21622,N_15220,N_14225);
or U21623 (N_21623,N_18646,N_13208);
or U21624 (N_21624,N_16721,N_13965);
and U21625 (N_21625,N_15831,N_15659);
nor U21626 (N_21626,N_14869,N_18421);
and U21627 (N_21627,N_17478,N_13526);
nor U21628 (N_21628,N_14914,N_13379);
or U21629 (N_21629,N_13845,N_17838);
or U21630 (N_21630,N_13226,N_14314);
and U21631 (N_21631,N_15131,N_14586);
xnor U21632 (N_21632,N_16749,N_13943);
or U21633 (N_21633,N_13084,N_18572);
nor U21634 (N_21634,N_17275,N_14830);
nor U21635 (N_21635,N_17191,N_13214);
xnor U21636 (N_21636,N_16895,N_12646);
xor U21637 (N_21637,N_12854,N_18229);
or U21638 (N_21638,N_14209,N_14461);
nand U21639 (N_21639,N_14853,N_12800);
or U21640 (N_21640,N_14995,N_16646);
nand U21641 (N_21641,N_18003,N_12860);
nor U21642 (N_21642,N_17885,N_15114);
xnor U21643 (N_21643,N_15771,N_15535);
nand U21644 (N_21644,N_16764,N_14259);
nor U21645 (N_21645,N_17162,N_15152);
or U21646 (N_21646,N_16551,N_13023);
nor U21647 (N_21647,N_12735,N_13014);
nand U21648 (N_21648,N_14213,N_13501);
nor U21649 (N_21649,N_12775,N_14341);
xor U21650 (N_21650,N_17410,N_16483);
xnor U21651 (N_21651,N_13072,N_14000);
xnor U21652 (N_21652,N_14929,N_15872);
or U21653 (N_21653,N_13650,N_17934);
xnor U21654 (N_21654,N_16475,N_14531);
and U21655 (N_21655,N_17508,N_17922);
and U21656 (N_21656,N_17338,N_14987);
nor U21657 (N_21657,N_14802,N_17655);
nor U21658 (N_21658,N_15645,N_15962);
nand U21659 (N_21659,N_18040,N_13426);
nor U21660 (N_21660,N_13638,N_17173);
or U21661 (N_21661,N_17863,N_14185);
and U21662 (N_21662,N_17026,N_18205);
and U21663 (N_21663,N_18289,N_13910);
nor U21664 (N_21664,N_15233,N_14858);
or U21665 (N_21665,N_16313,N_17203);
nor U21666 (N_21666,N_14483,N_13278);
nand U21667 (N_21667,N_18071,N_18043);
nand U21668 (N_21668,N_17706,N_17797);
and U21669 (N_21669,N_18525,N_18276);
and U21670 (N_21670,N_18008,N_17483);
or U21671 (N_21671,N_18368,N_14532);
nand U21672 (N_21672,N_12987,N_16383);
and U21673 (N_21673,N_16284,N_16859);
xnor U21674 (N_21674,N_16761,N_17307);
xnor U21675 (N_21675,N_14653,N_17851);
xor U21676 (N_21676,N_12881,N_18477);
nor U21677 (N_21677,N_16321,N_17633);
nor U21678 (N_21678,N_17984,N_14855);
nor U21679 (N_21679,N_17960,N_17891);
xnor U21680 (N_21680,N_13826,N_15001);
and U21681 (N_21681,N_16850,N_13421);
nand U21682 (N_21682,N_13069,N_14877);
nor U21683 (N_21683,N_15861,N_12831);
xor U21684 (N_21684,N_16022,N_15894);
nand U21685 (N_21685,N_17195,N_18116);
nor U21686 (N_21686,N_12971,N_17821);
xnor U21687 (N_21687,N_15781,N_17218);
xor U21688 (N_21688,N_13787,N_16863);
and U21689 (N_21689,N_15679,N_16262);
xor U21690 (N_21690,N_18354,N_18290);
xnor U21691 (N_21691,N_12515,N_15786);
nand U21692 (N_21692,N_15676,N_12658);
or U21693 (N_21693,N_14625,N_17682);
nor U21694 (N_21694,N_14257,N_16066);
and U21695 (N_21695,N_12677,N_13967);
nor U21696 (N_21696,N_17011,N_13858);
nand U21697 (N_21697,N_15142,N_17519);
nor U21698 (N_21698,N_14761,N_14800);
and U21699 (N_21699,N_14979,N_15902);
and U21700 (N_21700,N_16282,N_15295);
nand U21701 (N_21701,N_13652,N_14223);
nor U21702 (N_21702,N_13123,N_15791);
nand U21703 (N_21703,N_15813,N_18115);
and U21704 (N_21704,N_18195,N_18046);
or U21705 (N_21705,N_17105,N_17692);
xor U21706 (N_21706,N_17292,N_17571);
and U21707 (N_21707,N_17688,N_16219);
and U21708 (N_21708,N_13064,N_16194);
xor U21709 (N_21709,N_16947,N_13049);
and U21710 (N_21710,N_16913,N_16271);
nand U21711 (N_21711,N_16435,N_16508);
nor U21712 (N_21712,N_15222,N_14812);
xnor U21713 (N_21713,N_18702,N_14128);
nand U21714 (N_21714,N_14663,N_13776);
nand U21715 (N_21715,N_15930,N_16824);
xor U21716 (N_21716,N_13549,N_14479);
and U21717 (N_21717,N_16517,N_14465);
xnor U21718 (N_21718,N_17860,N_13723);
xor U21719 (N_21719,N_17341,N_12962);
xnor U21720 (N_21720,N_17078,N_18407);
nand U21721 (N_21721,N_16614,N_14493);
and U21722 (N_21722,N_14390,N_14876);
nor U21723 (N_21723,N_17890,N_13695);
or U21724 (N_21724,N_18744,N_13658);
xor U21725 (N_21725,N_17647,N_15660);
and U21726 (N_21726,N_13984,N_12749);
and U21727 (N_21727,N_13707,N_16033);
or U21728 (N_21728,N_14955,N_13020);
xor U21729 (N_21729,N_16482,N_17856);
or U21730 (N_21730,N_18573,N_12782);
and U21731 (N_21731,N_13464,N_18561);
nand U21732 (N_21732,N_15275,N_14892);
xor U21733 (N_21733,N_15086,N_12589);
xor U21734 (N_21734,N_12635,N_14616);
nor U21735 (N_21735,N_16292,N_13332);
nand U21736 (N_21736,N_14737,N_16056);
nand U21737 (N_21737,N_15526,N_17619);
and U21738 (N_21738,N_16618,N_18599);
and U21739 (N_21739,N_17506,N_12733);
nand U21740 (N_21740,N_15585,N_16993);
nor U21741 (N_21741,N_12833,N_18616);
xnor U21742 (N_21742,N_12777,N_15003);
nand U21743 (N_21743,N_17383,N_13908);
xnor U21744 (N_21744,N_18485,N_13112);
nand U21745 (N_21745,N_13269,N_17405);
nor U21746 (N_21746,N_17981,N_18568);
nor U21747 (N_21747,N_12706,N_15928);
nand U21748 (N_21748,N_14095,N_13622);
nand U21749 (N_21749,N_17357,N_16442);
or U21750 (N_21750,N_13817,N_17776);
and U21751 (N_21751,N_17316,N_17081);
or U21752 (N_21752,N_16460,N_17879);
nand U21753 (N_21753,N_14935,N_13710);
or U21754 (N_21754,N_18199,N_15175);
and U21755 (N_21755,N_17392,N_13586);
xnor U21756 (N_21756,N_15899,N_12900);
or U21757 (N_21757,N_16370,N_12956);
nor U21758 (N_21758,N_13371,N_15442);
xor U21759 (N_21759,N_16714,N_17016);
and U21760 (N_21760,N_13400,N_18608);
nor U21761 (N_21761,N_18611,N_16446);
or U21762 (N_21762,N_17671,N_14851);
and U21763 (N_21763,N_12976,N_14329);
nand U21764 (N_21764,N_16111,N_17291);
and U21765 (N_21765,N_14774,N_17210);
xor U21766 (N_21766,N_13906,N_16231);
or U21767 (N_21767,N_13599,N_13405);
nor U21768 (N_21768,N_17169,N_13103);
xor U21769 (N_21769,N_15283,N_18566);
and U21770 (N_21770,N_13894,N_13329);
nor U21771 (N_21771,N_16490,N_16599);
and U21772 (N_21772,N_17260,N_17120);
or U21773 (N_21773,N_17115,N_12783);
or U21774 (N_21774,N_17119,N_14403);
and U21775 (N_21775,N_15286,N_16728);
xnor U21776 (N_21776,N_18739,N_14588);
xor U21777 (N_21777,N_16307,N_17982);
nand U21778 (N_21778,N_15572,N_16404);
xnor U21779 (N_21779,N_14312,N_17915);
nor U21780 (N_21780,N_14299,N_16884);
xnor U21781 (N_21781,N_14570,N_15576);
nand U21782 (N_21782,N_13960,N_12595);
nor U21783 (N_21783,N_16727,N_17347);
xor U21784 (N_21784,N_13512,N_18513);
and U21785 (N_21785,N_12789,N_15682);
and U21786 (N_21786,N_14907,N_15420);
nor U21787 (N_21787,N_17342,N_17812);
nand U21788 (N_21788,N_13659,N_14071);
and U21789 (N_21789,N_13644,N_13368);
or U21790 (N_21790,N_18157,N_17179);
or U21791 (N_21791,N_18490,N_15937);
or U21792 (N_21792,N_15796,N_14485);
nor U21793 (N_21793,N_14034,N_13878);
nand U21794 (N_21794,N_12704,N_14913);
nor U21795 (N_21795,N_13430,N_16498);
or U21796 (N_21796,N_17419,N_16513);
or U21797 (N_21797,N_15503,N_14920);
and U21798 (N_21798,N_14113,N_16885);
or U21799 (N_21799,N_18686,N_14174);
and U21800 (N_21800,N_18506,N_18124);
or U21801 (N_21801,N_14710,N_15332);
nand U21802 (N_21802,N_12922,N_18082);
xnor U21803 (N_21803,N_17444,N_16555);
nor U21804 (N_21804,N_18565,N_13220);
and U21805 (N_21805,N_13438,N_17501);
nand U21806 (N_21806,N_15686,N_17174);
nand U21807 (N_21807,N_13235,N_17097);
nor U21808 (N_21808,N_15714,N_18682);
or U21809 (N_21809,N_16087,N_12695);
nand U21810 (N_21810,N_12734,N_14963);
xnor U21811 (N_21811,N_17804,N_17282);
or U21812 (N_21812,N_14353,N_17144);
nor U21813 (N_21813,N_16829,N_16397);
nor U21814 (N_21814,N_18615,N_14409);
and U21815 (N_21815,N_15154,N_14408);
xnor U21816 (N_21816,N_12899,N_18574);
xnor U21817 (N_21817,N_16587,N_13895);
xor U21818 (N_21818,N_16502,N_16339);
xnor U21819 (N_21819,N_14513,N_18610);
xor U21820 (N_21820,N_15556,N_15896);
nand U21821 (N_21821,N_18642,N_18110);
nand U21822 (N_21822,N_18664,N_15959);
xnor U21823 (N_21823,N_18602,N_17490);
or U21824 (N_21824,N_12951,N_15362);
nand U21825 (N_21825,N_12573,N_16221);
and U21826 (N_21826,N_17717,N_16441);
nor U21827 (N_21827,N_16982,N_14728);
xor U21828 (N_21828,N_14845,N_15241);
xor U21829 (N_21829,N_15268,N_13567);
or U21830 (N_21830,N_14747,N_17217);
nand U21831 (N_21831,N_18416,N_15935);
xnor U21832 (N_21832,N_17628,N_17964);
or U21833 (N_21833,N_16119,N_12715);
nor U21834 (N_21834,N_14614,N_15448);
nand U21835 (N_21835,N_14642,N_13174);
nor U21836 (N_21836,N_18679,N_13678);
or U21837 (N_21837,N_17959,N_18560);
nand U21838 (N_21838,N_17789,N_17793);
nor U21839 (N_21839,N_18278,N_15511);
nand U21840 (N_21840,N_18211,N_13417);
or U21841 (N_21841,N_18588,N_13544);
nand U21842 (N_21842,N_14523,N_18531);
and U21843 (N_21843,N_17904,N_17069);
nand U21844 (N_21844,N_16261,N_16415);
or U21845 (N_21845,N_17731,N_12835);
and U21846 (N_21846,N_14207,N_16057);
xor U21847 (N_21847,N_13192,N_17284);
nor U21848 (N_21848,N_14292,N_17945);
nor U21849 (N_21849,N_12566,N_17014);
nor U21850 (N_21850,N_15611,N_16923);
nand U21851 (N_21851,N_18448,N_13433);
and U21852 (N_21852,N_12918,N_18665);
or U21853 (N_21853,N_17456,N_13498);
and U21854 (N_21854,N_13714,N_17710);
or U21855 (N_21855,N_17336,N_17745);
nand U21856 (N_21856,N_17137,N_15265);
and U21857 (N_21857,N_17767,N_15140);
nand U21858 (N_21858,N_13816,N_14789);
xor U21859 (N_21859,N_14457,N_15149);
and U21860 (N_21860,N_17800,N_13717);
xor U21861 (N_21861,N_18376,N_13998);
and U21862 (N_21862,N_13462,N_18549);
nand U21863 (N_21863,N_17364,N_15706);
and U21864 (N_21864,N_14031,N_14901);
xor U21865 (N_21865,N_13563,N_13736);
and U21866 (N_21866,N_14274,N_16463);
xnor U21867 (N_21867,N_17881,N_12627);
and U21868 (N_21868,N_14349,N_14499);
or U21869 (N_21869,N_12978,N_12642);
nand U21870 (N_21870,N_13337,N_13803);
or U21871 (N_21871,N_16052,N_16700);
nand U21872 (N_21872,N_13633,N_14712);
nor U21873 (N_21873,N_17106,N_13674);
nor U21874 (N_21874,N_18053,N_16237);
or U21875 (N_21875,N_14990,N_17191);
or U21876 (N_21876,N_17138,N_16627);
nor U21877 (N_21877,N_16264,N_12849);
xor U21878 (N_21878,N_16786,N_14168);
xnor U21879 (N_21879,N_15744,N_17865);
or U21880 (N_21880,N_15657,N_15836);
xor U21881 (N_21881,N_16164,N_17174);
and U21882 (N_21882,N_16993,N_14605);
and U21883 (N_21883,N_17874,N_15447);
nor U21884 (N_21884,N_12831,N_15228);
and U21885 (N_21885,N_18651,N_14067);
or U21886 (N_21886,N_14092,N_13948);
and U21887 (N_21887,N_12902,N_15087);
xor U21888 (N_21888,N_17173,N_16824);
or U21889 (N_21889,N_17104,N_17075);
nand U21890 (N_21890,N_13773,N_12679);
and U21891 (N_21891,N_15940,N_17498);
nor U21892 (N_21892,N_13150,N_17758);
xnor U21893 (N_21893,N_14216,N_15355);
nor U21894 (N_21894,N_15348,N_12921);
nand U21895 (N_21895,N_15027,N_13926);
nor U21896 (N_21896,N_12903,N_16845);
nand U21897 (N_21897,N_16786,N_16788);
nand U21898 (N_21898,N_13197,N_18666);
and U21899 (N_21899,N_14922,N_17926);
xor U21900 (N_21900,N_14360,N_13432);
xor U21901 (N_21901,N_16375,N_15642);
nor U21902 (N_21902,N_14237,N_13276);
nand U21903 (N_21903,N_17708,N_13231);
xor U21904 (N_21904,N_14061,N_16944);
or U21905 (N_21905,N_12564,N_16673);
nor U21906 (N_21906,N_16763,N_14311);
xnor U21907 (N_21907,N_16047,N_17014);
nand U21908 (N_21908,N_15265,N_17281);
xor U21909 (N_21909,N_13062,N_16067);
or U21910 (N_21910,N_18009,N_15658);
nand U21911 (N_21911,N_17245,N_15152);
and U21912 (N_21912,N_17495,N_15006);
nor U21913 (N_21913,N_14121,N_15078);
nand U21914 (N_21914,N_18637,N_15781);
nand U21915 (N_21915,N_15723,N_17563);
xnor U21916 (N_21916,N_12565,N_14828);
and U21917 (N_21917,N_12902,N_13463);
and U21918 (N_21918,N_17245,N_13891);
xor U21919 (N_21919,N_17809,N_15459);
nor U21920 (N_21920,N_14251,N_13266);
xor U21921 (N_21921,N_17169,N_16768);
and U21922 (N_21922,N_14877,N_12741);
or U21923 (N_21923,N_16494,N_14670);
and U21924 (N_21924,N_12766,N_14232);
and U21925 (N_21925,N_16519,N_15333);
nor U21926 (N_21926,N_18139,N_18579);
nor U21927 (N_21927,N_16808,N_17655);
or U21928 (N_21928,N_12560,N_16314);
nand U21929 (N_21929,N_16077,N_16519);
nand U21930 (N_21930,N_13104,N_17253);
nor U21931 (N_21931,N_15799,N_14485);
xor U21932 (N_21932,N_12918,N_14522);
xor U21933 (N_21933,N_17114,N_17529);
and U21934 (N_21934,N_13843,N_15126);
and U21935 (N_21935,N_18334,N_16960);
nor U21936 (N_21936,N_15131,N_15816);
and U21937 (N_21937,N_13841,N_14450);
nand U21938 (N_21938,N_15439,N_16814);
and U21939 (N_21939,N_17886,N_18032);
and U21940 (N_21940,N_16546,N_18366);
xor U21941 (N_21941,N_18111,N_18498);
xor U21942 (N_21942,N_13929,N_12587);
nor U21943 (N_21943,N_18363,N_17003);
nor U21944 (N_21944,N_16512,N_14594);
nand U21945 (N_21945,N_17383,N_14811);
xor U21946 (N_21946,N_17740,N_15857);
and U21947 (N_21947,N_16317,N_17067);
xnor U21948 (N_21948,N_17762,N_14465);
or U21949 (N_21949,N_18266,N_17348);
nor U21950 (N_21950,N_17862,N_16582);
or U21951 (N_21951,N_18731,N_17838);
xnor U21952 (N_21952,N_16242,N_14914);
or U21953 (N_21953,N_15195,N_17330);
and U21954 (N_21954,N_14934,N_12812);
and U21955 (N_21955,N_16810,N_17123);
nor U21956 (N_21956,N_17181,N_14569);
nand U21957 (N_21957,N_18608,N_14871);
xnor U21958 (N_21958,N_17170,N_16398);
or U21959 (N_21959,N_14298,N_18693);
nor U21960 (N_21960,N_16711,N_17126);
or U21961 (N_21961,N_12765,N_17536);
and U21962 (N_21962,N_16368,N_18119);
and U21963 (N_21963,N_12848,N_15340);
nor U21964 (N_21964,N_12968,N_17214);
and U21965 (N_21965,N_15120,N_15493);
nand U21966 (N_21966,N_14736,N_15177);
nor U21967 (N_21967,N_18293,N_15028);
or U21968 (N_21968,N_17503,N_17632);
nand U21969 (N_21969,N_18737,N_15125);
nor U21970 (N_21970,N_14779,N_14353);
or U21971 (N_21971,N_15934,N_13907);
xnor U21972 (N_21972,N_15221,N_14482);
or U21973 (N_21973,N_13803,N_14755);
nand U21974 (N_21974,N_17969,N_14366);
or U21975 (N_21975,N_17693,N_17719);
and U21976 (N_21976,N_15898,N_17127);
or U21977 (N_21977,N_18006,N_15641);
and U21978 (N_21978,N_12851,N_16087);
nor U21979 (N_21979,N_16782,N_17345);
or U21980 (N_21980,N_13491,N_15505);
or U21981 (N_21981,N_18377,N_13038);
and U21982 (N_21982,N_14362,N_14911);
or U21983 (N_21983,N_13485,N_17603);
and U21984 (N_21984,N_13510,N_16872);
nand U21985 (N_21985,N_17351,N_13672);
nor U21986 (N_21986,N_18349,N_14191);
nor U21987 (N_21987,N_14941,N_13887);
or U21988 (N_21988,N_17864,N_18360);
and U21989 (N_21989,N_14511,N_15021);
nor U21990 (N_21990,N_16950,N_18238);
nor U21991 (N_21991,N_18058,N_13777);
or U21992 (N_21992,N_18256,N_17435);
nand U21993 (N_21993,N_12832,N_15485);
nor U21994 (N_21994,N_13290,N_17370);
or U21995 (N_21995,N_13518,N_13120);
nand U21996 (N_21996,N_17785,N_16457);
nor U21997 (N_21997,N_15448,N_17323);
nand U21998 (N_21998,N_13492,N_13660);
nor U21999 (N_21999,N_16917,N_17533);
nand U22000 (N_22000,N_18111,N_17179);
or U22001 (N_22001,N_18557,N_16559);
or U22002 (N_22002,N_12842,N_13287);
nand U22003 (N_22003,N_12617,N_13139);
or U22004 (N_22004,N_13006,N_16303);
xnor U22005 (N_22005,N_14853,N_18245);
nand U22006 (N_22006,N_14954,N_15773);
nor U22007 (N_22007,N_13897,N_17275);
or U22008 (N_22008,N_15814,N_13138);
xor U22009 (N_22009,N_17180,N_18143);
nor U22010 (N_22010,N_13118,N_12846);
and U22011 (N_22011,N_15605,N_17629);
nor U22012 (N_22012,N_14363,N_16252);
nand U22013 (N_22013,N_14867,N_15500);
or U22014 (N_22014,N_16020,N_17305);
xnor U22015 (N_22015,N_17544,N_14127);
nor U22016 (N_22016,N_12693,N_12552);
and U22017 (N_22017,N_15677,N_16512);
or U22018 (N_22018,N_14093,N_16661);
nor U22019 (N_22019,N_15086,N_15583);
or U22020 (N_22020,N_18730,N_18118);
or U22021 (N_22021,N_18256,N_15501);
xor U22022 (N_22022,N_16811,N_13006);
xnor U22023 (N_22023,N_16370,N_15442);
and U22024 (N_22024,N_16384,N_15286);
or U22025 (N_22025,N_17775,N_15664);
or U22026 (N_22026,N_14498,N_18478);
xor U22027 (N_22027,N_15054,N_15378);
nand U22028 (N_22028,N_15667,N_14615);
and U22029 (N_22029,N_14860,N_16834);
and U22030 (N_22030,N_18412,N_16126);
xnor U22031 (N_22031,N_12764,N_14258);
nand U22032 (N_22032,N_18097,N_16741);
nor U22033 (N_22033,N_17619,N_17704);
xor U22034 (N_22034,N_16250,N_15906);
and U22035 (N_22035,N_18447,N_15609);
or U22036 (N_22036,N_17276,N_12804);
nor U22037 (N_22037,N_13348,N_18126);
xnor U22038 (N_22038,N_16979,N_17625);
nand U22039 (N_22039,N_18693,N_14567);
nor U22040 (N_22040,N_16687,N_17774);
nor U22041 (N_22041,N_15607,N_17900);
nor U22042 (N_22042,N_14099,N_17690);
nand U22043 (N_22043,N_16225,N_14006);
nor U22044 (N_22044,N_12697,N_15013);
nor U22045 (N_22045,N_17470,N_15910);
xnor U22046 (N_22046,N_18032,N_15383);
xnor U22047 (N_22047,N_16172,N_18507);
or U22048 (N_22048,N_13033,N_12983);
and U22049 (N_22049,N_12963,N_14371);
or U22050 (N_22050,N_16896,N_18549);
nor U22051 (N_22051,N_14959,N_18542);
xnor U22052 (N_22052,N_16338,N_18365);
nor U22053 (N_22053,N_14880,N_13372);
nor U22054 (N_22054,N_12574,N_16806);
and U22055 (N_22055,N_13029,N_15910);
or U22056 (N_22056,N_15908,N_16752);
nand U22057 (N_22057,N_17098,N_13954);
nor U22058 (N_22058,N_15405,N_12545);
nor U22059 (N_22059,N_18026,N_12925);
nor U22060 (N_22060,N_14138,N_18082);
and U22061 (N_22061,N_15372,N_18719);
or U22062 (N_22062,N_13306,N_14331);
or U22063 (N_22063,N_16698,N_16516);
and U22064 (N_22064,N_12877,N_16707);
nand U22065 (N_22065,N_16747,N_16515);
and U22066 (N_22066,N_16077,N_15121);
nand U22067 (N_22067,N_17431,N_12774);
nand U22068 (N_22068,N_16885,N_18406);
and U22069 (N_22069,N_17081,N_15097);
nor U22070 (N_22070,N_14219,N_14380);
nor U22071 (N_22071,N_13343,N_15004);
nor U22072 (N_22072,N_14542,N_18107);
and U22073 (N_22073,N_13264,N_17701);
xnor U22074 (N_22074,N_14043,N_13880);
nand U22075 (N_22075,N_12925,N_13739);
nand U22076 (N_22076,N_15790,N_17272);
xnor U22077 (N_22077,N_14784,N_14558);
nand U22078 (N_22078,N_12666,N_16687);
nor U22079 (N_22079,N_14763,N_12906);
and U22080 (N_22080,N_13988,N_17238);
and U22081 (N_22081,N_18588,N_14785);
or U22082 (N_22082,N_15011,N_17882);
xnor U22083 (N_22083,N_14539,N_18696);
xor U22084 (N_22084,N_16657,N_12861);
xnor U22085 (N_22085,N_13445,N_12886);
nor U22086 (N_22086,N_15015,N_16042);
xor U22087 (N_22087,N_13624,N_14989);
nand U22088 (N_22088,N_12556,N_13057);
nand U22089 (N_22089,N_12756,N_17690);
and U22090 (N_22090,N_16589,N_13443);
nand U22091 (N_22091,N_18748,N_14243);
xor U22092 (N_22092,N_16670,N_12613);
and U22093 (N_22093,N_14685,N_13447);
and U22094 (N_22094,N_14434,N_13892);
nand U22095 (N_22095,N_13853,N_12881);
and U22096 (N_22096,N_17874,N_17355);
nor U22097 (N_22097,N_18580,N_12878);
nand U22098 (N_22098,N_17870,N_12914);
nor U22099 (N_22099,N_17503,N_13075);
or U22100 (N_22100,N_18488,N_16971);
nor U22101 (N_22101,N_13597,N_18600);
or U22102 (N_22102,N_15443,N_15738);
or U22103 (N_22103,N_17133,N_12999);
or U22104 (N_22104,N_14665,N_15754);
and U22105 (N_22105,N_18531,N_15404);
or U22106 (N_22106,N_17109,N_15910);
nand U22107 (N_22107,N_14312,N_15148);
nand U22108 (N_22108,N_18419,N_15590);
nor U22109 (N_22109,N_17313,N_17129);
and U22110 (N_22110,N_13878,N_13698);
and U22111 (N_22111,N_12530,N_13749);
or U22112 (N_22112,N_16788,N_14929);
nor U22113 (N_22113,N_15942,N_16791);
nand U22114 (N_22114,N_17436,N_17252);
or U22115 (N_22115,N_15665,N_15203);
nor U22116 (N_22116,N_16902,N_14579);
or U22117 (N_22117,N_14460,N_14842);
nor U22118 (N_22118,N_13421,N_17561);
or U22119 (N_22119,N_15615,N_17256);
xor U22120 (N_22120,N_15364,N_13401);
or U22121 (N_22121,N_14332,N_14466);
nor U22122 (N_22122,N_13820,N_15305);
nand U22123 (N_22123,N_17696,N_17454);
nor U22124 (N_22124,N_18501,N_16462);
and U22125 (N_22125,N_12849,N_17836);
nand U22126 (N_22126,N_17157,N_14718);
nor U22127 (N_22127,N_14445,N_16140);
xor U22128 (N_22128,N_14797,N_15742);
xnor U22129 (N_22129,N_17323,N_16225);
nor U22130 (N_22130,N_16768,N_16763);
nand U22131 (N_22131,N_17892,N_13737);
nor U22132 (N_22132,N_15372,N_13462);
or U22133 (N_22133,N_16519,N_13304);
or U22134 (N_22134,N_14514,N_16238);
and U22135 (N_22135,N_18310,N_14666);
nand U22136 (N_22136,N_14581,N_12812);
or U22137 (N_22137,N_15279,N_13758);
nor U22138 (N_22138,N_12885,N_17162);
nand U22139 (N_22139,N_14925,N_15246);
or U22140 (N_22140,N_13959,N_13426);
xor U22141 (N_22141,N_14014,N_16596);
nand U22142 (N_22142,N_17266,N_18547);
nand U22143 (N_22143,N_16707,N_16633);
and U22144 (N_22144,N_18445,N_16139);
or U22145 (N_22145,N_16702,N_12514);
or U22146 (N_22146,N_14511,N_12555);
nor U22147 (N_22147,N_17138,N_14642);
nor U22148 (N_22148,N_17086,N_16604);
xnor U22149 (N_22149,N_17249,N_14030);
nor U22150 (N_22150,N_13386,N_18546);
nand U22151 (N_22151,N_16205,N_13435);
and U22152 (N_22152,N_12801,N_13359);
xnor U22153 (N_22153,N_18272,N_12657);
xnor U22154 (N_22154,N_15496,N_16618);
and U22155 (N_22155,N_16082,N_15417);
nand U22156 (N_22156,N_14640,N_14674);
or U22157 (N_22157,N_13174,N_14921);
nand U22158 (N_22158,N_13010,N_17899);
nand U22159 (N_22159,N_17561,N_15445);
or U22160 (N_22160,N_16799,N_14213);
nand U22161 (N_22161,N_13799,N_14573);
nand U22162 (N_22162,N_15044,N_13629);
nor U22163 (N_22163,N_15514,N_14565);
or U22164 (N_22164,N_12793,N_13471);
or U22165 (N_22165,N_15322,N_15145);
nor U22166 (N_22166,N_16597,N_12674);
and U22167 (N_22167,N_16625,N_12830);
and U22168 (N_22168,N_13782,N_17960);
or U22169 (N_22169,N_16505,N_16370);
nand U22170 (N_22170,N_17819,N_15851);
xor U22171 (N_22171,N_16758,N_15192);
nand U22172 (N_22172,N_15949,N_16336);
or U22173 (N_22173,N_16406,N_14636);
nor U22174 (N_22174,N_13150,N_15860);
xnor U22175 (N_22175,N_17779,N_12964);
nand U22176 (N_22176,N_13128,N_14993);
nand U22177 (N_22177,N_13172,N_16361);
nor U22178 (N_22178,N_16485,N_15026);
or U22179 (N_22179,N_15817,N_17688);
or U22180 (N_22180,N_12758,N_13177);
xor U22181 (N_22181,N_14887,N_14128);
nand U22182 (N_22182,N_13900,N_12951);
or U22183 (N_22183,N_16532,N_12886);
nand U22184 (N_22184,N_12798,N_18597);
xnor U22185 (N_22185,N_15001,N_13297);
nand U22186 (N_22186,N_12529,N_15436);
or U22187 (N_22187,N_17143,N_15740);
xor U22188 (N_22188,N_16459,N_15572);
xnor U22189 (N_22189,N_15454,N_14076);
nand U22190 (N_22190,N_14036,N_15557);
nor U22191 (N_22191,N_15756,N_13805);
or U22192 (N_22192,N_15982,N_15977);
xnor U22193 (N_22193,N_15646,N_18165);
nand U22194 (N_22194,N_17644,N_16028);
xor U22195 (N_22195,N_14209,N_17376);
xor U22196 (N_22196,N_14570,N_15552);
or U22197 (N_22197,N_13425,N_14992);
and U22198 (N_22198,N_18277,N_15786);
and U22199 (N_22199,N_14846,N_13922);
xor U22200 (N_22200,N_16002,N_16267);
and U22201 (N_22201,N_15302,N_17235);
nor U22202 (N_22202,N_17167,N_15383);
or U22203 (N_22203,N_18078,N_16323);
or U22204 (N_22204,N_12518,N_14886);
or U22205 (N_22205,N_15774,N_17277);
and U22206 (N_22206,N_16569,N_17956);
xor U22207 (N_22207,N_14538,N_14242);
nand U22208 (N_22208,N_15576,N_12966);
nand U22209 (N_22209,N_16662,N_17472);
or U22210 (N_22210,N_17298,N_18427);
nor U22211 (N_22211,N_16489,N_17155);
nor U22212 (N_22212,N_18660,N_14581);
or U22213 (N_22213,N_17934,N_16219);
nor U22214 (N_22214,N_13600,N_17832);
nand U22215 (N_22215,N_12742,N_13973);
and U22216 (N_22216,N_14276,N_13246);
or U22217 (N_22217,N_13259,N_16993);
or U22218 (N_22218,N_13106,N_15083);
xnor U22219 (N_22219,N_14385,N_15486);
nor U22220 (N_22220,N_16083,N_15285);
nor U22221 (N_22221,N_13985,N_16008);
nand U22222 (N_22222,N_14972,N_13401);
nand U22223 (N_22223,N_15116,N_15145);
nand U22224 (N_22224,N_13210,N_12774);
and U22225 (N_22225,N_17945,N_13470);
nor U22226 (N_22226,N_13636,N_12590);
xnor U22227 (N_22227,N_18192,N_16086);
xor U22228 (N_22228,N_13053,N_18617);
and U22229 (N_22229,N_18584,N_15470);
and U22230 (N_22230,N_18698,N_18236);
xnor U22231 (N_22231,N_14038,N_15513);
xor U22232 (N_22232,N_13018,N_15574);
nor U22233 (N_22233,N_16880,N_17067);
or U22234 (N_22234,N_15618,N_18515);
nor U22235 (N_22235,N_18254,N_17536);
nor U22236 (N_22236,N_18557,N_15757);
and U22237 (N_22237,N_18574,N_14799);
and U22238 (N_22238,N_12577,N_17809);
nand U22239 (N_22239,N_12671,N_12962);
xnor U22240 (N_22240,N_13069,N_14614);
nor U22241 (N_22241,N_17436,N_12539);
nor U22242 (N_22242,N_16043,N_17693);
xor U22243 (N_22243,N_16553,N_12804);
xnor U22244 (N_22244,N_15326,N_13981);
xor U22245 (N_22245,N_16720,N_16885);
and U22246 (N_22246,N_12605,N_17662);
nor U22247 (N_22247,N_15781,N_15107);
or U22248 (N_22248,N_13077,N_13498);
and U22249 (N_22249,N_16659,N_16406);
xor U22250 (N_22250,N_18057,N_16275);
nor U22251 (N_22251,N_16294,N_18217);
or U22252 (N_22252,N_18080,N_16212);
or U22253 (N_22253,N_16678,N_13216);
and U22254 (N_22254,N_18383,N_12794);
nor U22255 (N_22255,N_15264,N_15504);
nand U22256 (N_22256,N_12821,N_13219);
and U22257 (N_22257,N_17431,N_13177);
and U22258 (N_22258,N_17255,N_18056);
nand U22259 (N_22259,N_17344,N_14529);
nor U22260 (N_22260,N_14567,N_16167);
xor U22261 (N_22261,N_15612,N_17280);
or U22262 (N_22262,N_12572,N_15651);
nor U22263 (N_22263,N_15566,N_13493);
nor U22264 (N_22264,N_17807,N_16973);
nand U22265 (N_22265,N_14588,N_18035);
xnor U22266 (N_22266,N_12575,N_16811);
xnor U22267 (N_22267,N_13909,N_18228);
or U22268 (N_22268,N_13873,N_14773);
or U22269 (N_22269,N_17782,N_13603);
nor U22270 (N_22270,N_16128,N_17408);
or U22271 (N_22271,N_17244,N_15264);
and U22272 (N_22272,N_17243,N_12614);
and U22273 (N_22273,N_15392,N_15229);
and U22274 (N_22274,N_14174,N_12741);
xnor U22275 (N_22275,N_12618,N_17448);
and U22276 (N_22276,N_16172,N_12736);
xor U22277 (N_22277,N_13591,N_15067);
xnor U22278 (N_22278,N_13111,N_13893);
or U22279 (N_22279,N_13292,N_16678);
xor U22280 (N_22280,N_13736,N_17659);
nor U22281 (N_22281,N_15875,N_14213);
nand U22282 (N_22282,N_12839,N_16196);
and U22283 (N_22283,N_15944,N_18624);
and U22284 (N_22284,N_15312,N_13673);
or U22285 (N_22285,N_15291,N_15449);
xnor U22286 (N_22286,N_14205,N_14133);
nor U22287 (N_22287,N_14784,N_16461);
and U22288 (N_22288,N_16783,N_17909);
or U22289 (N_22289,N_13742,N_16366);
nand U22290 (N_22290,N_17522,N_13176);
nand U22291 (N_22291,N_17076,N_16190);
xnor U22292 (N_22292,N_13831,N_12936);
nand U22293 (N_22293,N_17009,N_17044);
nand U22294 (N_22294,N_18499,N_13546);
or U22295 (N_22295,N_18176,N_17474);
and U22296 (N_22296,N_17552,N_14137);
and U22297 (N_22297,N_12805,N_12919);
xnor U22298 (N_22298,N_13040,N_18743);
and U22299 (N_22299,N_15776,N_16084);
and U22300 (N_22300,N_14926,N_14025);
or U22301 (N_22301,N_16480,N_15820);
xor U22302 (N_22302,N_14961,N_15796);
xor U22303 (N_22303,N_13570,N_13637);
or U22304 (N_22304,N_14963,N_17156);
and U22305 (N_22305,N_12907,N_17621);
nand U22306 (N_22306,N_13271,N_17565);
or U22307 (N_22307,N_13189,N_12702);
and U22308 (N_22308,N_17404,N_16239);
nand U22309 (N_22309,N_13557,N_13145);
xnor U22310 (N_22310,N_13670,N_16302);
and U22311 (N_22311,N_13710,N_15501);
or U22312 (N_22312,N_14087,N_15805);
or U22313 (N_22313,N_18518,N_16253);
and U22314 (N_22314,N_17551,N_15403);
and U22315 (N_22315,N_16798,N_18228);
and U22316 (N_22316,N_15761,N_13062);
xor U22317 (N_22317,N_12929,N_13114);
or U22318 (N_22318,N_13445,N_16577);
and U22319 (N_22319,N_17832,N_13400);
nor U22320 (N_22320,N_14761,N_13614);
xnor U22321 (N_22321,N_14746,N_13358);
xnor U22322 (N_22322,N_14211,N_17633);
nand U22323 (N_22323,N_12939,N_15059);
and U22324 (N_22324,N_16154,N_14817);
xor U22325 (N_22325,N_17395,N_17388);
xor U22326 (N_22326,N_16881,N_14603);
and U22327 (N_22327,N_16356,N_14187);
xor U22328 (N_22328,N_18734,N_16543);
nand U22329 (N_22329,N_15530,N_15776);
nor U22330 (N_22330,N_13664,N_13751);
nand U22331 (N_22331,N_18015,N_17305);
nor U22332 (N_22332,N_17266,N_12651);
or U22333 (N_22333,N_12620,N_15294);
nand U22334 (N_22334,N_17838,N_14345);
xnor U22335 (N_22335,N_18041,N_13952);
and U22336 (N_22336,N_13553,N_16170);
xnor U22337 (N_22337,N_15662,N_16768);
nor U22338 (N_22338,N_13092,N_18193);
nor U22339 (N_22339,N_18467,N_14345);
or U22340 (N_22340,N_18083,N_14779);
and U22341 (N_22341,N_18389,N_18511);
xor U22342 (N_22342,N_16166,N_14413);
xor U22343 (N_22343,N_12736,N_18285);
nor U22344 (N_22344,N_15049,N_17235);
nand U22345 (N_22345,N_12545,N_18567);
nand U22346 (N_22346,N_15788,N_16433);
and U22347 (N_22347,N_14492,N_16461);
and U22348 (N_22348,N_17673,N_15970);
nand U22349 (N_22349,N_17126,N_17623);
or U22350 (N_22350,N_17888,N_17384);
xor U22351 (N_22351,N_15438,N_17653);
or U22352 (N_22352,N_14040,N_16593);
and U22353 (N_22353,N_13282,N_17732);
xor U22354 (N_22354,N_17593,N_14100);
and U22355 (N_22355,N_17705,N_17998);
or U22356 (N_22356,N_12592,N_15412);
nor U22357 (N_22357,N_13758,N_18058);
and U22358 (N_22358,N_18473,N_13830);
nor U22359 (N_22359,N_15443,N_16337);
xnor U22360 (N_22360,N_12690,N_12792);
nand U22361 (N_22361,N_17102,N_15561);
nand U22362 (N_22362,N_16034,N_13046);
or U22363 (N_22363,N_13556,N_13229);
and U22364 (N_22364,N_15156,N_14200);
nor U22365 (N_22365,N_12948,N_12525);
and U22366 (N_22366,N_15589,N_14932);
or U22367 (N_22367,N_12924,N_17451);
or U22368 (N_22368,N_14092,N_12819);
xor U22369 (N_22369,N_16500,N_13725);
xor U22370 (N_22370,N_14277,N_13160);
and U22371 (N_22371,N_15274,N_15659);
or U22372 (N_22372,N_13474,N_18735);
nor U22373 (N_22373,N_13339,N_12938);
xnor U22374 (N_22374,N_18250,N_14517);
or U22375 (N_22375,N_17267,N_16197);
xor U22376 (N_22376,N_13379,N_15315);
xor U22377 (N_22377,N_16214,N_17644);
or U22378 (N_22378,N_18685,N_15822);
xnor U22379 (N_22379,N_13814,N_16969);
nor U22380 (N_22380,N_16363,N_15518);
and U22381 (N_22381,N_16571,N_13457);
and U22382 (N_22382,N_13217,N_13139);
nor U22383 (N_22383,N_14765,N_15593);
or U22384 (N_22384,N_14088,N_13934);
nand U22385 (N_22385,N_13476,N_15623);
or U22386 (N_22386,N_16662,N_15739);
and U22387 (N_22387,N_13379,N_14837);
nor U22388 (N_22388,N_14857,N_17345);
nand U22389 (N_22389,N_16277,N_17702);
nor U22390 (N_22390,N_17074,N_17895);
xnor U22391 (N_22391,N_17640,N_12647);
nor U22392 (N_22392,N_14090,N_14166);
or U22393 (N_22393,N_16684,N_12673);
or U22394 (N_22394,N_13326,N_13047);
or U22395 (N_22395,N_16576,N_16640);
and U22396 (N_22396,N_15874,N_15052);
and U22397 (N_22397,N_17329,N_17143);
or U22398 (N_22398,N_13714,N_13409);
or U22399 (N_22399,N_16732,N_14880);
nand U22400 (N_22400,N_18333,N_16762);
and U22401 (N_22401,N_15443,N_15104);
xnor U22402 (N_22402,N_16103,N_14543);
xnor U22403 (N_22403,N_12761,N_14744);
nor U22404 (N_22404,N_16393,N_12768);
nor U22405 (N_22405,N_17674,N_18481);
or U22406 (N_22406,N_18297,N_13372);
xnor U22407 (N_22407,N_14800,N_13768);
or U22408 (N_22408,N_12702,N_16174);
nor U22409 (N_22409,N_17386,N_15843);
or U22410 (N_22410,N_14725,N_13208);
nor U22411 (N_22411,N_13832,N_13932);
or U22412 (N_22412,N_18589,N_17124);
xnor U22413 (N_22413,N_13755,N_17608);
and U22414 (N_22414,N_14456,N_15386);
xnor U22415 (N_22415,N_13101,N_13535);
nand U22416 (N_22416,N_18681,N_14695);
xor U22417 (N_22417,N_16952,N_18010);
nor U22418 (N_22418,N_16090,N_14671);
or U22419 (N_22419,N_16905,N_17817);
or U22420 (N_22420,N_17777,N_13550);
xor U22421 (N_22421,N_14493,N_17950);
or U22422 (N_22422,N_15441,N_18698);
nor U22423 (N_22423,N_12584,N_13587);
nand U22424 (N_22424,N_17734,N_13086);
or U22425 (N_22425,N_17149,N_15057);
nor U22426 (N_22426,N_14818,N_17452);
nor U22427 (N_22427,N_14018,N_17749);
and U22428 (N_22428,N_17694,N_13753);
and U22429 (N_22429,N_14580,N_13106);
and U22430 (N_22430,N_15480,N_15360);
nor U22431 (N_22431,N_14558,N_16022);
or U22432 (N_22432,N_16751,N_15146);
nand U22433 (N_22433,N_13237,N_13983);
or U22434 (N_22434,N_14252,N_15679);
xor U22435 (N_22435,N_13585,N_17110);
and U22436 (N_22436,N_12790,N_18644);
xnor U22437 (N_22437,N_13255,N_17129);
nand U22438 (N_22438,N_14380,N_15143);
or U22439 (N_22439,N_13700,N_16662);
nand U22440 (N_22440,N_16130,N_17479);
nor U22441 (N_22441,N_13435,N_14242);
or U22442 (N_22442,N_14954,N_18426);
nor U22443 (N_22443,N_13468,N_18138);
xor U22444 (N_22444,N_16919,N_14096);
nor U22445 (N_22445,N_13041,N_17160);
xnor U22446 (N_22446,N_13317,N_16534);
or U22447 (N_22447,N_14420,N_18664);
or U22448 (N_22448,N_18421,N_17999);
or U22449 (N_22449,N_15851,N_14371);
xnor U22450 (N_22450,N_14300,N_14792);
and U22451 (N_22451,N_13759,N_18146);
nand U22452 (N_22452,N_13273,N_16631);
or U22453 (N_22453,N_15685,N_13805);
xor U22454 (N_22454,N_16912,N_13325);
nor U22455 (N_22455,N_14624,N_16967);
or U22456 (N_22456,N_14742,N_14239);
and U22457 (N_22457,N_17594,N_16278);
nand U22458 (N_22458,N_12714,N_14265);
and U22459 (N_22459,N_13599,N_12641);
nand U22460 (N_22460,N_15047,N_16878);
or U22461 (N_22461,N_17342,N_14245);
nand U22462 (N_22462,N_16934,N_16184);
nand U22463 (N_22463,N_15953,N_17431);
and U22464 (N_22464,N_16955,N_16445);
nor U22465 (N_22465,N_18704,N_14543);
nor U22466 (N_22466,N_13574,N_16757);
and U22467 (N_22467,N_18238,N_16902);
xnor U22468 (N_22468,N_14943,N_16133);
nand U22469 (N_22469,N_18630,N_13801);
nor U22470 (N_22470,N_17519,N_16528);
nor U22471 (N_22471,N_17191,N_13893);
xor U22472 (N_22472,N_16299,N_13033);
nand U22473 (N_22473,N_13350,N_13373);
nor U22474 (N_22474,N_16597,N_16344);
and U22475 (N_22475,N_17435,N_13319);
nand U22476 (N_22476,N_18575,N_14372);
or U22477 (N_22477,N_18212,N_17865);
nor U22478 (N_22478,N_14552,N_18494);
and U22479 (N_22479,N_15930,N_13355);
nor U22480 (N_22480,N_16469,N_14159);
nand U22481 (N_22481,N_16294,N_17441);
nor U22482 (N_22482,N_13182,N_17912);
nor U22483 (N_22483,N_17805,N_14155);
or U22484 (N_22484,N_17897,N_13683);
xor U22485 (N_22485,N_13610,N_17669);
and U22486 (N_22486,N_16488,N_14144);
and U22487 (N_22487,N_16715,N_13163);
nand U22488 (N_22488,N_17366,N_16556);
and U22489 (N_22489,N_14001,N_13006);
or U22490 (N_22490,N_17682,N_14620);
and U22491 (N_22491,N_14128,N_18051);
nor U22492 (N_22492,N_18403,N_12543);
nor U22493 (N_22493,N_15744,N_18170);
nor U22494 (N_22494,N_16247,N_13639);
xor U22495 (N_22495,N_15525,N_12698);
xnor U22496 (N_22496,N_14057,N_15157);
or U22497 (N_22497,N_16113,N_13203);
xor U22498 (N_22498,N_18209,N_16873);
xnor U22499 (N_22499,N_13125,N_16210);
or U22500 (N_22500,N_14948,N_18680);
nor U22501 (N_22501,N_12924,N_15024);
and U22502 (N_22502,N_15036,N_14240);
nor U22503 (N_22503,N_16812,N_15541);
nor U22504 (N_22504,N_16498,N_18005);
or U22505 (N_22505,N_18553,N_18476);
nand U22506 (N_22506,N_18054,N_14916);
and U22507 (N_22507,N_13851,N_15610);
and U22508 (N_22508,N_13907,N_15999);
nor U22509 (N_22509,N_12833,N_13593);
or U22510 (N_22510,N_16266,N_14032);
or U22511 (N_22511,N_15731,N_17790);
nor U22512 (N_22512,N_12961,N_12592);
and U22513 (N_22513,N_15696,N_14264);
nor U22514 (N_22514,N_16933,N_18326);
nand U22515 (N_22515,N_18692,N_13726);
xor U22516 (N_22516,N_14269,N_18691);
xnor U22517 (N_22517,N_13181,N_12787);
nand U22518 (N_22518,N_15582,N_16333);
nand U22519 (N_22519,N_15302,N_14338);
xor U22520 (N_22520,N_13906,N_18456);
and U22521 (N_22521,N_18314,N_16573);
and U22522 (N_22522,N_15841,N_15157);
xnor U22523 (N_22523,N_15067,N_18476);
nor U22524 (N_22524,N_16257,N_14852);
and U22525 (N_22525,N_15957,N_14281);
nand U22526 (N_22526,N_12585,N_16431);
and U22527 (N_22527,N_13840,N_18349);
nand U22528 (N_22528,N_16433,N_12975);
or U22529 (N_22529,N_18085,N_13917);
xnor U22530 (N_22530,N_15942,N_15813);
nand U22531 (N_22531,N_13831,N_13948);
nor U22532 (N_22532,N_17986,N_15840);
nor U22533 (N_22533,N_14556,N_14527);
nor U22534 (N_22534,N_16368,N_13026);
xnor U22535 (N_22535,N_16718,N_18049);
nand U22536 (N_22536,N_16709,N_12664);
xnor U22537 (N_22537,N_16897,N_14783);
or U22538 (N_22538,N_13895,N_16929);
and U22539 (N_22539,N_14920,N_15194);
nor U22540 (N_22540,N_12762,N_15892);
nand U22541 (N_22541,N_13380,N_17692);
nand U22542 (N_22542,N_17912,N_15738);
or U22543 (N_22543,N_14340,N_13297);
or U22544 (N_22544,N_14132,N_14454);
or U22545 (N_22545,N_14538,N_15993);
nor U22546 (N_22546,N_16649,N_18253);
and U22547 (N_22547,N_17157,N_16097);
or U22548 (N_22548,N_16781,N_12517);
nand U22549 (N_22549,N_13667,N_15448);
nor U22550 (N_22550,N_16279,N_18743);
xnor U22551 (N_22551,N_14488,N_15854);
and U22552 (N_22552,N_16767,N_17187);
nand U22553 (N_22553,N_15176,N_14200);
nand U22554 (N_22554,N_15629,N_18229);
and U22555 (N_22555,N_15659,N_18136);
nor U22556 (N_22556,N_14396,N_18185);
xor U22557 (N_22557,N_12516,N_17372);
nand U22558 (N_22558,N_13029,N_18131);
nor U22559 (N_22559,N_13164,N_12781);
xnor U22560 (N_22560,N_13913,N_14766);
nor U22561 (N_22561,N_18172,N_13895);
nor U22562 (N_22562,N_16486,N_17158);
xnor U22563 (N_22563,N_16861,N_18231);
nand U22564 (N_22564,N_14180,N_15881);
and U22565 (N_22565,N_15559,N_12982);
xor U22566 (N_22566,N_15450,N_14951);
xor U22567 (N_22567,N_16455,N_13856);
and U22568 (N_22568,N_15754,N_17324);
nor U22569 (N_22569,N_15537,N_15883);
nand U22570 (N_22570,N_15974,N_13244);
or U22571 (N_22571,N_17930,N_17751);
or U22572 (N_22572,N_16148,N_17561);
nand U22573 (N_22573,N_17685,N_18349);
xnor U22574 (N_22574,N_17363,N_17504);
and U22575 (N_22575,N_13494,N_18103);
nand U22576 (N_22576,N_17718,N_15972);
or U22577 (N_22577,N_15703,N_16769);
nor U22578 (N_22578,N_18409,N_13505);
and U22579 (N_22579,N_15024,N_15942);
xnor U22580 (N_22580,N_14845,N_16433);
nand U22581 (N_22581,N_17707,N_13749);
xor U22582 (N_22582,N_13863,N_12570);
nand U22583 (N_22583,N_16566,N_17866);
nand U22584 (N_22584,N_17831,N_14471);
or U22585 (N_22585,N_17307,N_15987);
or U22586 (N_22586,N_12849,N_15742);
or U22587 (N_22587,N_16014,N_13651);
nor U22588 (N_22588,N_15978,N_13279);
and U22589 (N_22589,N_17151,N_14449);
and U22590 (N_22590,N_12765,N_12827);
xnor U22591 (N_22591,N_13564,N_13883);
nand U22592 (N_22592,N_17607,N_16815);
xor U22593 (N_22593,N_14824,N_14002);
and U22594 (N_22594,N_18458,N_16611);
nand U22595 (N_22595,N_16008,N_18564);
or U22596 (N_22596,N_18684,N_14742);
nor U22597 (N_22597,N_17720,N_16980);
xnor U22598 (N_22598,N_14220,N_16025);
and U22599 (N_22599,N_13230,N_15299);
and U22600 (N_22600,N_18447,N_12989);
or U22601 (N_22601,N_16966,N_17983);
xnor U22602 (N_22602,N_17288,N_16838);
xor U22603 (N_22603,N_17793,N_16072);
and U22604 (N_22604,N_17640,N_12931);
or U22605 (N_22605,N_18646,N_16893);
nand U22606 (N_22606,N_13153,N_12864);
nor U22607 (N_22607,N_15128,N_15858);
xor U22608 (N_22608,N_13829,N_13910);
and U22609 (N_22609,N_16632,N_15727);
xor U22610 (N_22610,N_18061,N_14900);
nor U22611 (N_22611,N_16704,N_15664);
nand U22612 (N_22612,N_17248,N_16955);
xnor U22613 (N_22613,N_17690,N_13317);
or U22614 (N_22614,N_13313,N_13487);
or U22615 (N_22615,N_18564,N_17916);
and U22616 (N_22616,N_12617,N_16099);
or U22617 (N_22617,N_16535,N_15548);
and U22618 (N_22618,N_17629,N_18595);
nor U22619 (N_22619,N_13934,N_16259);
nor U22620 (N_22620,N_14071,N_16753);
or U22621 (N_22621,N_16503,N_15710);
xnor U22622 (N_22622,N_15990,N_15474);
and U22623 (N_22623,N_15781,N_17160);
nor U22624 (N_22624,N_17544,N_13038);
nor U22625 (N_22625,N_14194,N_12875);
nor U22626 (N_22626,N_14257,N_17070);
and U22627 (N_22627,N_14939,N_13154);
nand U22628 (N_22628,N_13645,N_17763);
or U22629 (N_22629,N_13008,N_13153);
or U22630 (N_22630,N_18426,N_17069);
or U22631 (N_22631,N_17074,N_12560);
and U22632 (N_22632,N_15496,N_17388);
xnor U22633 (N_22633,N_13188,N_18057);
or U22634 (N_22634,N_15957,N_16693);
xor U22635 (N_22635,N_13357,N_16075);
or U22636 (N_22636,N_16455,N_16469);
or U22637 (N_22637,N_14363,N_15966);
xnor U22638 (N_22638,N_18138,N_17617);
xnor U22639 (N_22639,N_17168,N_17468);
nand U22640 (N_22640,N_13913,N_18477);
and U22641 (N_22641,N_15511,N_17122);
nor U22642 (N_22642,N_18478,N_17564);
nand U22643 (N_22643,N_16960,N_14133);
xnor U22644 (N_22644,N_12642,N_18712);
xnor U22645 (N_22645,N_18514,N_18398);
xor U22646 (N_22646,N_15944,N_17227);
nand U22647 (N_22647,N_13971,N_13209);
and U22648 (N_22648,N_15211,N_14986);
and U22649 (N_22649,N_14140,N_17633);
nor U22650 (N_22650,N_14721,N_15196);
xnor U22651 (N_22651,N_18619,N_13189);
or U22652 (N_22652,N_14748,N_14384);
xnor U22653 (N_22653,N_14697,N_13255);
and U22654 (N_22654,N_13643,N_16955);
nor U22655 (N_22655,N_14521,N_17754);
xnor U22656 (N_22656,N_15786,N_15494);
nand U22657 (N_22657,N_16263,N_17042);
nor U22658 (N_22658,N_18326,N_17303);
or U22659 (N_22659,N_12582,N_16743);
and U22660 (N_22660,N_17175,N_14181);
and U22661 (N_22661,N_17742,N_13233);
and U22662 (N_22662,N_13978,N_15591);
nand U22663 (N_22663,N_14901,N_15699);
xnor U22664 (N_22664,N_17329,N_12789);
and U22665 (N_22665,N_14780,N_13720);
nor U22666 (N_22666,N_16796,N_18468);
and U22667 (N_22667,N_13618,N_15252);
nor U22668 (N_22668,N_13091,N_15891);
and U22669 (N_22669,N_17869,N_14384);
and U22670 (N_22670,N_16120,N_15903);
or U22671 (N_22671,N_13772,N_17039);
nand U22672 (N_22672,N_17824,N_12995);
nor U22673 (N_22673,N_13281,N_18619);
and U22674 (N_22674,N_15461,N_12948);
nor U22675 (N_22675,N_17939,N_13996);
nor U22676 (N_22676,N_17311,N_15453);
nor U22677 (N_22677,N_14955,N_12910);
and U22678 (N_22678,N_16862,N_16708);
and U22679 (N_22679,N_15786,N_15357);
or U22680 (N_22680,N_16308,N_15094);
nand U22681 (N_22681,N_16879,N_16618);
or U22682 (N_22682,N_14391,N_14890);
nand U22683 (N_22683,N_16916,N_13637);
nand U22684 (N_22684,N_14510,N_12890);
nand U22685 (N_22685,N_16512,N_17792);
and U22686 (N_22686,N_17727,N_16834);
nor U22687 (N_22687,N_15124,N_16949);
and U22688 (N_22688,N_17595,N_16593);
and U22689 (N_22689,N_13006,N_18496);
nor U22690 (N_22690,N_18670,N_14824);
xnor U22691 (N_22691,N_18658,N_15214);
xnor U22692 (N_22692,N_15619,N_16662);
nand U22693 (N_22693,N_14605,N_15331);
and U22694 (N_22694,N_13553,N_17498);
xor U22695 (N_22695,N_14013,N_15216);
or U22696 (N_22696,N_17977,N_12709);
xor U22697 (N_22697,N_15549,N_14647);
nor U22698 (N_22698,N_14283,N_14892);
or U22699 (N_22699,N_16747,N_13884);
nand U22700 (N_22700,N_18162,N_18012);
or U22701 (N_22701,N_18496,N_15709);
nand U22702 (N_22702,N_14157,N_12799);
nor U22703 (N_22703,N_13665,N_13063);
or U22704 (N_22704,N_13682,N_14359);
xnor U22705 (N_22705,N_18470,N_14623);
and U22706 (N_22706,N_13333,N_14350);
xor U22707 (N_22707,N_14984,N_17532);
xnor U22708 (N_22708,N_12954,N_14696);
and U22709 (N_22709,N_12689,N_14466);
or U22710 (N_22710,N_15607,N_12558);
xor U22711 (N_22711,N_13205,N_13118);
or U22712 (N_22712,N_13387,N_13215);
and U22713 (N_22713,N_15534,N_16984);
xnor U22714 (N_22714,N_18569,N_18659);
nand U22715 (N_22715,N_16865,N_17024);
and U22716 (N_22716,N_15965,N_17145);
or U22717 (N_22717,N_14293,N_13075);
nand U22718 (N_22718,N_13463,N_18535);
and U22719 (N_22719,N_14515,N_15461);
nand U22720 (N_22720,N_14367,N_16879);
xnor U22721 (N_22721,N_14092,N_17566);
nor U22722 (N_22722,N_16115,N_17340);
nand U22723 (N_22723,N_15999,N_16800);
nor U22724 (N_22724,N_18175,N_12678);
nand U22725 (N_22725,N_14861,N_16490);
nand U22726 (N_22726,N_18308,N_14322);
xnor U22727 (N_22727,N_15575,N_13392);
xor U22728 (N_22728,N_18688,N_13893);
nor U22729 (N_22729,N_13237,N_18335);
xor U22730 (N_22730,N_17691,N_16373);
nor U22731 (N_22731,N_14234,N_14362);
nand U22732 (N_22732,N_13284,N_15336);
or U22733 (N_22733,N_13456,N_15609);
and U22734 (N_22734,N_15014,N_13245);
xor U22735 (N_22735,N_16352,N_17845);
nand U22736 (N_22736,N_18156,N_14836);
and U22737 (N_22737,N_15864,N_16207);
and U22738 (N_22738,N_14663,N_18367);
and U22739 (N_22739,N_13232,N_16999);
nand U22740 (N_22740,N_13289,N_18654);
nor U22741 (N_22741,N_17657,N_17781);
nor U22742 (N_22742,N_14684,N_15026);
or U22743 (N_22743,N_14616,N_13029);
and U22744 (N_22744,N_16159,N_13231);
nor U22745 (N_22745,N_14499,N_15206);
or U22746 (N_22746,N_14024,N_15078);
and U22747 (N_22747,N_18386,N_17056);
or U22748 (N_22748,N_14812,N_14049);
nor U22749 (N_22749,N_15609,N_17304);
and U22750 (N_22750,N_12721,N_16248);
xnor U22751 (N_22751,N_17296,N_14753);
or U22752 (N_22752,N_18043,N_15278);
nor U22753 (N_22753,N_17742,N_16701);
nand U22754 (N_22754,N_16523,N_16813);
nand U22755 (N_22755,N_16392,N_14579);
xor U22756 (N_22756,N_13390,N_18316);
or U22757 (N_22757,N_15101,N_13288);
nor U22758 (N_22758,N_17395,N_18708);
and U22759 (N_22759,N_14833,N_18484);
nand U22760 (N_22760,N_15988,N_14501);
and U22761 (N_22761,N_13423,N_12605);
nor U22762 (N_22762,N_14392,N_16692);
or U22763 (N_22763,N_14843,N_15536);
xor U22764 (N_22764,N_13607,N_14325);
or U22765 (N_22765,N_16185,N_15610);
xor U22766 (N_22766,N_14424,N_18284);
or U22767 (N_22767,N_16159,N_18707);
or U22768 (N_22768,N_18283,N_17064);
xor U22769 (N_22769,N_13756,N_15672);
nand U22770 (N_22770,N_13486,N_14348);
nor U22771 (N_22771,N_17831,N_16006);
nand U22772 (N_22772,N_14606,N_13728);
and U22773 (N_22773,N_16090,N_15153);
xor U22774 (N_22774,N_15237,N_12925);
or U22775 (N_22775,N_17395,N_14242);
xnor U22776 (N_22776,N_17522,N_12838);
and U22777 (N_22777,N_15720,N_15117);
and U22778 (N_22778,N_15912,N_13554);
nor U22779 (N_22779,N_13121,N_14805);
nand U22780 (N_22780,N_15669,N_17633);
or U22781 (N_22781,N_13540,N_17415);
and U22782 (N_22782,N_12674,N_17422);
xnor U22783 (N_22783,N_16191,N_14994);
and U22784 (N_22784,N_12972,N_16960);
nor U22785 (N_22785,N_15062,N_13477);
nand U22786 (N_22786,N_18680,N_12537);
and U22787 (N_22787,N_12992,N_15553);
or U22788 (N_22788,N_14264,N_16538);
xnor U22789 (N_22789,N_15645,N_13998);
and U22790 (N_22790,N_17399,N_18527);
or U22791 (N_22791,N_12775,N_14466);
nand U22792 (N_22792,N_13428,N_12507);
nor U22793 (N_22793,N_13001,N_18230);
nand U22794 (N_22794,N_12615,N_17737);
nand U22795 (N_22795,N_18333,N_13561);
nand U22796 (N_22796,N_18483,N_13792);
xnor U22797 (N_22797,N_16237,N_17984);
xnor U22798 (N_22798,N_14791,N_13336);
nand U22799 (N_22799,N_16899,N_16086);
nor U22800 (N_22800,N_15528,N_12693);
xnor U22801 (N_22801,N_15523,N_13811);
nor U22802 (N_22802,N_16047,N_17573);
or U22803 (N_22803,N_13289,N_14168);
and U22804 (N_22804,N_17609,N_13729);
xnor U22805 (N_22805,N_18411,N_17796);
xor U22806 (N_22806,N_13927,N_13160);
nand U22807 (N_22807,N_13377,N_16725);
xnor U22808 (N_22808,N_14030,N_14333);
nand U22809 (N_22809,N_14980,N_14315);
and U22810 (N_22810,N_12707,N_13923);
nor U22811 (N_22811,N_16127,N_18011);
nand U22812 (N_22812,N_16516,N_18318);
nand U22813 (N_22813,N_12664,N_18736);
nor U22814 (N_22814,N_14799,N_13697);
or U22815 (N_22815,N_17018,N_18550);
xnor U22816 (N_22816,N_17537,N_18186);
nor U22817 (N_22817,N_15917,N_17325);
and U22818 (N_22818,N_15474,N_15960);
nand U22819 (N_22819,N_14303,N_12706);
and U22820 (N_22820,N_18004,N_13546);
xor U22821 (N_22821,N_18251,N_12755);
xnor U22822 (N_22822,N_17692,N_13566);
nand U22823 (N_22823,N_13803,N_13286);
xnor U22824 (N_22824,N_18672,N_15585);
xnor U22825 (N_22825,N_16619,N_13385);
and U22826 (N_22826,N_13221,N_14462);
or U22827 (N_22827,N_12504,N_15910);
or U22828 (N_22828,N_15805,N_14201);
xor U22829 (N_22829,N_17479,N_14635);
and U22830 (N_22830,N_15035,N_15740);
and U22831 (N_22831,N_16307,N_16526);
and U22832 (N_22832,N_14182,N_14344);
xor U22833 (N_22833,N_14718,N_16103);
nand U22834 (N_22834,N_12939,N_17086);
or U22835 (N_22835,N_12858,N_16447);
and U22836 (N_22836,N_17524,N_15269);
nand U22837 (N_22837,N_18703,N_13912);
nor U22838 (N_22838,N_13088,N_13767);
nand U22839 (N_22839,N_13176,N_17113);
nand U22840 (N_22840,N_12705,N_13248);
nand U22841 (N_22841,N_17547,N_17907);
and U22842 (N_22842,N_14379,N_14214);
or U22843 (N_22843,N_12909,N_12694);
and U22844 (N_22844,N_18382,N_17367);
xnor U22845 (N_22845,N_13790,N_18731);
or U22846 (N_22846,N_16775,N_15991);
nand U22847 (N_22847,N_18548,N_13948);
xnor U22848 (N_22848,N_14531,N_14976);
nand U22849 (N_22849,N_17900,N_12999);
and U22850 (N_22850,N_15366,N_14386);
nand U22851 (N_22851,N_15895,N_15948);
or U22852 (N_22852,N_17816,N_13269);
and U22853 (N_22853,N_14353,N_16143);
nor U22854 (N_22854,N_18485,N_15475);
and U22855 (N_22855,N_12756,N_14224);
nand U22856 (N_22856,N_18154,N_13331);
and U22857 (N_22857,N_16227,N_12642);
and U22858 (N_22858,N_14076,N_14811);
and U22859 (N_22859,N_17538,N_17653);
xor U22860 (N_22860,N_18692,N_14901);
and U22861 (N_22861,N_15650,N_15449);
xnor U22862 (N_22862,N_16669,N_12940);
and U22863 (N_22863,N_18448,N_17228);
and U22864 (N_22864,N_14648,N_13318);
nor U22865 (N_22865,N_12905,N_13642);
nor U22866 (N_22866,N_17381,N_16146);
nor U22867 (N_22867,N_13993,N_16157);
or U22868 (N_22868,N_12751,N_13039);
and U22869 (N_22869,N_18391,N_14390);
or U22870 (N_22870,N_16087,N_12714);
nand U22871 (N_22871,N_15699,N_15514);
and U22872 (N_22872,N_18249,N_16000);
nor U22873 (N_22873,N_15978,N_14720);
or U22874 (N_22874,N_16904,N_13012);
nand U22875 (N_22875,N_13268,N_18742);
xnor U22876 (N_22876,N_13545,N_14952);
xnor U22877 (N_22877,N_12541,N_13585);
or U22878 (N_22878,N_15399,N_13840);
xor U22879 (N_22879,N_15109,N_18059);
nor U22880 (N_22880,N_18345,N_17158);
or U22881 (N_22881,N_16232,N_17057);
nor U22882 (N_22882,N_13068,N_16379);
xor U22883 (N_22883,N_12713,N_18165);
and U22884 (N_22884,N_16472,N_12846);
xor U22885 (N_22885,N_14399,N_15336);
nand U22886 (N_22886,N_18148,N_13446);
and U22887 (N_22887,N_14556,N_13230);
xor U22888 (N_22888,N_17275,N_18401);
nand U22889 (N_22889,N_18475,N_14622);
nand U22890 (N_22890,N_15865,N_15886);
and U22891 (N_22891,N_15239,N_17498);
or U22892 (N_22892,N_13270,N_13728);
and U22893 (N_22893,N_15000,N_13662);
and U22894 (N_22894,N_18397,N_14560);
xor U22895 (N_22895,N_15683,N_14342);
xor U22896 (N_22896,N_18190,N_16946);
nand U22897 (N_22897,N_15921,N_15051);
nor U22898 (N_22898,N_18463,N_16070);
nand U22899 (N_22899,N_14012,N_17247);
xor U22900 (N_22900,N_14232,N_15438);
nor U22901 (N_22901,N_14069,N_17568);
and U22902 (N_22902,N_18306,N_17312);
nor U22903 (N_22903,N_13346,N_15854);
and U22904 (N_22904,N_16151,N_15786);
nor U22905 (N_22905,N_18656,N_14517);
xor U22906 (N_22906,N_13799,N_12601);
nor U22907 (N_22907,N_16316,N_13303);
or U22908 (N_22908,N_13030,N_15164);
and U22909 (N_22909,N_13072,N_17279);
nand U22910 (N_22910,N_17908,N_14835);
nand U22911 (N_22911,N_14600,N_12573);
or U22912 (N_22912,N_12572,N_15881);
nor U22913 (N_22913,N_17805,N_16174);
and U22914 (N_22914,N_12863,N_18197);
nor U22915 (N_22915,N_17833,N_13527);
and U22916 (N_22916,N_14240,N_18291);
xnor U22917 (N_22917,N_13541,N_14320);
and U22918 (N_22918,N_12608,N_18114);
or U22919 (N_22919,N_18218,N_15802);
nor U22920 (N_22920,N_15886,N_18737);
or U22921 (N_22921,N_15918,N_14585);
and U22922 (N_22922,N_16883,N_12654);
and U22923 (N_22923,N_16698,N_12712);
nor U22924 (N_22924,N_13332,N_16336);
nand U22925 (N_22925,N_12690,N_13015);
xnor U22926 (N_22926,N_15450,N_14025);
nand U22927 (N_22927,N_14254,N_15833);
or U22928 (N_22928,N_17987,N_13840);
and U22929 (N_22929,N_15378,N_16166);
or U22930 (N_22930,N_16593,N_15496);
nor U22931 (N_22931,N_15890,N_14613);
or U22932 (N_22932,N_18194,N_12587);
and U22933 (N_22933,N_15976,N_14781);
nand U22934 (N_22934,N_18729,N_18671);
nor U22935 (N_22935,N_18309,N_17125);
and U22936 (N_22936,N_16570,N_14941);
nor U22937 (N_22937,N_18019,N_13463);
and U22938 (N_22938,N_16544,N_18337);
or U22939 (N_22939,N_15799,N_14576);
xnor U22940 (N_22940,N_16150,N_13793);
nor U22941 (N_22941,N_15247,N_17741);
nand U22942 (N_22942,N_15619,N_16316);
and U22943 (N_22943,N_18011,N_15938);
nor U22944 (N_22944,N_18133,N_15341);
and U22945 (N_22945,N_13261,N_17617);
and U22946 (N_22946,N_16050,N_13119);
or U22947 (N_22947,N_16560,N_13167);
xor U22948 (N_22948,N_16403,N_18531);
and U22949 (N_22949,N_15269,N_16309);
nand U22950 (N_22950,N_12930,N_16485);
or U22951 (N_22951,N_16004,N_13378);
and U22952 (N_22952,N_13096,N_16190);
nand U22953 (N_22953,N_17567,N_18721);
or U22954 (N_22954,N_13678,N_17679);
nor U22955 (N_22955,N_18064,N_17060);
and U22956 (N_22956,N_14529,N_12784);
or U22957 (N_22957,N_15217,N_15641);
nand U22958 (N_22958,N_17227,N_18683);
xnor U22959 (N_22959,N_16219,N_16475);
nor U22960 (N_22960,N_14305,N_18455);
or U22961 (N_22961,N_16309,N_12941);
xor U22962 (N_22962,N_16594,N_15080);
and U22963 (N_22963,N_13644,N_15841);
xor U22964 (N_22964,N_16722,N_16225);
nor U22965 (N_22965,N_13416,N_18514);
nor U22966 (N_22966,N_13551,N_15928);
nor U22967 (N_22967,N_18368,N_13757);
xor U22968 (N_22968,N_15037,N_15492);
and U22969 (N_22969,N_18532,N_18006);
xnor U22970 (N_22970,N_12779,N_13594);
nor U22971 (N_22971,N_16838,N_13699);
and U22972 (N_22972,N_17257,N_18490);
nand U22973 (N_22973,N_16018,N_18668);
nor U22974 (N_22974,N_15968,N_18077);
and U22975 (N_22975,N_18439,N_16390);
xor U22976 (N_22976,N_15159,N_17873);
and U22977 (N_22977,N_15915,N_15060);
or U22978 (N_22978,N_18556,N_13016);
xnor U22979 (N_22979,N_18695,N_17099);
nand U22980 (N_22980,N_12928,N_14284);
nand U22981 (N_22981,N_14564,N_15811);
nand U22982 (N_22982,N_17455,N_14765);
xnor U22983 (N_22983,N_14204,N_17734);
nor U22984 (N_22984,N_13454,N_16798);
nand U22985 (N_22985,N_18502,N_17310);
xor U22986 (N_22986,N_14877,N_13603);
or U22987 (N_22987,N_16003,N_18130);
and U22988 (N_22988,N_12614,N_13448);
nor U22989 (N_22989,N_13987,N_13671);
nand U22990 (N_22990,N_14381,N_13118);
or U22991 (N_22991,N_18296,N_17378);
xor U22992 (N_22992,N_17330,N_12660);
and U22993 (N_22993,N_12607,N_13609);
and U22994 (N_22994,N_14806,N_15024);
or U22995 (N_22995,N_16432,N_14715);
nand U22996 (N_22996,N_12805,N_15409);
or U22997 (N_22997,N_16249,N_18748);
and U22998 (N_22998,N_12948,N_17583);
and U22999 (N_22999,N_14653,N_14274);
xnor U23000 (N_23000,N_17351,N_16080);
nor U23001 (N_23001,N_16281,N_14057);
and U23002 (N_23002,N_18593,N_13721);
or U23003 (N_23003,N_18208,N_18739);
or U23004 (N_23004,N_18159,N_16399);
nand U23005 (N_23005,N_16174,N_14020);
or U23006 (N_23006,N_17567,N_13550);
nand U23007 (N_23007,N_12862,N_13841);
xnor U23008 (N_23008,N_12983,N_16480);
and U23009 (N_23009,N_12926,N_16400);
nor U23010 (N_23010,N_18089,N_18328);
xor U23011 (N_23011,N_13092,N_17729);
xnor U23012 (N_23012,N_18023,N_17282);
nor U23013 (N_23013,N_17625,N_17159);
or U23014 (N_23014,N_17232,N_12747);
xor U23015 (N_23015,N_15778,N_13941);
or U23016 (N_23016,N_13017,N_14587);
xor U23017 (N_23017,N_17696,N_13455);
nor U23018 (N_23018,N_16032,N_18001);
nand U23019 (N_23019,N_14069,N_15915);
nor U23020 (N_23020,N_15926,N_18435);
nor U23021 (N_23021,N_17906,N_12708);
nor U23022 (N_23022,N_14762,N_16280);
nor U23023 (N_23023,N_18154,N_14440);
xor U23024 (N_23024,N_16947,N_13326);
xnor U23025 (N_23025,N_15940,N_17334);
xor U23026 (N_23026,N_17823,N_17301);
nor U23027 (N_23027,N_16345,N_18096);
nand U23028 (N_23028,N_18499,N_15568);
and U23029 (N_23029,N_13014,N_14318);
nor U23030 (N_23030,N_18490,N_15633);
and U23031 (N_23031,N_12664,N_18013);
nor U23032 (N_23032,N_14958,N_15347);
and U23033 (N_23033,N_17685,N_17012);
nor U23034 (N_23034,N_14486,N_17904);
nand U23035 (N_23035,N_13566,N_15177);
nor U23036 (N_23036,N_18073,N_12969);
and U23037 (N_23037,N_16179,N_15689);
xor U23038 (N_23038,N_15532,N_16593);
or U23039 (N_23039,N_16203,N_18245);
xnor U23040 (N_23040,N_13888,N_12988);
xor U23041 (N_23041,N_14663,N_17184);
nand U23042 (N_23042,N_12665,N_14126);
xnor U23043 (N_23043,N_12592,N_15242);
nor U23044 (N_23044,N_17413,N_16846);
xnor U23045 (N_23045,N_16244,N_12874);
or U23046 (N_23046,N_14828,N_18485);
or U23047 (N_23047,N_16491,N_17595);
nor U23048 (N_23048,N_16976,N_16809);
or U23049 (N_23049,N_14558,N_15725);
or U23050 (N_23050,N_15715,N_16297);
or U23051 (N_23051,N_18667,N_15111);
xor U23052 (N_23052,N_13435,N_17721);
nand U23053 (N_23053,N_17769,N_14702);
nand U23054 (N_23054,N_14764,N_14840);
nor U23055 (N_23055,N_14160,N_18377);
nand U23056 (N_23056,N_14828,N_16664);
nor U23057 (N_23057,N_13934,N_16707);
nor U23058 (N_23058,N_15907,N_15415);
and U23059 (N_23059,N_14373,N_14549);
or U23060 (N_23060,N_14979,N_17130);
or U23061 (N_23061,N_12701,N_14106);
nand U23062 (N_23062,N_17261,N_15585);
and U23063 (N_23063,N_16296,N_17460);
or U23064 (N_23064,N_14929,N_12610);
nor U23065 (N_23065,N_15953,N_14138);
xnor U23066 (N_23066,N_14040,N_13322);
nand U23067 (N_23067,N_14922,N_12696);
and U23068 (N_23068,N_18087,N_13961);
nand U23069 (N_23069,N_17451,N_12516);
nand U23070 (N_23070,N_16840,N_13659);
nor U23071 (N_23071,N_17048,N_17287);
xor U23072 (N_23072,N_15527,N_12610);
or U23073 (N_23073,N_17412,N_18388);
and U23074 (N_23074,N_17255,N_16332);
and U23075 (N_23075,N_17533,N_12569);
and U23076 (N_23076,N_13233,N_16515);
nor U23077 (N_23077,N_15364,N_13659);
xnor U23078 (N_23078,N_14465,N_18126);
xor U23079 (N_23079,N_16510,N_13782);
xnor U23080 (N_23080,N_13392,N_12762);
xor U23081 (N_23081,N_13423,N_18483);
or U23082 (N_23082,N_12740,N_18164);
xor U23083 (N_23083,N_16136,N_14000);
or U23084 (N_23084,N_14160,N_13996);
and U23085 (N_23085,N_17309,N_14845);
xor U23086 (N_23086,N_13099,N_18040);
nor U23087 (N_23087,N_17355,N_16425);
xor U23088 (N_23088,N_14127,N_17975);
xnor U23089 (N_23089,N_14251,N_13625);
nor U23090 (N_23090,N_17240,N_14054);
nor U23091 (N_23091,N_15796,N_13107);
xor U23092 (N_23092,N_17377,N_14783);
xor U23093 (N_23093,N_18661,N_17476);
xnor U23094 (N_23094,N_18395,N_13344);
and U23095 (N_23095,N_13326,N_15967);
and U23096 (N_23096,N_16750,N_17577);
or U23097 (N_23097,N_18331,N_14885);
xor U23098 (N_23098,N_15863,N_14906);
nor U23099 (N_23099,N_17560,N_14276);
and U23100 (N_23100,N_17641,N_17256);
xnor U23101 (N_23101,N_14425,N_15107);
nand U23102 (N_23102,N_13660,N_15106);
nand U23103 (N_23103,N_13786,N_17492);
and U23104 (N_23104,N_18480,N_16718);
xnor U23105 (N_23105,N_16385,N_15083);
nand U23106 (N_23106,N_15129,N_16724);
and U23107 (N_23107,N_15612,N_13255);
xor U23108 (N_23108,N_15525,N_15706);
xnor U23109 (N_23109,N_13887,N_13043);
xor U23110 (N_23110,N_15793,N_17481);
or U23111 (N_23111,N_17968,N_18199);
and U23112 (N_23112,N_18714,N_15417);
nand U23113 (N_23113,N_16248,N_15256);
or U23114 (N_23114,N_18084,N_13036);
xnor U23115 (N_23115,N_12711,N_13244);
nor U23116 (N_23116,N_13473,N_18411);
nor U23117 (N_23117,N_16670,N_16317);
or U23118 (N_23118,N_18037,N_15396);
xor U23119 (N_23119,N_15894,N_13056);
and U23120 (N_23120,N_15192,N_18000);
xor U23121 (N_23121,N_17655,N_16037);
and U23122 (N_23122,N_16263,N_17034);
nor U23123 (N_23123,N_16671,N_17497);
nand U23124 (N_23124,N_15853,N_12950);
nor U23125 (N_23125,N_16861,N_17170);
xor U23126 (N_23126,N_13784,N_16583);
and U23127 (N_23127,N_17754,N_17468);
and U23128 (N_23128,N_14349,N_14904);
nor U23129 (N_23129,N_13850,N_14117);
xor U23130 (N_23130,N_14258,N_13612);
nand U23131 (N_23131,N_12896,N_16129);
xnor U23132 (N_23132,N_15019,N_14545);
xor U23133 (N_23133,N_18442,N_15279);
nand U23134 (N_23134,N_12931,N_13624);
xnor U23135 (N_23135,N_14430,N_17107);
xor U23136 (N_23136,N_17623,N_14942);
nor U23137 (N_23137,N_13484,N_16250);
or U23138 (N_23138,N_15060,N_12639);
or U23139 (N_23139,N_12662,N_16320);
nand U23140 (N_23140,N_13173,N_14663);
or U23141 (N_23141,N_12676,N_16590);
and U23142 (N_23142,N_18457,N_13102);
nor U23143 (N_23143,N_13816,N_16729);
nor U23144 (N_23144,N_16988,N_15300);
nor U23145 (N_23145,N_13748,N_13317);
and U23146 (N_23146,N_13611,N_15264);
or U23147 (N_23147,N_13224,N_18321);
nand U23148 (N_23148,N_15419,N_18266);
or U23149 (N_23149,N_13579,N_18321);
or U23150 (N_23150,N_16953,N_12944);
and U23151 (N_23151,N_13369,N_16216);
xor U23152 (N_23152,N_17776,N_15928);
or U23153 (N_23153,N_14887,N_18056);
or U23154 (N_23154,N_16520,N_14299);
and U23155 (N_23155,N_16646,N_16309);
nor U23156 (N_23156,N_14949,N_17084);
xnor U23157 (N_23157,N_17829,N_17436);
and U23158 (N_23158,N_18710,N_17102);
or U23159 (N_23159,N_15852,N_18138);
or U23160 (N_23160,N_17243,N_14402);
nand U23161 (N_23161,N_16357,N_14211);
and U23162 (N_23162,N_15055,N_13987);
nand U23163 (N_23163,N_17402,N_17170);
nand U23164 (N_23164,N_13501,N_18177);
and U23165 (N_23165,N_17446,N_15777);
nor U23166 (N_23166,N_17845,N_14770);
xor U23167 (N_23167,N_12544,N_12944);
or U23168 (N_23168,N_16137,N_18513);
and U23169 (N_23169,N_14407,N_15610);
nand U23170 (N_23170,N_16181,N_16997);
nand U23171 (N_23171,N_12657,N_18118);
nor U23172 (N_23172,N_14298,N_16469);
nand U23173 (N_23173,N_12535,N_13407);
nor U23174 (N_23174,N_12818,N_17752);
nand U23175 (N_23175,N_16340,N_18055);
nand U23176 (N_23176,N_17855,N_18600);
or U23177 (N_23177,N_13331,N_15488);
or U23178 (N_23178,N_14407,N_13225);
nand U23179 (N_23179,N_12689,N_16017);
or U23180 (N_23180,N_17374,N_14599);
nand U23181 (N_23181,N_16549,N_15252);
or U23182 (N_23182,N_16697,N_13892);
nor U23183 (N_23183,N_18254,N_14087);
or U23184 (N_23184,N_17843,N_15389);
nand U23185 (N_23185,N_16019,N_14723);
and U23186 (N_23186,N_16971,N_13228);
xnor U23187 (N_23187,N_15273,N_14083);
xor U23188 (N_23188,N_15694,N_16908);
or U23189 (N_23189,N_17898,N_16404);
or U23190 (N_23190,N_15593,N_16578);
xnor U23191 (N_23191,N_18489,N_14578);
nand U23192 (N_23192,N_14403,N_12819);
nand U23193 (N_23193,N_18062,N_12582);
and U23194 (N_23194,N_18084,N_17081);
or U23195 (N_23195,N_13321,N_14244);
xor U23196 (N_23196,N_15422,N_15888);
and U23197 (N_23197,N_14504,N_18301);
or U23198 (N_23198,N_16212,N_18442);
and U23199 (N_23199,N_16400,N_17393);
nand U23200 (N_23200,N_15503,N_17889);
nor U23201 (N_23201,N_14475,N_14381);
or U23202 (N_23202,N_15363,N_15292);
xor U23203 (N_23203,N_14672,N_13068);
nand U23204 (N_23204,N_13510,N_13427);
and U23205 (N_23205,N_12589,N_17008);
or U23206 (N_23206,N_16832,N_16854);
nor U23207 (N_23207,N_15041,N_12574);
or U23208 (N_23208,N_14615,N_15219);
xor U23209 (N_23209,N_16653,N_13787);
xor U23210 (N_23210,N_12504,N_16324);
nand U23211 (N_23211,N_14107,N_18296);
nor U23212 (N_23212,N_16083,N_15945);
nor U23213 (N_23213,N_18702,N_18442);
nand U23214 (N_23214,N_17457,N_13396);
nand U23215 (N_23215,N_12726,N_15425);
xor U23216 (N_23216,N_13898,N_15718);
xnor U23217 (N_23217,N_16595,N_18621);
and U23218 (N_23218,N_17300,N_15358);
and U23219 (N_23219,N_17647,N_17209);
nand U23220 (N_23220,N_15853,N_16861);
nor U23221 (N_23221,N_17249,N_13692);
nor U23222 (N_23222,N_18522,N_13006);
and U23223 (N_23223,N_17494,N_15132);
and U23224 (N_23224,N_16882,N_15230);
and U23225 (N_23225,N_18590,N_17313);
and U23226 (N_23226,N_18261,N_13442);
nand U23227 (N_23227,N_17336,N_12785);
nand U23228 (N_23228,N_14357,N_13388);
xnor U23229 (N_23229,N_12905,N_16317);
and U23230 (N_23230,N_18543,N_14026);
or U23231 (N_23231,N_14736,N_17847);
and U23232 (N_23232,N_18113,N_13099);
or U23233 (N_23233,N_12576,N_16252);
or U23234 (N_23234,N_16120,N_17557);
nor U23235 (N_23235,N_14197,N_13238);
and U23236 (N_23236,N_14508,N_15971);
or U23237 (N_23237,N_17506,N_12843);
xnor U23238 (N_23238,N_13062,N_14747);
nand U23239 (N_23239,N_17818,N_14732);
nor U23240 (N_23240,N_14754,N_16864);
nand U23241 (N_23241,N_12602,N_15173);
and U23242 (N_23242,N_17621,N_15875);
xor U23243 (N_23243,N_17795,N_14437);
and U23244 (N_23244,N_17952,N_13087);
and U23245 (N_23245,N_13589,N_17937);
and U23246 (N_23246,N_13174,N_12785);
and U23247 (N_23247,N_15513,N_15589);
xor U23248 (N_23248,N_17903,N_18701);
nand U23249 (N_23249,N_17198,N_16378);
or U23250 (N_23250,N_17472,N_17140);
or U23251 (N_23251,N_14469,N_14159);
or U23252 (N_23252,N_13982,N_15770);
xnor U23253 (N_23253,N_18079,N_12975);
and U23254 (N_23254,N_14475,N_14533);
or U23255 (N_23255,N_16438,N_13381);
nor U23256 (N_23256,N_12586,N_16325);
or U23257 (N_23257,N_13998,N_13809);
nor U23258 (N_23258,N_13674,N_14319);
nand U23259 (N_23259,N_14780,N_13292);
and U23260 (N_23260,N_16354,N_12681);
xor U23261 (N_23261,N_18385,N_17454);
and U23262 (N_23262,N_15907,N_18587);
xnor U23263 (N_23263,N_16814,N_18121);
or U23264 (N_23264,N_14579,N_13040);
and U23265 (N_23265,N_13757,N_17844);
nand U23266 (N_23266,N_13347,N_15137);
or U23267 (N_23267,N_17248,N_14830);
nor U23268 (N_23268,N_17243,N_18634);
or U23269 (N_23269,N_14119,N_17070);
or U23270 (N_23270,N_15689,N_18262);
or U23271 (N_23271,N_14014,N_12655);
nor U23272 (N_23272,N_16280,N_18573);
nand U23273 (N_23273,N_14159,N_15054);
and U23274 (N_23274,N_15947,N_13673);
nor U23275 (N_23275,N_14961,N_17354);
nor U23276 (N_23276,N_17859,N_14904);
nor U23277 (N_23277,N_15099,N_12619);
nand U23278 (N_23278,N_16382,N_18648);
or U23279 (N_23279,N_17201,N_13574);
and U23280 (N_23280,N_12901,N_17147);
nand U23281 (N_23281,N_16304,N_18525);
xor U23282 (N_23282,N_17310,N_15006);
or U23283 (N_23283,N_14689,N_15295);
nand U23284 (N_23284,N_12818,N_13525);
and U23285 (N_23285,N_15188,N_16995);
nor U23286 (N_23286,N_14054,N_16433);
and U23287 (N_23287,N_12712,N_16671);
xor U23288 (N_23288,N_13567,N_13346);
xnor U23289 (N_23289,N_13666,N_17877);
or U23290 (N_23290,N_13139,N_14534);
nand U23291 (N_23291,N_13491,N_17030);
and U23292 (N_23292,N_18064,N_14680);
nor U23293 (N_23293,N_17947,N_18166);
nand U23294 (N_23294,N_16305,N_18136);
and U23295 (N_23295,N_13489,N_14139);
xor U23296 (N_23296,N_15227,N_16608);
xnor U23297 (N_23297,N_15538,N_15506);
nand U23298 (N_23298,N_14058,N_15975);
and U23299 (N_23299,N_16198,N_17412);
and U23300 (N_23300,N_12723,N_15215);
nand U23301 (N_23301,N_14809,N_13129);
and U23302 (N_23302,N_13744,N_14002);
nor U23303 (N_23303,N_14612,N_16861);
nor U23304 (N_23304,N_17549,N_18483);
or U23305 (N_23305,N_16503,N_17806);
xor U23306 (N_23306,N_17348,N_17086);
nand U23307 (N_23307,N_14069,N_16715);
xor U23308 (N_23308,N_13041,N_15653);
nand U23309 (N_23309,N_16141,N_15423);
and U23310 (N_23310,N_15812,N_12545);
xor U23311 (N_23311,N_14636,N_13323);
nor U23312 (N_23312,N_18196,N_18170);
or U23313 (N_23313,N_13331,N_13955);
xor U23314 (N_23314,N_12639,N_15251);
or U23315 (N_23315,N_12845,N_16279);
nor U23316 (N_23316,N_17270,N_14782);
nand U23317 (N_23317,N_18481,N_16102);
or U23318 (N_23318,N_17744,N_13264);
nand U23319 (N_23319,N_13037,N_13732);
or U23320 (N_23320,N_13259,N_15000);
nand U23321 (N_23321,N_16227,N_13289);
or U23322 (N_23322,N_13255,N_17409);
or U23323 (N_23323,N_13328,N_14861);
nand U23324 (N_23324,N_13682,N_18105);
or U23325 (N_23325,N_14460,N_16653);
and U23326 (N_23326,N_14116,N_17915);
nor U23327 (N_23327,N_15806,N_13526);
nor U23328 (N_23328,N_12505,N_17389);
or U23329 (N_23329,N_16797,N_15607);
nand U23330 (N_23330,N_14944,N_16610);
nand U23331 (N_23331,N_13497,N_16582);
nor U23332 (N_23332,N_15265,N_16471);
or U23333 (N_23333,N_13887,N_13422);
xor U23334 (N_23334,N_15799,N_14344);
or U23335 (N_23335,N_14291,N_15806);
and U23336 (N_23336,N_12527,N_16347);
and U23337 (N_23337,N_16362,N_14977);
xor U23338 (N_23338,N_14231,N_17415);
nand U23339 (N_23339,N_18535,N_17546);
and U23340 (N_23340,N_18371,N_18413);
xor U23341 (N_23341,N_17058,N_13199);
nand U23342 (N_23342,N_14287,N_13169);
nand U23343 (N_23343,N_18716,N_17382);
xnor U23344 (N_23344,N_14862,N_15290);
nor U23345 (N_23345,N_13809,N_15671);
nand U23346 (N_23346,N_13636,N_16657);
or U23347 (N_23347,N_15279,N_18041);
and U23348 (N_23348,N_15518,N_12865);
nand U23349 (N_23349,N_18676,N_14485);
or U23350 (N_23350,N_17847,N_15259);
and U23351 (N_23351,N_16386,N_17363);
or U23352 (N_23352,N_13121,N_18073);
and U23353 (N_23353,N_16656,N_14251);
nand U23354 (N_23354,N_16565,N_18207);
xor U23355 (N_23355,N_18561,N_16784);
xnor U23356 (N_23356,N_15393,N_12744);
xnor U23357 (N_23357,N_13440,N_13136);
xor U23358 (N_23358,N_12540,N_14798);
nor U23359 (N_23359,N_15051,N_18614);
and U23360 (N_23360,N_13517,N_17477);
nand U23361 (N_23361,N_14583,N_18352);
xor U23362 (N_23362,N_16305,N_18427);
and U23363 (N_23363,N_16963,N_18220);
nand U23364 (N_23364,N_15735,N_13115);
or U23365 (N_23365,N_13345,N_13551);
xor U23366 (N_23366,N_17523,N_15450);
nor U23367 (N_23367,N_16286,N_13807);
or U23368 (N_23368,N_16401,N_16330);
nand U23369 (N_23369,N_18184,N_18269);
nand U23370 (N_23370,N_17420,N_12689);
and U23371 (N_23371,N_16148,N_12828);
or U23372 (N_23372,N_15508,N_13122);
xnor U23373 (N_23373,N_15753,N_13629);
nand U23374 (N_23374,N_15101,N_14905);
or U23375 (N_23375,N_17632,N_17449);
nand U23376 (N_23376,N_12589,N_18117);
nor U23377 (N_23377,N_14448,N_13691);
xor U23378 (N_23378,N_17096,N_15674);
or U23379 (N_23379,N_16964,N_14723);
and U23380 (N_23380,N_15865,N_15876);
nand U23381 (N_23381,N_15699,N_17094);
or U23382 (N_23382,N_14081,N_14091);
xnor U23383 (N_23383,N_16434,N_17093);
or U23384 (N_23384,N_13870,N_14001);
xor U23385 (N_23385,N_17814,N_17676);
nand U23386 (N_23386,N_12730,N_17923);
or U23387 (N_23387,N_15872,N_17135);
or U23388 (N_23388,N_13202,N_16895);
nand U23389 (N_23389,N_15062,N_12777);
nand U23390 (N_23390,N_18459,N_18422);
and U23391 (N_23391,N_14005,N_13794);
and U23392 (N_23392,N_17276,N_18614);
nor U23393 (N_23393,N_12976,N_16558);
or U23394 (N_23394,N_13879,N_13694);
xnor U23395 (N_23395,N_15174,N_14131);
nand U23396 (N_23396,N_12714,N_14975);
nand U23397 (N_23397,N_18179,N_14765);
and U23398 (N_23398,N_13625,N_18218);
and U23399 (N_23399,N_18048,N_17901);
nand U23400 (N_23400,N_15584,N_13203);
and U23401 (N_23401,N_15239,N_12878);
nand U23402 (N_23402,N_14316,N_17896);
and U23403 (N_23403,N_17875,N_13652);
xnor U23404 (N_23404,N_15001,N_18453);
xor U23405 (N_23405,N_18202,N_18634);
or U23406 (N_23406,N_13074,N_16213);
nand U23407 (N_23407,N_15363,N_16110);
nand U23408 (N_23408,N_18510,N_17645);
xor U23409 (N_23409,N_14901,N_16971);
nand U23410 (N_23410,N_13306,N_17809);
xnor U23411 (N_23411,N_18692,N_17556);
nor U23412 (N_23412,N_17958,N_16647);
and U23413 (N_23413,N_17795,N_15462);
xnor U23414 (N_23414,N_14156,N_13017);
nand U23415 (N_23415,N_18280,N_18257);
xnor U23416 (N_23416,N_12534,N_14207);
nand U23417 (N_23417,N_18139,N_18680);
nor U23418 (N_23418,N_16726,N_18516);
or U23419 (N_23419,N_13869,N_16419);
nand U23420 (N_23420,N_13133,N_12898);
and U23421 (N_23421,N_17524,N_14797);
nor U23422 (N_23422,N_16938,N_13690);
and U23423 (N_23423,N_17883,N_16028);
and U23424 (N_23424,N_12665,N_17513);
nor U23425 (N_23425,N_18343,N_14423);
xor U23426 (N_23426,N_15675,N_12518);
and U23427 (N_23427,N_12559,N_13570);
and U23428 (N_23428,N_16480,N_17058);
or U23429 (N_23429,N_15211,N_14580);
xor U23430 (N_23430,N_15816,N_17929);
nor U23431 (N_23431,N_13955,N_13608);
nor U23432 (N_23432,N_16745,N_12835);
or U23433 (N_23433,N_13995,N_15517);
or U23434 (N_23434,N_18677,N_16629);
xor U23435 (N_23435,N_14888,N_13712);
or U23436 (N_23436,N_16344,N_16083);
nand U23437 (N_23437,N_15788,N_14055);
and U23438 (N_23438,N_18466,N_14105);
or U23439 (N_23439,N_16698,N_12884);
nand U23440 (N_23440,N_18069,N_16795);
xnor U23441 (N_23441,N_17733,N_13214);
nand U23442 (N_23442,N_15992,N_18454);
nand U23443 (N_23443,N_18407,N_13894);
or U23444 (N_23444,N_13074,N_16842);
and U23445 (N_23445,N_16368,N_16482);
xor U23446 (N_23446,N_13149,N_13640);
or U23447 (N_23447,N_14811,N_13659);
and U23448 (N_23448,N_18076,N_15101);
nand U23449 (N_23449,N_13662,N_16246);
nand U23450 (N_23450,N_13373,N_13348);
and U23451 (N_23451,N_17057,N_15262);
or U23452 (N_23452,N_13124,N_15475);
nand U23453 (N_23453,N_18385,N_13787);
or U23454 (N_23454,N_15652,N_17892);
nor U23455 (N_23455,N_12683,N_18123);
xor U23456 (N_23456,N_15582,N_12721);
nand U23457 (N_23457,N_18245,N_12992);
xnor U23458 (N_23458,N_18171,N_13118);
and U23459 (N_23459,N_13914,N_13152);
or U23460 (N_23460,N_17021,N_17319);
and U23461 (N_23461,N_15565,N_16680);
or U23462 (N_23462,N_17485,N_13289);
nor U23463 (N_23463,N_16784,N_13626);
nor U23464 (N_23464,N_17056,N_16971);
xor U23465 (N_23465,N_14100,N_15455);
or U23466 (N_23466,N_16940,N_17153);
xnor U23467 (N_23467,N_13540,N_14167);
nor U23468 (N_23468,N_13091,N_17373);
or U23469 (N_23469,N_13122,N_18501);
xnor U23470 (N_23470,N_16184,N_18645);
nand U23471 (N_23471,N_17859,N_14269);
and U23472 (N_23472,N_16758,N_13864);
and U23473 (N_23473,N_13872,N_17158);
xnor U23474 (N_23474,N_15878,N_15715);
xor U23475 (N_23475,N_14617,N_16523);
and U23476 (N_23476,N_12932,N_14030);
nor U23477 (N_23477,N_12616,N_17322);
and U23478 (N_23478,N_17062,N_17926);
nand U23479 (N_23479,N_15563,N_18483);
nand U23480 (N_23480,N_13601,N_17416);
xor U23481 (N_23481,N_13195,N_15616);
and U23482 (N_23482,N_14764,N_14800);
nand U23483 (N_23483,N_15202,N_16404);
nor U23484 (N_23484,N_12951,N_14713);
xnor U23485 (N_23485,N_13851,N_17762);
nand U23486 (N_23486,N_16600,N_18650);
or U23487 (N_23487,N_15193,N_18683);
xor U23488 (N_23488,N_18117,N_15335);
and U23489 (N_23489,N_14445,N_16338);
and U23490 (N_23490,N_14054,N_12634);
or U23491 (N_23491,N_13748,N_17539);
xor U23492 (N_23492,N_17811,N_13447);
xor U23493 (N_23493,N_15367,N_15051);
or U23494 (N_23494,N_14573,N_12578);
xor U23495 (N_23495,N_17133,N_17937);
or U23496 (N_23496,N_12505,N_13591);
xor U23497 (N_23497,N_16623,N_18159);
and U23498 (N_23498,N_17646,N_13694);
and U23499 (N_23499,N_17876,N_15645);
or U23500 (N_23500,N_16971,N_14494);
and U23501 (N_23501,N_12881,N_15559);
nor U23502 (N_23502,N_13507,N_14652);
nand U23503 (N_23503,N_13838,N_16668);
nand U23504 (N_23504,N_16404,N_16153);
xor U23505 (N_23505,N_17104,N_18168);
xor U23506 (N_23506,N_15467,N_13442);
and U23507 (N_23507,N_16263,N_17938);
nor U23508 (N_23508,N_17867,N_12857);
nand U23509 (N_23509,N_15392,N_17599);
xor U23510 (N_23510,N_16197,N_15682);
nor U23511 (N_23511,N_13728,N_15743);
and U23512 (N_23512,N_16565,N_13383);
nor U23513 (N_23513,N_16253,N_17219);
nor U23514 (N_23514,N_12593,N_14750);
and U23515 (N_23515,N_18574,N_15147);
xnor U23516 (N_23516,N_15781,N_15003);
nor U23517 (N_23517,N_14537,N_14063);
nand U23518 (N_23518,N_13591,N_15008);
or U23519 (N_23519,N_14359,N_13539);
nand U23520 (N_23520,N_18083,N_18225);
xor U23521 (N_23521,N_17908,N_17457);
nor U23522 (N_23522,N_14115,N_14842);
nand U23523 (N_23523,N_14279,N_15713);
xor U23524 (N_23524,N_13955,N_16913);
nand U23525 (N_23525,N_13901,N_17191);
nand U23526 (N_23526,N_18451,N_15115);
xnor U23527 (N_23527,N_14510,N_15148);
nand U23528 (N_23528,N_14377,N_14066);
or U23529 (N_23529,N_17089,N_16084);
and U23530 (N_23530,N_12584,N_18726);
nor U23531 (N_23531,N_18554,N_12968);
nand U23532 (N_23532,N_14910,N_18348);
or U23533 (N_23533,N_17890,N_15924);
nand U23534 (N_23534,N_17902,N_14442);
xor U23535 (N_23535,N_15942,N_18671);
and U23536 (N_23536,N_15679,N_14501);
or U23537 (N_23537,N_15693,N_14759);
or U23538 (N_23538,N_15327,N_13949);
nor U23539 (N_23539,N_14694,N_13304);
nor U23540 (N_23540,N_14212,N_18500);
and U23541 (N_23541,N_16421,N_14267);
or U23542 (N_23542,N_15616,N_17253);
nor U23543 (N_23543,N_16185,N_17440);
and U23544 (N_23544,N_14047,N_14521);
nand U23545 (N_23545,N_16075,N_13193);
and U23546 (N_23546,N_17126,N_12772);
nor U23547 (N_23547,N_13225,N_16645);
xnor U23548 (N_23548,N_15348,N_13189);
and U23549 (N_23549,N_16264,N_14899);
xor U23550 (N_23550,N_13864,N_16498);
nor U23551 (N_23551,N_16247,N_17400);
or U23552 (N_23552,N_13511,N_15405);
nand U23553 (N_23553,N_15126,N_13425);
and U23554 (N_23554,N_15191,N_12702);
and U23555 (N_23555,N_15928,N_17666);
xnor U23556 (N_23556,N_18061,N_13964);
or U23557 (N_23557,N_16998,N_15123);
nor U23558 (N_23558,N_18364,N_15475);
or U23559 (N_23559,N_13589,N_18551);
and U23560 (N_23560,N_13469,N_12704);
xor U23561 (N_23561,N_15608,N_16178);
nor U23562 (N_23562,N_17351,N_17010);
and U23563 (N_23563,N_17734,N_14986);
or U23564 (N_23564,N_13468,N_15102);
or U23565 (N_23565,N_17889,N_17285);
xnor U23566 (N_23566,N_18525,N_13706);
nor U23567 (N_23567,N_12834,N_17804);
or U23568 (N_23568,N_14462,N_15026);
nor U23569 (N_23569,N_13167,N_15134);
or U23570 (N_23570,N_18414,N_12980);
nand U23571 (N_23571,N_14850,N_15252);
nand U23572 (N_23572,N_15229,N_14948);
xnor U23573 (N_23573,N_18563,N_14330);
and U23574 (N_23574,N_14811,N_16890);
nand U23575 (N_23575,N_12977,N_12961);
nor U23576 (N_23576,N_16731,N_16665);
nand U23577 (N_23577,N_17684,N_15803);
or U23578 (N_23578,N_12596,N_15996);
or U23579 (N_23579,N_18116,N_14090);
and U23580 (N_23580,N_13716,N_12875);
nor U23581 (N_23581,N_16446,N_14640);
or U23582 (N_23582,N_13610,N_15473);
xor U23583 (N_23583,N_16969,N_13436);
nand U23584 (N_23584,N_12685,N_16830);
nor U23585 (N_23585,N_16642,N_14462);
or U23586 (N_23586,N_14503,N_13638);
or U23587 (N_23587,N_13753,N_16084);
xnor U23588 (N_23588,N_18255,N_15290);
or U23589 (N_23589,N_15523,N_16573);
nand U23590 (N_23590,N_12773,N_16891);
xor U23591 (N_23591,N_16905,N_18590);
and U23592 (N_23592,N_18315,N_18397);
nor U23593 (N_23593,N_15781,N_18508);
or U23594 (N_23594,N_16711,N_17292);
nor U23595 (N_23595,N_15324,N_18746);
nand U23596 (N_23596,N_15691,N_12859);
or U23597 (N_23597,N_17752,N_17623);
nand U23598 (N_23598,N_18333,N_13818);
or U23599 (N_23599,N_15912,N_18537);
xnor U23600 (N_23600,N_15850,N_15306);
xor U23601 (N_23601,N_13565,N_17683);
nor U23602 (N_23602,N_16325,N_14775);
nand U23603 (N_23603,N_16055,N_17500);
nand U23604 (N_23604,N_13939,N_13303);
nor U23605 (N_23605,N_14635,N_18653);
nand U23606 (N_23606,N_16832,N_13308);
nand U23607 (N_23607,N_13831,N_16501);
nand U23608 (N_23608,N_13477,N_17131);
or U23609 (N_23609,N_14791,N_12633);
nand U23610 (N_23610,N_16375,N_14977);
nor U23611 (N_23611,N_14376,N_18627);
xor U23612 (N_23612,N_14041,N_15439);
and U23613 (N_23613,N_12521,N_16919);
or U23614 (N_23614,N_17090,N_16763);
or U23615 (N_23615,N_16212,N_15920);
nor U23616 (N_23616,N_17727,N_14528);
xnor U23617 (N_23617,N_15170,N_12628);
and U23618 (N_23618,N_18749,N_14634);
nor U23619 (N_23619,N_14085,N_15171);
xor U23620 (N_23620,N_15536,N_14748);
nand U23621 (N_23621,N_12708,N_16560);
nor U23622 (N_23622,N_14914,N_12846);
nand U23623 (N_23623,N_15683,N_16861);
nand U23624 (N_23624,N_17703,N_16643);
or U23625 (N_23625,N_13593,N_16046);
or U23626 (N_23626,N_18528,N_15386);
xnor U23627 (N_23627,N_16521,N_12673);
or U23628 (N_23628,N_12887,N_12801);
or U23629 (N_23629,N_14931,N_13838);
nor U23630 (N_23630,N_17920,N_18193);
and U23631 (N_23631,N_14043,N_18536);
nand U23632 (N_23632,N_16442,N_13660);
xor U23633 (N_23633,N_15943,N_13407);
and U23634 (N_23634,N_13821,N_15952);
nor U23635 (N_23635,N_18454,N_16721);
nor U23636 (N_23636,N_17512,N_13875);
nand U23637 (N_23637,N_13170,N_14641);
nand U23638 (N_23638,N_18071,N_15335);
or U23639 (N_23639,N_14489,N_13775);
and U23640 (N_23640,N_13885,N_15818);
or U23641 (N_23641,N_16078,N_14315);
xnor U23642 (N_23642,N_16789,N_15393);
or U23643 (N_23643,N_15215,N_12946);
nand U23644 (N_23644,N_18314,N_13659);
and U23645 (N_23645,N_12668,N_15549);
nand U23646 (N_23646,N_17680,N_14501);
or U23647 (N_23647,N_17466,N_14413);
or U23648 (N_23648,N_17004,N_18416);
nand U23649 (N_23649,N_16751,N_12757);
and U23650 (N_23650,N_15998,N_13862);
or U23651 (N_23651,N_12845,N_12815);
or U23652 (N_23652,N_16372,N_13140);
xor U23653 (N_23653,N_14930,N_16226);
nand U23654 (N_23654,N_13674,N_13855);
xnor U23655 (N_23655,N_16750,N_12973);
xor U23656 (N_23656,N_16949,N_15257);
nand U23657 (N_23657,N_15698,N_15650);
nor U23658 (N_23658,N_17494,N_17013);
and U23659 (N_23659,N_15675,N_14341);
nor U23660 (N_23660,N_15119,N_17883);
and U23661 (N_23661,N_17001,N_16770);
xor U23662 (N_23662,N_17622,N_16725);
nor U23663 (N_23663,N_14489,N_15792);
or U23664 (N_23664,N_15539,N_18006);
and U23665 (N_23665,N_17533,N_16179);
nor U23666 (N_23666,N_12787,N_16438);
and U23667 (N_23667,N_16026,N_13317);
nor U23668 (N_23668,N_13628,N_16557);
nor U23669 (N_23669,N_18196,N_14624);
xor U23670 (N_23670,N_17426,N_18646);
nor U23671 (N_23671,N_13141,N_16373);
and U23672 (N_23672,N_15712,N_16293);
nand U23673 (N_23673,N_13743,N_15288);
nor U23674 (N_23674,N_13867,N_13790);
xnor U23675 (N_23675,N_15772,N_13868);
or U23676 (N_23676,N_12873,N_18030);
or U23677 (N_23677,N_15973,N_13340);
or U23678 (N_23678,N_12538,N_15660);
nor U23679 (N_23679,N_17224,N_18056);
or U23680 (N_23680,N_17878,N_16509);
nand U23681 (N_23681,N_18428,N_14262);
and U23682 (N_23682,N_15847,N_14153);
xor U23683 (N_23683,N_18184,N_14312);
nor U23684 (N_23684,N_17122,N_18403);
xnor U23685 (N_23685,N_15054,N_13277);
and U23686 (N_23686,N_16520,N_13454);
or U23687 (N_23687,N_16507,N_15392);
xnor U23688 (N_23688,N_18719,N_13791);
and U23689 (N_23689,N_18632,N_13201);
nand U23690 (N_23690,N_17211,N_16859);
nand U23691 (N_23691,N_13228,N_15116);
nor U23692 (N_23692,N_12515,N_17381);
nand U23693 (N_23693,N_12662,N_13626);
xnor U23694 (N_23694,N_17050,N_16130);
nor U23695 (N_23695,N_16156,N_16324);
nor U23696 (N_23696,N_12927,N_17595);
nand U23697 (N_23697,N_16447,N_15884);
nor U23698 (N_23698,N_16850,N_18277);
nand U23699 (N_23699,N_13198,N_16698);
or U23700 (N_23700,N_18122,N_18496);
or U23701 (N_23701,N_16955,N_13695);
nand U23702 (N_23702,N_16002,N_13779);
or U23703 (N_23703,N_18118,N_17420);
xor U23704 (N_23704,N_13981,N_14592);
xnor U23705 (N_23705,N_12941,N_17751);
nor U23706 (N_23706,N_16488,N_18440);
or U23707 (N_23707,N_15825,N_16309);
nor U23708 (N_23708,N_17240,N_14735);
nand U23709 (N_23709,N_17837,N_16352);
nor U23710 (N_23710,N_15061,N_14519);
nor U23711 (N_23711,N_13160,N_16532);
nand U23712 (N_23712,N_17009,N_14419);
or U23713 (N_23713,N_16001,N_14610);
nor U23714 (N_23714,N_14221,N_18054);
nand U23715 (N_23715,N_18426,N_16338);
and U23716 (N_23716,N_14764,N_14167);
or U23717 (N_23717,N_17488,N_16109);
nor U23718 (N_23718,N_15744,N_17006);
nor U23719 (N_23719,N_15599,N_14726);
or U23720 (N_23720,N_13756,N_14372);
nand U23721 (N_23721,N_16119,N_16997);
xnor U23722 (N_23722,N_16383,N_17385);
and U23723 (N_23723,N_17073,N_12647);
and U23724 (N_23724,N_17802,N_14920);
nor U23725 (N_23725,N_17888,N_17876);
or U23726 (N_23726,N_14006,N_16341);
xor U23727 (N_23727,N_15417,N_16162);
nor U23728 (N_23728,N_12913,N_14168);
xnor U23729 (N_23729,N_14423,N_13265);
or U23730 (N_23730,N_15024,N_14258);
and U23731 (N_23731,N_17574,N_18596);
nor U23732 (N_23732,N_14083,N_15893);
nand U23733 (N_23733,N_12737,N_17566);
xor U23734 (N_23734,N_18734,N_13814);
or U23735 (N_23735,N_18612,N_14383);
and U23736 (N_23736,N_12788,N_13878);
or U23737 (N_23737,N_15933,N_13926);
xnor U23738 (N_23738,N_17161,N_16737);
or U23739 (N_23739,N_16239,N_17935);
nor U23740 (N_23740,N_16642,N_13260);
xor U23741 (N_23741,N_16814,N_12702);
xnor U23742 (N_23742,N_16167,N_16506);
nand U23743 (N_23743,N_16726,N_18035);
nand U23744 (N_23744,N_17506,N_18189);
and U23745 (N_23745,N_17146,N_14278);
nand U23746 (N_23746,N_13325,N_14915);
or U23747 (N_23747,N_15784,N_15151);
or U23748 (N_23748,N_14222,N_15994);
and U23749 (N_23749,N_12972,N_16834);
and U23750 (N_23750,N_13856,N_15494);
nor U23751 (N_23751,N_14209,N_16177);
nor U23752 (N_23752,N_17350,N_17195);
nand U23753 (N_23753,N_16591,N_15919);
nor U23754 (N_23754,N_15681,N_14697);
nor U23755 (N_23755,N_12521,N_13544);
nor U23756 (N_23756,N_18643,N_16126);
nor U23757 (N_23757,N_12980,N_16026);
and U23758 (N_23758,N_13733,N_16581);
nor U23759 (N_23759,N_14265,N_15243);
or U23760 (N_23760,N_13904,N_14497);
nand U23761 (N_23761,N_17695,N_14120);
xnor U23762 (N_23762,N_14255,N_13986);
xor U23763 (N_23763,N_16525,N_14182);
xnor U23764 (N_23764,N_15675,N_18264);
xor U23765 (N_23765,N_16301,N_15103);
xor U23766 (N_23766,N_14777,N_14310);
and U23767 (N_23767,N_15964,N_16548);
nor U23768 (N_23768,N_18309,N_17053);
xnor U23769 (N_23769,N_16529,N_13242);
nand U23770 (N_23770,N_16961,N_14124);
nand U23771 (N_23771,N_16943,N_18711);
xor U23772 (N_23772,N_18021,N_14020);
xor U23773 (N_23773,N_14069,N_17680);
and U23774 (N_23774,N_16882,N_16230);
xnor U23775 (N_23775,N_17650,N_13077);
nand U23776 (N_23776,N_18465,N_15468);
and U23777 (N_23777,N_15696,N_13015);
nor U23778 (N_23778,N_14270,N_13169);
xnor U23779 (N_23779,N_18250,N_14183);
or U23780 (N_23780,N_15414,N_15691);
nand U23781 (N_23781,N_14858,N_13309);
and U23782 (N_23782,N_18618,N_18621);
or U23783 (N_23783,N_12673,N_12589);
nor U23784 (N_23784,N_12770,N_13965);
and U23785 (N_23785,N_16610,N_14734);
nor U23786 (N_23786,N_18020,N_16437);
nand U23787 (N_23787,N_18433,N_14946);
xnor U23788 (N_23788,N_13171,N_15762);
nand U23789 (N_23789,N_15300,N_17143);
nand U23790 (N_23790,N_15824,N_16777);
or U23791 (N_23791,N_14428,N_16602);
xnor U23792 (N_23792,N_13250,N_15308);
nand U23793 (N_23793,N_14226,N_15342);
and U23794 (N_23794,N_15355,N_17330);
or U23795 (N_23795,N_16789,N_13240);
or U23796 (N_23796,N_15598,N_17357);
or U23797 (N_23797,N_13314,N_18064);
nand U23798 (N_23798,N_16708,N_13797);
nor U23799 (N_23799,N_15248,N_15805);
xnor U23800 (N_23800,N_15109,N_17170);
nor U23801 (N_23801,N_16397,N_18724);
nor U23802 (N_23802,N_13902,N_16508);
nor U23803 (N_23803,N_15281,N_12692);
nand U23804 (N_23804,N_17378,N_16807);
xnor U23805 (N_23805,N_12538,N_17845);
nor U23806 (N_23806,N_16318,N_14724);
xor U23807 (N_23807,N_13459,N_12574);
nor U23808 (N_23808,N_13997,N_16867);
nand U23809 (N_23809,N_12552,N_17578);
xor U23810 (N_23810,N_18350,N_13500);
or U23811 (N_23811,N_13608,N_14493);
nor U23812 (N_23812,N_17609,N_15370);
and U23813 (N_23813,N_12825,N_15111);
nand U23814 (N_23814,N_14137,N_13195);
nand U23815 (N_23815,N_18367,N_17184);
or U23816 (N_23816,N_14655,N_15090);
nor U23817 (N_23817,N_15950,N_13863);
xnor U23818 (N_23818,N_17181,N_13029);
nand U23819 (N_23819,N_13552,N_18303);
xor U23820 (N_23820,N_17813,N_14951);
xor U23821 (N_23821,N_16361,N_15903);
or U23822 (N_23822,N_12850,N_15126);
xnor U23823 (N_23823,N_17415,N_12608);
nor U23824 (N_23824,N_18044,N_17723);
and U23825 (N_23825,N_18018,N_15980);
xor U23826 (N_23826,N_18183,N_12757);
xnor U23827 (N_23827,N_12724,N_16461);
nand U23828 (N_23828,N_15488,N_15074);
xnor U23829 (N_23829,N_15389,N_17379);
nand U23830 (N_23830,N_14601,N_14408);
xor U23831 (N_23831,N_13529,N_18473);
nor U23832 (N_23832,N_13485,N_15081);
xnor U23833 (N_23833,N_18611,N_13894);
or U23834 (N_23834,N_15242,N_18499);
xor U23835 (N_23835,N_14020,N_15897);
xnor U23836 (N_23836,N_18175,N_18141);
nand U23837 (N_23837,N_17323,N_15866);
and U23838 (N_23838,N_14556,N_17442);
nand U23839 (N_23839,N_17140,N_17874);
nand U23840 (N_23840,N_18703,N_14230);
and U23841 (N_23841,N_13732,N_14307);
nand U23842 (N_23842,N_16336,N_15179);
or U23843 (N_23843,N_15004,N_18482);
or U23844 (N_23844,N_17376,N_17149);
or U23845 (N_23845,N_15495,N_17142);
nand U23846 (N_23846,N_12571,N_16261);
xor U23847 (N_23847,N_18304,N_16883);
nor U23848 (N_23848,N_17892,N_13370);
nor U23849 (N_23849,N_13404,N_13527);
or U23850 (N_23850,N_15991,N_12903);
and U23851 (N_23851,N_13162,N_17701);
nor U23852 (N_23852,N_15126,N_14956);
nor U23853 (N_23853,N_16095,N_16069);
nand U23854 (N_23854,N_16060,N_18276);
or U23855 (N_23855,N_16109,N_13333);
nor U23856 (N_23856,N_14176,N_12880);
or U23857 (N_23857,N_17503,N_16699);
and U23858 (N_23858,N_12794,N_12762);
and U23859 (N_23859,N_16880,N_16419);
or U23860 (N_23860,N_14600,N_18044);
xnor U23861 (N_23861,N_17941,N_13342);
nand U23862 (N_23862,N_18659,N_18513);
nand U23863 (N_23863,N_18747,N_13301);
xnor U23864 (N_23864,N_14291,N_18388);
and U23865 (N_23865,N_16179,N_18252);
nand U23866 (N_23866,N_17548,N_13080);
and U23867 (N_23867,N_13501,N_14665);
nand U23868 (N_23868,N_18334,N_16703);
nand U23869 (N_23869,N_15030,N_16055);
nor U23870 (N_23870,N_13635,N_15111);
nand U23871 (N_23871,N_18188,N_17250);
xnor U23872 (N_23872,N_17502,N_15514);
nor U23873 (N_23873,N_12806,N_17502);
and U23874 (N_23874,N_14312,N_17419);
nand U23875 (N_23875,N_13468,N_18054);
nand U23876 (N_23876,N_18538,N_15043);
and U23877 (N_23877,N_14698,N_17583);
xnor U23878 (N_23878,N_13642,N_16077);
nor U23879 (N_23879,N_16589,N_14589);
xnor U23880 (N_23880,N_17964,N_16437);
nor U23881 (N_23881,N_12976,N_17333);
and U23882 (N_23882,N_13846,N_14316);
or U23883 (N_23883,N_17300,N_15229);
nand U23884 (N_23884,N_12973,N_16664);
xor U23885 (N_23885,N_15078,N_17895);
nand U23886 (N_23886,N_16647,N_14232);
and U23887 (N_23887,N_15273,N_15250);
nand U23888 (N_23888,N_14611,N_14753);
or U23889 (N_23889,N_17676,N_13743);
xnor U23890 (N_23890,N_15647,N_15186);
nor U23891 (N_23891,N_17396,N_14370);
nand U23892 (N_23892,N_17051,N_18021);
nor U23893 (N_23893,N_16212,N_15199);
xor U23894 (N_23894,N_18245,N_14310);
or U23895 (N_23895,N_14749,N_16988);
nand U23896 (N_23896,N_14838,N_16751);
and U23897 (N_23897,N_15658,N_17356);
or U23898 (N_23898,N_13987,N_18227);
nor U23899 (N_23899,N_14481,N_18601);
nor U23900 (N_23900,N_15788,N_15754);
or U23901 (N_23901,N_18033,N_17799);
nand U23902 (N_23902,N_13474,N_15920);
nor U23903 (N_23903,N_13961,N_16651);
and U23904 (N_23904,N_18717,N_17921);
and U23905 (N_23905,N_16751,N_12705);
nor U23906 (N_23906,N_14518,N_16220);
xnor U23907 (N_23907,N_17472,N_17023);
or U23908 (N_23908,N_12606,N_13196);
or U23909 (N_23909,N_17674,N_16579);
and U23910 (N_23910,N_14754,N_16536);
nor U23911 (N_23911,N_14739,N_16972);
and U23912 (N_23912,N_17131,N_16604);
or U23913 (N_23913,N_15911,N_14629);
and U23914 (N_23914,N_15619,N_12534);
or U23915 (N_23915,N_18693,N_16932);
nor U23916 (N_23916,N_13931,N_14758);
nand U23917 (N_23917,N_17062,N_15255);
xor U23918 (N_23918,N_16146,N_13769);
nor U23919 (N_23919,N_15752,N_14859);
nand U23920 (N_23920,N_18598,N_18649);
xnor U23921 (N_23921,N_16671,N_17107);
nand U23922 (N_23922,N_13398,N_16024);
and U23923 (N_23923,N_18547,N_14215);
and U23924 (N_23924,N_14116,N_18256);
or U23925 (N_23925,N_13085,N_17127);
nor U23926 (N_23926,N_13690,N_13047);
xnor U23927 (N_23927,N_17776,N_12737);
and U23928 (N_23928,N_15119,N_17559);
and U23929 (N_23929,N_18023,N_13173);
nor U23930 (N_23930,N_15702,N_13870);
nor U23931 (N_23931,N_18178,N_17436);
nand U23932 (N_23932,N_16017,N_12742);
and U23933 (N_23933,N_18401,N_16592);
nand U23934 (N_23934,N_13849,N_15445);
nor U23935 (N_23935,N_14533,N_16563);
or U23936 (N_23936,N_17672,N_15777);
or U23937 (N_23937,N_16285,N_13115);
or U23938 (N_23938,N_17098,N_12526);
nand U23939 (N_23939,N_18299,N_17166);
nor U23940 (N_23940,N_15288,N_17750);
nand U23941 (N_23941,N_17947,N_12873);
nor U23942 (N_23942,N_16173,N_17153);
and U23943 (N_23943,N_17700,N_18360);
xnor U23944 (N_23944,N_14302,N_15756);
nand U23945 (N_23945,N_16567,N_18189);
and U23946 (N_23946,N_16885,N_14837);
or U23947 (N_23947,N_15209,N_13172);
nor U23948 (N_23948,N_14342,N_18693);
nor U23949 (N_23949,N_15377,N_13505);
nand U23950 (N_23950,N_15033,N_13735);
nand U23951 (N_23951,N_13248,N_14419);
nor U23952 (N_23952,N_16308,N_16195);
nor U23953 (N_23953,N_15580,N_18206);
nand U23954 (N_23954,N_15219,N_16563);
xor U23955 (N_23955,N_15764,N_15015);
nor U23956 (N_23956,N_16472,N_16812);
and U23957 (N_23957,N_17840,N_15703);
and U23958 (N_23958,N_15378,N_17897);
and U23959 (N_23959,N_13279,N_13228);
or U23960 (N_23960,N_17176,N_17236);
nor U23961 (N_23961,N_14170,N_17172);
nor U23962 (N_23962,N_12541,N_14010);
nor U23963 (N_23963,N_16535,N_15085);
xor U23964 (N_23964,N_17282,N_17744);
xor U23965 (N_23965,N_12565,N_14667);
nor U23966 (N_23966,N_16549,N_12679);
xor U23967 (N_23967,N_12990,N_18125);
nand U23968 (N_23968,N_18059,N_13254);
or U23969 (N_23969,N_16708,N_16812);
nor U23970 (N_23970,N_18220,N_17991);
and U23971 (N_23971,N_16155,N_14516);
or U23972 (N_23972,N_18459,N_16391);
and U23973 (N_23973,N_13393,N_17621);
nand U23974 (N_23974,N_17258,N_14259);
and U23975 (N_23975,N_14366,N_12879);
nand U23976 (N_23976,N_16665,N_17383);
nand U23977 (N_23977,N_17185,N_17819);
nor U23978 (N_23978,N_18731,N_18246);
xnor U23979 (N_23979,N_17348,N_16612);
or U23980 (N_23980,N_14811,N_16659);
nor U23981 (N_23981,N_17985,N_17138);
nand U23982 (N_23982,N_16258,N_15945);
nand U23983 (N_23983,N_12995,N_18486);
xnor U23984 (N_23984,N_12862,N_16541);
or U23985 (N_23985,N_12918,N_15123);
or U23986 (N_23986,N_14680,N_13986);
or U23987 (N_23987,N_17237,N_17529);
nor U23988 (N_23988,N_18382,N_14326);
or U23989 (N_23989,N_13033,N_17508);
or U23990 (N_23990,N_16770,N_13356);
nand U23991 (N_23991,N_15741,N_16581);
or U23992 (N_23992,N_14691,N_18292);
nand U23993 (N_23993,N_18138,N_16952);
xnor U23994 (N_23994,N_17756,N_18486);
nand U23995 (N_23995,N_18271,N_18532);
xnor U23996 (N_23996,N_15302,N_13073);
nor U23997 (N_23997,N_14670,N_15807);
xnor U23998 (N_23998,N_17926,N_15884);
nand U23999 (N_23999,N_14079,N_16606);
or U24000 (N_24000,N_15575,N_18203);
nand U24001 (N_24001,N_16174,N_18160);
nand U24002 (N_24002,N_18679,N_13487);
xnor U24003 (N_24003,N_15636,N_16006);
xor U24004 (N_24004,N_12624,N_16088);
or U24005 (N_24005,N_18633,N_17255);
nand U24006 (N_24006,N_13579,N_16525);
xor U24007 (N_24007,N_14971,N_16011);
and U24008 (N_24008,N_15011,N_16679);
and U24009 (N_24009,N_18302,N_13597);
nand U24010 (N_24010,N_17534,N_15756);
nor U24011 (N_24011,N_14913,N_13366);
xor U24012 (N_24012,N_16173,N_13066);
and U24013 (N_24013,N_14303,N_16463);
xnor U24014 (N_24014,N_17980,N_17732);
xnor U24015 (N_24015,N_18278,N_13144);
xor U24016 (N_24016,N_17358,N_17353);
nand U24017 (N_24017,N_13621,N_13900);
nor U24018 (N_24018,N_13068,N_18243);
xor U24019 (N_24019,N_18028,N_14347);
nor U24020 (N_24020,N_13120,N_17666);
or U24021 (N_24021,N_16739,N_12924);
nand U24022 (N_24022,N_16805,N_13587);
nor U24023 (N_24023,N_14133,N_16611);
xor U24024 (N_24024,N_18630,N_16384);
nand U24025 (N_24025,N_14716,N_16995);
and U24026 (N_24026,N_15427,N_15882);
and U24027 (N_24027,N_17053,N_17262);
and U24028 (N_24028,N_13936,N_13445);
and U24029 (N_24029,N_12827,N_17247);
and U24030 (N_24030,N_13745,N_13031);
nand U24031 (N_24031,N_16539,N_17079);
nor U24032 (N_24032,N_15263,N_13344);
nor U24033 (N_24033,N_13632,N_16319);
nand U24034 (N_24034,N_15735,N_18365);
nor U24035 (N_24035,N_13291,N_14790);
or U24036 (N_24036,N_17960,N_14035);
and U24037 (N_24037,N_13769,N_16879);
nand U24038 (N_24038,N_16918,N_14797);
or U24039 (N_24039,N_18171,N_18358);
xnor U24040 (N_24040,N_17359,N_13322);
or U24041 (N_24041,N_15603,N_16507);
xor U24042 (N_24042,N_12665,N_14423);
nand U24043 (N_24043,N_15967,N_13573);
or U24044 (N_24044,N_13859,N_17646);
and U24045 (N_24045,N_18415,N_13047);
xor U24046 (N_24046,N_18125,N_14993);
nand U24047 (N_24047,N_15027,N_17168);
and U24048 (N_24048,N_14496,N_18193);
xor U24049 (N_24049,N_14820,N_14936);
or U24050 (N_24050,N_12916,N_18117);
nand U24051 (N_24051,N_17916,N_16742);
nand U24052 (N_24052,N_17063,N_12586);
or U24053 (N_24053,N_12858,N_13700);
xor U24054 (N_24054,N_14136,N_16937);
or U24055 (N_24055,N_14846,N_15392);
xor U24056 (N_24056,N_16656,N_18020);
xnor U24057 (N_24057,N_15530,N_18246);
xnor U24058 (N_24058,N_18438,N_12944);
nor U24059 (N_24059,N_12521,N_12715);
nand U24060 (N_24060,N_15540,N_17796);
nand U24061 (N_24061,N_15834,N_12910);
nand U24062 (N_24062,N_13068,N_14096);
nor U24063 (N_24063,N_18379,N_14024);
nand U24064 (N_24064,N_17469,N_14877);
nand U24065 (N_24065,N_16470,N_14572);
xor U24066 (N_24066,N_13537,N_16957);
nor U24067 (N_24067,N_14911,N_13433);
xnor U24068 (N_24068,N_15019,N_15198);
or U24069 (N_24069,N_17891,N_15435);
xnor U24070 (N_24070,N_14398,N_18017);
or U24071 (N_24071,N_15164,N_17542);
nand U24072 (N_24072,N_15877,N_14473);
or U24073 (N_24073,N_13348,N_14764);
nor U24074 (N_24074,N_13206,N_16444);
xnor U24075 (N_24075,N_16729,N_15833);
xnor U24076 (N_24076,N_13523,N_16353);
or U24077 (N_24077,N_13949,N_15106);
xnor U24078 (N_24078,N_18092,N_13549);
nand U24079 (N_24079,N_16476,N_13043);
nor U24080 (N_24080,N_15896,N_18715);
or U24081 (N_24081,N_17999,N_18518);
and U24082 (N_24082,N_13245,N_12635);
or U24083 (N_24083,N_13261,N_18719);
and U24084 (N_24084,N_18210,N_15207);
and U24085 (N_24085,N_17744,N_18703);
nand U24086 (N_24086,N_18747,N_17580);
nand U24087 (N_24087,N_16113,N_13308);
nor U24088 (N_24088,N_15999,N_16646);
nand U24089 (N_24089,N_13234,N_12808);
xor U24090 (N_24090,N_15466,N_15271);
nor U24091 (N_24091,N_15599,N_16826);
and U24092 (N_24092,N_14758,N_18605);
nand U24093 (N_24093,N_16902,N_16209);
or U24094 (N_24094,N_16651,N_15671);
and U24095 (N_24095,N_15904,N_12602);
or U24096 (N_24096,N_15985,N_13805);
and U24097 (N_24097,N_16314,N_18665);
nand U24098 (N_24098,N_16063,N_15991);
xnor U24099 (N_24099,N_15783,N_13049);
nor U24100 (N_24100,N_15066,N_17106);
nand U24101 (N_24101,N_16399,N_17332);
nand U24102 (N_24102,N_14227,N_15098);
nand U24103 (N_24103,N_13000,N_15953);
or U24104 (N_24104,N_17132,N_17437);
and U24105 (N_24105,N_13183,N_14024);
nand U24106 (N_24106,N_14928,N_16731);
xor U24107 (N_24107,N_12889,N_16963);
and U24108 (N_24108,N_13886,N_18420);
or U24109 (N_24109,N_18611,N_15455);
nand U24110 (N_24110,N_14960,N_15074);
or U24111 (N_24111,N_18092,N_14547);
xnor U24112 (N_24112,N_15217,N_15827);
nand U24113 (N_24113,N_18471,N_17644);
xor U24114 (N_24114,N_15192,N_16084);
nor U24115 (N_24115,N_14199,N_15513);
xnor U24116 (N_24116,N_18304,N_15195);
and U24117 (N_24117,N_17473,N_12533);
or U24118 (N_24118,N_17698,N_13496);
nor U24119 (N_24119,N_15609,N_13430);
nand U24120 (N_24120,N_13786,N_17478);
or U24121 (N_24121,N_15179,N_17946);
or U24122 (N_24122,N_15967,N_18724);
or U24123 (N_24123,N_18448,N_14028);
or U24124 (N_24124,N_17747,N_13990);
xnor U24125 (N_24125,N_18213,N_18673);
nor U24126 (N_24126,N_15494,N_12860);
nand U24127 (N_24127,N_14763,N_14331);
xnor U24128 (N_24128,N_15541,N_17933);
or U24129 (N_24129,N_15815,N_15467);
and U24130 (N_24130,N_12509,N_15468);
and U24131 (N_24131,N_14814,N_14142);
xor U24132 (N_24132,N_16271,N_14611);
nor U24133 (N_24133,N_14113,N_14616);
or U24134 (N_24134,N_13869,N_14131);
nand U24135 (N_24135,N_14465,N_14555);
nor U24136 (N_24136,N_18004,N_14736);
or U24137 (N_24137,N_16192,N_12622);
and U24138 (N_24138,N_16162,N_13602);
or U24139 (N_24139,N_13873,N_16377);
or U24140 (N_24140,N_16973,N_16913);
and U24141 (N_24141,N_17780,N_17129);
xnor U24142 (N_24142,N_17327,N_14443);
and U24143 (N_24143,N_18273,N_17032);
and U24144 (N_24144,N_17130,N_13128);
and U24145 (N_24145,N_12957,N_15066);
xnor U24146 (N_24146,N_16964,N_17046);
nor U24147 (N_24147,N_17595,N_15476);
xor U24148 (N_24148,N_13019,N_18248);
nor U24149 (N_24149,N_14274,N_14516);
nand U24150 (N_24150,N_17329,N_16908);
nor U24151 (N_24151,N_13291,N_16138);
nor U24152 (N_24152,N_13699,N_18161);
nor U24153 (N_24153,N_17657,N_13509);
and U24154 (N_24154,N_15765,N_13949);
xor U24155 (N_24155,N_14864,N_13315);
xor U24156 (N_24156,N_17571,N_18562);
nand U24157 (N_24157,N_13078,N_15922);
nor U24158 (N_24158,N_15861,N_15588);
nand U24159 (N_24159,N_14427,N_13973);
xor U24160 (N_24160,N_18391,N_17268);
or U24161 (N_24161,N_14429,N_17722);
xor U24162 (N_24162,N_15342,N_14995);
and U24163 (N_24163,N_16184,N_14709);
and U24164 (N_24164,N_18513,N_13610);
nor U24165 (N_24165,N_17228,N_14322);
and U24166 (N_24166,N_13362,N_15001);
or U24167 (N_24167,N_13273,N_15227);
xnor U24168 (N_24168,N_16353,N_18408);
or U24169 (N_24169,N_13927,N_13227);
and U24170 (N_24170,N_12576,N_18736);
nand U24171 (N_24171,N_13136,N_13366);
xor U24172 (N_24172,N_12558,N_15484);
xnor U24173 (N_24173,N_16043,N_17504);
nand U24174 (N_24174,N_16651,N_15273);
and U24175 (N_24175,N_13296,N_15484);
or U24176 (N_24176,N_18254,N_14700);
xnor U24177 (N_24177,N_12941,N_13516);
and U24178 (N_24178,N_14121,N_12797);
xor U24179 (N_24179,N_15693,N_17324);
or U24180 (N_24180,N_13319,N_18259);
nor U24181 (N_24181,N_17356,N_18690);
nand U24182 (N_24182,N_17648,N_15654);
and U24183 (N_24183,N_15178,N_14751);
or U24184 (N_24184,N_15232,N_13282);
nor U24185 (N_24185,N_15976,N_17661);
or U24186 (N_24186,N_18525,N_12782);
nor U24187 (N_24187,N_13882,N_13321);
and U24188 (N_24188,N_16650,N_12830);
nand U24189 (N_24189,N_16795,N_14142);
nand U24190 (N_24190,N_14263,N_17143);
nor U24191 (N_24191,N_17818,N_12895);
xnor U24192 (N_24192,N_17426,N_14729);
nor U24193 (N_24193,N_13374,N_15016);
and U24194 (N_24194,N_17891,N_18485);
or U24195 (N_24195,N_13853,N_12517);
and U24196 (N_24196,N_17644,N_15539);
and U24197 (N_24197,N_17215,N_15802);
xnor U24198 (N_24198,N_17462,N_16546);
nor U24199 (N_24199,N_17211,N_17866);
or U24200 (N_24200,N_15260,N_13629);
or U24201 (N_24201,N_16807,N_18478);
and U24202 (N_24202,N_17157,N_16455);
and U24203 (N_24203,N_14961,N_14128);
nand U24204 (N_24204,N_13298,N_14669);
nor U24205 (N_24205,N_15468,N_18540);
nand U24206 (N_24206,N_16015,N_13510);
nand U24207 (N_24207,N_15464,N_13451);
nand U24208 (N_24208,N_16238,N_15874);
or U24209 (N_24209,N_16536,N_16428);
or U24210 (N_24210,N_18193,N_14172);
xor U24211 (N_24211,N_17685,N_15952);
xor U24212 (N_24212,N_17468,N_17083);
xnor U24213 (N_24213,N_16430,N_17942);
nand U24214 (N_24214,N_13339,N_13089);
nor U24215 (N_24215,N_16149,N_14109);
xor U24216 (N_24216,N_15534,N_15312);
nor U24217 (N_24217,N_16379,N_14612);
nor U24218 (N_24218,N_13928,N_15027);
nand U24219 (N_24219,N_14303,N_18613);
nand U24220 (N_24220,N_14963,N_17504);
xor U24221 (N_24221,N_13891,N_15155);
and U24222 (N_24222,N_16966,N_15068);
nor U24223 (N_24223,N_17672,N_15356);
or U24224 (N_24224,N_13430,N_17950);
nor U24225 (N_24225,N_17115,N_14426);
and U24226 (N_24226,N_17129,N_17636);
and U24227 (N_24227,N_12608,N_18724);
xnor U24228 (N_24228,N_17671,N_15775);
or U24229 (N_24229,N_18240,N_13865);
and U24230 (N_24230,N_12915,N_16113);
xnor U24231 (N_24231,N_15175,N_14627);
nand U24232 (N_24232,N_12753,N_13499);
and U24233 (N_24233,N_18243,N_18693);
and U24234 (N_24234,N_13950,N_13114);
nand U24235 (N_24235,N_18664,N_17576);
xnor U24236 (N_24236,N_15888,N_16405);
and U24237 (N_24237,N_12854,N_17625);
nor U24238 (N_24238,N_17884,N_14786);
nor U24239 (N_24239,N_14721,N_18122);
and U24240 (N_24240,N_15823,N_18547);
or U24241 (N_24241,N_17306,N_15218);
nand U24242 (N_24242,N_13135,N_16635);
and U24243 (N_24243,N_12836,N_16416);
nand U24244 (N_24244,N_16968,N_13942);
and U24245 (N_24245,N_16813,N_15712);
or U24246 (N_24246,N_16427,N_16543);
nor U24247 (N_24247,N_16966,N_18670);
and U24248 (N_24248,N_12724,N_17716);
nor U24249 (N_24249,N_13416,N_15175);
and U24250 (N_24250,N_17202,N_13433);
nand U24251 (N_24251,N_13057,N_14408);
nor U24252 (N_24252,N_14083,N_18016);
nor U24253 (N_24253,N_16176,N_18032);
nor U24254 (N_24254,N_18189,N_18327);
nor U24255 (N_24255,N_17687,N_17010);
and U24256 (N_24256,N_15677,N_15179);
or U24257 (N_24257,N_17049,N_17842);
nand U24258 (N_24258,N_16604,N_18003);
nand U24259 (N_24259,N_12582,N_14751);
nand U24260 (N_24260,N_14192,N_16412);
and U24261 (N_24261,N_13468,N_17886);
nor U24262 (N_24262,N_15419,N_17795);
or U24263 (N_24263,N_17072,N_12714);
nor U24264 (N_24264,N_16142,N_17144);
xor U24265 (N_24265,N_15751,N_16321);
nor U24266 (N_24266,N_16044,N_13055);
nand U24267 (N_24267,N_14467,N_16840);
nor U24268 (N_24268,N_16347,N_15740);
nand U24269 (N_24269,N_13243,N_14649);
nand U24270 (N_24270,N_12568,N_16330);
nor U24271 (N_24271,N_17925,N_17011);
nand U24272 (N_24272,N_18736,N_17702);
nand U24273 (N_24273,N_12645,N_16957);
xnor U24274 (N_24274,N_15408,N_18696);
nor U24275 (N_24275,N_17878,N_14409);
nor U24276 (N_24276,N_18083,N_14788);
or U24277 (N_24277,N_18253,N_15857);
nand U24278 (N_24278,N_17488,N_17976);
xor U24279 (N_24279,N_15431,N_14606);
nand U24280 (N_24280,N_13380,N_14532);
and U24281 (N_24281,N_16248,N_18517);
nand U24282 (N_24282,N_12941,N_16202);
nand U24283 (N_24283,N_17378,N_17719);
nand U24284 (N_24284,N_15469,N_17057);
nor U24285 (N_24285,N_17489,N_15206);
nand U24286 (N_24286,N_17370,N_15842);
nor U24287 (N_24287,N_12655,N_13610);
nand U24288 (N_24288,N_14574,N_16839);
or U24289 (N_24289,N_17286,N_13150);
nor U24290 (N_24290,N_12773,N_14461);
nor U24291 (N_24291,N_14727,N_13143);
and U24292 (N_24292,N_14999,N_14737);
and U24293 (N_24293,N_16279,N_13237);
nor U24294 (N_24294,N_18425,N_14833);
xor U24295 (N_24295,N_15106,N_17322);
nand U24296 (N_24296,N_18196,N_16276);
nor U24297 (N_24297,N_14737,N_15247);
or U24298 (N_24298,N_18183,N_14277);
nor U24299 (N_24299,N_16059,N_14840);
nand U24300 (N_24300,N_16848,N_18543);
nand U24301 (N_24301,N_13527,N_15088);
and U24302 (N_24302,N_18258,N_13050);
xnor U24303 (N_24303,N_13332,N_12617);
nand U24304 (N_24304,N_15799,N_13006);
xor U24305 (N_24305,N_17971,N_12505);
nand U24306 (N_24306,N_16400,N_15408);
nor U24307 (N_24307,N_16387,N_15540);
and U24308 (N_24308,N_14505,N_13408);
and U24309 (N_24309,N_13931,N_13523);
nand U24310 (N_24310,N_12994,N_15250);
nor U24311 (N_24311,N_18708,N_14124);
xor U24312 (N_24312,N_17017,N_18662);
xnor U24313 (N_24313,N_18284,N_13228);
xor U24314 (N_24314,N_16401,N_14114);
or U24315 (N_24315,N_12995,N_15816);
or U24316 (N_24316,N_12973,N_15243);
or U24317 (N_24317,N_18030,N_15359);
nor U24318 (N_24318,N_12962,N_15386);
nor U24319 (N_24319,N_17660,N_14679);
and U24320 (N_24320,N_14875,N_16016);
nand U24321 (N_24321,N_12718,N_18253);
and U24322 (N_24322,N_16193,N_16728);
nor U24323 (N_24323,N_13448,N_17337);
or U24324 (N_24324,N_18068,N_14019);
and U24325 (N_24325,N_17149,N_15868);
nor U24326 (N_24326,N_16600,N_18058);
and U24327 (N_24327,N_16793,N_16293);
xor U24328 (N_24328,N_14308,N_15447);
or U24329 (N_24329,N_14350,N_14288);
nor U24330 (N_24330,N_12937,N_12856);
xor U24331 (N_24331,N_17373,N_14462);
or U24332 (N_24332,N_17470,N_14630);
and U24333 (N_24333,N_16543,N_14064);
nor U24334 (N_24334,N_15082,N_17159);
nor U24335 (N_24335,N_12743,N_15130);
nand U24336 (N_24336,N_15674,N_17740);
nand U24337 (N_24337,N_15178,N_15892);
nor U24338 (N_24338,N_16024,N_18738);
nand U24339 (N_24339,N_17228,N_16135);
xor U24340 (N_24340,N_12765,N_18328);
and U24341 (N_24341,N_18469,N_16695);
and U24342 (N_24342,N_13189,N_16798);
nand U24343 (N_24343,N_14109,N_18136);
or U24344 (N_24344,N_12617,N_14698);
xnor U24345 (N_24345,N_17682,N_14684);
xor U24346 (N_24346,N_17528,N_13101);
or U24347 (N_24347,N_13909,N_13934);
and U24348 (N_24348,N_17753,N_15551);
nor U24349 (N_24349,N_17913,N_17409);
and U24350 (N_24350,N_13277,N_17206);
nand U24351 (N_24351,N_14555,N_16500);
nand U24352 (N_24352,N_12930,N_18417);
nand U24353 (N_24353,N_15171,N_17167);
nand U24354 (N_24354,N_16085,N_13578);
and U24355 (N_24355,N_15333,N_14905);
and U24356 (N_24356,N_17323,N_13712);
nand U24357 (N_24357,N_13125,N_18511);
and U24358 (N_24358,N_14719,N_18546);
xnor U24359 (N_24359,N_17552,N_14840);
or U24360 (N_24360,N_16786,N_15855);
xnor U24361 (N_24361,N_17674,N_14210);
nand U24362 (N_24362,N_18723,N_16793);
and U24363 (N_24363,N_13420,N_17349);
nor U24364 (N_24364,N_14436,N_14338);
or U24365 (N_24365,N_13481,N_14863);
and U24366 (N_24366,N_17234,N_17978);
or U24367 (N_24367,N_12501,N_16729);
nor U24368 (N_24368,N_17225,N_15608);
or U24369 (N_24369,N_17358,N_12947);
or U24370 (N_24370,N_14973,N_17455);
nand U24371 (N_24371,N_12819,N_15011);
or U24372 (N_24372,N_15378,N_14924);
nor U24373 (N_24373,N_12622,N_17583);
nand U24374 (N_24374,N_12601,N_14410);
xor U24375 (N_24375,N_15211,N_18383);
and U24376 (N_24376,N_13300,N_17149);
and U24377 (N_24377,N_17721,N_13940);
or U24378 (N_24378,N_15796,N_13219);
or U24379 (N_24379,N_17785,N_13401);
nand U24380 (N_24380,N_17792,N_18029);
nor U24381 (N_24381,N_12639,N_14314);
xor U24382 (N_24382,N_14770,N_15195);
nor U24383 (N_24383,N_14204,N_16477);
or U24384 (N_24384,N_17090,N_15604);
nor U24385 (N_24385,N_15530,N_17389);
nand U24386 (N_24386,N_17485,N_18172);
or U24387 (N_24387,N_13163,N_16176);
nand U24388 (N_24388,N_17449,N_16159);
and U24389 (N_24389,N_15543,N_13665);
nand U24390 (N_24390,N_18452,N_17291);
and U24391 (N_24391,N_17773,N_14787);
nor U24392 (N_24392,N_18209,N_17923);
xor U24393 (N_24393,N_17426,N_17078);
and U24394 (N_24394,N_18434,N_15422);
and U24395 (N_24395,N_16092,N_17949);
nor U24396 (N_24396,N_15205,N_13783);
nor U24397 (N_24397,N_18414,N_14668);
or U24398 (N_24398,N_13880,N_14156);
or U24399 (N_24399,N_16500,N_14497);
nor U24400 (N_24400,N_15995,N_17858);
nand U24401 (N_24401,N_13065,N_15379);
and U24402 (N_24402,N_15444,N_14091);
nand U24403 (N_24403,N_18611,N_14594);
nand U24404 (N_24404,N_18084,N_16745);
nor U24405 (N_24405,N_16827,N_18010);
or U24406 (N_24406,N_18647,N_12897);
nand U24407 (N_24407,N_13613,N_13396);
and U24408 (N_24408,N_15492,N_16670);
nor U24409 (N_24409,N_14625,N_17746);
or U24410 (N_24410,N_18464,N_12911);
and U24411 (N_24411,N_16410,N_16052);
nand U24412 (N_24412,N_12602,N_14209);
or U24413 (N_24413,N_18672,N_17862);
and U24414 (N_24414,N_14172,N_18278);
or U24415 (N_24415,N_13648,N_12993);
nor U24416 (N_24416,N_12895,N_17148);
xor U24417 (N_24417,N_14927,N_17021);
or U24418 (N_24418,N_12970,N_15304);
nand U24419 (N_24419,N_13878,N_15621);
nor U24420 (N_24420,N_15250,N_16426);
or U24421 (N_24421,N_16279,N_18053);
xnor U24422 (N_24422,N_14663,N_14938);
or U24423 (N_24423,N_14540,N_13632);
or U24424 (N_24424,N_16165,N_16419);
or U24425 (N_24425,N_15815,N_13842);
nand U24426 (N_24426,N_14085,N_17553);
or U24427 (N_24427,N_14361,N_14424);
or U24428 (N_24428,N_15337,N_12890);
and U24429 (N_24429,N_14734,N_15530);
xor U24430 (N_24430,N_17048,N_17853);
nand U24431 (N_24431,N_14574,N_16483);
xor U24432 (N_24432,N_13360,N_13405);
nand U24433 (N_24433,N_13741,N_17230);
and U24434 (N_24434,N_16131,N_15970);
or U24435 (N_24435,N_15968,N_14182);
nor U24436 (N_24436,N_15278,N_15844);
xor U24437 (N_24437,N_13024,N_18440);
or U24438 (N_24438,N_13109,N_13800);
xnor U24439 (N_24439,N_12801,N_14017);
xnor U24440 (N_24440,N_17803,N_16647);
nor U24441 (N_24441,N_17385,N_13450);
xor U24442 (N_24442,N_18580,N_15810);
nand U24443 (N_24443,N_16767,N_17086);
nand U24444 (N_24444,N_15526,N_17147);
nor U24445 (N_24445,N_15202,N_12732);
or U24446 (N_24446,N_14735,N_14780);
or U24447 (N_24447,N_16860,N_14616);
xnor U24448 (N_24448,N_18070,N_17767);
and U24449 (N_24449,N_15029,N_16807);
nand U24450 (N_24450,N_14610,N_14831);
xnor U24451 (N_24451,N_18148,N_13601);
and U24452 (N_24452,N_14324,N_18256);
xor U24453 (N_24453,N_18356,N_17023);
or U24454 (N_24454,N_14990,N_18441);
nor U24455 (N_24455,N_17692,N_15433);
xor U24456 (N_24456,N_18663,N_13143);
nand U24457 (N_24457,N_14407,N_15112);
nor U24458 (N_24458,N_15575,N_13275);
nor U24459 (N_24459,N_13290,N_14802);
and U24460 (N_24460,N_16968,N_15308);
and U24461 (N_24461,N_17929,N_16940);
nand U24462 (N_24462,N_17550,N_12984);
and U24463 (N_24463,N_12894,N_17078);
or U24464 (N_24464,N_14549,N_16525);
and U24465 (N_24465,N_18246,N_17715);
nand U24466 (N_24466,N_13064,N_13963);
or U24467 (N_24467,N_14166,N_15437);
nor U24468 (N_24468,N_12970,N_16366);
nor U24469 (N_24469,N_17396,N_14057);
xor U24470 (N_24470,N_16146,N_16393);
xor U24471 (N_24471,N_14818,N_16430);
nand U24472 (N_24472,N_14779,N_16003);
nand U24473 (N_24473,N_16844,N_15346);
nor U24474 (N_24474,N_12963,N_16911);
nor U24475 (N_24475,N_16921,N_15704);
and U24476 (N_24476,N_14565,N_13469);
xor U24477 (N_24477,N_13900,N_15906);
nand U24478 (N_24478,N_16680,N_13560);
nand U24479 (N_24479,N_13879,N_18553);
nand U24480 (N_24480,N_18613,N_16689);
xor U24481 (N_24481,N_13524,N_12880);
and U24482 (N_24482,N_16079,N_14071);
nor U24483 (N_24483,N_13047,N_14796);
nor U24484 (N_24484,N_16433,N_18033);
and U24485 (N_24485,N_17225,N_13663);
or U24486 (N_24486,N_12858,N_12986);
nor U24487 (N_24487,N_16586,N_15810);
nand U24488 (N_24488,N_16912,N_13337);
and U24489 (N_24489,N_12512,N_17602);
xor U24490 (N_24490,N_16713,N_13356);
nor U24491 (N_24491,N_15653,N_14641);
nand U24492 (N_24492,N_13104,N_16795);
or U24493 (N_24493,N_13374,N_15636);
nand U24494 (N_24494,N_13035,N_15089);
nand U24495 (N_24495,N_12943,N_13593);
or U24496 (N_24496,N_14142,N_16430);
nand U24497 (N_24497,N_13520,N_15892);
nor U24498 (N_24498,N_18644,N_16126);
nand U24499 (N_24499,N_12704,N_16952);
nand U24500 (N_24500,N_16104,N_16806);
nand U24501 (N_24501,N_15844,N_18427);
or U24502 (N_24502,N_17145,N_13605);
nand U24503 (N_24503,N_16209,N_14722);
nor U24504 (N_24504,N_14182,N_18485);
or U24505 (N_24505,N_17883,N_13864);
or U24506 (N_24506,N_16735,N_15812);
nand U24507 (N_24507,N_15306,N_18270);
nand U24508 (N_24508,N_14637,N_15241);
or U24509 (N_24509,N_17200,N_13261);
nand U24510 (N_24510,N_13136,N_13603);
nor U24511 (N_24511,N_14087,N_15993);
and U24512 (N_24512,N_18119,N_16135);
or U24513 (N_24513,N_15988,N_14444);
nor U24514 (N_24514,N_13005,N_13587);
or U24515 (N_24515,N_17843,N_14670);
and U24516 (N_24516,N_18474,N_14925);
nand U24517 (N_24517,N_14122,N_14711);
xnor U24518 (N_24518,N_16873,N_17066);
or U24519 (N_24519,N_15557,N_17131);
or U24520 (N_24520,N_14859,N_13735);
and U24521 (N_24521,N_17594,N_14650);
xnor U24522 (N_24522,N_14542,N_18219);
nand U24523 (N_24523,N_17886,N_12832);
or U24524 (N_24524,N_17144,N_16327);
nor U24525 (N_24525,N_18488,N_17248);
nand U24526 (N_24526,N_12838,N_14043);
or U24527 (N_24527,N_15789,N_15778);
or U24528 (N_24528,N_15401,N_15749);
and U24529 (N_24529,N_15814,N_14999);
xor U24530 (N_24530,N_13906,N_15252);
xor U24531 (N_24531,N_13285,N_16334);
xor U24532 (N_24532,N_16799,N_17139);
xnor U24533 (N_24533,N_17930,N_16862);
and U24534 (N_24534,N_12985,N_15044);
or U24535 (N_24535,N_14075,N_15239);
and U24536 (N_24536,N_14367,N_18033);
nor U24537 (N_24537,N_12793,N_15915);
or U24538 (N_24538,N_14796,N_16795);
nor U24539 (N_24539,N_16125,N_14401);
nand U24540 (N_24540,N_17203,N_14120);
nand U24541 (N_24541,N_15091,N_12721);
or U24542 (N_24542,N_17234,N_12912);
xor U24543 (N_24543,N_18596,N_15966);
xor U24544 (N_24544,N_17473,N_13579);
nand U24545 (N_24545,N_17884,N_18069);
nor U24546 (N_24546,N_17493,N_14275);
xor U24547 (N_24547,N_14956,N_13067);
and U24548 (N_24548,N_15737,N_18143);
xor U24549 (N_24549,N_15464,N_18674);
nor U24550 (N_24550,N_14665,N_17944);
nand U24551 (N_24551,N_17050,N_18494);
xnor U24552 (N_24552,N_12954,N_12599);
and U24553 (N_24553,N_17860,N_16183);
nor U24554 (N_24554,N_15370,N_14087);
and U24555 (N_24555,N_14218,N_16132);
and U24556 (N_24556,N_14221,N_17364);
or U24557 (N_24557,N_18187,N_14580);
or U24558 (N_24558,N_16248,N_16893);
or U24559 (N_24559,N_15941,N_18205);
or U24560 (N_24560,N_12544,N_13400);
nor U24561 (N_24561,N_15088,N_16920);
xnor U24562 (N_24562,N_15715,N_17434);
or U24563 (N_24563,N_18691,N_14080);
and U24564 (N_24564,N_16271,N_17412);
xor U24565 (N_24565,N_18113,N_16662);
xor U24566 (N_24566,N_15286,N_12845);
xnor U24567 (N_24567,N_13855,N_14727);
or U24568 (N_24568,N_13791,N_13579);
xnor U24569 (N_24569,N_18389,N_16195);
nor U24570 (N_24570,N_18150,N_14384);
xnor U24571 (N_24571,N_15290,N_18139);
and U24572 (N_24572,N_17584,N_18322);
and U24573 (N_24573,N_16016,N_16808);
and U24574 (N_24574,N_12656,N_17743);
nor U24575 (N_24575,N_15214,N_13570);
or U24576 (N_24576,N_17289,N_12525);
or U24577 (N_24577,N_14098,N_17791);
and U24578 (N_24578,N_15185,N_15563);
and U24579 (N_24579,N_17932,N_13754);
or U24580 (N_24580,N_15360,N_17818);
nand U24581 (N_24581,N_13660,N_16492);
or U24582 (N_24582,N_13338,N_13839);
nor U24583 (N_24583,N_18037,N_12964);
nor U24584 (N_24584,N_18178,N_16135);
nand U24585 (N_24585,N_14673,N_16905);
nor U24586 (N_24586,N_16127,N_12992);
nor U24587 (N_24587,N_17641,N_17350);
nor U24588 (N_24588,N_16992,N_14366);
and U24589 (N_24589,N_14869,N_14531);
nand U24590 (N_24590,N_13170,N_13823);
and U24591 (N_24591,N_17805,N_14183);
or U24592 (N_24592,N_16772,N_15754);
xnor U24593 (N_24593,N_17887,N_14559);
xnor U24594 (N_24594,N_17750,N_12647);
nor U24595 (N_24595,N_15390,N_14782);
nand U24596 (N_24596,N_15942,N_13128);
nor U24597 (N_24597,N_14582,N_12564);
nor U24598 (N_24598,N_16923,N_17539);
nor U24599 (N_24599,N_17613,N_14341);
xnor U24600 (N_24600,N_14975,N_16952);
xnor U24601 (N_24601,N_15058,N_17604);
xor U24602 (N_24602,N_16989,N_17621);
and U24603 (N_24603,N_13258,N_15159);
nand U24604 (N_24604,N_17442,N_18706);
nor U24605 (N_24605,N_14698,N_15287);
or U24606 (N_24606,N_16815,N_13549);
nor U24607 (N_24607,N_18586,N_14041);
or U24608 (N_24608,N_14439,N_15765);
or U24609 (N_24609,N_14431,N_18446);
nand U24610 (N_24610,N_15687,N_15078);
nand U24611 (N_24611,N_14329,N_14472);
nor U24612 (N_24612,N_15342,N_18539);
xor U24613 (N_24613,N_14711,N_13914);
or U24614 (N_24614,N_17455,N_15634);
nor U24615 (N_24615,N_16310,N_17745);
nor U24616 (N_24616,N_14562,N_14383);
xor U24617 (N_24617,N_17662,N_15465);
and U24618 (N_24618,N_15792,N_16807);
nand U24619 (N_24619,N_17326,N_13585);
xor U24620 (N_24620,N_13842,N_14194);
nor U24621 (N_24621,N_12576,N_16995);
and U24622 (N_24622,N_13578,N_17167);
xnor U24623 (N_24623,N_13110,N_17256);
or U24624 (N_24624,N_14069,N_15075);
or U24625 (N_24625,N_13540,N_17174);
nand U24626 (N_24626,N_14890,N_13305);
nand U24627 (N_24627,N_18542,N_14371);
nand U24628 (N_24628,N_16425,N_13574);
nor U24629 (N_24629,N_17771,N_17579);
or U24630 (N_24630,N_17491,N_14483);
xor U24631 (N_24631,N_15904,N_12529);
nor U24632 (N_24632,N_14177,N_15692);
and U24633 (N_24633,N_17356,N_13446);
and U24634 (N_24634,N_16735,N_14395);
or U24635 (N_24635,N_17156,N_14292);
nand U24636 (N_24636,N_18687,N_15118);
or U24637 (N_24637,N_15326,N_18290);
or U24638 (N_24638,N_12522,N_16235);
xnor U24639 (N_24639,N_15764,N_16987);
xnor U24640 (N_24640,N_14649,N_18031);
nand U24641 (N_24641,N_14753,N_18748);
or U24642 (N_24642,N_14913,N_15232);
nor U24643 (N_24643,N_13985,N_13905);
xor U24644 (N_24644,N_16417,N_16952);
xor U24645 (N_24645,N_15700,N_17409);
or U24646 (N_24646,N_15453,N_15488);
nand U24647 (N_24647,N_17396,N_16606);
nor U24648 (N_24648,N_12992,N_17358);
xnor U24649 (N_24649,N_12720,N_12930);
xnor U24650 (N_24650,N_12802,N_17998);
nor U24651 (N_24651,N_14244,N_13891);
and U24652 (N_24652,N_17386,N_17538);
and U24653 (N_24653,N_15011,N_12894);
or U24654 (N_24654,N_15039,N_12957);
nor U24655 (N_24655,N_13543,N_13655);
xnor U24656 (N_24656,N_16368,N_13665);
nor U24657 (N_24657,N_14353,N_14096);
nand U24658 (N_24658,N_17704,N_16867);
xnor U24659 (N_24659,N_16865,N_15921);
and U24660 (N_24660,N_16340,N_17335);
and U24661 (N_24661,N_12873,N_12924);
nor U24662 (N_24662,N_17885,N_17546);
nand U24663 (N_24663,N_18712,N_17707);
nor U24664 (N_24664,N_15874,N_18236);
and U24665 (N_24665,N_14946,N_13866);
nand U24666 (N_24666,N_16239,N_14589);
nor U24667 (N_24667,N_15371,N_12760);
xor U24668 (N_24668,N_17705,N_17848);
or U24669 (N_24669,N_15601,N_18054);
and U24670 (N_24670,N_15032,N_14206);
and U24671 (N_24671,N_16383,N_12901);
or U24672 (N_24672,N_14501,N_13888);
nand U24673 (N_24673,N_18499,N_15708);
nor U24674 (N_24674,N_13814,N_12792);
nand U24675 (N_24675,N_17178,N_17205);
and U24676 (N_24676,N_15914,N_18186);
or U24677 (N_24677,N_13690,N_17799);
and U24678 (N_24678,N_13102,N_13095);
and U24679 (N_24679,N_14763,N_14231);
and U24680 (N_24680,N_17402,N_12580);
or U24681 (N_24681,N_17406,N_15192);
and U24682 (N_24682,N_16486,N_18508);
nor U24683 (N_24683,N_16831,N_17110);
xor U24684 (N_24684,N_14347,N_17326);
xnor U24685 (N_24685,N_16438,N_18261);
or U24686 (N_24686,N_15406,N_15533);
and U24687 (N_24687,N_14666,N_14987);
xnor U24688 (N_24688,N_15167,N_13912);
nand U24689 (N_24689,N_18151,N_15726);
and U24690 (N_24690,N_14868,N_17023);
xnor U24691 (N_24691,N_13071,N_12970);
nand U24692 (N_24692,N_14928,N_15550);
and U24693 (N_24693,N_15484,N_15641);
nand U24694 (N_24694,N_15485,N_16124);
and U24695 (N_24695,N_12530,N_15646);
nand U24696 (N_24696,N_17438,N_18333);
nor U24697 (N_24697,N_12697,N_15345);
and U24698 (N_24698,N_18056,N_17300);
xor U24699 (N_24699,N_12735,N_17008);
and U24700 (N_24700,N_15993,N_17489);
nand U24701 (N_24701,N_13735,N_12613);
xnor U24702 (N_24702,N_18384,N_15744);
and U24703 (N_24703,N_16094,N_16349);
nor U24704 (N_24704,N_17838,N_14644);
and U24705 (N_24705,N_13139,N_15807);
and U24706 (N_24706,N_18677,N_17601);
nand U24707 (N_24707,N_14562,N_13495);
nand U24708 (N_24708,N_18643,N_12778);
nand U24709 (N_24709,N_18639,N_17885);
nand U24710 (N_24710,N_13980,N_16404);
and U24711 (N_24711,N_17481,N_16368);
or U24712 (N_24712,N_16699,N_17685);
nor U24713 (N_24713,N_17617,N_12539);
nand U24714 (N_24714,N_16529,N_15650);
xnor U24715 (N_24715,N_15112,N_16579);
nor U24716 (N_24716,N_17342,N_18299);
xnor U24717 (N_24717,N_18663,N_17080);
xnor U24718 (N_24718,N_12671,N_15444);
nor U24719 (N_24719,N_13411,N_15389);
xor U24720 (N_24720,N_14390,N_15243);
or U24721 (N_24721,N_17529,N_12898);
nand U24722 (N_24722,N_14219,N_12870);
nor U24723 (N_24723,N_16530,N_16722);
nor U24724 (N_24724,N_13425,N_15854);
nand U24725 (N_24725,N_18442,N_14214);
or U24726 (N_24726,N_16784,N_16654);
xnor U24727 (N_24727,N_15721,N_14302);
and U24728 (N_24728,N_15539,N_16394);
xnor U24729 (N_24729,N_14004,N_16982);
nand U24730 (N_24730,N_18330,N_17546);
nand U24731 (N_24731,N_12501,N_18725);
and U24732 (N_24732,N_16544,N_16389);
and U24733 (N_24733,N_14949,N_14307);
xor U24734 (N_24734,N_16373,N_12665);
xnor U24735 (N_24735,N_18120,N_14329);
and U24736 (N_24736,N_17694,N_17321);
and U24737 (N_24737,N_15393,N_14712);
and U24738 (N_24738,N_15274,N_13675);
xor U24739 (N_24739,N_14978,N_14429);
nor U24740 (N_24740,N_18501,N_17951);
xor U24741 (N_24741,N_17584,N_16878);
and U24742 (N_24742,N_17859,N_17619);
and U24743 (N_24743,N_12810,N_15214);
nand U24744 (N_24744,N_14203,N_16823);
or U24745 (N_24745,N_16996,N_17272);
xnor U24746 (N_24746,N_15390,N_16507);
xnor U24747 (N_24747,N_15127,N_16418);
nand U24748 (N_24748,N_13850,N_18278);
and U24749 (N_24749,N_16022,N_17000);
or U24750 (N_24750,N_13127,N_17406);
nand U24751 (N_24751,N_13118,N_17968);
xor U24752 (N_24752,N_14078,N_14989);
nor U24753 (N_24753,N_16767,N_17243);
nand U24754 (N_24754,N_17536,N_17118);
xor U24755 (N_24755,N_14681,N_12573);
nor U24756 (N_24756,N_17756,N_17017);
or U24757 (N_24757,N_13176,N_17016);
nand U24758 (N_24758,N_12614,N_17187);
xor U24759 (N_24759,N_14240,N_16319);
nand U24760 (N_24760,N_13662,N_17868);
nor U24761 (N_24761,N_12615,N_17516);
xnor U24762 (N_24762,N_16885,N_18339);
nand U24763 (N_24763,N_17693,N_13639);
nand U24764 (N_24764,N_12843,N_17791);
nor U24765 (N_24765,N_14707,N_14976);
and U24766 (N_24766,N_16472,N_14508);
xnor U24767 (N_24767,N_13559,N_12731);
nand U24768 (N_24768,N_16395,N_17013);
xor U24769 (N_24769,N_14158,N_17608);
or U24770 (N_24770,N_17836,N_16095);
nor U24771 (N_24771,N_15853,N_18486);
or U24772 (N_24772,N_12947,N_14233);
nor U24773 (N_24773,N_14390,N_14343);
xnor U24774 (N_24774,N_17039,N_14059);
or U24775 (N_24775,N_15502,N_17167);
nand U24776 (N_24776,N_12578,N_18069);
or U24777 (N_24777,N_18116,N_15051);
or U24778 (N_24778,N_16694,N_16663);
nor U24779 (N_24779,N_16019,N_16751);
or U24780 (N_24780,N_17945,N_12769);
or U24781 (N_24781,N_18153,N_16000);
and U24782 (N_24782,N_17421,N_15349);
nor U24783 (N_24783,N_18380,N_16663);
nor U24784 (N_24784,N_15581,N_15116);
or U24785 (N_24785,N_14513,N_18591);
nor U24786 (N_24786,N_13850,N_12916);
and U24787 (N_24787,N_13579,N_16785);
or U24788 (N_24788,N_13082,N_16921);
and U24789 (N_24789,N_13710,N_13990);
and U24790 (N_24790,N_12653,N_17008);
and U24791 (N_24791,N_18561,N_17552);
and U24792 (N_24792,N_14166,N_13633);
xnor U24793 (N_24793,N_17921,N_15157);
nand U24794 (N_24794,N_17400,N_17952);
or U24795 (N_24795,N_14214,N_13469);
nand U24796 (N_24796,N_15769,N_15415);
nor U24797 (N_24797,N_16226,N_16885);
and U24798 (N_24798,N_13936,N_13125);
or U24799 (N_24799,N_15216,N_17118);
nand U24800 (N_24800,N_18479,N_17630);
or U24801 (N_24801,N_15921,N_17021);
and U24802 (N_24802,N_15583,N_15150);
nand U24803 (N_24803,N_12512,N_18430);
xnor U24804 (N_24804,N_13779,N_13796);
nand U24805 (N_24805,N_18589,N_12664);
nand U24806 (N_24806,N_16407,N_15435);
and U24807 (N_24807,N_12688,N_18081);
or U24808 (N_24808,N_17843,N_15996);
and U24809 (N_24809,N_17349,N_17430);
and U24810 (N_24810,N_13092,N_18749);
nand U24811 (N_24811,N_13489,N_14283);
and U24812 (N_24812,N_18015,N_13892);
and U24813 (N_24813,N_16717,N_17308);
nor U24814 (N_24814,N_17515,N_12893);
xor U24815 (N_24815,N_17533,N_17540);
xor U24816 (N_24816,N_16306,N_18389);
or U24817 (N_24817,N_17518,N_16800);
nor U24818 (N_24818,N_13620,N_18652);
nor U24819 (N_24819,N_17419,N_18051);
xnor U24820 (N_24820,N_15499,N_16653);
xor U24821 (N_24821,N_15780,N_14110);
or U24822 (N_24822,N_17230,N_18242);
nor U24823 (N_24823,N_14048,N_18129);
xnor U24824 (N_24824,N_16502,N_12905);
xnor U24825 (N_24825,N_16806,N_17164);
nand U24826 (N_24826,N_16466,N_14267);
or U24827 (N_24827,N_13116,N_17075);
xor U24828 (N_24828,N_16210,N_12705);
xor U24829 (N_24829,N_13954,N_14939);
or U24830 (N_24830,N_14524,N_17416);
xnor U24831 (N_24831,N_12827,N_16177);
xnor U24832 (N_24832,N_13015,N_17718);
or U24833 (N_24833,N_13987,N_17751);
xor U24834 (N_24834,N_14622,N_14999);
nand U24835 (N_24835,N_14510,N_16370);
nand U24836 (N_24836,N_14038,N_12731);
nor U24837 (N_24837,N_17998,N_17317);
nor U24838 (N_24838,N_15262,N_13158);
nor U24839 (N_24839,N_16185,N_14648);
or U24840 (N_24840,N_17932,N_17302);
and U24841 (N_24841,N_16589,N_16019);
nor U24842 (N_24842,N_16825,N_16813);
nor U24843 (N_24843,N_13206,N_17913);
or U24844 (N_24844,N_13272,N_12563);
and U24845 (N_24845,N_14883,N_18319);
xor U24846 (N_24846,N_18660,N_15982);
nor U24847 (N_24847,N_15402,N_15513);
nand U24848 (N_24848,N_18678,N_15043);
or U24849 (N_24849,N_13966,N_15784);
or U24850 (N_24850,N_17964,N_14145);
or U24851 (N_24851,N_14917,N_17035);
xnor U24852 (N_24852,N_13548,N_13729);
nor U24853 (N_24853,N_15101,N_18192);
nor U24854 (N_24854,N_13144,N_14931);
or U24855 (N_24855,N_15198,N_17754);
and U24856 (N_24856,N_15985,N_12650);
xnor U24857 (N_24857,N_17125,N_14463);
and U24858 (N_24858,N_14416,N_14893);
and U24859 (N_24859,N_17863,N_17276);
and U24860 (N_24860,N_13858,N_12729);
and U24861 (N_24861,N_14778,N_12911);
or U24862 (N_24862,N_18412,N_14625);
nor U24863 (N_24863,N_16585,N_17765);
xnor U24864 (N_24864,N_15103,N_15191);
and U24865 (N_24865,N_15332,N_15989);
and U24866 (N_24866,N_12513,N_14685);
xnor U24867 (N_24867,N_15904,N_18329);
nand U24868 (N_24868,N_18465,N_17738);
and U24869 (N_24869,N_16323,N_18694);
or U24870 (N_24870,N_12767,N_16529);
nand U24871 (N_24871,N_14385,N_17777);
nor U24872 (N_24872,N_15269,N_15577);
nor U24873 (N_24873,N_16774,N_15494);
nand U24874 (N_24874,N_14927,N_17630);
xor U24875 (N_24875,N_12985,N_13868);
and U24876 (N_24876,N_12684,N_18432);
nor U24877 (N_24877,N_14739,N_12884);
nor U24878 (N_24878,N_14884,N_13311);
or U24879 (N_24879,N_16387,N_13435);
xnor U24880 (N_24880,N_17164,N_17394);
xnor U24881 (N_24881,N_16740,N_15062);
nor U24882 (N_24882,N_17855,N_18603);
xor U24883 (N_24883,N_13194,N_15474);
and U24884 (N_24884,N_18274,N_12696);
nor U24885 (N_24885,N_17165,N_14110);
nand U24886 (N_24886,N_16179,N_15213);
or U24887 (N_24887,N_15087,N_14390);
nand U24888 (N_24888,N_18087,N_17343);
nand U24889 (N_24889,N_14836,N_12977);
nor U24890 (N_24890,N_17863,N_17368);
nor U24891 (N_24891,N_14746,N_13821);
or U24892 (N_24892,N_14002,N_18626);
or U24893 (N_24893,N_12580,N_15578);
xnor U24894 (N_24894,N_17516,N_15070);
and U24895 (N_24895,N_15782,N_17163);
nand U24896 (N_24896,N_18243,N_18416);
or U24897 (N_24897,N_12915,N_14259);
and U24898 (N_24898,N_12601,N_13126);
or U24899 (N_24899,N_15436,N_14742);
or U24900 (N_24900,N_15706,N_15457);
xor U24901 (N_24901,N_14822,N_12559);
and U24902 (N_24902,N_13508,N_16951);
nor U24903 (N_24903,N_14344,N_12511);
xor U24904 (N_24904,N_13242,N_17886);
nand U24905 (N_24905,N_17574,N_16537);
and U24906 (N_24906,N_17669,N_14141);
xor U24907 (N_24907,N_15510,N_18473);
nand U24908 (N_24908,N_14136,N_15540);
xor U24909 (N_24909,N_17208,N_13199);
or U24910 (N_24910,N_16514,N_17715);
nand U24911 (N_24911,N_17974,N_12898);
or U24912 (N_24912,N_14642,N_17091);
nor U24913 (N_24913,N_18574,N_18096);
and U24914 (N_24914,N_13649,N_12547);
and U24915 (N_24915,N_13660,N_18126);
nand U24916 (N_24916,N_18018,N_13139);
and U24917 (N_24917,N_16836,N_17869);
nor U24918 (N_24918,N_16511,N_14528);
or U24919 (N_24919,N_15928,N_16177);
nor U24920 (N_24920,N_16976,N_12612);
nor U24921 (N_24921,N_14046,N_13395);
xor U24922 (N_24922,N_18474,N_16199);
and U24923 (N_24923,N_16399,N_15634);
and U24924 (N_24924,N_17260,N_15506);
or U24925 (N_24925,N_14800,N_12902);
xor U24926 (N_24926,N_15836,N_15838);
nor U24927 (N_24927,N_16496,N_15594);
and U24928 (N_24928,N_13492,N_14262);
nor U24929 (N_24929,N_14064,N_13738);
or U24930 (N_24930,N_18194,N_12767);
nor U24931 (N_24931,N_18548,N_17568);
xor U24932 (N_24932,N_17278,N_16604);
nand U24933 (N_24933,N_14105,N_13922);
xor U24934 (N_24934,N_12967,N_18356);
and U24935 (N_24935,N_18744,N_17860);
xor U24936 (N_24936,N_12664,N_14226);
xor U24937 (N_24937,N_17248,N_16360);
nand U24938 (N_24938,N_17227,N_16191);
or U24939 (N_24939,N_13544,N_12687);
xnor U24940 (N_24940,N_18596,N_15669);
xor U24941 (N_24941,N_15777,N_13390);
and U24942 (N_24942,N_16315,N_17899);
or U24943 (N_24943,N_16458,N_18152);
nor U24944 (N_24944,N_15704,N_14051);
nand U24945 (N_24945,N_16949,N_15182);
xor U24946 (N_24946,N_12514,N_15075);
nor U24947 (N_24947,N_17195,N_17715);
and U24948 (N_24948,N_14544,N_16937);
xnor U24949 (N_24949,N_14327,N_13975);
or U24950 (N_24950,N_17018,N_15753);
nand U24951 (N_24951,N_18148,N_12510);
nand U24952 (N_24952,N_18434,N_16487);
nand U24953 (N_24953,N_13068,N_18278);
nand U24954 (N_24954,N_17608,N_18733);
nor U24955 (N_24955,N_18680,N_15152);
xor U24956 (N_24956,N_17113,N_15158);
or U24957 (N_24957,N_15457,N_12712);
xor U24958 (N_24958,N_12700,N_15316);
and U24959 (N_24959,N_15912,N_16637);
nor U24960 (N_24960,N_14432,N_15532);
xor U24961 (N_24961,N_13898,N_15419);
nor U24962 (N_24962,N_13297,N_18556);
xor U24963 (N_24963,N_18047,N_16037);
or U24964 (N_24964,N_12609,N_16059);
xor U24965 (N_24965,N_13504,N_13477);
nand U24966 (N_24966,N_18025,N_18194);
and U24967 (N_24967,N_13755,N_18206);
xor U24968 (N_24968,N_13231,N_15904);
nand U24969 (N_24969,N_12666,N_15282);
nor U24970 (N_24970,N_13066,N_13444);
xnor U24971 (N_24971,N_14842,N_15827);
nor U24972 (N_24972,N_13222,N_15742);
xor U24973 (N_24973,N_15672,N_18708);
or U24974 (N_24974,N_13438,N_15476);
or U24975 (N_24975,N_12769,N_17486);
nor U24976 (N_24976,N_12891,N_14340);
or U24977 (N_24977,N_16082,N_17627);
nor U24978 (N_24978,N_15808,N_17192);
or U24979 (N_24979,N_14365,N_15994);
xor U24980 (N_24980,N_13201,N_18256);
and U24981 (N_24981,N_13618,N_13800);
xnor U24982 (N_24982,N_16297,N_13903);
nand U24983 (N_24983,N_18588,N_12725);
and U24984 (N_24984,N_12920,N_14410);
and U24985 (N_24985,N_15257,N_17546);
and U24986 (N_24986,N_16090,N_16656);
xnor U24987 (N_24987,N_14414,N_18486);
and U24988 (N_24988,N_14223,N_18062);
or U24989 (N_24989,N_13759,N_14321);
xor U24990 (N_24990,N_16372,N_18533);
or U24991 (N_24991,N_14931,N_18537);
and U24992 (N_24992,N_14413,N_14269);
or U24993 (N_24993,N_13160,N_16599);
xor U24994 (N_24994,N_15067,N_13002);
and U24995 (N_24995,N_15672,N_18485);
xnor U24996 (N_24996,N_18337,N_17281);
and U24997 (N_24997,N_16450,N_16565);
nor U24998 (N_24998,N_15349,N_15938);
xor U24999 (N_24999,N_13724,N_12822);
nand UO_0 (O_0,N_24264,N_21999);
or UO_1 (O_1,N_19945,N_19259);
nand UO_2 (O_2,N_22518,N_24784);
or UO_3 (O_3,N_23944,N_22362);
and UO_4 (O_4,N_20148,N_20097);
nand UO_5 (O_5,N_23092,N_21690);
or UO_6 (O_6,N_21704,N_22567);
and UO_7 (O_7,N_21971,N_23212);
and UO_8 (O_8,N_21524,N_21674);
nor UO_9 (O_9,N_23912,N_23647);
nor UO_10 (O_10,N_22712,N_19626);
and UO_11 (O_11,N_22405,N_24935);
nor UO_12 (O_12,N_23239,N_21217);
xnor UO_13 (O_13,N_24757,N_19023);
and UO_14 (O_14,N_20152,N_22602);
and UO_15 (O_15,N_23030,N_19197);
nor UO_16 (O_16,N_23392,N_22551);
or UO_17 (O_17,N_19838,N_21309);
and UO_18 (O_18,N_21799,N_22107);
or UO_19 (O_19,N_19534,N_20965);
xor UO_20 (O_20,N_20651,N_23098);
and UO_21 (O_21,N_19428,N_23524);
nor UO_22 (O_22,N_19607,N_22773);
nor UO_23 (O_23,N_21884,N_20857);
nor UO_24 (O_24,N_22461,N_22009);
nand UO_25 (O_25,N_24581,N_19910);
nor UO_26 (O_26,N_23410,N_20584);
nor UO_27 (O_27,N_22149,N_18790);
nand UO_28 (O_28,N_20568,N_22744);
xor UO_29 (O_29,N_20736,N_21509);
nor UO_30 (O_30,N_19163,N_21223);
and UO_31 (O_31,N_18832,N_20223);
and UO_32 (O_32,N_21439,N_23135);
xnor UO_33 (O_33,N_19931,N_19084);
or UO_34 (O_34,N_20942,N_19759);
nand UO_35 (O_35,N_19106,N_20566);
xnor UO_36 (O_36,N_22341,N_21399);
or UO_37 (O_37,N_20534,N_21206);
xnor UO_38 (O_38,N_20463,N_23445);
and UO_39 (O_39,N_19145,N_21843);
nand UO_40 (O_40,N_23115,N_21355);
nand UO_41 (O_41,N_20944,N_20507);
or UO_42 (O_42,N_22636,N_22704);
nand UO_43 (O_43,N_19615,N_23126);
and UO_44 (O_44,N_22080,N_24197);
nor UO_45 (O_45,N_24016,N_21541);
nor UO_46 (O_46,N_19898,N_19899);
xor UO_47 (O_47,N_20428,N_24573);
nand UO_48 (O_48,N_21129,N_18809);
and UO_49 (O_49,N_19577,N_23731);
and UO_50 (O_50,N_22964,N_21059);
nand UO_51 (O_51,N_19734,N_22464);
nand UO_52 (O_52,N_23626,N_21721);
nor UO_53 (O_53,N_22365,N_22971);
and UO_54 (O_54,N_21087,N_19194);
nor UO_55 (O_55,N_23309,N_19047);
nand UO_56 (O_56,N_21047,N_21154);
xor UO_57 (O_57,N_22136,N_24751);
xor UO_58 (O_58,N_23621,N_22643);
xor UO_59 (O_59,N_21640,N_23110);
and UO_60 (O_60,N_22309,N_19420);
nor UO_61 (O_61,N_19599,N_23151);
nand UO_62 (O_62,N_23259,N_20078);
xor UO_63 (O_63,N_22391,N_20861);
nor UO_64 (O_64,N_24919,N_19202);
xor UO_65 (O_65,N_21603,N_20635);
or UO_66 (O_66,N_22846,N_19268);
xor UO_67 (O_67,N_23946,N_24021);
nor UO_68 (O_68,N_19887,N_24647);
nor UO_69 (O_69,N_24672,N_24825);
or UO_70 (O_70,N_20472,N_22446);
nand UO_71 (O_71,N_21708,N_18857);
nand UO_72 (O_72,N_20918,N_23032);
nor UO_73 (O_73,N_22796,N_21761);
xnor UO_74 (O_74,N_21646,N_22538);
and UO_75 (O_75,N_18964,N_23982);
or UO_76 (O_76,N_23646,N_21289);
nor UO_77 (O_77,N_19060,N_24462);
and UO_78 (O_78,N_19390,N_22211);
or UO_79 (O_79,N_20200,N_20423);
xor UO_80 (O_80,N_22992,N_19854);
and UO_81 (O_81,N_22652,N_22326);
nor UO_82 (O_82,N_22085,N_21575);
xnor UO_83 (O_83,N_19857,N_19940);
nor UO_84 (O_84,N_18975,N_21747);
nor UO_85 (O_85,N_21307,N_20885);
xor UO_86 (O_86,N_21095,N_23473);
or UO_87 (O_87,N_21490,N_21769);
xnor UO_88 (O_88,N_19653,N_22675);
nor UO_89 (O_89,N_22465,N_22916);
and UO_90 (O_90,N_23661,N_19487);
or UO_91 (O_91,N_23291,N_24137);
nor UO_92 (O_92,N_23520,N_19966);
nor UO_93 (O_93,N_24775,N_21876);
nor UO_94 (O_94,N_19529,N_20840);
and UO_95 (O_95,N_19647,N_22479);
nor UO_96 (O_96,N_19422,N_24731);
or UO_97 (O_97,N_21466,N_19355);
xor UO_98 (O_98,N_23539,N_24830);
or UO_99 (O_99,N_21369,N_19425);
xor UO_100 (O_100,N_22584,N_19446);
xnor UO_101 (O_101,N_23750,N_22889);
nor UO_102 (O_102,N_20000,N_23562);
xnor UO_103 (O_103,N_19370,N_19474);
or UO_104 (O_104,N_24285,N_18982);
nor UO_105 (O_105,N_23889,N_20034);
xnor UO_106 (O_106,N_21513,N_19712);
nor UO_107 (O_107,N_21498,N_22590);
xor UO_108 (O_108,N_21684,N_23699);
nand UO_109 (O_109,N_21290,N_20720);
or UO_110 (O_110,N_20661,N_21112);
xnor UO_111 (O_111,N_22497,N_23512);
nand UO_112 (O_112,N_21548,N_19770);
xnor UO_113 (O_113,N_23854,N_24044);
xnor UO_114 (O_114,N_19188,N_24798);
xnor UO_115 (O_115,N_20043,N_19120);
and UO_116 (O_116,N_19150,N_21121);
nand UO_117 (O_117,N_24539,N_23173);
nor UO_118 (O_118,N_22789,N_24867);
or UO_119 (O_119,N_22027,N_24811);
nand UO_120 (O_120,N_20754,N_24135);
nor UO_121 (O_121,N_22170,N_24275);
and UO_122 (O_122,N_20216,N_23303);
or UO_123 (O_123,N_23070,N_19609);
nand UO_124 (O_124,N_19637,N_21225);
nor UO_125 (O_125,N_24450,N_23448);
nor UO_126 (O_126,N_21109,N_20979);
or UO_127 (O_127,N_23142,N_19782);
nand UO_128 (O_128,N_22867,N_21350);
xor UO_129 (O_129,N_20529,N_21032);
nand UO_130 (O_130,N_19462,N_21444);
nor UO_131 (O_131,N_23915,N_19727);
xnor UO_132 (O_132,N_21797,N_20949);
nand UO_133 (O_133,N_19318,N_18897);
or UO_134 (O_134,N_23736,N_19121);
nor UO_135 (O_135,N_21322,N_23163);
nand UO_136 (O_136,N_21858,N_21072);
nand UO_137 (O_137,N_24330,N_23877);
nand UO_138 (O_138,N_22904,N_23614);
nand UO_139 (O_139,N_20275,N_20518);
and UO_140 (O_140,N_20176,N_24478);
or UO_141 (O_141,N_21919,N_21991);
nand UO_142 (O_142,N_22310,N_22190);
nand UO_143 (O_143,N_22022,N_23475);
nand UO_144 (O_144,N_19287,N_23814);
nand UO_145 (O_145,N_24753,N_20737);
xor UO_146 (O_146,N_21897,N_19969);
nand UO_147 (O_147,N_19872,N_24957);
and UO_148 (O_148,N_19654,N_24054);
nor UO_149 (O_149,N_19600,N_22532);
nand UO_150 (O_150,N_24587,N_24964);
nand UO_151 (O_151,N_24903,N_23454);
nor UO_152 (O_152,N_22577,N_19914);
nand UO_153 (O_153,N_20978,N_24040);
nand UO_154 (O_154,N_22018,N_20970);
nor UO_155 (O_155,N_21330,N_22220);
or UO_156 (O_156,N_21437,N_19745);
xnor UO_157 (O_157,N_20118,N_20386);
or UO_158 (O_158,N_21910,N_23033);
nor UO_159 (O_159,N_20186,N_24405);
xnor UO_160 (O_160,N_24008,N_20930);
nor UO_161 (O_161,N_21004,N_24748);
or UO_162 (O_162,N_20811,N_21807);
and UO_163 (O_163,N_20788,N_23093);
xor UO_164 (O_164,N_19317,N_21683);
or UO_165 (O_165,N_21793,N_24041);
and UO_166 (O_166,N_18924,N_19291);
and UO_167 (O_167,N_24737,N_23930);
or UO_168 (O_168,N_23997,N_22760);
or UO_169 (O_169,N_22963,N_22345);
xnor UO_170 (O_170,N_21782,N_22657);
and UO_171 (O_171,N_22293,N_20286);
nor UO_172 (O_172,N_22694,N_24743);
xnor UO_173 (O_173,N_23594,N_20458);
nand UO_174 (O_174,N_21600,N_18847);
nand UO_175 (O_175,N_22677,N_22986);
and UO_176 (O_176,N_19398,N_24723);
xnor UO_177 (O_177,N_19808,N_21015);
nand UO_178 (O_178,N_22624,N_21478);
nand UO_179 (O_179,N_20555,N_19724);
xor UO_180 (O_180,N_22687,N_23490);
nand UO_181 (O_181,N_19307,N_23109);
nand UO_182 (O_182,N_18759,N_24296);
xor UO_183 (O_183,N_22113,N_22762);
xnor UO_184 (O_184,N_21311,N_20452);
and UO_185 (O_185,N_22952,N_19869);
or UO_186 (O_186,N_19911,N_20672);
nand UO_187 (O_187,N_21804,N_24902);
xnor UO_188 (O_188,N_19074,N_22161);
nand UO_189 (O_189,N_19913,N_23097);
nor UO_190 (O_190,N_22241,N_23394);
nor UO_191 (O_191,N_19042,N_22861);
and UO_192 (O_192,N_23607,N_21891);
and UO_193 (O_193,N_24501,N_18991);
nand UO_194 (O_194,N_18801,N_22234);
xor UO_195 (O_195,N_19924,N_23738);
and UO_196 (O_196,N_22797,N_20415);
nor UO_197 (O_197,N_18981,N_22934);
xor UO_198 (O_198,N_19226,N_24271);
or UO_199 (O_199,N_23991,N_19744);
and UO_200 (O_200,N_19840,N_21984);
nand UO_201 (O_201,N_21409,N_23245);
nor UO_202 (O_202,N_23044,N_20863);
or UO_203 (O_203,N_23100,N_24231);
or UO_204 (O_204,N_24949,N_21756);
nor UO_205 (O_205,N_19056,N_22219);
or UO_206 (O_206,N_23174,N_24590);
or UO_207 (O_207,N_20947,N_23304);
xnor UO_208 (O_208,N_22360,N_23408);
or UO_209 (O_209,N_20704,N_21762);
nand UO_210 (O_210,N_19246,N_23101);
nand UO_211 (O_211,N_22856,N_20786);
and UO_212 (O_212,N_22500,N_21652);
and UO_213 (O_213,N_24878,N_21040);
xor UO_214 (O_214,N_23599,N_23271);
and UO_215 (O_215,N_21609,N_20189);
nand UO_216 (O_216,N_18978,N_23516);
nand UO_217 (O_217,N_19172,N_18922);
xor UO_218 (O_218,N_19295,N_19697);
xnor UO_219 (O_219,N_22598,N_19382);
and UO_220 (O_220,N_24490,N_19820);
nand UO_221 (O_221,N_21483,N_24159);
nor UO_222 (O_222,N_23747,N_22776);
or UO_223 (O_223,N_20929,N_22553);
nand UO_224 (O_224,N_23210,N_24451);
nand UO_225 (O_225,N_24864,N_23324);
nand UO_226 (O_226,N_21382,N_24497);
or UO_227 (O_227,N_23083,N_21363);
and UO_228 (O_228,N_21617,N_20860);
or UO_229 (O_229,N_20416,N_22945);
and UO_230 (O_230,N_20309,N_22150);
xnor UO_231 (O_231,N_22718,N_24627);
and UO_232 (O_232,N_20351,N_20207);
or UO_233 (O_233,N_19363,N_24065);
nor UO_234 (O_234,N_23327,N_19706);
and UO_235 (O_235,N_21394,N_22033);
nor UO_236 (O_236,N_20036,N_22357);
xnor UO_237 (O_237,N_22116,N_24629);
and UO_238 (O_238,N_24172,N_24715);
xnor UO_239 (O_239,N_22530,N_22880);
nor UO_240 (O_240,N_24885,N_22906);
xor UO_241 (O_241,N_22226,N_21859);
and UO_242 (O_242,N_21120,N_20089);
xor UO_243 (O_243,N_20859,N_21140);
xnor UO_244 (O_244,N_20898,N_23065);
xor UO_245 (O_245,N_21750,N_21806);
xnor UO_246 (O_246,N_23632,N_19799);
or UO_247 (O_247,N_23132,N_19339);
nand UO_248 (O_248,N_24786,N_23479);
nand UO_249 (O_249,N_23179,N_21631);
xnor UO_250 (O_250,N_21268,N_22647);
nor UO_251 (O_251,N_19029,N_19257);
and UO_252 (O_252,N_20264,N_24165);
xor UO_253 (O_253,N_21123,N_21751);
and UO_254 (O_254,N_20958,N_23375);
nor UO_255 (O_255,N_18833,N_23859);
nand UO_256 (O_256,N_19443,N_22995);
nand UO_257 (O_257,N_20065,N_21563);
or UO_258 (O_258,N_23315,N_23809);
xor UO_259 (O_259,N_19488,N_19305);
and UO_260 (O_260,N_24153,N_18974);
nand UO_261 (O_261,N_24302,N_23251);
or UO_262 (O_262,N_21519,N_22680);
xnor UO_263 (O_263,N_22338,N_21632);
and UO_264 (O_264,N_22879,N_19538);
or UO_265 (O_265,N_22402,N_24310);
or UO_266 (O_266,N_24063,N_20547);
xnor UO_267 (O_267,N_23892,N_19008);
xnor UO_268 (O_268,N_19619,N_20825);
and UO_269 (O_269,N_19376,N_21488);
and UO_270 (O_270,N_20009,N_24123);
nand UO_271 (O_271,N_23140,N_24236);
nand UO_272 (O_272,N_23671,N_19592);
or UO_273 (O_273,N_24609,N_19650);
xnor UO_274 (O_274,N_21990,N_21176);
and UO_275 (O_275,N_22614,N_20732);
nor UO_276 (O_276,N_23684,N_24525);
xor UO_277 (O_277,N_22303,N_22185);
or UO_278 (O_278,N_22258,N_24158);
nor UO_279 (O_279,N_19932,N_19930);
nor UO_280 (O_280,N_21758,N_19523);
nand UO_281 (O_281,N_24116,N_23393);
and UO_282 (O_282,N_24245,N_24362);
nand UO_283 (O_283,N_23609,N_23222);
xnor UO_284 (O_284,N_21879,N_18856);
and UO_285 (O_285,N_21787,N_19496);
xor UO_286 (O_286,N_20470,N_20308);
or UO_287 (O_287,N_19812,N_20134);
xnor UO_288 (O_288,N_19602,N_23356);
and UO_289 (O_289,N_23633,N_21183);
or UO_290 (O_290,N_23095,N_19183);
xnor UO_291 (O_291,N_20374,N_22327);
nor UO_292 (O_292,N_21801,N_21726);
nor UO_293 (O_293,N_24771,N_24071);
or UO_294 (O_294,N_21832,N_22571);
xnor UO_295 (O_295,N_23124,N_19664);
or UO_296 (O_296,N_21452,N_21484);
xor UO_297 (O_297,N_20935,N_24541);
or UO_298 (O_298,N_19053,N_20364);
xnor UO_299 (O_299,N_20653,N_22753);
and UO_300 (O_300,N_23219,N_23885);
xnor UO_301 (O_301,N_22317,N_19865);
nand UO_302 (O_302,N_23968,N_23102);
nand UO_303 (O_303,N_23637,N_22540);
xnor UO_304 (O_304,N_22407,N_24473);
or UO_305 (O_305,N_23342,N_21349);
xnor UO_306 (O_306,N_23592,N_22173);
nand UO_307 (O_307,N_20199,N_22582);
or UO_308 (O_308,N_18937,N_24600);
and UO_309 (O_309,N_24712,N_21987);
and UO_310 (O_310,N_21127,N_23740);
xor UO_311 (O_311,N_21300,N_19974);
or UO_312 (O_312,N_24918,N_24481);
nor UO_313 (O_313,N_24641,N_22557);
nand UO_314 (O_314,N_23279,N_23498);
xor UO_315 (O_315,N_23723,N_21555);
and UO_316 (O_316,N_22253,N_22991);
nor UO_317 (O_317,N_24717,N_19206);
nand UO_318 (O_318,N_24424,N_21174);
and UO_319 (O_319,N_22940,N_18789);
or UO_320 (O_320,N_22300,N_23893);
nand UO_321 (O_321,N_19776,N_24214);
and UO_322 (O_322,N_24711,N_22823);
or UO_323 (O_323,N_22871,N_22489);
nand UO_324 (O_324,N_18878,N_23751);
xnor UO_325 (O_325,N_20710,N_19722);
and UO_326 (O_326,N_19320,N_22117);
nor UO_327 (O_327,N_24239,N_18992);
nand UO_328 (O_328,N_22573,N_20143);
nand UO_329 (O_329,N_20375,N_24968);
nor UO_330 (O_330,N_19248,N_23326);
and UO_331 (O_331,N_24487,N_24227);
or UO_332 (O_332,N_24531,N_22307);
xnor UO_333 (O_333,N_21427,N_18934);
nor UO_334 (O_334,N_24169,N_20129);
xor UO_335 (O_335,N_23269,N_19521);
nor UO_336 (O_336,N_21024,N_19742);
nor UO_337 (O_337,N_19601,N_22717);
or UO_338 (O_338,N_19442,N_21189);
or UO_339 (O_339,N_24536,N_19823);
or UO_340 (O_340,N_24216,N_19294);
nor UO_341 (O_341,N_23246,N_21297);
and UO_342 (O_342,N_23668,N_21224);
nor UO_343 (O_343,N_23909,N_21267);
and UO_344 (O_344,N_24913,N_22834);
nor UO_345 (O_345,N_20535,N_20320);
or UO_346 (O_346,N_20440,N_20832);
xnor UO_347 (O_347,N_19325,N_24502);
nand UO_348 (O_348,N_20538,N_23852);
nand UO_349 (O_349,N_21035,N_23346);
nand UO_350 (O_350,N_20580,N_23069);
nor UO_351 (O_351,N_19164,N_22828);
or UO_352 (O_352,N_19131,N_20936);
or UO_353 (O_353,N_22422,N_19586);
or UO_354 (O_354,N_24097,N_24974);
and UO_355 (O_355,N_22028,N_19277);
or UO_356 (O_356,N_22900,N_21082);
and UO_357 (O_357,N_21917,N_20522);
xor UO_358 (O_358,N_20248,N_22390);
and UO_359 (O_359,N_22695,N_19009);
xor UO_360 (O_360,N_23357,N_20781);
and UO_361 (O_361,N_20873,N_20201);
or UO_362 (O_362,N_22209,N_23182);
nand UO_363 (O_363,N_21443,N_20062);
xnor UO_364 (O_364,N_23037,N_24985);
or UO_365 (O_365,N_24822,N_22936);
and UO_366 (O_366,N_23153,N_21668);
xnor UO_367 (O_367,N_23470,N_19110);
or UO_368 (O_368,N_20084,N_22648);
or UO_369 (O_369,N_21871,N_24560);
and UO_370 (O_370,N_24185,N_19683);
or UO_371 (O_371,N_22783,N_23417);
or UO_372 (O_372,N_23391,N_18908);
or UO_373 (O_373,N_22152,N_22070);
nor UO_374 (O_374,N_22466,N_19322);
and UO_375 (O_375,N_20544,N_22174);
nor UO_376 (O_376,N_20562,N_20981);
nand UO_377 (O_377,N_22325,N_23672);
or UO_378 (O_378,N_23420,N_23819);
and UO_379 (O_379,N_24327,N_23020);
xor UO_380 (O_380,N_20412,N_19736);
nor UO_381 (O_381,N_19168,N_19691);
nor UO_382 (O_382,N_19105,N_24925);
or UO_383 (O_383,N_21187,N_23497);
nand UO_384 (O_384,N_23482,N_23587);
nor UO_385 (O_385,N_20693,N_20344);
nor UO_386 (O_386,N_18923,N_20837);
or UO_387 (O_387,N_22385,N_23709);
nand UO_388 (O_388,N_22137,N_24209);
nor UO_389 (O_389,N_21781,N_21836);
xnor UO_390 (O_390,N_19587,N_22699);
and UO_391 (O_391,N_23334,N_20038);
nand UO_392 (O_392,N_20110,N_23242);
or UO_393 (O_393,N_20896,N_21020);
xnor UO_394 (O_394,N_20763,N_23973);
nand UO_395 (O_395,N_24666,N_21587);
and UO_396 (O_396,N_24709,N_24276);
and UO_397 (O_397,N_19616,N_24309);
and UO_398 (O_398,N_18807,N_23074);
nor UO_399 (O_399,N_23270,N_19375);
nor UO_400 (O_400,N_20776,N_23006);
nor UO_401 (O_401,N_20365,N_23111);
or UO_402 (O_402,N_21114,N_19517);
or UO_403 (O_403,N_20255,N_18965);
xnor UO_404 (O_404,N_19173,N_22359);
or UO_405 (O_405,N_24244,N_22721);
xor UO_406 (O_406,N_21146,N_18766);
or UO_407 (O_407,N_21141,N_21687);
nand UO_408 (O_408,N_20623,N_21457);
and UO_409 (O_409,N_20677,N_23519);
xnor UO_410 (O_410,N_20473,N_24059);
and UO_411 (O_411,N_18911,N_22741);
nand UO_412 (O_412,N_20471,N_23419);
nand UO_413 (O_413,N_20424,N_20597);
nor UO_414 (O_414,N_22725,N_22589);
nand UO_415 (O_415,N_20325,N_19681);
xor UO_416 (O_416,N_24544,N_23007);
xnor UO_417 (O_417,N_19374,N_18850);
xor UO_418 (O_418,N_22962,N_24503);
nor UO_419 (O_419,N_24367,N_18968);
or UO_420 (O_420,N_22514,N_22469);
nor UO_421 (O_421,N_23068,N_20486);
and UO_422 (O_422,N_21299,N_22888);
nand UO_423 (O_423,N_23550,N_19472);
nor UO_424 (O_424,N_24943,N_22673);
nand UO_425 (O_425,N_23344,N_22752);
xor UO_426 (O_426,N_21381,N_22012);
nor UO_427 (O_427,N_24515,N_19450);
or UO_428 (O_428,N_22382,N_22318);
and UO_429 (O_429,N_23481,N_20770);
nand UO_430 (O_430,N_23667,N_20019);
nor UO_431 (O_431,N_22662,N_20551);
nor UO_432 (O_432,N_24548,N_24472);
xor UO_433 (O_433,N_23989,N_22651);
or UO_434 (O_434,N_24942,N_22486);
or UO_435 (O_435,N_21021,N_24851);
xnor UO_436 (O_436,N_22286,N_20531);
xnor UO_437 (O_437,N_20133,N_19825);
xor UO_438 (O_438,N_21686,N_22284);
or UO_439 (O_439,N_23561,N_23706);
xnor UO_440 (O_440,N_24713,N_19635);
and UO_441 (O_441,N_24181,N_23285);
nor UO_442 (O_442,N_23588,N_23252);
or UO_443 (O_443,N_22110,N_22772);
nor UO_444 (O_444,N_20790,N_22572);
nor UO_445 (O_445,N_21822,N_20705);
or UO_446 (O_446,N_19296,N_22740);
nand UO_447 (O_447,N_20679,N_19253);
or UO_448 (O_448,N_23129,N_19617);
nand UO_449 (O_449,N_24635,N_22355);
xnor UO_450 (O_450,N_21111,N_22426);
and UO_451 (O_451,N_23737,N_24891);
and UO_452 (O_452,N_20330,N_20871);
and UO_453 (O_453,N_20109,N_23653);
and UO_454 (O_454,N_21557,N_20050);
and UO_455 (O_455,N_23778,N_20210);
nor UO_456 (O_456,N_19464,N_20479);
nor UO_457 (O_457,N_20571,N_24828);
nor UO_458 (O_458,N_21558,N_20229);
xnor UO_459 (O_459,N_22377,N_19814);
and UO_460 (O_460,N_24170,N_19806);
nand UO_461 (O_461,N_23422,N_20132);
nand UO_462 (O_462,N_19580,N_18913);
or UO_463 (O_463,N_22749,N_22696);
nor UO_464 (O_464,N_22984,N_21261);
nor UO_465 (O_465,N_24180,N_21579);
nand UO_466 (O_466,N_20456,N_18993);
nand UO_467 (O_467,N_22344,N_19493);
and UO_468 (O_468,N_21106,N_18765);
xnor UO_469 (O_469,N_22162,N_22366);
or UO_470 (O_470,N_19332,N_21277);
and UO_471 (O_471,N_20636,N_22646);
nor UO_472 (O_472,N_19153,N_19882);
nor UO_473 (O_473,N_22496,N_23213);
nand UO_474 (O_474,N_21063,N_23434);
or UO_475 (O_475,N_23012,N_20155);
or UO_476 (O_476,N_19666,N_22835);
nor UO_477 (O_477,N_18824,N_23679);
nand UO_478 (O_478,N_22658,N_22755);
or UO_479 (O_479,N_23954,N_19588);
nand UO_480 (O_480,N_22035,N_23043);
or UO_481 (O_481,N_18845,N_21264);
nand UO_482 (O_482,N_22690,N_20574);
nand UO_483 (O_483,N_24745,N_19978);
nand UO_484 (O_484,N_18960,N_22095);
and UO_485 (O_485,N_20439,N_24002);
xor UO_486 (O_486,N_19804,N_20596);
and UO_487 (O_487,N_24118,N_22931);
or UO_488 (O_488,N_24897,N_20835);
and UO_489 (O_489,N_24077,N_20616);
nor UO_490 (O_490,N_22508,N_21882);
nor UO_491 (O_491,N_19936,N_20261);
nor UO_492 (O_492,N_20406,N_22837);
nor UO_493 (O_493,N_18976,N_21645);
or UO_494 (O_494,N_23586,N_24603);
or UO_495 (O_495,N_24331,N_21025);
or UO_496 (O_496,N_23829,N_23322);
or UO_497 (O_497,N_24970,N_24762);
xnor UO_498 (O_498,N_20310,N_19585);
and UO_499 (O_499,N_24623,N_22683);
nand UO_500 (O_500,N_21837,N_19667);
xnor UO_501 (O_501,N_24317,N_19096);
xor UO_502 (O_502,N_24371,N_24094);
xnor UO_503 (O_503,N_21156,N_22290);
nand UO_504 (O_504,N_19893,N_19757);
or UO_505 (O_505,N_20818,N_21003);
nor UO_506 (O_506,N_24446,N_20711);
nor UO_507 (O_507,N_22779,N_21041);
and UO_508 (O_508,N_21468,N_20652);
nor UO_509 (O_509,N_19591,N_24601);
nor UO_510 (O_510,N_22519,N_19249);
nor UO_511 (O_511,N_24333,N_22665);
xnor UO_512 (O_512,N_22961,N_24184);
nor UO_513 (O_513,N_19710,N_22639);
nand UO_514 (O_514,N_23923,N_23217);
xnor UO_515 (O_515,N_21592,N_21353);
xor UO_516 (O_516,N_24735,N_19122);
and UO_517 (O_517,N_19200,N_20485);
nor UO_518 (O_518,N_21993,N_21680);
or UO_519 (O_519,N_21108,N_20560);
and UO_520 (O_520,N_24485,N_24674);
nand UO_521 (O_521,N_21074,N_23268);
and UO_522 (O_522,N_20077,N_19896);
nor UO_523 (O_523,N_20015,N_19660);
and UO_524 (O_524,N_23683,N_22853);
nand UO_525 (O_525,N_22334,N_18788);
and UO_526 (O_526,N_20508,N_20866);
or UO_527 (O_527,N_21662,N_21593);
xnor UO_528 (O_528,N_22802,N_23860);
or UO_529 (O_529,N_21691,N_18842);
nor UO_530 (O_530,N_20916,N_24756);
and UO_531 (O_531,N_18777,N_23943);
or UO_532 (O_532,N_22138,N_22010);
xnor UO_533 (O_533,N_20864,N_19645);
nand UO_534 (O_534,N_19477,N_23501);
nand UO_535 (O_535,N_20893,N_21936);
nand UO_536 (O_536,N_20336,N_22884);
xor UO_537 (O_537,N_24358,N_22438);
or UO_538 (O_538,N_21388,N_21002);
and UO_539 (O_539,N_19801,N_20459);
or UO_540 (O_540,N_24779,N_21157);
or UO_541 (O_541,N_24564,N_22886);
nor UO_542 (O_542,N_21234,N_21046);
or UO_543 (O_543,N_21571,N_24625);
nand UO_544 (O_544,N_23049,N_23527);
nand UO_545 (O_545,N_23638,N_20335);
or UO_546 (O_546,N_20158,N_20096);
or UO_547 (O_547,N_20662,N_24457);
and UO_548 (O_548,N_20606,N_22758);
and UO_549 (O_549,N_22930,N_19036);
nor UO_550 (O_550,N_20738,N_24308);
or UO_551 (O_551,N_24025,N_21066);
nand UO_552 (O_552,N_23639,N_21184);
or UO_553 (O_553,N_20668,N_22993);
nand UO_554 (O_554,N_23801,N_18944);
or UO_555 (O_555,N_22100,N_21278);
or UO_556 (O_556,N_20150,N_21453);
or UO_557 (O_557,N_21682,N_23214);
nor UO_558 (O_558,N_21461,N_20085);
and UO_559 (O_559,N_22291,N_23415);
xor UO_560 (O_560,N_20124,N_24592);
xor UO_561 (O_561,N_21681,N_24837);
xnor UO_562 (O_562,N_23403,N_24556);
nand UO_563 (O_563,N_19184,N_20103);
nor UO_564 (O_564,N_19261,N_20919);
nor UO_565 (O_565,N_24932,N_21233);
nand UO_566 (O_566,N_21357,N_20285);
and UO_567 (O_567,N_23312,N_20627);
and UO_568 (O_568,N_18950,N_23756);
nand UO_569 (O_569,N_23590,N_23247);
xnor UO_570 (O_570,N_22064,N_24012);
and UO_571 (O_571,N_19711,N_21899);
nor UO_572 (O_572,N_22467,N_22957);
or UO_573 (O_573,N_19352,N_19419);
nor UO_574 (O_574,N_21507,N_24896);
nor UO_575 (O_575,N_24476,N_24785);
and UO_576 (O_576,N_21878,N_19649);
nor UO_577 (O_577,N_21754,N_21870);
xor UO_578 (O_578,N_24937,N_19473);
xor UO_579 (O_579,N_22075,N_19423);
or UO_580 (O_580,N_24223,N_21414);
and UO_581 (O_581,N_24334,N_22259);
or UO_582 (O_582,N_22094,N_19237);
nand UO_583 (O_583,N_21892,N_19429);
and UO_584 (O_584,N_24313,N_23496);
nor UO_585 (O_585,N_24017,N_19080);
and UO_586 (O_586,N_24127,N_23837);
xor UO_587 (O_587,N_22733,N_21016);
and UO_588 (O_588,N_19178,N_24098);
nand UO_589 (O_589,N_21505,N_19644);
or UO_590 (O_590,N_20206,N_24606);
and UO_591 (O_591,N_24687,N_20829);
nand UO_592 (O_592,N_23597,N_19623);
and UO_593 (O_593,N_19424,N_21338);
nand UO_594 (O_594,N_23378,N_21697);
nand UO_595 (O_595,N_21677,N_23963);
and UO_596 (O_596,N_22672,N_20912);
or UO_597 (O_597,N_21707,N_19437);
or UO_598 (O_598,N_20315,N_19947);
or UO_599 (O_599,N_20833,N_24795);
xor UO_600 (O_600,N_20277,N_20235);
nor UO_601 (O_601,N_19963,N_19004);
or UO_602 (O_602,N_23557,N_23538);
or UO_603 (O_603,N_20372,N_22860);
xnor UO_604 (O_604,N_24277,N_21411);
nand UO_605 (O_605,N_22419,N_19765);
and UO_606 (O_606,N_23890,N_20174);
nand UO_607 (O_607,N_21659,N_21522);
nand UO_608 (O_608,N_20505,N_22023);
nor UO_609 (O_609,N_20639,N_20957);
xor UO_610 (O_610,N_24215,N_23634);
or UO_611 (O_611,N_20012,N_23583);
xor UO_612 (O_612,N_21616,N_21005);
xnor UO_613 (O_613,N_23071,N_23461);
xor UO_614 (O_614,N_21834,N_22208);
and UO_615 (O_615,N_23872,N_19394);
or UO_616 (O_616,N_22275,N_19377);
xor UO_617 (O_617,N_18755,N_24703);
or UO_618 (O_618,N_21308,N_23185);
nor UO_619 (O_619,N_21086,N_23674);
xor UO_620 (O_620,N_20069,N_20988);
xnor UO_621 (O_621,N_23052,N_23521);
or UO_622 (O_622,N_19965,N_20796);
or UO_623 (O_623,N_19467,N_22298);
or UO_624 (O_624,N_20400,N_24363);
nand UO_625 (O_625,N_23458,N_23894);
nor UO_626 (O_626,N_19949,N_21845);
xnor UO_627 (O_627,N_20076,N_19457);
and UO_628 (O_628,N_21354,N_24730);
xor UO_629 (O_629,N_22048,N_24408);
xnor UO_630 (O_630,N_23769,N_23645);
or UO_631 (O_631,N_24020,N_23385);
nand UO_632 (O_632,N_21026,N_22457);
and UO_633 (O_633,N_20903,N_24788);
or UO_634 (O_634,N_22370,N_22785);
or UO_635 (O_635,N_24962,N_24742);
xnor UO_636 (O_636,N_19072,N_20986);
or UO_637 (O_637,N_24945,N_21075);
nand UO_638 (O_638,N_18818,N_23460);
xor UO_639 (O_639,N_19392,N_23301);
and UO_640 (O_640,N_22304,N_19803);
or UO_641 (O_641,N_19014,N_21445);
nand UO_642 (O_642,N_24024,N_23551);
and UO_643 (O_643,N_22045,N_19571);
nand UO_644 (O_644,N_22270,N_24005);
and UO_645 (O_645,N_23526,N_23624);
xnor UO_646 (O_646,N_23388,N_20523);
and UO_647 (O_647,N_24526,N_23746);
nand UO_648 (O_648,N_22411,N_20217);
and UO_649 (O_649,N_24722,N_23985);
and UO_650 (O_650,N_23858,N_21050);
and UO_651 (O_651,N_24877,N_20013);
nor UO_652 (O_652,N_24954,N_23221);
or UO_653 (O_653,N_20022,N_24946);
nand UO_654 (O_654,N_24880,N_19844);
xor UO_655 (O_655,N_23028,N_19598);
xnor UO_656 (O_656,N_21618,N_23341);
and UO_657 (O_657,N_20197,N_21544);
or UO_658 (O_658,N_22821,N_22849);
or UO_659 (O_659,N_22922,N_24866);
nand UO_660 (O_660,N_19605,N_23721);
nand UO_661 (O_661,N_21569,N_24643);
xnor UO_662 (O_662,N_20690,N_21514);
xnor UO_663 (O_663,N_22156,N_18836);
nor UO_664 (O_664,N_22596,N_20442);
or UO_665 (O_665,N_21281,N_21436);
xor UO_666 (O_666,N_20901,N_23772);
nand UO_667 (O_667,N_19408,N_20391);
xnor UO_668 (O_668,N_24619,N_22047);
or UO_669 (O_669,N_23106,N_21192);
xnor UO_670 (O_670,N_22401,N_24350);
xnor UO_671 (O_671,N_19098,N_22492);
and UO_672 (O_672,N_23995,N_24610);
nor UO_673 (O_673,N_23386,N_19695);
or UO_674 (O_674,N_21883,N_19732);
or UO_675 (O_675,N_19285,N_19448);
and UO_676 (O_676,N_19211,N_24238);
xnor UO_677 (O_677,N_19479,N_21283);
xnor UO_678 (O_678,N_21417,N_21092);
xor UO_679 (O_679,N_19858,N_21038);
or UO_680 (O_680,N_22509,N_24781);
or UO_681 (O_681,N_18770,N_23659);
and UO_682 (O_682,N_24732,N_21595);
or UO_683 (O_683,N_19676,N_24489);
xnor UO_684 (O_684,N_23146,N_23436);
or UO_685 (O_685,N_18912,N_21511);
or UO_686 (O_686,N_19328,N_23438);
and UO_687 (O_687,N_22759,N_19315);
and UO_688 (O_688,N_19010,N_23361);
nor UO_689 (O_689,N_20107,N_18771);
nand UO_690 (O_690,N_22533,N_21780);
nand UO_691 (O_691,N_23313,N_20208);
or UO_692 (O_692,N_24591,N_20180);
xor UO_693 (O_693,N_23990,N_24022);
xor UO_694 (O_694,N_18890,N_21862);
nor UO_695 (O_695,N_24253,N_22480);
nor UO_696 (O_696,N_24959,N_21405);
xnor UO_697 (O_697,N_20650,N_21532);
and UO_698 (O_698,N_22630,N_24874);
nor UO_699 (O_699,N_22937,N_20480);
nor UO_700 (O_700,N_20469,N_23118);
nand UO_701 (O_701,N_21788,N_21364);
and UO_702 (O_702,N_24995,N_21732);
nand UO_703 (O_703,N_24311,N_22081);
nor UO_704 (O_704,N_23673,N_21191);
nor UO_705 (O_705,N_20079,N_19957);
nand UO_706 (O_706,N_23319,N_23072);
or UO_707 (O_707,N_22975,N_23666);
nand UO_708 (O_708,N_24865,N_22693);
or UO_709 (O_709,N_21116,N_20082);
xor UO_710 (O_710,N_22640,N_21554);
nor UO_711 (O_711,N_19378,N_20170);
nor UO_712 (O_712,N_18887,N_23399);
xnor UO_713 (O_713,N_22720,N_24341);
or UO_714 (O_714,N_22714,N_24144);
nor UO_715 (O_715,N_19017,N_20115);
xnor UO_716 (O_716,N_23310,N_20610);
xor UO_717 (O_717,N_23591,N_20474);
and UO_718 (O_718,N_19123,N_20941);
nor UO_719 (O_719,N_23412,N_21499);
nor UO_720 (O_720,N_23613,N_21545);
xor UO_721 (O_721,N_19003,N_19409);
nor UO_722 (O_722,N_23949,N_21348);
nand UO_723 (O_723,N_19212,N_20801);
nand UO_724 (O_724,N_19435,N_21729);
xor UO_725 (O_725,N_19684,N_19701);
xor UO_726 (O_726,N_20074,N_20080);
nand UO_727 (O_727,N_21084,N_23433);
nor UO_728 (O_728,N_23845,N_18998);
nor UO_729 (O_729,N_22512,N_23542);
nand UO_730 (O_730,N_19077,N_20033);
and UO_731 (O_731,N_22669,N_20006);
nor UO_732 (O_732,N_20269,N_19465);
or UO_733 (O_733,N_24765,N_23477);
and UO_734 (O_734,N_24175,N_23256);
xnor UO_735 (O_735,N_21389,N_19441);
or UO_736 (O_736,N_20268,N_21347);
and UO_737 (O_737,N_20477,N_21916);
nor UO_738 (O_738,N_19547,N_19725);
nand UO_739 (O_739,N_21247,N_22336);
xor UO_740 (O_740,N_24390,N_20671);
nand UO_741 (O_741,N_24114,N_20615);
xnor UO_742 (O_742,N_22038,N_23121);
nor UO_743 (O_743,N_24204,N_19867);
xor UO_744 (O_744,N_20305,N_21213);
nand UO_745 (O_745,N_21226,N_24840);
nand UO_746 (O_746,N_20756,N_24566);
and UO_747 (O_747,N_20068,N_23732);
or UO_748 (O_748,N_21573,N_24930);
and UO_749 (O_749,N_23870,N_23295);
and UO_750 (O_750,N_24076,N_22848);
nand UO_751 (O_751,N_19541,N_20585);
or UO_752 (O_752,N_20600,N_21927);
nor UO_753 (O_753,N_24186,N_21670);
nor UO_754 (O_754,N_21255,N_24028);
nand UO_755 (O_755,N_21236,N_20702);
or UO_756 (O_756,N_22408,N_24561);
xor UO_757 (O_757,N_24189,N_19786);
nor UO_758 (O_758,N_22769,N_19079);
nor UO_759 (O_759,N_22340,N_19875);
or UO_760 (O_760,N_20729,N_24728);
nand UO_761 (O_761,N_19883,N_24369);
or UO_762 (O_762,N_22999,N_19749);
nand UO_763 (O_763,N_19922,N_24876);
xor UO_764 (O_764,N_23863,N_23064);
nor UO_765 (O_765,N_22463,N_21815);
and UO_766 (O_766,N_23194,N_24938);
or UO_767 (O_767,N_21853,N_20991);
or UO_768 (O_768,N_19245,N_21679);
or UO_769 (O_769,N_24449,N_20141);
nand UO_770 (O_770,N_22960,N_21286);
and UO_771 (O_771,N_22800,N_19233);
or UO_772 (O_772,N_19572,N_20667);
or UO_773 (O_773,N_24815,N_20127);
and UO_774 (O_774,N_24431,N_19846);
and UO_775 (O_775,N_24247,N_21676);
and UO_776 (O_776,N_23716,N_18889);
nand UO_777 (O_777,N_19549,N_24988);
nand UO_778 (O_778,N_22967,N_24057);
xor UO_779 (O_779,N_23282,N_21830);
and UO_780 (O_780,N_23241,N_23082);
nor UO_781 (O_781,N_18843,N_19848);
xor UO_782 (O_782,N_24043,N_21186);
xor UO_783 (O_783,N_23339,N_23956);
nand UO_784 (O_784,N_22175,N_21506);
nand UO_785 (O_785,N_24766,N_23215);
nand UO_786 (O_786,N_24667,N_23321);
or UO_787 (O_787,N_19758,N_24651);
or UO_788 (O_788,N_24774,N_24381);
and UO_789 (O_789,N_20520,N_21517);
nand UO_790 (O_790,N_20165,N_19905);
and UO_791 (O_791,N_24151,N_23752);
or UO_792 (O_792,N_21045,N_21122);
or UO_793 (O_793,N_20302,N_20517);
or UO_794 (O_794,N_23895,N_21901);
xor UO_795 (O_795,N_23585,N_20447);
nor UO_796 (O_796,N_20094,N_19270);
and UO_797 (O_797,N_23042,N_24255);
xor UO_798 (O_798,N_21928,N_19810);
and UO_799 (O_799,N_21044,N_19620);
and UO_800 (O_800,N_22210,N_22536);
nor UO_801 (O_801,N_20880,N_24770);
xor UO_802 (O_802,N_22932,N_19421);
or UO_803 (O_803,N_20583,N_23827);
xor UO_804 (O_804,N_23843,N_24755);
nand UO_805 (O_805,N_24099,N_24553);
nor UO_806 (O_806,N_21886,N_23166);
and UO_807 (O_807,N_21985,N_22655);
nor UO_808 (O_808,N_21027,N_22086);
xnor UO_809 (O_809,N_19800,N_20617);
xnor UO_810 (O_810,N_24504,N_18863);
nor UO_811 (O_811,N_21387,N_23418);
or UO_812 (O_812,N_20812,N_23902);
nand UO_813 (O_813,N_20484,N_18956);
or UO_814 (O_814,N_19950,N_19819);
nor UO_815 (O_815,N_23116,N_23760);
nor UO_816 (O_816,N_21340,N_21472);
nand UO_817 (O_817,N_18900,N_18943);
and UO_818 (O_818,N_18969,N_20577);
nor UO_819 (O_819,N_24578,N_23423);
nor UO_820 (O_820,N_20701,N_19346);
and UO_821 (O_821,N_22372,N_24557);
nand UO_822 (O_822,N_19447,N_19502);
nand UO_823 (O_823,N_21315,N_24412);
or UO_824 (O_824,N_20343,N_23472);
or UO_825 (O_825,N_21337,N_24168);
and UO_826 (O_826,N_22872,N_19192);
or UO_827 (O_827,N_18980,N_19781);
and UO_828 (O_828,N_23776,N_23701);
nor UO_829 (O_829,N_19514,N_22685);
nor UO_830 (O_830,N_21475,N_23058);
or UO_831 (O_831,N_23886,N_22109);
xor UO_832 (O_832,N_23964,N_24736);
and UO_833 (O_833,N_24680,N_21734);
nand UO_834 (O_834,N_21864,N_22148);
nand UO_835 (O_835,N_24103,N_20299);
nand UO_836 (O_836,N_24048,N_22580);
xnor UO_837 (O_837,N_20163,N_20301);
xnor UO_838 (O_838,N_18873,N_21896);
nor UO_839 (O_839,N_23904,N_21067);
xnor UO_840 (O_840,N_24488,N_22606);
nor UO_841 (O_841,N_20973,N_19929);
nand UO_842 (O_842,N_20984,N_20620);
or UO_843 (O_843,N_20824,N_18758);
nand UO_844 (O_844,N_20095,N_19995);
and UO_845 (O_845,N_20145,N_19536);
and UO_846 (O_846,N_22819,N_24861);
nor UO_847 (O_847,N_22062,N_23096);
nand UO_848 (O_848,N_24554,N_20892);
nor UO_849 (O_849,N_24414,N_22410);
or UO_850 (O_850,N_23950,N_21689);
nor UO_851 (O_851,N_19044,N_22956);
xnor UO_852 (O_852,N_19368,N_20826);
and UO_853 (O_853,N_19218,N_23786);
or UO_854 (O_854,N_24582,N_19302);
and UO_855 (O_855,N_22863,N_20581);
or UO_856 (O_856,N_21585,N_22968);
xnor UO_857 (O_857,N_21314,N_24383);
or UO_858 (O_858,N_24477,N_22432);
or UO_859 (O_859,N_22034,N_20717);
nand UO_860 (O_860,N_19915,N_19624);
xor UO_861 (O_861,N_22706,N_18917);
or UO_862 (O_862,N_18997,N_20188);
and UO_863 (O_863,N_20073,N_23733);
nand UO_864 (O_864,N_24507,N_24700);
and UO_865 (O_865,N_20026,N_21458);
and UO_866 (O_866,N_22927,N_24439);
nor UO_867 (O_867,N_19584,N_19530);
and UO_868 (O_868,N_18955,N_23136);
and UO_869 (O_869,N_21574,N_24343);
or UO_870 (O_870,N_21518,N_23262);
nor UO_871 (O_871,N_18971,N_20245);
nor UO_872 (O_872,N_20595,N_21765);
and UO_873 (O_873,N_19890,N_19030);
or UO_874 (O_874,N_21844,N_20806);
nor UO_875 (O_875,N_20676,N_22798);
nor UO_876 (O_876,N_18989,N_19527);
nor UO_877 (O_877,N_24329,N_18776);
or UO_878 (O_878,N_23926,N_24740);
nand UO_879 (O_879,N_20769,N_21395);
nor UO_880 (O_880,N_20153,N_19578);
nand UO_881 (O_881,N_21403,N_22249);
or UO_882 (O_882,N_19690,N_21947);
nor UO_883 (O_883,N_19657,N_24657);
and UO_884 (O_884,N_20779,N_23265);
xor UO_885 (O_885,N_24527,N_21102);
and UO_886 (O_886,N_22575,N_21193);
or UO_887 (O_887,N_21007,N_24484);
nor UO_888 (O_888,N_22159,N_23348);
nand UO_889 (O_889,N_19632,N_21565);
nor UO_890 (O_890,N_20950,N_23207);
nand UO_891 (O_891,N_23935,N_23696);
and UO_892 (O_892,N_24430,N_19094);
nand UO_893 (O_893,N_20187,N_24324);
nand UO_894 (O_894,N_21974,N_18879);
nand UO_895 (O_895,N_20695,N_22947);
nor UO_896 (O_896,N_20764,N_20931);
xnor UO_897 (O_897,N_24816,N_18948);
nor UO_898 (O_898,N_21178,N_24538);
nor UO_899 (O_899,N_24519,N_22490);
xor UO_900 (O_900,N_22398,N_21373);
xor UO_901 (O_901,N_22133,N_21150);
and UO_902 (O_902,N_23289,N_19216);
nor UO_903 (O_903,N_22181,N_22314);
nor UO_904 (O_904,N_20121,N_21132);
nor UO_905 (O_905,N_20834,N_22282);
and UO_906 (O_906,N_23744,N_24790);
nand UO_907 (O_907,N_22187,N_19537);
nor UO_908 (O_908,N_22564,N_19603);
nor UO_909 (O_909,N_24436,N_19528);
or UO_910 (O_910,N_23084,N_20246);
or UO_911 (O_911,N_23984,N_21313);
xnor UO_912 (O_912,N_23514,N_21438);
or UO_913 (O_913,N_19391,N_22256);
and UO_914 (O_914,N_21966,N_19871);
nor UO_915 (O_915,N_19693,N_21949);
xor UO_916 (O_916,N_22448,N_23790);
nor UO_917 (O_917,N_23180,N_23495);
or UO_918 (O_918,N_24989,N_24972);
nor UO_919 (O_919,N_22066,N_23307);
and UO_920 (O_920,N_19468,N_19853);
xor UO_921 (O_921,N_22132,N_21279);
nand UO_922 (O_922,N_23227,N_23449);
xor UO_923 (O_923,N_24055,N_24233);
nand UO_924 (O_924,N_21898,N_20113);
or UO_925 (O_925,N_24997,N_18782);
nand UO_926 (O_926,N_24620,N_18754);
and UO_927 (O_927,N_21071,N_21253);
nand UO_928 (O_928,N_21164,N_20850);
and UO_929 (O_929,N_22494,N_23952);
xnor UO_930 (O_930,N_22083,N_22387);
nand UO_931 (O_931,N_21502,N_18808);
and UO_932 (O_932,N_21635,N_20852);
nor UO_933 (O_933,N_20593,N_22566);
and UO_934 (O_934,N_19807,N_22039);
xor UO_935 (O_935,N_19916,N_22233);
xnor UO_936 (O_936,N_21269,N_19794);
nor UO_937 (O_937,N_22168,N_24178);
or UO_938 (O_938,N_21562,N_20014);
xor UO_939 (O_939,N_24219,N_24993);
and UO_940 (O_940,N_23311,N_22668);
nor UO_941 (O_941,N_20211,N_24939);
nand UO_942 (O_942,N_21553,N_23148);
xnor UO_943 (O_943,N_19445,N_21070);
or UO_944 (O_944,N_19276,N_20055);
or UO_945 (O_945,N_21752,N_19852);
nor UO_946 (O_946,N_20039,N_22225);
and UO_947 (O_947,N_21520,N_21265);
nand UO_948 (O_948,N_18867,N_22921);
nor UO_949 (O_949,N_20347,N_22439);
nand UO_950 (O_950,N_19921,N_21934);
or UO_951 (O_951,N_23755,N_19019);
or UO_952 (O_952,N_20644,N_23815);
xnor UO_953 (O_953,N_24407,N_22212);
xor UO_954 (O_954,N_23491,N_24268);
nand UO_955 (O_955,N_19596,N_18829);
or UO_956 (O_956,N_21702,N_24070);
and UO_957 (O_957,N_23630,N_19373);
nor UO_958 (O_958,N_22349,N_23836);
nand UO_959 (O_959,N_19777,N_19519);
or UO_960 (O_960,N_20476,N_23233);
and UO_961 (O_961,N_22025,N_20787);
nand UO_962 (O_962,N_20051,N_24193);
and UO_963 (O_963,N_23425,N_21200);
or UO_964 (O_964,N_21924,N_22654);
xor UO_965 (O_965,N_19764,N_19750);
or UO_966 (O_966,N_18835,N_22379);
nor UO_967 (O_967,N_21851,N_21133);
and UO_968 (O_968,N_23169,N_22363);
or UO_969 (O_969,N_20219,N_20098);
nand UO_970 (O_970,N_20232,N_22537);
xor UO_971 (O_971,N_21867,N_19469);
and UO_972 (O_972,N_24252,N_21407);
and UO_973 (O_973,N_24626,N_23913);
and UO_974 (O_974,N_20175,N_21341);
and UO_975 (O_975,N_22491,N_21449);
nor UO_976 (O_976,N_24498,N_24924);
or UO_977 (O_977,N_24973,N_21077);
or UO_978 (O_978,N_23781,N_24471);
nor UO_979 (O_979,N_23023,N_22715);
nor UO_980 (O_980,N_24266,N_22333);
or UO_981 (O_981,N_24029,N_24777);
xor UO_982 (O_982,N_23619,N_20353);
nor UO_983 (O_983,N_23631,N_22134);
nor UO_984 (O_984,N_24571,N_19515);
xor UO_985 (O_985,N_23288,N_23120);
nor UO_986 (O_986,N_22196,N_24250);
or UO_987 (O_987,N_20099,N_22194);
nor UO_988 (O_988,N_20766,N_22612);
and UO_989 (O_989,N_21602,N_22264);
and UO_990 (O_990,N_22565,N_19399);
and UO_991 (O_991,N_24119,N_21813);
or UO_992 (O_992,N_24796,N_22114);
nand UO_993 (O_993,N_24257,N_19863);
or UO_994 (O_994,N_19772,N_20377);
or UO_995 (O_995,N_22625,N_22051);
xor UO_996 (O_996,N_20540,N_19215);
nor UO_997 (O_997,N_23704,N_20848);
nor UO_998 (O_998,N_18881,N_24279);
nand UO_999 (O_999,N_24494,N_19885);
or UO_1000 (O_1000,N_21215,N_18907);
nand UO_1001 (O_1001,N_20977,N_24648);
or UO_1002 (O_1002,N_19522,N_19239);
nor UO_1003 (O_1003,N_21828,N_19763);
or UO_1004 (O_1004,N_19050,N_21245);
xor UO_1005 (O_1005,N_23799,N_21811);
and UO_1006 (O_1006,N_19719,N_24389);
nor UO_1007 (O_1007,N_24294,N_23831);
or UO_1008 (O_1008,N_19114,N_19180);
xnor UO_1009 (O_1009,N_23525,N_21607);
or UO_1010 (O_1010,N_21329,N_22232);
and UO_1011 (O_1011,N_22915,N_24747);
nand UO_1012 (O_1012,N_21921,N_19752);
nand UO_1013 (O_1013,N_18796,N_19709);
nor UO_1014 (O_1014,N_23038,N_24394);
nand UO_1015 (O_1015,N_22339,N_22709);
nand UO_1016 (O_1016,N_20126,N_23087);
and UO_1017 (O_1017,N_24887,N_21800);
xor UO_1018 (O_1018,N_22104,N_23925);
xnor UO_1019 (O_1019,N_23338,N_24148);
nor UO_1020 (O_1020,N_21295,N_20252);
xnor UO_1021 (O_1021,N_24614,N_19327);
nand UO_1022 (O_1022,N_21017,N_21970);
and UO_1023 (O_1023,N_18972,N_20854);
nand UO_1024 (O_1024,N_22004,N_18858);
and UO_1025 (O_1025,N_21775,N_19730);
nor UO_1026 (O_1026,N_23767,N_23431);
and UO_1027 (O_1027,N_20478,N_22420);
xor UO_1028 (O_1028,N_19702,N_20119);
xnor UO_1029 (O_1029,N_24570,N_23998);
nand UO_1030 (O_1030,N_20827,N_22925);
xnor UO_1031 (O_1031,N_24106,N_24342);
nor UO_1032 (O_1032,N_21989,N_18892);
and UO_1033 (O_1033,N_20510,N_21079);
or UO_1034 (O_1034,N_19051,N_19043);
nand UO_1035 (O_1035,N_18802,N_21292);
nor UO_1036 (O_1036,N_23377,N_23560);
nor UO_1037 (O_1037,N_24353,N_19985);
or UO_1038 (O_1038,N_24671,N_18762);
or UO_1039 (O_1039,N_19525,N_24456);
nor UO_1040 (O_1040,N_23283,N_20340);
xnor UO_1041 (O_1041,N_19265,N_23257);
and UO_1042 (O_1042,N_23364,N_23960);
nor UO_1043 (O_1043,N_22090,N_24352);
and UO_1044 (O_1044,N_20001,N_20911);
or UO_1045 (O_1045,N_24206,N_23605);
or UO_1046 (O_1046,N_22737,N_20225);
and UO_1047 (O_1047,N_24088,N_24998);
xnor UO_1048 (O_1048,N_20321,N_20546);
xnor UO_1049 (O_1049,N_21510,N_23443);
nor UO_1050 (O_1050,N_21637,N_19142);
nand UO_1051 (O_1051,N_18834,N_21408);
nand UO_1052 (O_1052,N_21818,N_21527);
and UO_1053 (O_1053,N_20382,N_24810);
nand UO_1054 (O_1054,N_21596,N_22547);
xor UO_1055 (O_1055,N_19126,N_22179);
or UO_1056 (O_1056,N_20982,N_22549);
nor UO_1057 (O_1057,N_19417,N_23818);
xnor UO_1058 (O_1058,N_23474,N_21792);
xor UO_1059 (O_1059,N_22851,N_18946);
nor UO_1060 (O_1060,N_21849,N_20663);
nor UO_1061 (O_1061,N_24034,N_24208);
and UO_1062 (O_1062,N_19532,N_21763);
and UO_1063 (O_1063,N_21298,N_18861);
nor UO_1064 (O_1064,N_23478,N_20432);
nand UO_1065 (O_1065,N_23779,N_19073);
xor UO_1066 (O_1066,N_21435,N_22734);
nor UO_1067 (O_1067,N_19411,N_22829);
xnor UO_1068 (O_1068,N_24195,N_21238);
nor UO_1069 (O_1069,N_21372,N_24373);
nand UO_1070 (O_1070,N_24467,N_20292);
or UO_1071 (O_1071,N_23359,N_22204);
nor UO_1072 (O_1072,N_22901,N_20909);
nor UO_1073 (O_1073,N_23547,N_24653);
xor UO_1074 (O_1074,N_20974,N_20645);
xor UO_1075 (O_1075,N_22358,N_19707);
and UO_1076 (O_1076,N_24616,N_20604);
or UO_1077 (O_1077,N_24461,N_24909);
nor UO_1078 (O_1078,N_23483,N_23170);
nand UO_1079 (O_1079,N_20122,N_23891);
and UO_1080 (O_1080,N_21019,N_18904);
and UO_1081 (O_1081,N_23421,N_22483);
and UO_1082 (O_1082,N_20405,N_24848);
and UO_1083 (O_1083,N_23405,N_19260);
nor UO_1084 (O_1084,N_23903,N_20847);
nand UO_1085 (O_1085,N_20169,N_23155);
or UO_1086 (O_1086,N_22431,N_24975);
and UO_1087 (O_1087,N_19563,N_20403);
nand UO_1088 (O_1088,N_22814,N_21235);
nor UO_1089 (O_1089,N_22394,N_20749);
xnor UO_1090 (O_1090,N_24642,N_23506);
xnor UO_1091 (O_1091,N_19127,N_20171);
or UO_1092 (O_1092,N_21933,N_22429);
nand UO_1093 (O_1093,N_18898,N_21561);
and UO_1094 (O_1094,N_19880,N_22058);
and UO_1095 (O_1095,N_23444,N_22621);
and UO_1096 (O_1096,N_20727,N_22531);
or UO_1097 (O_1097,N_20920,N_23029);
and UO_1098 (O_1098,N_21248,N_21287);
or UO_1099 (O_1099,N_20939,N_22056);
nand UO_1100 (O_1100,N_23874,N_19300);
nor UO_1101 (O_1101,N_20179,N_20139);
nand UO_1102 (O_1102,N_20280,N_23413);
nand UO_1103 (O_1103,N_19228,N_22442);
xnor UO_1104 (O_1104,N_24234,N_19780);
or UO_1105 (O_1105,N_22801,N_21366);
nor UO_1106 (O_1106,N_19000,N_20281);
and UO_1107 (O_1107,N_24332,N_22101);
nand UO_1108 (O_1108,N_19027,N_20841);
and UO_1109 (O_1109,N_18932,N_22084);
nand UO_1110 (O_1110,N_23416,N_23191);
xor UO_1111 (O_1111,N_22074,N_24441);
and UO_1112 (O_1112,N_20369,N_21638);
nor UO_1113 (O_1113,N_23176,N_24349);
nor UO_1114 (O_1114,N_23664,N_22841);
xor UO_1115 (O_1115,N_18885,N_23853);
nor UO_1116 (O_1116,N_22869,N_21712);
xnor UO_1117 (O_1117,N_20521,N_24994);
xnor UO_1118 (O_1118,N_24923,N_19881);
nor UO_1119 (O_1119,N_23523,N_23486);
nor UO_1120 (O_1120,N_23842,N_24589);
nor UO_1121 (O_1121,N_21542,N_22585);
or UO_1122 (O_1122,N_19349,N_21526);
xnor UO_1123 (O_1123,N_23152,N_20493);
xor UO_1124 (O_1124,N_24996,N_19746);
or UO_1125 (O_1125,N_21211,N_24718);
xor UO_1126 (O_1126,N_22726,N_18906);
or UO_1127 (O_1127,N_22428,N_19505);
nand UO_1128 (O_1128,N_22044,N_21393);
nor UO_1129 (O_1129,N_18995,N_22453);
nor UO_1130 (O_1130,N_18999,N_20184);
and UO_1131 (O_1131,N_22082,N_20791);
and UO_1132 (O_1132,N_23264,N_22375);
xnor UO_1133 (O_1133,N_23828,N_21675);
or UO_1134 (O_1134,N_20925,N_21604);
or UO_1135 (O_1135,N_19198,N_23376);
nand UO_1136 (O_1136,N_19231,N_19638);
and UO_1137 (O_1137,N_20244,N_18819);
and UO_1138 (O_1138,N_20943,N_21250);
nand UO_1139 (O_1139,N_22030,N_22724);
xor UO_1140 (O_1140,N_21209,N_21426);
and UO_1141 (O_1141,N_21523,N_20409);
nor UO_1142 (O_1142,N_23226,N_24145);
nand UO_1143 (O_1143,N_22273,N_21052);
nor UO_1144 (O_1144,N_20159,N_20397);
or UO_1145 (O_1145,N_20287,N_19546);
or UO_1146 (O_1146,N_19284,N_21487);
and UO_1147 (O_1147,N_20233,N_21422);
nand UO_1148 (O_1148,N_23505,N_20753);
nor UO_1149 (O_1149,N_23518,N_24171);
or UO_1150 (O_1150,N_24388,N_24892);
or UO_1151 (O_1151,N_19484,N_21240);
xor UO_1152 (O_1152,N_20956,N_20782);
xnor UO_1153 (O_1153,N_24534,N_20018);
and UO_1154 (O_1154,N_20249,N_22781);
and UO_1155 (O_1155,N_23138,N_20816);
or UO_1156 (O_1156,N_18838,N_20955);
and UO_1157 (O_1157,N_22988,N_24857);
nand UO_1158 (O_1158,N_20140,N_23759);
or UO_1159 (O_1159,N_21188,N_21658);
xnor UO_1160 (O_1160,N_22099,N_19912);
xor UO_1161 (O_1161,N_18927,N_24221);
nor UO_1162 (O_1162,N_21920,N_22831);
nand UO_1163 (O_1163,N_21643,N_22242);
xnor UO_1164 (O_1164,N_23272,N_19024);
and UO_1165 (O_1165,N_20785,N_21716);
nor UO_1166 (O_1166,N_22550,N_20657);
and UO_1167 (O_1167,N_20220,N_20436);
xnor UO_1168 (O_1168,N_19510,N_19130);
nand UO_1169 (O_1169,N_19093,N_23880);
nor UO_1170 (O_1170,N_20881,N_24621);
nand UO_1171 (O_1171,N_22641,N_19430);
nor UO_1172 (O_1172,N_21275,N_23203);
or UO_1173 (O_1173,N_19927,N_20994);
or UO_1174 (O_1174,N_23001,N_19551);
or UO_1175 (O_1175,N_22807,N_23318);
nand UO_1176 (O_1176,N_20462,N_24776);
xnor UO_1177 (O_1177,N_23618,N_19083);
or UO_1178 (O_1178,N_21594,N_20063);
nor UO_1179 (O_1179,N_19359,N_21566);
nand UO_1180 (O_1180,N_24510,N_20731);
nand UO_1181 (O_1181,N_22982,N_24940);
nand UO_1182 (O_1182,N_24161,N_23367);
and UO_1183 (O_1183,N_22913,N_24631);
nor UO_1184 (O_1184,N_22615,N_22306);
or UO_1185 (O_1185,N_21455,N_20963);
nand UO_1186 (O_1186,N_20260,N_22766);
xor UO_1187 (O_1187,N_21180,N_22719);
nand UO_1188 (O_1188,N_20708,N_21535);
nand UO_1189 (O_1189,N_24655,N_21693);
xor UO_1190 (O_1190,N_21959,N_21302);
xnor UO_1191 (O_1191,N_24241,N_23566);
nand UO_1192 (O_1192,N_21379,N_19809);
and UO_1193 (O_1193,N_23996,N_23615);
or UO_1194 (O_1194,N_23040,N_22858);
nor UO_1195 (O_1195,N_22331,N_23933);
nor UO_1196 (O_1196,N_22268,N_24288);
nand UO_1197 (O_1197,N_20359,N_22414);
or UO_1198 (O_1198,N_18837,N_20317);
or UO_1199 (O_1199,N_22476,N_24386);
nand UO_1200 (O_1200,N_18778,N_20706);
xnor UO_1201 (O_1201,N_20262,N_22729);
xor UO_1202 (O_1202,N_20185,N_21718);
or UO_1203 (O_1203,N_20609,N_22197);
nand UO_1204 (O_1204,N_23820,N_24920);
nor UO_1205 (O_1205,N_19459,N_24326);
and UO_1206 (O_1206,N_21599,N_22061);
and UO_1207 (O_1207,N_22434,N_19426);
or UO_1208 (O_1208,N_19313,N_21301);
nor UO_1209 (O_1209,N_22745,N_23797);
xor UO_1210 (O_1210,N_24495,N_23143);
or UO_1211 (O_1211,N_23675,N_23838);
xor UO_1212 (O_1212,N_23901,N_24969);
or UO_1213 (O_1213,N_19652,N_21979);
nand UO_1214 (O_1214,N_23384,N_21241);
nand UO_1215 (O_1215,N_23932,N_21796);
nand UO_1216 (O_1216,N_20843,N_21644);
nand UO_1217 (O_1217,N_19267,N_22838);
xnor UO_1218 (O_1218,N_23515,N_23016);
nand UO_1219 (O_1219,N_22369,N_18828);
nor UO_1220 (O_1220,N_20144,N_22705);
nand UO_1221 (O_1221,N_19062,N_21730);
or UO_1222 (O_1222,N_21695,N_18864);
nor UO_1223 (O_1223,N_19242,N_22526);
or UO_1224 (O_1224,N_21723,N_21983);
or UO_1225 (O_1225,N_20037,N_24190);
nor UO_1226 (O_1226,N_21386,N_22343);
nor UO_1227 (O_1227,N_24921,N_21055);
and UO_1228 (O_1228,N_24915,N_22896);
nor UO_1229 (O_1229,N_20709,N_20318);
nand UO_1230 (O_1230,N_23184,N_19960);
xor UO_1231 (O_1231,N_19119,N_20745);
nor UO_1232 (O_1232,N_20603,N_21260);
and UO_1233 (O_1233,N_19851,N_20998);
nor UO_1234 (O_1234,N_21816,N_18852);
and UO_1235 (O_1235,N_24267,N_23372);
or UO_1236 (O_1236,N_21477,N_20023);
nand UO_1237 (O_1237,N_22650,N_23868);
nor UO_1238 (O_1238,N_20611,N_19039);
xnor UO_1239 (O_1239,N_18977,N_20205);
nand UO_1240 (O_1240,N_19941,N_23186);
nor UO_1241 (O_1241,N_21220,N_24907);
or UO_1242 (O_1242,N_21331,N_19095);
nand UO_1243 (O_1243,N_23517,N_21319);
nor UO_1244 (O_1244,N_23939,N_23112);
nand UO_1245 (O_1245,N_21034,N_23374);
nand UO_1246 (O_1246,N_23480,N_22645);
and UO_1247 (O_1247,N_24085,N_22671);
xor UO_1248 (O_1248,N_22072,N_21946);
and UO_1249 (O_1249,N_18841,N_19874);
nor UO_1250 (O_1250,N_22451,N_24112);
xor UO_1251 (O_1251,N_23232,N_23817);
xor UO_1252 (O_1252,N_23456,N_19400);
and UO_1253 (O_1253,N_18938,N_23465);
nand UO_1254 (O_1254,N_24862,N_22180);
xnor UO_1255 (O_1255,N_24149,N_19544);
or UO_1256 (O_1256,N_21181,N_23195);
nor UO_1257 (O_1257,N_20579,N_23455);
nand UO_1258 (O_1258,N_21722,N_20300);
nor UO_1259 (O_1259,N_19169,N_19864);
and UO_1260 (O_1260,N_21303,N_19543);
nor UO_1261 (O_1261,N_21713,N_22261);
nand UO_1262 (O_1262,N_22546,N_23536);
and UO_1263 (O_1263,N_22329,N_20276);
and UO_1264 (O_1264,N_20041,N_21100);
nand UO_1265 (O_1265,N_22812,N_24400);
nor UO_1266 (O_1266,N_20227,N_20550);
or UO_1267 (O_1267,N_20542,N_22381);
and UO_1268 (O_1268,N_19329,N_24832);
and UO_1269 (O_1269,N_23305,N_19508);
xnor UO_1270 (O_1270,N_19822,N_22545);
and UO_1271 (O_1271,N_19193,N_19055);
xor UO_1272 (O_1272,N_23439,N_20061);
or UO_1273 (O_1273,N_19630,N_19942);
and UO_1274 (O_1274,N_24087,N_23336);
and UO_1275 (O_1275,N_19224,N_19877);
xnor UO_1276 (O_1276,N_22295,N_22485);
nand UO_1277 (O_1277,N_22865,N_20648);
or UO_1278 (O_1278,N_22525,N_19983);
and UO_1279 (O_1279,N_24320,N_21296);
or UO_1280 (O_1280,N_23382,N_24003);
and UO_1281 (O_1281,N_22929,N_24200);
nor UO_1282 (O_1282,N_21054,N_23165);
nand UO_1283 (O_1283,N_24458,N_19975);
nor UO_1284 (O_1284,N_19656,N_23154);
xnor UO_1285 (O_1285,N_24177,N_18935);
and UO_1286 (O_1286,N_18899,N_23022);
and UO_1287 (O_1287,N_23596,N_24049);
and UO_1288 (O_1288,N_20539,N_21113);
nand UO_1289 (O_1289,N_19717,N_22803);
and UO_1290 (O_1290,N_24792,N_20557);
and UO_1291 (O_1291,N_19312,N_22102);
nand UO_1292 (O_1292,N_22165,N_19988);
nand UO_1293 (O_1293,N_21784,N_21493);
nor UO_1294 (O_1294,N_24243,N_23691);
or UO_1295 (O_1295,N_21190,N_23002);
or UO_1296 (O_1296,N_23383,N_22356);
and UO_1297 (O_1297,N_19463,N_24522);
nor UO_1298 (O_1298,N_22813,N_20803);
nor UO_1299 (O_1299,N_24427,N_23015);
nand UO_1300 (O_1300,N_20467,N_22143);
xor UO_1301 (O_1301,N_20324,N_22057);
or UO_1302 (O_1302,N_24708,N_23844);
nand UO_1303 (O_1303,N_24281,N_24051);
nor UO_1304 (O_1304,N_24415,N_22788);
nand UO_1305 (O_1305,N_22308,N_22633);
nor UO_1306 (O_1306,N_18985,N_21939);
xnor UO_1307 (O_1307,N_24124,N_20327);
nor UO_1308 (O_1308,N_22471,N_19685);
nand UO_1309 (O_1309,N_22498,N_20100);
nand UO_1310 (O_1310,N_22949,N_24899);
and UO_1311 (O_1311,N_24660,N_19579);
nor UO_1312 (O_1312,N_20890,N_21463);
or UO_1313 (O_1313,N_24251,N_19132);
or UO_1314 (O_1314,N_19161,N_21374);
or UO_1315 (O_1315,N_23725,N_20563);
and UO_1316 (O_1316,N_24611,N_22599);
nor UO_1317 (O_1317,N_18823,N_23718);
nor UO_1318 (O_1318,N_21433,N_20800);
xor UO_1319 (O_1319,N_18750,N_21809);
nor UO_1320 (O_1320,N_23775,N_24729);
nor UO_1321 (O_1321,N_22323,N_19340);
nand UO_1322 (O_1322,N_18886,N_22878);
nand UO_1323 (O_1323,N_21634,N_21590);
or UO_1324 (O_1324,N_19860,N_20605);
and UO_1325 (O_1325,N_23652,N_19148);
or UO_1326 (O_1326,N_23934,N_19737);
or UO_1327 (O_1327,N_24726,N_23063);
or UO_1328 (O_1328,N_19227,N_22437);
nand UO_1329 (O_1329,N_23573,N_24174);
or UO_1330 (O_1330,N_20914,N_24305);
and UO_1331 (O_1331,N_22315,N_22707);
nor UO_1332 (O_1332,N_19903,N_20195);
xor UO_1333 (O_1333,N_24120,N_19494);
or UO_1334 (O_1334,N_21115,N_21888);
nand UO_1335 (O_1335,N_22563,N_22855);
xor UO_1336 (O_1336,N_22918,N_20972);
and UO_1337 (O_1337,N_24807,N_22793);
xor UO_1338 (O_1338,N_23598,N_19937);
or UO_1339 (O_1339,N_22637,N_21464);
or UO_1340 (O_1340,N_23821,N_21152);
nand UO_1341 (O_1341,N_19733,N_22222);
nor UO_1342 (O_1342,N_20441,N_22678);
and UO_1343 (O_1343,N_18784,N_20937);
or UO_1344 (O_1344,N_23442,N_24568);
nor UO_1345 (O_1345,N_23061,N_23979);
and UO_1346 (O_1346,N_23848,N_19048);
xnor UO_1347 (O_1347,N_19567,N_20830);
and UO_1348 (O_1348,N_22423,N_23274);
or UO_1349 (O_1349,N_20498,N_22541);
nand UO_1350 (O_1350,N_20713,N_23178);
or UO_1351 (O_1351,N_24142,N_21536);
nor UO_1352 (O_1352,N_22368,N_19485);
xor UO_1353 (O_1353,N_19389,N_20497);
or UO_1354 (O_1354,N_24752,N_20874);
nand UO_1355 (O_1355,N_19321,N_18958);
xor UO_1356 (O_1356,N_21492,N_24594);
and UO_1357 (O_1357,N_20853,N_22444);
nor UO_1358 (O_1358,N_20501,N_24404);
xor UO_1359 (O_1359,N_23856,N_22236);
and UO_1360 (O_1360,N_19308,N_19028);
xnor UO_1361 (O_1361,N_18827,N_22367);
or UO_1362 (O_1362,N_19263,N_24679);
xor UO_1363 (O_1363,N_22610,N_21777);
or UO_1364 (O_1364,N_20283,N_19238);
xnor UO_1365 (O_1365,N_19884,N_23826);
nor UO_1366 (O_1366,N_24058,N_22939);
and UO_1367 (O_1367,N_24900,N_23187);
xor UO_1368 (O_1368,N_19569,N_21869);
and UO_1369 (O_1369,N_23234,N_22757);
nand UO_1370 (O_1370,N_21450,N_22322);
or UO_1371 (O_1371,N_24452,N_21808);
xnor UO_1372 (O_1372,N_22750,N_19976);
xnor UO_1373 (O_1373,N_22424,N_23358);
nor UO_1374 (O_1374,N_22818,N_18767);
and UO_1375 (O_1375,N_24298,N_22958);
xor UO_1376 (O_1376,N_24440,N_19997);
nand UO_1377 (O_1377,N_20985,N_23198);
and UO_1378 (O_1378,N_22700,N_23441);
nand UO_1379 (O_1379,N_22007,N_19679);
nor UO_1380 (O_1380,N_21649,N_20136);
and UO_1381 (O_1381,N_24273,N_20784);
or UO_1382 (O_1382,N_21906,N_23114);
xor UO_1383 (O_1383,N_23878,N_18926);
xnor UO_1384 (O_1384,N_24663,N_22708);
and UO_1385 (O_1385,N_23676,N_20910);
nor UO_1386 (O_1386,N_21194,N_19826);
xor UO_1387 (O_1387,N_24081,N_22535);
nor UO_1388 (O_1388,N_20345,N_22332);
and UO_1389 (O_1389,N_19167,N_21961);
xor UO_1390 (O_1390,N_23488,N_24354);
nor UO_1391 (O_1391,N_21401,N_19064);
or UO_1392 (O_1392,N_20429,N_24287);
nor UO_1393 (O_1393,N_22415,N_20434);
xnor UO_1394 (O_1394,N_24417,N_19251);
nor UO_1395 (O_1395,N_19959,N_24056);
and UO_1396 (O_1396,N_23822,N_22634);
xnor UO_1397 (O_1397,N_20524,N_23582);
or UO_1398 (O_1398,N_21969,N_24901);
or UO_1399 (O_1399,N_20081,N_23616);
and UO_1400 (O_1400,N_21471,N_23530);
or UO_1401 (O_1401,N_23728,N_21932);
nand UO_1402 (O_1402,N_19593,N_21817);
and UO_1403 (O_1403,N_21814,N_23158);
nor UO_1404 (O_1404,N_19894,N_21673);
and UO_1405 (O_1405,N_21089,N_20291);
nand UO_1406 (O_1406,N_24237,N_24319);
nand UO_1407 (O_1407,N_23019,N_18942);
xor UO_1408 (O_1408,N_20656,N_20586);
xnor UO_1409 (O_1409,N_19767,N_21628);
nor UO_1410 (O_1410,N_22396,N_22231);
nand UO_1411 (O_1411,N_19539,N_24809);
nor UO_1412 (O_1412,N_19518,N_22684);
or UO_1413 (O_1413,N_23081,N_20070);
nor UO_1414 (O_1414,N_22026,N_19134);
nor UO_1415 (O_1415,N_24284,N_22552);
nand UO_1416 (O_1416,N_24622,N_19855);
and UO_1417 (O_1417,N_23041,N_22763);
nor UO_1418 (O_1418,N_22893,N_24963);
xnor UO_1419 (O_1419,N_19336,N_23986);
nor UO_1420 (O_1420,N_21430,N_24514);
nor UO_1421 (O_1421,N_23469,N_22416);
or UO_1422 (O_1422,N_19836,N_18979);
nor UO_1423 (O_1423,N_22515,N_19908);
or UO_1424 (O_1424,N_19670,N_19892);
and UO_1425 (O_1425,N_20228,N_20509);
nor UO_1426 (O_1426,N_18909,N_21840);
nand UO_1427 (O_1427,N_19303,N_19061);
nor UO_1428 (O_1428,N_24739,N_19661);
or UO_1429 (O_1429,N_24727,N_20514);
xnor UO_1430 (O_1430,N_19678,N_20573);
or UO_1431 (O_1431,N_20357,N_23788);
nor UO_1432 (O_1432,N_22527,N_22587);
or UO_1433 (O_1433,N_20527,N_20021);
or UO_1434 (O_1434,N_19991,N_23839);
nand UO_1435 (O_1435,N_24261,N_18756);
and UO_1436 (O_1436,N_19636,N_21165);
nor UO_1437 (O_1437,N_22579,N_22374);
nor UO_1438 (O_1438,N_19861,N_21719);
nand UO_1439 (O_1439,N_24833,N_19689);
xnor UO_1440 (O_1440,N_22421,N_23741);
nor UO_1441 (O_1441,N_22560,N_20461);
nor UO_1442 (O_1442,N_21727,N_20674);
nand UO_1443 (O_1443,N_19662,N_24289);
xnor UO_1444 (O_1444,N_23499,N_22723);
or UO_1445 (O_1445,N_22822,N_18799);
and UO_1446 (O_1446,N_22944,N_18840);
nor UO_1447 (O_1447,N_22845,N_24376);
and UO_1448 (O_1448,N_23091,N_20504);
nand UO_1449 (O_1449,N_23796,N_19805);
or UO_1450 (O_1450,N_22663,N_24509);
or UO_1451 (O_1451,N_20969,N_21273);
xor UO_1452 (O_1452,N_19498,N_24443);
nand UO_1453 (O_1453,N_19639,N_24009);
xnor UO_1454 (O_1454,N_23079,N_21119);
and UO_1455 (O_1455,N_21043,N_19262);
and UO_1456 (O_1456,N_22014,N_23128);
xnor UO_1457 (O_1457,N_21909,N_21306);
nand UO_1458 (O_1458,N_23919,N_22255);
nor UO_1459 (O_1459,N_21855,N_19868);
nand UO_1460 (O_1460,N_20851,N_24694);
or UO_1461 (O_1461,N_21564,N_18764);
or UO_1462 (O_1462,N_23739,N_23463);
and UO_1463 (O_1463,N_19611,N_21672);
nor UO_1464 (O_1464,N_22053,N_19031);
xnor UO_1465 (O_1465,N_23623,N_24420);
nand UO_1466 (O_1466,N_23608,N_23485);
and UO_1467 (O_1467,N_18954,N_20238);
nand UO_1468 (O_1468,N_19606,N_24941);
or UO_1469 (O_1469,N_24321,N_19229);
nor UO_1470 (O_1470,N_19367,N_21724);
nor UO_1471 (O_1471,N_21117,N_21251);
xnor UO_1472 (O_1472,N_24508,N_20913);
nor UO_1473 (O_1473,N_24633,N_24664);
or UO_1474 (O_1474,N_24520,N_22502);
nor UO_1475 (O_1475,N_21440,N_23369);
nand UO_1476 (O_1476,N_20734,N_24337);
and UO_1477 (O_1477,N_22235,N_21144);
xnor UO_1478 (O_1478,N_19504,N_24649);
nand UO_1479 (O_1479,N_21451,N_19876);
and UO_1480 (O_1480,N_24089,N_20154);
nand UO_1481 (O_1481,N_22487,N_23172);
nand UO_1482 (O_1482,N_19558,N_19069);
nand UO_1483 (O_1483,N_21343,N_21624);
xnor UO_1484 (O_1484,N_23869,N_19090);
nor UO_1485 (O_1485,N_18945,N_24615);
and UO_1486 (O_1486,N_20856,N_22430);
nor UO_1487 (O_1487,N_21383,N_22735);
or UO_1488 (O_1488,N_20162,N_20263);
or UO_1489 (O_1489,N_21229,N_23761);
nand UO_1490 (O_1490,N_23452,N_23953);
or UO_1491 (O_1491,N_19692,N_19199);
xor UO_1492 (O_1492,N_24167,N_24391);
xnor UO_1493 (O_1493,N_24905,N_19557);
xor UO_1494 (O_1494,N_20758,N_22301);
nor UO_1495 (O_1495,N_23278,N_22371);
and UO_1496 (O_1496,N_22096,N_20466);
or UO_1497 (O_1497,N_20156,N_23824);
nor UO_1498 (O_1498,N_24339,N_19680);
nand UO_1499 (O_1499,N_21481,N_22972);
xor UO_1500 (O_1500,N_20895,N_22032);
and UO_1501 (O_1501,N_19628,N_21547);
nor UO_1502 (O_1502,N_21327,N_23075);
nand UO_1503 (O_1503,N_19380,N_22019);
nand UO_1504 (O_1504,N_20105,N_20054);
and UO_1505 (O_1505,N_24829,N_24421);
and UO_1506 (O_1506,N_21420,N_23105);
nand UO_1507 (O_1507,N_19280,N_20319);
and UO_1508 (O_1508,N_22049,N_23951);
or UO_1509 (O_1509,N_22743,N_23500);
nor UO_1510 (O_1510,N_22898,N_23793);
nor UO_1511 (O_1511,N_20951,N_22278);
nor UO_1512 (O_1512,N_18779,N_22910);
nor UO_1513 (O_1513,N_23813,N_21696);
xnor UO_1514 (O_1514,N_22607,N_23663);
or UO_1515 (O_1515,N_24910,N_18791);
or UO_1516 (O_1516,N_21586,N_22427);
nand UO_1517 (O_1517,N_23223,N_23009);
or UO_1518 (O_1518,N_21872,N_20876);
nor UO_1519 (O_1519,N_21580,N_22795);
and UO_1520 (O_1520,N_23085,N_19642);
nand UO_1521 (O_1521,N_23576,N_24661);
or UO_1522 (O_1522,N_24368,N_22254);
nand UO_1523 (O_1523,N_19135,N_23381);
xor UO_1524 (O_1524,N_21733,N_23464);
nand UO_1525 (O_1525,N_21641,N_21706);
nand UO_1526 (O_1526,N_19128,N_22911);
xnor UO_1527 (O_1527,N_18757,N_21914);
and UO_1528 (O_1528,N_24397,N_20995);
and UO_1529 (O_1529,N_21731,N_23175);
or UO_1530 (O_1530,N_24202,N_24883);
and UO_1531 (O_1531,N_24068,N_24702);
or UO_1532 (O_1532,N_21495,N_19101);
xnor UO_1533 (O_1533,N_18817,N_21207);
nor UO_1534 (O_1534,N_22413,N_24050);
and UO_1535 (O_1535,N_20502,N_23350);
nand UO_1536 (O_1536,N_21392,N_23908);
and UO_1537 (O_1537,N_20191,N_20621);
or UO_1538 (O_1538,N_23726,N_20046);
nand UO_1539 (O_1539,N_21196,N_18810);
nand UO_1540 (O_1540,N_22462,N_22833);
and UO_1541 (O_1541,N_20487,N_18812);
nor UO_1542 (O_1542,N_24460,N_22335);
and UO_1543 (O_1543,N_19271,N_23657);
nor UO_1544 (O_1544,N_20193,N_23593);
and UO_1545 (O_1545,N_24506,N_23658);
xnor UO_1546 (O_1546,N_22716,N_24393);
xor UO_1547 (O_1547,N_23387,N_20515);
or UO_1548 (O_1548,N_23190,N_21826);
xnor UO_1549 (O_1549,N_23035,N_20198);
and UO_1550 (O_1550,N_18816,N_21941);
nor UO_1551 (O_1551,N_24799,N_20295);
or UO_1552 (O_1552,N_22513,N_19788);
xor UO_1553 (O_1553,N_20025,N_20256);
nand UO_1554 (O_1554,N_24764,N_20565);
xnor UO_1555 (O_1555,N_19082,N_23297);
xor UO_1556 (O_1556,N_19545,N_24966);
nand UO_1557 (O_1557,N_20303,N_21744);
nor UO_1558 (O_1558,N_22129,N_24220);
or UO_1559 (O_1559,N_19956,N_24513);
nand UO_1560 (O_1560,N_19556,N_21246);
nand UO_1561 (O_1561,N_22842,N_19646);
nand UO_1562 (O_1562,N_24991,N_22948);
and UO_1563 (O_1563,N_23181,N_24293);
xor UO_1564 (O_1564,N_19490,N_23149);
xor UO_1565 (O_1565,N_20768,N_20407);
and UO_1566 (O_1566,N_21105,N_20443);
nand UO_1567 (O_1567,N_21549,N_19946);
and UO_1568 (O_1568,N_19962,N_24567);
nor UO_1569 (O_1569,N_19286,N_21351);
nand UO_1570 (O_1570,N_19497,N_22468);
nand UO_1571 (O_1571,N_21922,N_21352);
nor UO_1572 (O_1572,N_19057,N_20091);
xnor UO_1573 (O_1573,N_23611,N_22979);
nor UO_1574 (O_1574,N_20537,N_20196);
or UO_1575 (O_1575,N_22441,N_22978);
or UO_1576 (O_1576,N_21759,N_19713);
and UO_1577 (O_1577,N_21486,N_20402);
xor UO_1578 (O_1578,N_23703,N_21023);
xnor UO_1579 (O_1579,N_22811,N_22542);
or UO_1580 (O_1580,N_20237,N_22046);
or UO_1581 (O_1581,N_23014,N_21945);
nor UO_1582 (O_1582,N_24835,N_24977);
xnor UO_1583 (O_1583,N_19564,N_20990);
xnor UO_1584 (O_1584,N_23978,N_22216);
xnor UO_1585 (O_1585,N_20437,N_21534);
nor UO_1586 (O_1586,N_19843,N_18919);
and UO_1587 (O_1587,N_20658,N_20813);
nor UO_1588 (O_1588,N_19356,N_19902);
nor UO_1589 (O_1589,N_20243,N_24377);
or UO_1590 (O_1590,N_21064,N_21062);
xnor UO_1591 (O_1591,N_22844,N_18941);
and UO_1592 (O_1592,N_24654,N_19136);
and UO_1593 (O_1593,N_20664,N_18970);
xor UO_1594 (O_1594,N_21530,N_18952);
or UO_1595 (O_1595,N_24677,N_20355);
nor UO_1596 (O_1596,N_20057,N_19343);
or UO_1597 (O_1597,N_21182,N_20793);
and UO_1598 (O_1598,N_21323,N_20680);
xor UO_1599 (O_1599,N_19659,N_21208);
or UO_1600 (O_1600,N_22877,N_20842);
or UO_1601 (O_1601,N_19561,N_22177);
nor UO_1602 (O_1602,N_24014,N_22203);
nor UO_1603 (O_1603,N_24203,N_24976);
nand UO_1604 (O_1604,N_21825,N_19386);
nand UO_1605 (O_1605,N_23777,N_23380);
and UO_1606 (O_1606,N_21345,N_20213);
or UO_1607 (O_1607,N_24272,N_23328);
nor UO_1608 (O_1608,N_20454,N_22054);
and UO_1609 (O_1609,N_20297,N_24248);
nor UO_1610 (O_1610,N_19432,N_24346);
nand UO_1611 (O_1611,N_23711,N_22383);
nand UO_1612 (O_1612,N_22230,N_23802);
or UO_1613 (O_1613,N_23462,N_23089);
nor UO_1614 (O_1614,N_20932,N_21655);
or UO_1615 (O_1615,N_23017,N_19495);
and UO_1616 (O_1616,N_23734,N_24297);
xnor UO_1617 (O_1617,N_24162,N_23906);
or UO_1618 (O_1618,N_24027,N_19540);
nor UO_1619 (O_1619,N_24881,N_24418);
and UO_1620 (O_1620,N_23535,N_20304);
or UO_1621 (O_1621,N_19618,N_23047);
nand UO_1622 (O_1622,N_21293,N_19006);
or UO_1623 (O_1623,N_21398,N_23161);
and UO_1624 (O_1624,N_19817,N_22666);
or UO_1625 (O_1625,N_20983,N_23051);
xnor UO_1626 (O_1626,N_21272,N_23308);
nor UO_1627 (O_1627,N_20767,N_19397);
or UO_1628 (O_1628,N_19984,N_20214);
and UO_1629 (O_1629,N_20900,N_24226);
or UO_1630 (O_1630,N_21835,N_22732);
or UO_1631 (O_1631,N_19243,N_22794);
xnor UO_1632 (O_1632,N_22881,N_19555);
nand UO_1633 (O_1633,N_19928,N_24069);
or UO_1634 (O_1634,N_21104,N_20821);
or UO_1635 (O_1635,N_22321,N_20748);
and UO_1636 (O_1636,N_23432,N_23625);
and UO_1637 (O_1637,N_23076,N_20686);
or UO_1638 (O_1638,N_19507,N_18994);
and UO_1639 (O_1639,N_19147,N_24624);
xor UO_1640 (O_1640,N_18896,N_23832);
nor UO_1641 (O_1641,N_18820,N_22731);
nor UO_1642 (O_1642,N_22043,N_23784);
or UO_1643 (O_1643,N_20311,N_18839);
xor UO_1644 (O_1644,N_21887,N_21185);
and UO_1645 (O_1645,N_20298,N_21489);
nand UO_1646 (O_1646,N_24192,N_19849);
nand UO_1647 (O_1647,N_24318,N_23712);
and UO_1648 (O_1648,N_21516,N_19920);
xor UO_1649 (O_1649,N_19830,N_19873);
or UO_1650 (O_1650,N_20356,N_21500);
xnor UO_1651 (O_1651,N_23335,N_24644);
xor UO_1652 (O_1652,N_24422,N_20341);
nor UO_1653 (O_1653,N_24429,N_21954);
nor UO_1654 (O_1654,N_23945,N_24826);
nand UO_1655 (O_1655,N_18811,N_19438);
nor UO_1656 (O_1656,N_24908,N_23745);
xnor UO_1657 (O_1657,N_19761,N_22257);
nand UO_1658 (O_1658,N_23546,N_21294);
nand UO_1659 (O_1659,N_22158,N_18866);
nor UO_1660 (O_1660,N_24984,N_20363);
nor UO_1661 (O_1661,N_23835,N_24357);
and UO_1662 (O_1662,N_23544,N_19499);
and UO_1663 (O_1663,N_19768,N_19934);
or UO_1664 (O_1664,N_24596,N_22594);
and UO_1665 (O_1665,N_20168,N_19235);
and UO_1666 (O_1666,N_19816,N_24147);
nand UO_1667 (O_1667,N_24218,N_23967);
and UO_1668 (O_1668,N_19583,N_22994);
or UO_1669 (O_1669,N_21935,N_22980);
nor UO_1670 (O_1670,N_23851,N_19802);
nand UO_1671 (O_1671,N_21494,N_19828);
nor UO_1672 (O_1672,N_21110,N_24758);
xnor UO_1673 (O_1673,N_22274,N_21029);
nand UO_1674 (O_1674,N_19152,N_21473);
nor UO_1675 (O_1675,N_21480,N_18868);
xnor UO_1676 (O_1676,N_21736,N_19723);
nand UO_1677 (O_1677,N_21540,N_20922);
and UO_1678 (O_1678,N_21753,N_21138);
xnor UO_1679 (O_1679,N_24072,N_23036);
nor UO_1680 (O_1680,N_20007,N_20624);
and UO_1681 (O_1681,N_21866,N_22920);
xnor UO_1682 (O_1682,N_20166,N_21531);
xnor UO_1683 (O_1683,N_23553,N_20775);
or UO_1684 (O_1684,N_22400,N_22603);
nand UO_1685 (O_1685,N_20747,N_19068);
or UO_1686 (O_1686,N_22280,N_21147);
or UO_1687 (O_1687,N_21948,N_21078);
nand UO_1688 (O_1688,N_24772,N_23768);
xor UO_1689 (O_1689,N_20819,N_19815);
and UO_1690 (O_1690,N_21550,N_23757);
xnor UO_1691 (O_1691,N_24291,N_23957);
or UO_1692 (O_1692,N_24146,N_19186);
or UO_1693 (O_1693,N_22691,N_21317);
and UO_1694 (O_1694,N_20449,N_19311);
nand UO_1695 (O_1695,N_20358,N_19015);
or UO_1696 (O_1696,N_23276,N_20167);
and UO_1697 (O_1697,N_23983,N_21705);
nand UO_1698 (O_1698,N_22250,N_24535);
nand UO_1699 (O_1699,N_21539,N_24474);
or UO_1700 (O_1700,N_21210,N_23635);
or UO_1701 (O_1701,N_20759,N_20883);
or UO_1702 (O_1702,N_20564,N_22534);
and UO_1703 (O_1703,N_21915,N_22908);
or UO_1704 (O_1704,N_20728,N_21326);
and UO_1705 (O_1705,N_22570,N_18893);
xor UO_1706 (O_1706,N_24030,N_22820);
or UO_1707 (O_1707,N_21755,N_20915);
or UO_1708 (O_1708,N_20215,N_19482);
or UO_1709 (O_1709,N_19866,N_22595);
nand UO_1710 (O_1710,N_19195,N_23062);
nor UO_1711 (O_1711,N_21432,N_21143);
and UO_1712 (O_1712,N_22458,N_20699);
nand UO_1713 (O_1713,N_21416,N_22144);
nand UO_1714 (O_1714,N_19720,N_20125);
nand UO_1715 (O_1715,N_24931,N_21097);
nor UO_1716 (O_1716,N_21648,N_22388);
nor UO_1717 (O_1717,N_20160,N_20862);
or UO_1718 (O_1718,N_19016,N_19182);
xnor UO_1719 (O_1719,N_19365,N_20755);
nand UO_1720 (O_1720,N_24670,N_23287);
nor UO_1721 (O_1721,N_19665,N_22998);
or UO_1722 (O_1722,N_20226,N_22569);
nand UO_1723 (O_1723,N_21018,N_19146);
and UO_1724 (O_1724,N_22141,N_18877);
xor UO_1725 (O_1725,N_23428,N_21359);
or UO_1726 (O_1726,N_19087,N_18815);
xor UO_1727 (O_1727,N_22393,N_22455);
or UO_1728 (O_1728,N_24366,N_23294);
and UO_1729 (O_1729,N_24141,N_20368);
nand UO_1730 (O_1730,N_20418,N_21710);
and UO_1731 (O_1731,N_20684,N_20719);
and UO_1732 (O_1732,N_23540,N_21161);
xor UO_1733 (O_1733,N_24378,N_20003);
nand UO_1734 (O_1734,N_20279,N_23355);
xor UO_1735 (O_1735,N_23922,N_20060);
nand UO_1736 (O_1736,N_24361,N_22926);
nor UO_1737 (O_1737,N_21423,N_24499);
nor UO_1738 (O_1738,N_23117,N_24160);
nor UO_1739 (O_1739,N_22205,N_19520);
and UO_1740 (O_1740,N_22350,N_18903);
or UO_1741 (O_1741,N_24122,N_22548);
and UO_1742 (O_1742,N_20601,N_24301);
nand UO_1743 (O_1743,N_24823,N_21742);
and UO_1744 (O_1744,N_19766,N_23936);
nand UO_1745 (O_1745,N_22816,N_23961);
nand UO_1746 (O_1746,N_19613,N_18825);
or UO_1747 (O_1747,N_22297,N_20052);
nor UO_1748 (O_1748,N_21058,N_21952);
or UO_1749 (O_1749,N_19085,N_21365);
xnor UO_1750 (O_1750,N_22088,N_19176);
and UO_1751 (O_1751,N_23139,N_24187);
nor UO_1752 (O_1752,N_22703,N_21581);
xor UO_1753 (O_1753,N_22765,N_23267);
and UO_1754 (O_1754,N_19842,N_24721);
or UO_1755 (O_1755,N_20448,N_20569);
and UO_1756 (O_1756,N_24406,N_24061);
nor UO_1757 (O_1757,N_23162,N_18803);
xnor UO_1758 (O_1758,N_20271,N_21567);
and UO_1759 (O_1759,N_23127,N_23762);
nand UO_1760 (O_1760,N_21981,N_19614);
xnor UO_1761 (O_1761,N_22627,N_21061);
nor UO_1762 (O_1762,N_19597,N_21663);
xnor UO_1763 (O_1763,N_23329,N_24039);
nor UO_1764 (O_1764,N_21610,N_24827);
or UO_1765 (O_1765,N_20807,N_19278);
nor UO_1766 (O_1766,N_23250,N_23337);
and UO_1767 (O_1767,N_23144,N_19444);
and UO_1768 (O_1768,N_21212,N_20496);
nor UO_1769 (O_1769,N_23899,N_20385);
xor UO_1770 (O_1770,N_23255,N_21131);
nand UO_1771 (O_1771,N_20290,N_24082);
xnor UO_1772 (O_1772,N_19909,N_23792);
nor UO_1773 (O_1773,N_19982,N_22126);
xor UO_1774 (O_1774,N_22895,N_19141);
xnor UO_1775 (O_1775,N_24961,N_24841);
or UO_1776 (O_1776,N_22440,N_20762);
xor UO_1777 (O_1777,N_19492,N_23937);
and UO_1778 (O_1778,N_22843,N_20475);
nand UO_1779 (O_1779,N_23261,N_18846);
nand UO_1780 (O_1780,N_24716,N_20798);
xnor UO_1781 (O_1781,N_22202,N_18805);
nor UO_1782 (O_1782,N_23424,N_22764);
nor UO_1783 (O_1783,N_22473,N_20017);
or UO_1784 (O_1784,N_24714,N_18787);
nor UO_1785 (O_1785,N_20465,N_22251);
xnor UO_1786 (O_1786,N_19273,N_19324);
xnor UO_1787 (O_1787,N_24659,N_22710);
xnor UO_1788 (O_1788,N_21160,N_24563);
or UO_1789 (O_1789,N_23157,N_23682);
or UO_1790 (O_1790,N_18959,N_19337);
nand UO_1791 (O_1791,N_21875,N_20258);
nor UO_1792 (O_1792,N_24448,N_24090);
or UO_1793 (O_1793,N_18763,N_22767);
or UO_1794 (O_1794,N_23078,N_22933);
xnor UO_1795 (O_1795,N_22121,N_24978);
nor UO_1796 (O_1796,N_21904,N_19574);
or UO_1797 (O_1797,N_19137,N_21447);
nor UO_1798 (O_1798,N_21739,N_24936);
nor UO_1799 (O_1799,N_19413,N_22020);
or UO_1800 (O_1800,N_23236,N_21149);
or UO_1801 (O_1801,N_21318,N_23211);
xnor UO_1802 (O_1802,N_19792,N_20810);
or UO_1803 (O_1803,N_21356,N_20040);
nor UO_1804 (O_1804,N_21885,N_23617);
and UO_1805 (O_1805,N_20735,N_23927);
and UO_1806 (O_1806,N_22730,N_24079);
or UO_1807 (O_1807,N_19046,N_20634);
nand UO_1808 (O_1808,N_20548,N_24138);
nand UO_1809 (O_1809,N_24432,N_21802);
nand UO_1810 (O_1810,N_21838,N_20906);
nor UO_1811 (O_1811,N_20420,N_22447);
xnor UO_1812 (O_1812,N_19850,N_24906);
and UO_1813 (O_1813,N_21810,N_22245);
nand UO_1814 (O_1814,N_21497,N_23905);
nor UO_1815 (O_1815,N_20591,N_24286);
and UO_1816 (O_1816,N_20590,N_23622);
and UO_1817 (O_1817,N_21042,N_21056);
nand UO_1818 (O_1818,N_24733,N_21893);
and UO_1819 (O_1819,N_22484,N_20946);
and UO_1820 (O_1820,N_24395,N_23275);
nor UO_1821 (O_1821,N_21694,N_20413);
or UO_1822 (O_1822,N_22106,N_24552);
and UO_1823 (O_1823,N_19796,N_22229);
xor UO_1824 (O_1824,N_24240,N_24818);
nand UO_1825 (O_1825,N_24469,N_21037);
nand UO_1826 (O_1826,N_20367,N_24782);
xor UO_1827 (O_1827,N_19348,N_20567);
nor UO_1828 (O_1828,N_24351,N_21779);
or UO_1829 (O_1829,N_22817,N_23003);
xnor UO_1830 (O_1830,N_23644,N_22139);
xor UO_1831 (O_1831,N_24306,N_20814);
xnor UO_1832 (O_1832,N_22874,N_23010);
nor UO_1833 (O_1833,N_24340,N_24023);
xor UO_1834 (O_1834,N_24805,N_20029);
nand UO_1835 (O_1835,N_24746,N_24413);
and UO_1836 (O_1836,N_21820,N_22965);
and UO_1837 (O_1837,N_19743,N_24521);
nand UO_1838 (O_1838,N_20379,N_20151);
nor UO_1839 (O_1839,N_19824,N_19641);
or UO_1840 (O_1840,N_23397,N_23708);
and UO_1841 (O_1841,N_19827,N_22445);
and UO_1842 (O_1842,N_21073,N_19025);
or UO_1843 (O_1843,N_21570,N_20541);
and UO_1844 (O_1844,N_22543,N_18939);
nor UO_1845 (O_1845,N_22864,N_20536);
xnor UO_1846 (O_1846,N_23133,N_23770);
xor UO_1847 (O_1847,N_22558,N_19964);
nor UO_1848 (O_1848,N_22746,N_20879);
nand UO_1849 (O_1849,N_19951,N_19754);
nand UO_1850 (O_1850,N_24934,N_23437);
nor UO_1851 (O_1851,N_22272,N_23783);
or UO_1852 (O_1852,N_23898,N_23537);
nor UO_1853 (O_1853,N_19269,N_20612);
and UO_1854 (O_1854,N_21474,N_24282);
and UO_1855 (O_1855,N_21441,N_24872);
xor UO_1856 (O_1856,N_22969,N_24207);
or UO_1857 (O_1857,N_21907,N_20687);
nor UO_1858 (O_1858,N_22005,N_19621);
xor UO_1859 (O_1859,N_20578,N_19175);
and UO_1860 (O_1860,N_23713,N_19798);
or UO_1861 (O_1861,N_22656,N_19612);
or UO_1862 (O_1862,N_20254,N_22395);
or UO_1863 (O_1863,N_23156,N_19999);
nand UO_1864 (O_1864,N_23992,N_19393);
or UO_1865 (O_1865,N_23218,N_21254);
nand UO_1866 (O_1866,N_23794,N_23508);
and UO_1867 (O_1867,N_20637,N_24675);
or UO_1868 (O_1868,N_21861,N_20976);
or UO_1869 (O_1869,N_19535,N_23131);
nand UO_1870 (O_1870,N_22617,N_24820);
nand UO_1871 (O_1871,N_24665,N_23791);
xnor UO_1872 (O_1872,N_18891,N_20654);
or UO_1873 (O_1873,N_24847,N_21559);
and UO_1874 (O_1874,N_24300,N_21214);
nand UO_1875 (O_1875,N_19509,N_21768);
xor UO_1876 (O_1876,N_20274,N_22951);
or UO_1877 (O_1877,N_19013,N_19005);
xor UO_1878 (O_1878,N_19948,N_23572);
xnor UO_1879 (O_1879,N_24447,N_20247);
or UO_1880 (O_1880,N_21485,N_23086);
or UO_1881 (O_1881,N_21406,N_19364);
and UO_1882 (O_1882,N_24410,N_18844);
and UO_1883 (O_1883,N_24365,N_22041);
and UO_1884 (O_1884,N_20500,N_22885);
nor UO_1885 (O_1885,N_22460,N_19952);
nand UO_1886 (O_1886,N_20388,N_21276);
xor UO_1887 (O_1887,N_23204,N_22342);
or UO_1888 (O_1888,N_21310,N_23349);
xnor UO_1889 (O_1889,N_21469,N_19402);
and UO_1890 (O_1890,N_22891,N_19967);
nor UO_1891 (O_1891,N_20945,N_22917);
or UO_1892 (O_1892,N_24710,N_19590);
nor UO_1893 (O_1893,N_22850,N_24249);
nor UO_1894 (O_1894,N_20455,N_21913);
xor UO_1895 (O_1895,N_24583,N_24328);
and UO_1896 (O_1896,N_22108,N_19566);
xor UO_1897 (O_1897,N_19347,N_21332);
and UO_1898 (O_1898,N_21911,N_20172);
nand UO_1899 (O_1899,N_22482,N_24933);
nand UO_1900 (O_1900,N_21172,N_21202);
or UO_1901 (O_1901,N_21069,N_22504);
xnor UO_1902 (O_1902,N_23670,N_23800);
nor UO_1903 (O_1903,N_20780,N_21656);
xor UO_1904 (O_1904,N_22215,N_21925);
nor UO_1905 (O_1905,N_24183,N_22686);
nor UO_1906 (O_1906,N_22516,N_20692);
xor UO_1907 (O_1907,N_18925,N_24630);
xor UO_1908 (O_1908,N_23053,N_20891);
nor UO_1909 (O_1909,N_19040,N_20804);
and UO_1910 (O_1910,N_22481,N_21938);
or UO_1911 (O_1911,N_23545,N_21263);
xor UO_1912 (O_1912,N_19351,N_20164);
nand UO_1913 (O_1913,N_19344,N_21145);
xor UO_1914 (O_1914,N_24211,N_19067);
nor UO_1915 (O_1915,N_19449,N_21621);
nand UO_1916 (O_1916,N_23402,N_19565);
nor UO_1917 (O_1917,N_22770,N_18947);
xor UO_1918 (O_1918,N_24385,N_24982);
xnor UO_1919 (O_1919,N_22942,N_23284);
nand UO_1920 (O_1920,N_22425,N_22130);
nand UO_1921 (O_1921,N_20730,N_19568);
and UO_1922 (O_1922,N_18928,N_21284);
and UO_1923 (O_1923,N_22983,N_21912);
nor UO_1924 (O_1924,N_20959,N_24401);
and UO_1925 (O_1925,N_19668,N_21833);
xor UO_1926 (O_1926,N_22011,N_23700);
nor UO_1927 (O_1927,N_21125,N_19099);
nor UO_1928 (O_1928,N_24364,N_20481);
and UO_1929 (O_1929,N_20682,N_24562);
and UO_1930 (O_1930,N_23921,N_23489);
and UO_1931 (O_1931,N_21926,N_21965);
xor UO_1932 (O_1932,N_22178,N_24559);
nand UO_1933 (O_1933,N_20751,N_24707);
nor UO_1934 (O_1934,N_23702,N_24944);
xor UO_1935 (O_1935,N_20966,N_23689);
nor UO_1936 (O_1936,N_22449,N_24259);
or UO_1937 (O_1937,N_22364,N_20494);
or UO_1938 (O_1938,N_18869,N_21446);
xor UO_1939 (O_1939,N_20707,N_23056);
and UO_1940 (O_1940,N_19918,N_24274);
or UO_1941 (O_1941,N_23680,N_21606);
nand UO_1942 (O_1942,N_20928,N_24372);
nor UO_1943 (O_1943,N_24882,N_22976);
nand UO_1944 (O_1944,N_20242,N_21142);
and UO_1945 (O_1945,N_18800,N_23280);
and UO_1946 (O_1946,N_21857,N_23717);
or UO_1947 (O_1947,N_22285,N_20629);
xor UO_1948 (O_1948,N_24928,N_22938);
nor UO_1949 (O_1949,N_21390,N_24091);
and UO_1950 (O_1950,N_19751,N_24741);
and UO_1951 (O_1951,N_24115,N_24392);
or UO_1952 (O_1952,N_24763,N_24425);
and UO_1953 (O_1953,N_23958,N_23325);
xor UO_1954 (O_1954,N_24884,N_20389);
or UO_1955 (O_1955,N_21865,N_20464);
nor UO_1956 (O_1956,N_24093,N_22172);
or UO_1957 (O_1957,N_20266,N_18849);
nand UO_1958 (O_1958,N_19220,N_22313);
and UO_1959 (O_1959,N_24047,N_24576);
nor UO_1960 (O_1960,N_24262,N_22001);
nand UO_1961 (O_1961,N_22191,N_20433);
or UO_1962 (O_1962,N_23864,N_18792);
nand UO_1963 (O_1963,N_19489,N_21943);
nor UO_1964 (O_1964,N_18769,N_20882);
and UO_1965 (O_1965,N_19288,N_24686);
xor UO_1966 (O_1966,N_23804,N_23628);
nor UO_1967 (O_1967,N_21992,N_19236);
xnor UO_1968 (O_1968,N_22622,N_22299);
or UO_1969 (O_1969,N_22501,N_23045);
or UO_1970 (O_1970,N_19506,N_22830);
nor UO_1971 (O_1971,N_20681,N_22638);
nor UO_1972 (O_1972,N_23244,N_22098);
xor UO_1973 (O_1973,N_19986,N_21367);
or UO_1974 (O_1974,N_24402,N_23220);
or UO_1975 (O_1975,N_20394,N_23555);
or UO_1976 (O_1976,N_22351,N_21101);
and UO_1977 (O_1977,N_21424,N_22328);
nand UO_1978 (O_1978,N_18760,N_22037);
nor UO_1979 (O_1979,N_22742,N_21877);
xor UO_1980 (O_1980,N_19625,N_19548);
and UO_1981 (O_1981,N_20265,N_22778);
or UO_1982 (O_1982,N_23263,N_24863);
nand UO_1983 (O_1983,N_24652,N_18895);
and UO_1984 (O_1984,N_22118,N_20491);
nand UO_1985 (O_1985,N_23057,N_22348);
nor UO_1986 (O_1986,N_24492,N_23534);
nor UO_1987 (O_1987,N_23698,N_24849);
xnor UO_1988 (O_1988,N_24986,N_23581);
nand UO_1989 (O_1989,N_23459,N_19879);
or UO_1990 (O_1990,N_19187,N_23812);
or UO_1991 (O_1991,N_20989,N_23730);
and UO_1992 (O_1992,N_18854,N_22810);
nor UO_1993 (O_1993,N_20934,N_19926);
nor UO_1994 (O_1994,N_20230,N_24283);
or UO_1995 (O_1995,N_24126,N_22403);
nor UO_1996 (O_1996,N_22008,N_22089);
or UO_1997 (O_1997,N_24705,N_21195);
and UO_1998 (O_1998,N_24483,N_18914);
and UO_1999 (O_1999,N_22780,N_19516);
nor UO_2000 (O_2000,N_21854,N_23401);
xor UO_2001 (O_2001,N_20503,N_19250);
nor UO_2002 (O_2002,N_19431,N_21789);
xor UO_2003 (O_2003,N_19981,N_23669);
or UO_2004 (O_2004,N_23249,N_22060);
and UO_2005 (O_2005,N_21929,N_24695);
nor UO_2006 (O_2006,N_22243,N_23225);
and UO_2007 (O_2007,N_23938,N_19088);
and UO_2008 (O_2008,N_20633,N_21669);
nor UO_2009 (O_2009,N_24083,N_23159);
nand UO_2010 (O_2010,N_23507,N_19847);
and UO_2011 (O_2011,N_21692,N_22664);
xor UO_2012 (O_2012,N_23196,N_23971);
or UO_2013 (O_2013,N_21103,N_23910);
and UO_2014 (O_2014,N_23206,N_24125);
nand UO_2015 (O_2015,N_24129,N_22905);
and UO_2016 (O_2016,N_20743,N_18797);
nand UO_2017 (O_2017,N_19032,N_20056);
or UO_2018 (O_2018,N_23947,N_24454);
nor UO_2019 (O_2019,N_22649,N_23021);
xor UO_2020 (O_2020,N_18894,N_18783);
or UO_2021 (O_2021,N_22079,N_20999);
or UO_2022 (O_2022,N_19111,N_24773);
xor UO_2023 (O_2023,N_21728,N_19513);
or UO_2024 (O_2024,N_20010,N_23649);
and UO_2025 (O_2025,N_19129,N_24791);
and UO_2026 (O_2026,N_20511,N_21476);
and UO_2027 (O_2027,N_24697,N_20902);
or UO_2028 (O_2028,N_20177,N_24006);
xor UO_2029 (O_2029,N_23994,N_20655);
and UO_2030 (O_2030,N_24537,N_22031);
nor UO_2031 (O_2031,N_20490,N_24546);
nor UO_2032 (O_2032,N_24011,N_19309);
and UO_2033 (O_2033,N_24426,N_19831);
and UO_2034 (O_2034,N_22892,N_20971);
nand UO_2035 (O_2035,N_23579,N_23293);
and UO_2036 (O_2036,N_19366,N_20408);
xnor UO_2037 (O_2037,N_23230,N_20795);
nand UO_2038 (O_2038,N_20799,N_24696);
nand UO_2039 (O_2039,N_24845,N_22092);
and UO_2040 (O_2040,N_24808,N_22417);
and UO_2041 (O_2041,N_21795,N_22063);
and UO_2042 (O_2042,N_18918,N_20721);
and UO_2043 (O_2043,N_18961,N_20750);
and UO_2044 (O_2044,N_19971,N_23722);
xnor UO_2045 (O_2045,N_23999,N_21324);
or UO_2046 (O_2046,N_20669,N_24468);
or UO_2047 (O_2047,N_23427,N_23533);
xnor UO_2048 (O_2048,N_20194,N_22263);
or UO_2049 (O_2049,N_23865,N_23202);
nor UO_2050 (O_2050,N_24951,N_19330);
nand UO_2051 (O_2051,N_21552,N_24761);
nor UO_2052 (O_2052,N_22875,N_20948);
nor UO_2053 (O_2053,N_21850,N_19582);
nor UO_2054 (O_2054,N_21612,N_19731);
nor UO_2055 (O_2055,N_23887,N_22799);
and UO_2056 (O_2056,N_21977,N_20917);
or UO_2057 (O_2057,N_21232,N_24886);
nor UO_2058 (O_2058,N_19672,N_20752);
or UO_2059 (O_2059,N_23855,N_23088);
and UO_2060 (O_2060,N_19475,N_19232);
and UO_2061 (O_2061,N_23685,N_23258);
and UO_2062 (O_2062,N_22164,N_20064);
xor UO_2063 (O_2063,N_22176,N_21748);
or UO_2064 (O_2064,N_19977,N_20888);
nor UO_2065 (O_2065,N_23450,N_21895);
xnor UO_2066 (O_2066,N_18830,N_24911);
and UO_2067 (O_2067,N_21262,N_23846);
nand UO_2068 (O_2068,N_19041,N_24475);
or UO_2069 (O_2069,N_19560,N_22689);
or UO_2070 (O_2070,N_21894,N_22123);
xor UO_2071 (O_2071,N_20250,N_22157);
nand UO_2072 (O_2072,N_24518,N_23867);
xnor UO_2073 (O_2073,N_20809,N_23371);
or UO_2074 (O_2074,N_21980,N_21525);
or UO_2075 (O_2075,N_24111,N_20071);
nor UO_2076 (O_2076,N_23970,N_20272);
and UO_2077 (O_2077,N_20002,N_24965);
or UO_2078 (O_2078,N_18880,N_24092);
xor UO_2079 (O_2079,N_20008,N_22632);
or UO_2080 (O_2080,N_19453,N_24873);
and UO_2081 (O_2081,N_24004,N_19961);
or UO_2082 (O_2082,N_24922,N_23931);
or UO_2083 (O_2083,N_24929,N_24585);
nand UO_2084 (O_2084,N_22240,N_22827);
nand UO_2085 (O_2085,N_24860,N_22935);
or UO_2086 (O_2086,N_21325,N_23900);
or UO_2087 (O_2087,N_21203,N_21699);
nor UO_2088 (O_2088,N_21266,N_22267);
or UO_2089 (O_2089,N_21151,N_19466);
xor UO_2090 (O_2090,N_19306,N_19177);
or UO_2091 (O_2091,N_23941,N_21128);
or UO_2092 (O_2092,N_24155,N_19214);
or UO_2093 (O_2093,N_18853,N_24706);
nor UO_2094 (O_2094,N_20328,N_22199);
or UO_2095 (O_2095,N_21344,N_20093);
nor UO_2096 (O_2096,N_19171,N_22380);
nor UO_2097 (O_2097,N_19160,N_20294);
nand UO_2098 (O_2098,N_20333,N_20222);
nor UO_2099 (O_2099,N_21304,N_20869);
and UO_2100 (O_2100,N_19149,N_23807);
nand UO_2101 (O_2101,N_18957,N_19151);
xnor UO_2102 (O_2102,N_23426,N_22825);
nand UO_2103 (O_2103,N_19381,N_23565);
nor UO_2104 (O_2104,N_21010,N_23942);
nand UO_2105 (O_2105,N_21470,N_18781);
and UO_2106 (O_2106,N_19189,N_21515);
or UO_2107 (O_2107,N_23753,N_24444);
xnor UO_2108 (O_2108,N_22873,N_20632);
xnor UO_2109 (O_2109,N_24074,N_24128);
nor UO_2110 (O_2110,N_20659,N_20513);
nor UO_2111 (O_2111,N_19608,N_19001);
or UO_2112 (O_2112,N_23201,N_19954);
xor UO_2113 (O_2113,N_23570,N_24769);
xnor UO_2114 (O_2114,N_22281,N_22676);
nand UO_2115 (O_2115,N_24701,N_21576);
and UO_2116 (O_2116,N_22472,N_24971);
xor UO_2117 (O_2117,N_22131,N_19066);
nand UO_2118 (O_2118,N_20938,N_20239);
and UO_2119 (O_2119,N_24579,N_20923);
xnor UO_2120 (O_2120,N_24102,N_19213);
and UO_2121 (O_2121,N_22153,N_20020);
nor UO_2122 (O_2122,N_22824,N_20778);
and UO_2123 (O_2123,N_19771,N_20877);
and UO_2124 (O_2124,N_23300,N_23823);
or UO_2125 (O_2125,N_22125,N_21305);
or UO_2126 (O_2126,N_19089,N_24398);
nand UO_2127 (O_2127,N_21218,N_23330);
or UO_2128 (O_2128,N_20558,N_23888);
and UO_2129 (O_2129,N_24260,N_23323);
nand UO_2130 (O_2130,N_23924,N_21376);
and UO_2131 (O_2131,N_22154,N_22970);
and UO_2132 (O_2132,N_18901,N_20618);
nand UO_2133 (O_2133,N_22626,N_20526);
nor UO_2134 (O_2134,N_24409,N_22914);
and UO_2135 (O_2135,N_23871,N_19821);
xnor UO_2136 (O_2136,N_20646,N_24500);
nor UO_2137 (O_2137,N_22977,N_19718);
xor UO_2138 (O_2138,N_24838,N_23558);
nand UO_2139 (O_2139,N_23145,N_22024);
nand UO_2140 (O_2140,N_19070,N_18876);
xor UO_2141 (O_2141,N_24356,N_19451);
and UO_2142 (O_2142,N_21137,N_24480);
nand UO_2143 (O_2143,N_21839,N_19832);
xnor UO_2144 (O_2144,N_21940,N_24073);
xor UO_2145 (O_2145,N_19501,N_22399);
or UO_2146 (O_2146,N_22748,N_21358);
nand UO_2147 (O_2147,N_21448,N_23197);
or UO_2148 (O_2148,N_23224,N_24323);
nand UO_2149 (O_2149,N_23965,N_20545);
or UO_2150 (O_2150,N_20553,N_24066);
nor UO_2151 (O_2151,N_19272,N_24095);
nor UO_2152 (O_2152,N_22955,N_19919);
nor UO_2153 (O_2153,N_21930,N_20314);
and UO_2154 (O_2154,N_23298,N_19154);
and UO_2155 (O_2155,N_24213,N_23509);
or UO_2156 (O_2156,N_22711,N_21378);
or UO_2157 (O_2157,N_24999,N_24853);
xnor UO_2158 (O_2158,N_23248,N_22897);
nor UO_2159 (O_2159,N_22620,N_22623);
nand UO_2160 (O_2160,N_24819,N_21766);
nand UO_2161 (O_2161,N_21591,N_19627);
nand UO_2162 (O_2162,N_20212,N_21413);
and UO_2163 (O_2163,N_20378,N_24814);
nand UO_2164 (O_2164,N_23916,N_22592);
and UO_2165 (O_2165,N_21798,N_22507);
nor UO_2166 (O_2166,N_22522,N_23005);
nor UO_2167 (O_2167,N_19092,N_21166);
nor UO_2168 (O_2168,N_19673,N_22228);
nand UO_2169 (O_2169,N_20889,N_21873);
nand UO_2170 (O_2170,N_21328,N_19107);
and UO_2171 (O_2171,N_19870,N_18773);
xor UO_2172 (O_2172,N_20108,N_20739);
and UO_2173 (O_2173,N_22200,N_20765);
and UO_2174 (O_2174,N_23504,N_21778);
and UO_2175 (O_2175,N_20867,N_22246);
and UO_2176 (O_2176,N_23798,N_21415);
and UO_2177 (O_2177,N_19369,N_19748);
nand UO_2178 (O_2178,N_24806,N_19222);
or UO_2179 (O_2179,N_19316,N_20926);
and UO_2180 (O_2180,N_23039,N_21321);
and UO_2181 (O_2181,N_20204,N_21760);
xnor UO_2182 (O_2182,N_24136,N_21698);
and UO_2183 (O_2183,N_20839,N_22002);
nor UO_2184 (O_2184,N_19456,N_23987);
or UO_2185 (O_2185,N_22266,N_23541);
and UO_2186 (O_2186,N_22189,N_19203);
and UO_2187 (O_2187,N_21582,N_20326);
nand UO_2188 (O_2188,N_24987,N_24844);
or UO_2189 (O_2189,N_24640,N_24533);
nor UO_2190 (O_2190,N_23253,N_21467);
xor UO_2191 (O_2191,N_20619,N_19714);
nand UO_2192 (O_2192,N_21153,N_19779);
and UO_2193 (O_2193,N_24010,N_24338);
or UO_2194 (O_2194,N_22902,N_24370);
or UO_2195 (O_2195,N_19018,N_19980);
and UO_2196 (O_2196,N_23200,N_22616);
nor UO_2197 (O_2197,N_19686,N_21627);
nor UO_2198 (O_2198,N_18986,N_20904);
nand UO_2199 (O_2199,N_19354,N_19886);
and UO_2200 (O_2200,N_20138,N_24100);
and UO_2201 (O_2201,N_21346,N_19406);
or UO_2202 (O_2202,N_21242,N_24511);
xnor UO_2203 (O_2203,N_23636,N_23059);
or UO_2204 (O_2204,N_20278,N_24685);
nand UO_2205 (O_2205,N_21419,N_19907);
and UO_2206 (O_2206,N_24569,N_22903);
or UO_2207 (O_2207,N_20532,N_22836);
nand UO_2208 (O_2208,N_24734,N_19503);
xnor UO_2209 (O_2209,N_22122,N_20673);
and UO_2210 (O_2210,N_18962,N_24898);
xnor UO_2211 (O_2211,N_24084,N_20446);
or UO_2212 (O_2212,N_24839,N_19170);
and UO_2213 (O_2213,N_23502,N_21139);
or UO_2214 (O_2214,N_23577,N_18804);
nand UO_2215 (O_2215,N_21543,N_20528);
nand UO_2216 (O_2216,N_20331,N_24032);
nor UO_2217 (O_2217,N_19471,N_23134);
xnor UO_2218 (O_2218,N_19835,N_23277);
or UO_2219 (O_2219,N_20582,N_24046);
nand UO_2220 (O_2220,N_24157,N_22608);
or UO_2221 (O_2221,N_24191,N_24947);
xor UO_2222 (O_2222,N_21819,N_21846);
nor UO_2223 (O_2223,N_21259,N_21391);
and UO_2224 (O_2224,N_20554,N_21661);
nor UO_2225 (O_2225,N_22660,N_21767);
xnor UO_2226 (O_2226,N_19595,N_22077);
xor UO_2227 (O_2227,N_20575,N_21667);
nand UO_2228 (O_2228,N_19091,N_23940);
or UO_2229 (O_2229,N_20221,N_20457);
nor UO_2230 (O_2230,N_22311,N_22237);
nor UO_2231 (O_2231,N_19405,N_20683);
or UO_2232 (O_2232,N_24698,N_20313);
xor UO_2233 (O_2233,N_22378,N_19075);
xor UO_2234 (O_2234,N_18884,N_24760);
and UO_2235 (O_2235,N_21053,N_20506);
xor UO_2236 (O_2236,N_20370,N_22119);
nand UO_2237 (O_2237,N_23273,N_19891);
nand UO_2238 (O_2238,N_24689,N_21080);
and UO_2239 (O_2239,N_20024,N_21385);
or UO_2240 (O_2240,N_19297,N_24850);
nand UO_2241 (O_2241,N_19416,N_21963);
nand UO_2242 (O_2242,N_23569,N_24540);
or UO_2243 (O_2243,N_20332,N_20488);
or UO_2244 (O_2244,N_21124,N_21396);
nand UO_2245 (O_2245,N_23396,N_23026);
and UO_2246 (O_2246,N_20427,N_19255);
xnor UO_2247 (O_2247,N_18902,N_24121);
nand UO_2248 (O_2248,N_19581,N_22768);
or UO_2249 (O_2249,N_20306,N_24958);
and UO_2250 (O_2250,N_22312,N_20855);
xnor UO_2251 (O_2251,N_24269,N_20426);
xor UO_2252 (O_2252,N_21821,N_19350);
or UO_2253 (O_2253,N_21890,N_21774);
and UO_2254 (O_2254,N_19797,N_21368);
xnor UO_2255 (O_2255,N_21937,N_22840);
or UO_2256 (O_2256,N_21456,N_19944);
nand UO_2257 (O_2257,N_20887,N_21642);
and UO_2258 (O_2258,N_18768,N_24593);
or UO_2259 (O_2259,N_24893,N_24290);
and UO_2260 (O_2260,N_21001,N_19594);
xor UO_2261 (O_2261,N_24411,N_23471);
nor UO_2262 (O_2262,N_24528,N_22477);
or UO_2263 (O_2263,N_19811,N_21588);
nand UO_2264 (O_2264,N_23578,N_20049);
and UO_2265 (O_2265,N_21918,N_20987);
and UO_2266 (O_2266,N_20058,N_23640);
xnor UO_2267 (O_2267,N_22883,N_24955);
xor UO_2268 (O_2268,N_20047,N_23929);
and UO_2269 (O_2269,N_23873,N_20587);
xor UO_2270 (O_2270,N_20387,N_23317);
or UO_2271 (O_2271,N_20718,N_18882);
and UO_2272 (O_2272,N_23168,N_20670);
or UO_2273 (O_2273,N_20181,N_23510);
xor UO_2274 (O_2274,N_24131,N_22470);
nor UO_2275 (O_2275,N_21031,N_22289);
xnor UO_2276 (O_2276,N_18973,N_18996);
nand UO_2277 (O_2277,N_20401,N_21770);
nand UO_2278 (O_2278,N_23137,N_20092);
or UO_2279 (O_2279,N_20628,N_19979);
nand UO_2280 (O_2280,N_24382,N_19140);
or UO_2281 (O_2281,N_19035,N_22568);
and UO_2282 (O_2282,N_24256,N_21216);
or UO_2283 (O_2283,N_24547,N_24465);
nand UO_2284 (O_2284,N_23238,N_21068);
or UO_2285 (O_2285,N_22052,N_23574);
nor UO_2286 (O_2286,N_24134,N_19669);
nand UO_2287 (O_2287,N_24198,N_21746);
and UO_2288 (O_2288,N_23080,N_24869);
nand UO_2289 (O_2289,N_19698,N_24442);
xor UO_2290 (O_2290,N_20789,N_22521);
xnor UO_2291 (O_2291,N_21709,N_20190);
nor UO_2292 (O_2292,N_21362,N_20772);
and UO_2293 (O_2293,N_24254,N_22127);
xnor UO_2294 (O_2294,N_20137,N_20004);
or UO_2295 (O_2295,N_20660,N_20516);
and UO_2296 (O_2296,N_24683,N_23849);
or UO_2297 (O_2297,N_23333,N_23686);
nor UO_2298 (O_2298,N_20733,N_20740);
nor UO_2299 (O_2299,N_21794,N_21975);
nand UO_2300 (O_2300,N_20273,N_21342);
nor UO_2301 (O_2301,N_19116,N_19384);
nor UO_2302 (O_2302,N_19100,N_22361);
or UO_2303 (O_2303,N_19775,N_19533);
nor UO_2304 (O_2304,N_21496,N_23332);
xnor UO_2305 (O_2305,N_24316,N_23787);
nor UO_2306 (O_2306,N_23795,N_23920);
and UO_2307 (O_2307,N_21096,N_24759);
or UO_2308 (O_2308,N_20533,N_21060);
nor UO_2309 (O_2309,N_21521,N_21923);
nor UO_2310 (O_2310,N_24550,N_18814);
xnor UO_2311 (O_2311,N_23917,N_20641);
xnor UO_2312 (O_2312,N_19304,N_22523);
or UO_2313 (O_2313,N_21972,N_22319);
nor UO_2314 (O_2314,N_23188,N_24646);
or UO_2315 (O_2315,N_23292,N_19274);
nor UO_2316 (O_2316,N_20622,N_22524);
or UO_2317 (O_2317,N_19531,N_20831);
and UO_2318 (O_2318,N_22135,N_23897);
and UO_2319 (O_2319,N_24981,N_23266);
xnor UO_2320 (O_2320,N_21512,N_19333);
and UO_2321 (O_2321,N_23806,N_21944);
nand UO_2322 (O_2322,N_24855,N_24516);
xor UO_2323 (O_2323,N_24019,N_21198);
or UO_2324 (O_2324,N_24229,N_21776);
or UO_2325 (O_2325,N_21665,N_24109);
nor UO_2326 (O_2326,N_24315,N_20032);
nor UO_2327 (O_2327,N_24035,N_19987);
nand UO_2328 (O_2328,N_21425,N_24524);
nor UO_2329 (O_2329,N_19388,N_21700);
and UO_2330 (O_2330,N_23366,N_18875);
nor UO_2331 (O_2331,N_22013,N_23345);
or UO_2332 (O_2332,N_23861,N_19204);
nor UO_2333 (O_2333,N_20954,N_24645);
nor UO_2334 (O_2334,N_23840,N_22692);
nand UO_2335 (O_2335,N_21772,N_22124);
and UO_2336 (O_2336,N_20312,N_19219);
or UO_2337 (O_2337,N_23988,N_20202);
nand UO_2338 (O_2338,N_21903,N_22981);
nand UO_2339 (O_2339,N_23024,N_24532);
nand UO_2340 (O_2340,N_19994,N_22059);
nand UO_2341 (O_2341,N_23094,N_21083);
nor UO_2342 (O_2342,N_24692,N_20373);
nand UO_2343 (O_2343,N_19856,N_19166);
or UO_2344 (O_2344,N_19726,N_24396);
nand UO_2345 (O_2345,N_21629,N_22928);
xnor UO_2346 (O_2346,N_22069,N_22826);
and UO_2347 (O_2347,N_22578,N_18859);
nand UO_2348 (O_2348,N_23763,N_21657);
and UO_2349 (O_2349,N_24086,N_19281);
nand UO_2350 (O_2350,N_18871,N_23365);
nand UO_2351 (O_2351,N_22384,N_22697);
and UO_2352 (O_2352,N_24523,N_23629);
nand UO_2353 (O_2353,N_24992,N_20642);
and UO_2354 (O_2354,N_20561,N_22890);
nand UO_2355 (O_2355,N_24295,N_20725);
xor UO_2356 (O_2356,N_23962,N_22593);
xor UO_2357 (O_2357,N_21847,N_18933);
nand UO_2358 (O_2358,N_20130,N_22499);
and UO_2359 (O_2359,N_20178,N_20209);
nand UO_2360 (O_2360,N_21577,N_20142);
nand UO_2361 (O_2361,N_22115,N_22198);
nand UO_2362 (O_2362,N_19103,N_21584);
or UO_2363 (O_2363,N_19165,N_21785);
xor UO_2364 (O_2364,N_21316,N_22539);
and UO_2365 (O_2365,N_21988,N_23803);
or UO_2366 (O_2366,N_23810,N_23907);
or UO_2367 (O_2367,N_23589,N_19335);
xor UO_2368 (O_2368,N_20339,N_19756);
or UO_2369 (O_2369,N_21764,N_19674);
nand UO_2370 (O_2370,N_19741,N_22887);
nand UO_2371 (O_2371,N_19326,N_22050);
or UO_2372 (O_2372,N_20576,N_20608);
nand UO_2373 (O_2373,N_23977,N_22105);
nand UO_2374 (O_2374,N_19862,N_22320);
nor UO_2375 (O_2375,N_20102,N_21491);
nor UO_2376 (O_2376,N_21968,N_22017);
nand UO_2377 (O_2377,N_20116,N_19418);
xnor UO_2378 (O_2378,N_20921,N_23554);
xnor UO_2379 (O_2379,N_23748,N_19139);
nand UO_2380 (O_2380,N_20149,N_20559);
xnor UO_2381 (O_2381,N_24875,N_19181);
or UO_2382 (O_2382,N_24470,N_21630);
xor UO_2383 (O_2383,N_24690,N_21334);
or UO_2384 (O_2384,N_19708,N_24632);
or UO_2385 (O_2385,N_18921,N_22412);
nor UO_2386 (O_2386,N_20282,N_23707);
xor UO_2387 (O_2387,N_22493,N_18774);
nor UO_2388 (O_2388,N_21222,N_22450);
or UO_2389 (O_2389,N_24225,N_21418);
and UO_2390 (O_2390,N_23825,N_21088);
nand UO_2391 (O_2391,N_20450,N_22223);
and UO_2392 (O_2392,N_19716,N_23692);
and UO_2393 (O_2393,N_24598,N_23883);
nor UO_2394 (O_2394,N_19387,N_24045);
nor UO_2395 (O_2395,N_22042,N_21288);
nand UO_2396 (O_2396,N_24639,N_24602);
and UO_2397 (O_2397,N_23974,N_21671);
or UO_2398 (O_2398,N_22324,N_21065);
nand UO_2399 (O_2399,N_21258,N_21973);
nand UO_2400 (O_2400,N_24824,N_20289);
xnor UO_2401 (O_2401,N_23447,N_23189);
and UO_2402 (O_2402,N_19696,N_20059);
xnor UO_2403 (O_2403,N_24555,N_19841);
xnor UO_2404 (O_2404,N_24780,N_22511);
nor UO_2405 (O_2405,N_23866,N_19063);
or UO_2406 (O_2406,N_22954,N_18936);
or UO_2407 (O_2407,N_19156,N_20794);
xnor UO_2408 (O_2408,N_24529,N_22352);
nor UO_2409 (O_2409,N_22581,N_18988);
xor UO_2410 (O_2410,N_20960,N_24143);
nor UO_2411 (O_2411,N_23018,N_19729);
xor UO_2412 (O_2412,N_24292,N_23193);
xnor UO_2413 (O_2413,N_22554,N_23620);
or UO_2414 (O_2414,N_19904,N_20131);
or UO_2415 (O_2415,N_24854,N_18855);
nand UO_2416 (O_2416,N_21749,N_24113);
and UO_2417 (O_2417,N_21623,N_21134);
xor UO_2418 (O_2418,N_18987,N_22628);
nand UO_2419 (O_2419,N_24926,N_21997);
nand UO_2420 (O_2420,N_19289,N_24586);
nor UO_2421 (O_2421,N_23678,N_22876);
xor UO_2422 (O_2422,N_20419,N_23727);
nor UO_2423 (O_2423,N_21889,N_24179);
or UO_2424 (O_2424,N_22832,N_18862);
and UO_2425 (O_2425,N_21501,N_24139);
and UO_2426 (O_2426,N_20614,N_18920);
and UO_2427 (O_2427,N_19813,N_23373);
and UO_2428 (O_2428,N_19360,N_24078);
or UO_2429 (O_2429,N_21291,N_20053);
or UO_2430 (O_2430,N_20792,N_20726);
or UO_2431 (O_2431,N_24312,N_24015);
and UO_2432 (O_2432,N_22815,N_24434);
xnor UO_2433 (O_2433,N_20715,N_21688);
nor UO_2434 (O_2434,N_20649,N_20135);
nand UO_2435 (O_2435,N_21783,N_22252);
nor UO_2436 (O_2436,N_22140,N_24416);
and UO_2437 (O_2437,N_19155,N_19412);
nor UO_2438 (O_2438,N_24399,N_24173);
xnor UO_2439 (O_2439,N_21036,N_23320);
xor UO_2440 (O_2440,N_19791,N_18798);
nor UO_2441 (O_2441,N_21057,N_19290);
and UO_2442 (O_2442,N_21274,N_19301);
or UO_2443 (O_2443,N_23435,N_20316);
nand UO_2444 (O_2444,N_23882,N_18966);
nand UO_2445 (O_2445,N_20495,N_23205);
or UO_2446 (O_2446,N_19738,N_20689);
nand UO_2447 (O_2447,N_22777,N_21081);
nor UO_2448 (O_2448,N_20631,N_19834);
or UO_2449 (O_2449,N_24375,N_24013);
nor UO_2450 (O_2450,N_23060,N_19996);
xnor UO_2451 (O_2451,N_23724,N_20549);
nor UO_2452 (O_2452,N_22574,N_24956);
xor UO_2453 (O_2453,N_21271,N_19818);
and UO_2454 (O_2454,N_21598,N_19524);
xor UO_2455 (O_2455,N_23693,N_23164);
nor UO_2456 (O_2456,N_19677,N_19889);
and UO_2457 (O_2457,N_24693,N_22619);
nor UO_2458 (O_2458,N_19385,N_23735);
xnor UO_2459 (O_2459,N_23108,N_22040);
nand UO_2460 (O_2460,N_20884,N_23351);
nand UO_2461 (O_2461,N_22073,N_22217);
nor UO_2462 (O_2462,N_24154,N_21842);
xnor UO_2463 (O_2463,N_20685,N_23150);
nor UO_2464 (O_2464,N_22806,N_24575);
or UO_2465 (O_2465,N_20016,N_24953);
nand UO_2466 (O_2466,N_20844,N_21022);
xor UO_2467 (O_2467,N_21994,N_19998);
nand UO_2468 (O_2468,N_19065,N_24750);
xnor UO_2469 (O_2469,N_20066,N_23969);
xnor UO_2470 (O_2470,N_19396,N_19439);
nand UO_2471 (O_2471,N_22183,N_24650);
nand UO_2472 (O_2472,N_20430,N_21982);
or UO_2473 (O_2473,N_19264,N_22899);
nor UO_2474 (O_2474,N_22702,N_19124);
and UO_2475 (O_2475,N_21546,N_23743);
and UO_2476 (O_2476,N_20027,N_24983);
or UO_2477 (O_2477,N_22727,N_23677);
and UO_2478 (O_2478,N_24230,N_22262);
nor UO_2479 (O_2479,N_21583,N_24280);
nor UO_2480 (O_2480,N_20797,N_20030);
xnor UO_2481 (O_2481,N_24754,N_18967);
xor UO_2482 (O_2482,N_19575,N_24360);
or UO_2483 (O_2483,N_20530,N_20381);
xor UO_2484 (O_2484,N_21905,N_21950);
xnor UO_2485 (O_2485,N_19319,N_19097);
nand UO_2486 (O_2486,N_23467,N_18990);
xnor UO_2487 (O_2487,N_24856,N_21168);
nor UO_2488 (O_2488,N_22354,N_19476);
nor UO_2489 (O_2489,N_20846,N_23125);
or UO_2490 (O_2490,N_19491,N_21465);
and UO_2491 (O_2491,N_19735,N_23414);
and UO_2492 (O_2492,N_22784,N_23862);
and UO_2493 (O_2493,N_20870,N_20241);
and UO_2494 (O_2494,N_20849,N_22924);
or UO_2495 (O_2495,N_20031,N_22188);
and UO_2496 (O_2496,N_24804,N_24505);
nand UO_2497 (O_2497,N_21285,N_20771);
nand UO_2498 (O_2498,N_21957,N_21098);
nor UO_2499 (O_2499,N_23451,N_20350);
nor UO_2500 (O_2500,N_22894,N_23568);
and UO_2501 (O_2501,N_22456,N_24325);
xor UO_2502 (O_2502,N_23066,N_24166);
and UO_2503 (O_2503,N_21094,N_19671);
nor UO_2504 (O_2504,N_23340,N_19901);
or UO_2505 (O_2505,N_22919,N_24307);
and UO_2506 (O_2506,N_18753,N_24595);
and UO_2507 (O_2507,N_19783,N_20643);
nor UO_2508 (O_2508,N_20512,N_22195);
nor UO_2509 (O_2509,N_23584,N_22182);
nor UO_2510 (O_2510,N_22775,N_24062);
nor UO_2511 (O_2511,N_21653,N_21421);
and UO_2512 (O_2512,N_19970,N_21205);
xor UO_2513 (O_2513,N_23466,N_22260);
nand UO_2514 (O_2514,N_23296,N_19012);
nand UO_2515 (O_2515,N_24662,N_23690);
nand UO_2516 (O_2516,N_20697,N_22604);
or UO_2517 (O_2517,N_23642,N_19454);
nand UO_2518 (O_2518,N_22859,N_19115);
xor UO_2519 (O_2519,N_21380,N_20961);
and UO_2520 (O_2520,N_20886,N_19897);
xor UO_2521 (O_2521,N_22373,N_19345);
xor UO_2522 (O_2522,N_23643,N_19225);
nand UO_2523 (O_2523,N_18915,N_24542);
nor UO_2524 (O_2524,N_24355,N_23243);
or UO_2525 (O_2525,N_22739,N_19755);
nand UO_2526 (O_2526,N_20362,N_24890);
nand UO_2527 (O_2527,N_22488,N_24637);
xor UO_2528 (O_2528,N_20975,N_21608);
and UO_2529 (O_2529,N_21227,N_19622);
xor UO_2530 (O_2530,N_20072,N_21239);
nand UO_2531 (O_2531,N_19458,N_24130);
nor UO_2532 (O_2532,N_24749,N_23600);
nand UO_2533 (O_2533,N_23559,N_21402);
nor UO_2534 (O_2534,N_21597,N_21824);
nor UO_2535 (O_2535,N_22021,N_24914);
nor UO_2536 (O_2536,N_23749,N_23122);
or UO_2537 (O_2537,N_21578,N_19210);
xnor UO_2538 (O_2538,N_19972,N_20411);
nor UO_2539 (O_2539,N_20630,N_19208);
nor UO_2540 (O_2540,N_21533,N_19404);
or UO_2541 (O_2541,N_21030,N_19703);
xor UO_2542 (O_2542,N_22959,N_20106);
nor UO_2543 (O_2543,N_23235,N_24007);
nand UO_2544 (O_2544,N_23955,N_23966);
xor UO_2545 (O_2545,N_24052,N_19002);
and UO_2546 (O_2546,N_18888,N_20647);
nor UO_2547 (O_2547,N_19159,N_21611);
xor UO_2548 (O_2548,N_23972,N_19049);
nand UO_2549 (O_2549,N_22941,N_23406);
and UO_2550 (O_2550,N_24545,N_19341);
xnor UO_2551 (O_2551,N_22674,N_23494);
or UO_2552 (O_2552,N_20307,N_21280);
nand UO_2553 (O_2553,N_20805,N_20161);
or UO_2554 (O_2554,N_24577,N_24801);
nor UO_2555 (O_2555,N_21508,N_22103);
or UO_2556 (O_2556,N_24950,N_24496);
or UO_2557 (O_2557,N_24802,N_24117);
or UO_2558 (O_2558,N_20417,N_19207);
nand UO_2559 (O_2559,N_19371,N_22386);
nand UO_2560 (O_2560,N_19955,N_20090);
nand UO_2561 (O_2561,N_23352,N_19113);
nor UO_2562 (O_2562,N_24379,N_24744);
xnor UO_2563 (O_2563,N_20716,N_20570);
and UO_2564 (O_2564,N_21375,N_21006);
or UO_2565 (O_2565,N_19104,N_19241);
or UO_2566 (O_2566,N_19773,N_22055);
nand UO_2567 (O_2567,N_19338,N_22003);
and UO_2568 (O_2568,N_19361,N_20589);
nand UO_2569 (O_2569,N_19993,N_23260);
nand UO_2570 (O_2570,N_24889,N_24656);
nor UO_2571 (O_2571,N_20722,N_22265);
nand UO_2572 (O_2572,N_23879,N_22224);
nand UO_2573 (O_2573,N_19125,N_23976);
or UO_2574 (O_2574,N_24000,N_22495);
and UO_2575 (O_2575,N_24196,N_24846);
nor UO_2576 (O_2576,N_24628,N_21737);
nor UO_2577 (O_2577,N_23531,N_24980);
and UO_2578 (O_2578,N_19923,N_23484);
or UO_2579 (O_2579,N_23660,N_20838);
or UO_2580 (O_2580,N_22376,N_19314);
or UO_2581 (O_2581,N_24990,N_19038);
nand UO_2582 (O_2582,N_21714,N_21049);
nor UO_2583 (O_2583,N_19196,N_19633);
and UO_2584 (O_2584,N_20323,N_24778);
and UO_2585 (O_2585,N_24235,N_19118);
xor UO_2586 (O_2586,N_22279,N_19117);
nor UO_2587 (O_2587,N_22852,N_23370);
nand UO_2588 (O_2588,N_21848,N_24960);
xor UO_2589 (O_2589,N_22653,N_22847);
xor UO_2590 (O_2590,N_24026,N_23013);
nor UO_2591 (O_2591,N_23758,N_23563);
nand UO_2592 (O_2592,N_19334,N_22642);
or UO_2593 (O_2593,N_24789,N_18949);
and UO_2594 (O_2594,N_22283,N_21745);
nor UO_2595 (O_2595,N_23453,N_19888);
xor UO_2596 (O_2596,N_19829,N_20878);
and UO_2597 (O_2597,N_23073,N_19395);
or UO_2598 (O_2598,N_22909,N_24486);
xor UO_2599 (O_2599,N_24917,N_21033);
nor UO_2600 (O_2600,N_23209,N_24842);
nand UO_2601 (O_2601,N_20640,N_19554);
nor UO_2602 (O_2602,N_24888,N_23119);
xor UO_2603 (O_2603,N_23850,N_24075);
xnor UO_2604 (O_2604,N_19256,N_23841);
and UO_2605 (O_2605,N_23720,N_24794);
nand UO_2606 (O_2606,N_23847,N_19785);
and UO_2607 (O_2607,N_19383,N_21336);
nand UO_2608 (O_2608,N_24725,N_22294);
xnor UO_2609 (O_2609,N_22155,N_19461);
nor UO_2610 (O_2610,N_24688,N_20438);
nor UO_2611 (O_2611,N_19990,N_20666);
nor UO_2612 (O_2612,N_23766,N_18910);
nand UO_2613 (O_2613,N_22316,N_19715);
or UO_2614 (O_2614,N_19144,N_20183);
nand UO_2615 (O_2615,N_20872,N_22221);
xnor UO_2616 (O_2616,N_23446,N_20592);
xnor UO_2617 (O_2617,N_24345,N_19434);
xor UO_2618 (O_2618,N_21162,N_21556);
nor UO_2619 (O_2619,N_20742,N_19682);
nand UO_2620 (O_2620,N_22151,N_23694);
nor UO_2621 (O_2621,N_23347,N_24800);
and UO_2622 (O_2622,N_19589,N_21158);
nand UO_2623 (O_2623,N_20224,N_19133);
xor UO_2624 (O_2624,N_20688,N_23228);
nand UO_2625 (O_2625,N_19191,N_20724);
nand UO_2626 (O_2626,N_19007,N_21000);
xor UO_2627 (O_2627,N_24242,N_21459);
xor UO_2628 (O_2628,N_24720,N_22389);
and UO_2629 (O_2629,N_19342,N_22433);
nand UO_2630 (O_2630,N_21572,N_19209);
and UO_2631 (O_2631,N_22093,N_23975);
xor UO_2632 (O_2632,N_24164,N_22271);
and UO_2633 (O_2633,N_21412,N_20822);
and UO_2634 (O_2634,N_23648,N_20468);
or UO_2635 (O_2635,N_21738,N_20218);
xor UO_2636 (O_2636,N_21237,N_23398);
or UO_2637 (O_2637,N_24793,N_23580);
nand UO_2638 (O_2638,N_22985,N_21159);
nand UO_2639 (O_2639,N_21201,N_23281);
nand UO_2640 (O_2640,N_23780,N_19217);
and UO_2641 (O_2641,N_21384,N_19793);
nand UO_2642 (O_2642,N_23395,N_23543);
and UO_2643 (O_2643,N_23314,N_19247);
and UO_2644 (O_2644,N_23754,N_19240);
nand UO_2645 (O_2645,N_20712,N_20777);
and UO_2646 (O_2646,N_18951,N_20543);
or UO_2647 (O_2647,N_20607,N_20296);
xor UO_2648 (O_2648,N_23881,N_22670);
and UO_2649 (O_2649,N_24435,N_21377);
nand UO_2650 (O_2650,N_22882,N_22186);
xnor UO_2651 (O_2651,N_20203,N_20005);
nand UO_2652 (O_2652,N_19562,N_22667);
or UO_2653 (O_2653,N_22738,N_24246);
or UO_2654 (O_2654,N_20451,N_24304);
and UO_2655 (O_2655,N_19784,N_24812);
nand UO_2656 (O_2656,N_24684,N_20044);
and UO_2657 (O_2657,N_19795,N_20952);
nand UO_2658 (O_2658,N_23407,N_19640);
or UO_2659 (O_2659,N_21051,N_22989);
and UO_2660 (O_2660,N_24212,N_24768);
nor UO_2661 (O_2661,N_21976,N_23687);
or UO_2662 (O_2662,N_22244,N_20897);
or UO_2663 (O_2663,N_22761,N_19470);
nand UO_2664 (O_2664,N_21479,N_23567);
xnor UO_2665 (O_2665,N_24270,N_21666);
xor UO_2666 (O_2666,N_20083,N_21460);
nand UO_2667 (O_2667,N_23354,N_23980);
and UO_2668 (O_2668,N_21256,N_22506);
and UO_2669 (O_2669,N_20899,N_18870);
or UO_2670 (O_2670,N_24967,N_24347);
and UO_2671 (O_2671,N_19576,N_20396);
nor UO_2672 (O_2672,N_19973,N_20380);
nor UO_2673 (O_2673,N_19704,N_19109);
and UO_2674 (O_2674,N_19252,N_19688);
xor UO_2675 (O_2675,N_21442,N_20980);
and UO_2676 (O_2676,N_24597,N_18761);
xor UO_2677 (O_2677,N_20823,N_20399);
and UO_2678 (O_2678,N_19143,N_24912);
or UO_2679 (O_2679,N_22145,N_22782);
nor UO_2680 (O_2680,N_20483,N_20384);
and UO_2681 (O_2681,N_24858,N_24558);
nor UO_2682 (O_2682,N_20953,N_19162);
nand UO_2683 (O_2683,N_20342,N_19483);
xnor UO_2684 (O_2684,N_19282,N_23055);
nand UO_2685 (O_2685,N_20322,N_24904);
nor UO_2686 (O_2686,N_23167,N_19323);
nand UO_2687 (O_2687,N_21090,N_19223);
nor UO_2688 (O_2688,N_23834,N_21651);
nand UO_2689 (O_2689,N_20270,N_24222);
nand UO_2690 (O_2690,N_24228,N_23641);
and UO_2691 (O_2691,N_24201,N_22854);
or UO_2692 (O_2692,N_21685,N_19021);
nand UO_2693 (O_2693,N_20182,N_20723);
nand UO_2694 (O_2694,N_21028,N_19655);
or UO_2695 (O_2695,N_24916,N_20499);
nand UO_2696 (O_2696,N_19033,N_24699);
or UO_2697 (O_2697,N_19917,N_23254);
and UO_2698 (O_2698,N_18780,N_22436);
xnor UO_2699 (O_2699,N_22681,N_24658);
xor UO_2700 (O_2700,N_18752,N_24618);
or UO_2701 (O_2701,N_19221,N_22087);
nand UO_2702 (O_2702,N_19651,N_22644);
and UO_2703 (O_2703,N_23511,N_20395);
xnor UO_2704 (O_2704,N_23729,N_19550);
and UO_2705 (O_2705,N_24232,N_21757);
xor UO_2706 (O_2706,N_21908,N_23123);
xor UO_2707 (O_2707,N_23389,N_22227);
and UO_2708 (O_2708,N_21703,N_23104);
xor UO_2709 (O_2709,N_20354,N_19526);
or UO_2710 (O_2710,N_23742,N_21678);
nand UO_2711 (O_2711,N_20817,N_21177);
and UO_2712 (O_2712,N_23552,N_22591);
nor UO_2713 (O_2713,N_23183,N_22635);
or UO_2714 (O_2714,N_18795,N_20120);
nor UO_2715 (O_2715,N_21009,N_22016);
and UO_2716 (O_2716,N_23107,N_20371);
xor UO_2717 (O_2717,N_20714,N_20783);
or UO_2718 (O_2718,N_18831,N_21228);
nor UO_2719 (O_2719,N_19943,N_22544);
or UO_2720 (O_2720,N_23896,N_19675);
and UO_2721 (O_2721,N_19992,N_24638);
and UO_2722 (O_2722,N_24831,N_19925);
xor UO_2723 (O_2723,N_19157,N_24682);
and UO_2724 (O_2724,N_20907,N_24258);
nor UO_2725 (O_2725,N_20525,N_22418);
or UO_2726 (O_2726,N_20157,N_22943);
nor UO_2727 (O_2727,N_19486,N_19769);
xnor UO_2728 (O_2728,N_21528,N_22213);
xor UO_2729 (O_2729,N_23360,N_19895);
nand UO_2730 (O_2730,N_21958,N_23918);
or UO_2731 (O_2731,N_23981,N_20087);
or UO_2732 (O_2732,N_24018,N_22305);
and UO_2733 (O_2733,N_21107,N_19939);
or UO_2734 (O_2734,N_23503,N_19279);
or UO_2735 (O_2735,N_21771,N_22091);
and UO_2736 (O_2736,N_22163,N_24445);
nand UO_2737 (O_2737,N_21429,N_18821);
nand UO_2738 (O_2738,N_19058,N_18940);
nor UO_2739 (O_2739,N_19293,N_19570);
nor UO_2740 (O_2740,N_20346,N_23808);
and UO_2741 (O_2741,N_21986,N_23884);
nand UO_2742 (O_2742,N_23522,N_23229);
nor UO_2743 (O_2743,N_19480,N_22503);
nand UO_2744 (O_2744,N_23771,N_22111);
or UO_2745 (O_2745,N_21482,N_20675);
and UO_2746 (O_2746,N_22166,N_22239);
nor UO_2747 (O_2747,N_23290,N_23411);
or UO_2748 (O_2748,N_21249,N_19112);
and UO_2749 (O_2749,N_21252,N_19205);
and UO_2750 (O_2750,N_24265,N_21130);
nor UO_2751 (O_2751,N_19648,N_21013);
or UO_2752 (O_2752,N_20352,N_19552);
nor UO_2753 (O_2753,N_20293,N_20117);
and UO_2754 (O_2754,N_19185,N_23549);
nand UO_2755 (O_2755,N_22870,N_21735);
and UO_2756 (O_2756,N_23782,N_21244);
nand UO_2757 (O_2757,N_19022,N_23316);
nor UO_2758 (O_2758,N_21230,N_18785);
nand UO_2759 (O_2759,N_19938,N_22907);
nand UO_2760 (O_2760,N_23457,N_24588);
nand UO_2761 (O_2761,N_24681,N_18874);
nor UO_2762 (O_2762,N_22015,N_19379);
nand UO_2763 (O_2763,N_21538,N_22974);
and UO_2764 (O_2764,N_20905,N_24031);
nand UO_2765 (O_2765,N_19362,N_24466);
or UO_2766 (O_2766,N_24783,N_19699);
nor UO_2767 (O_2767,N_21955,N_21361);
and UO_2768 (O_2768,N_23343,N_21099);
or UO_2769 (O_2769,N_22562,N_19900);
nor UO_2770 (O_2770,N_20147,N_24132);
or UO_2771 (O_2771,N_23231,N_18822);
or UO_2772 (O_2772,N_22120,N_19076);
and UO_2773 (O_2773,N_19837,N_22751);
xnor UO_2774 (O_2774,N_22192,N_21148);
xor UO_2775 (O_2775,N_20703,N_19778);
or UO_2776 (O_2776,N_21175,N_22409);
nand UO_2777 (O_2777,N_24543,N_24108);
or UO_2778 (O_2778,N_21169,N_18931);
nor UO_2779 (O_2779,N_20048,N_24380);
nor UO_2780 (O_2780,N_23719,N_24817);
or UO_2781 (O_2781,N_24852,N_21560);
xnor UO_2782 (O_2782,N_23548,N_21039);
nor UO_2783 (O_2783,N_21537,N_21221);
nor UO_2784 (O_2784,N_24979,N_19839);
or UO_2785 (O_2785,N_21805,N_24459);
nand UO_2786 (O_2786,N_22839,N_21093);
xnor UO_2787 (O_2787,N_23532,N_21243);
or UO_2788 (O_2788,N_22973,N_22528);
or UO_2789 (O_2789,N_18929,N_21155);
or UO_2790 (O_2790,N_21931,N_21360);
xor UO_2791 (O_2791,N_21197,N_19427);
and UO_2792 (O_2792,N_22097,N_24668);
nor UO_2793 (O_2793,N_19511,N_23000);
nor UO_2794 (O_2794,N_24423,N_22805);
xnor UO_2795 (O_2795,N_19634,N_21812);
nor UO_2796 (O_2796,N_21717,N_21967);
xor UO_2797 (O_2797,N_23715,N_23299);
nand UO_2798 (O_2798,N_19102,N_20908);
or UO_2799 (O_2799,N_24604,N_23216);
nand UO_2800 (O_2800,N_20192,N_22792);
and UO_2801 (O_2801,N_18883,N_20383);
xor UO_2802 (O_2802,N_22167,N_23199);
and UO_2803 (O_2803,N_19310,N_21664);
or UO_2804 (O_2804,N_22146,N_23302);
xor UO_2805 (O_2805,N_21626,N_24150);
and UO_2806 (O_2806,N_24859,N_21011);
and UO_2807 (O_2807,N_23785,N_21136);
or UO_2808 (O_2808,N_22078,N_18953);
or UO_2809 (O_2809,N_23656,N_20678);
or UO_2810 (O_2810,N_21633,N_19705);
nand UO_2811 (O_2811,N_24419,N_20253);
or UO_2812 (O_2812,N_21270,N_24096);
and UO_2813 (O_2813,N_19071,N_19372);
xor UO_2814 (O_2814,N_24803,N_23487);
xnor UO_2815 (O_2815,N_24303,N_22953);
and UO_2816 (O_2816,N_19790,N_19275);
nand UO_2817 (O_2817,N_23067,N_22169);
or UO_2818 (O_2818,N_23556,N_20996);
or UO_2819 (O_2819,N_19753,N_24464);
xnor UO_2820 (O_2820,N_23011,N_24605);
nor UO_2821 (O_2821,N_21135,N_24704);
nand UO_2822 (O_2822,N_19878,N_24491);
or UO_2823 (O_2823,N_24580,N_20392);
nand UO_2824 (O_2824,N_23595,N_20444);
and UO_2825 (O_2825,N_19403,N_20288);
or UO_2826 (O_2826,N_20086,N_21725);
nor UO_2827 (O_2827,N_22160,N_23603);
nor UO_2828 (O_2828,N_22337,N_19478);
nand UO_2829 (O_2829,N_20602,N_23141);
or UO_2830 (O_2830,N_22287,N_24205);
nor UO_2831 (O_2831,N_24156,N_22857);
or UO_2832 (O_2832,N_22248,N_19436);
or UO_2833 (O_2833,N_20348,N_20828);
or UO_2834 (O_2834,N_24676,N_21786);
and UO_2835 (O_2835,N_20594,N_23876);
nor UO_2836 (O_2836,N_22756,N_23306);
xor UO_2837 (O_2837,N_24403,N_21589);
or UO_2838 (O_2838,N_22736,N_20638);
nor UO_2839 (O_2839,N_18793,N_18794);
nand UO_2840 (O_2840,N_22701,N_21529);
and UO_2841 (O_2841,N_20492,N_24738);
xnor UO_2842 (O_2842,N_20865,N_19452);
nand UO_2843 (O_2843,N_24107,N_23571);
nor UO_2844 (O_2844,N_23575,N_22966);
and UO_2845 (O_2845,N_24176,N_20284);
or UO_2846 (O_2846,N_22559,N_20337);
nor UO_2847 (O_2847,N_22435,N_19604);
nand UO_2848 (O_2848,N_21008,N_24549);
nand UO_2849 (O_2849,N_21428,N_22618);
nor UO_2850 (O_2850,N_20741,N_22576);
or UO_2851 (O_2851,N_22698,N_19933);
nor UO_2852 (O_2852,N_20173,N_20101);
and UO_2853 (O_2853,N_20334,N_24152);
nand UO_2854 (O_2854,N_22296,N_23363);
and UO_2855 (O_2855,N_18983,N_20390);
xor UO_2856 (O_2856,N_19787,N_24787);
nor UO_2857 (O_2857,N_20338,N_24438);
xor UO_2858 (O_2858,N_21863,N_24724);
or UO_2859 (O_2859,N_22346,N_20240);
nor UO_2860 (O_2860,N_23171,N_22713);
and UO_2861 (O_2861,N_21860,N_24053);
and UO_2862 (O_2862,N_23409,N_21639);
or UO_2863 (O_2863,N_22193,N_23833);
and UO_2864 (O_2864,N_21167,N_23237);
nor UO_2865 (O_2865,N_22443,N_24433);
and UO_2866 (O_2866,N_22722,N_22659);
xnor UO_2867 (O_2867,N_19859,N_22946);
or UO_2868 (O_2868,N_22682,N_24033);
nor UO_2869 (O_2869,N_22600,N_20088);
and UO_2870 (O_2870,N_19401,N_23130);
xnor UO_2871 (O_2871,N_22147,N_19906);
nand UO_2872 (O_2872,N_19266,N_20556);
and UO_2873 (O_2873,N_19935,N_23025);
or UO_2874 (O_2874,N_23476,N_21740);
nand UO_2875 (O_2875,N_23048,N_21619);
nand UO_2876 (O_2876,N_19201,N_22529);
nand UO_2877 (O_2877,N_19739,N_20744);
or UO_2878 (O_2878,N_19953,N_23857);
or UO_2879 (O_2879,N_19059,N_22520);
and UO_2880 (O_2880,N_20552,N_23601);
or UO_2881 (O_2881,N_20234,N_24335);
nand UO_2882 (O_2882,N_22862,N_19845);
or UO_2883 (O_2883,N_20588,N_21503);
nor UO_2884 (O_2884,N_24359,N_21312);
nor UO_2885 (O_2885,N_24463,N_21996);
or UO_2886 (O_2886,N_23493,N_20858);
or UO_2887 (O_2887,N_23610,N_24344);
nor UO_2888 (O_2888,N_22353,N_20267);
and UO_2889 (O_2889,N_22288,N_22987);
and UO_2890 (O_2890,N_21404,N_20820);
or UO_2891 (O_2891,N_23911,N_18813);
nor UO_2892 (O_2892,N_19687,N_20366);
nor UO_2893 (O_2893,N_19629,N_22688);
and UO_2894 (O_2894,N_21650,N_20259);
nand UO_2895 (O_2895,N_20445,N_23714);
or UO_2896 (O_2896,N_19414,N_20940);
or UO_2897 (O_2897,N_18905,N_22006);
or UO_2898 (O_2898,N_23612,N_22950);
and UO_2899 (O_2899,N_24551,N_20360);
xor UO_2900 (O_2900,N_20414,N_22404);
or UO_2901 (O_2901,N_24767,N_23705);
and UO_2902 (O_2902,N_24482,N_24037);
or UO_2903 (O_2903,N_24322,N_20489);
nand UO_2904 (O_2904,N_24565,N_23774);
and UO_2905 (O_2905,N_24479,N_21605);
or UO_2906 (O_2906,N_21951,N_22597);
xnor UO_2907 (O_2907,N_23602,N_24530);
or UO_2908 (O_2908,N_21791,N_22990);
nor UO_2909 (O_2909,N_20128,N_23805);
or UO_2910 (O_2910,N_20694,N_19512);
or UO_2911 (O_2911,N_19433,N_22866);
or UO_2912 (O_2912,N_21431,N_21454);
xnor UO_2913 (O_2913,N_24834,N_22184);
nand UO_2914 (O_2914,N_22561,N_20700);
nand UO_2915 (O_2915,N_21654,N_22510);
and UO_2916 (O_2916,N_21410,N_24607);
xnor UO_2917 (O_2917,N_22076,N_23286);
xnor UO_2918 (O_2918,N_21660,N_21823);
nor UO_2919 (O_2919,N_20696,N_21962);
or UO_2920 (O_2920,N_24299,N_22631);
nand UO_2921 (O_2921,N_21960,N_20992);
or UO_2922 (O_2922,N_19138,N_20431);
nor UO_2923 (O_2923,N_21551,N_19833);
xnor UO_2924 (O_2924,N_24813,N_20815);
or UO_2925 (O_2925,N_23400,N_19078);
and UO_2926 (O_2926,N_21568,N_19234);
nand UO_2927 (O_2927,N_20460,N_24927);
xnor UO_2928 (O_2928,N_21741,N_22747);
nor UO_2929 (O_2929,N_24879,N_23928);
or UO_2930 (O_2930,N_24455,N_19694);
xnor UO_2931 (O_2931,N_21048,N_19011);
and UO_2932 (O_2932,N_21333,N_21219);
and UO_2933 (O_2933,N_22206,N_19721);
nand UO_2934 (O_2934,N_24453,N_23662);
nor UO_2935 (O_2935,N_24719,N_23440);
xor UO_2936 (O_2936,N_22238,N_22613);
and UO_2937 (O_2937,N_20964,N_21614);
or UO_2938 (O_2938,N_24673,N_23528);
nand UO_2939 (O_2939,N_24080,N_19026);
nand UO_2940 (O_2940,N_21964,N_24678);
or UO_2941 (O_2941,N_20665,N_20894);
xor UO_2942 (O_2942,N_23362,N_24036);
nand UO_2943 (O_2943,N_19610,N_20114);
or UO_2944 (O_2944,N_19045,N_21014);
or UO_2945 (O_2945,N_20927,N_21998);
nand UO_2946 (O_2946,N_21622,N_22207);
and UO_2947 (O_2947,N_20146,N_20933);
nor UO_2948 (O_2948,N_23606,N_23147);
nand UO_2949 (O_2949,N_22601,N_20997);
xnor UO_2950 (O_2950,N_24064,N_20746);
nand UO_2951 (O_2951,N_20042,N_19762);
or UO_2952 (O_2952,N_22392,N_18848);
and UO_2953 (O_2953,N_20421,N_24952);
nand UO_2954 (O_2954,N_21829,N_23034);
or UO_2955 (O_2955,N_21085,N_23811);
nor UO_2956 (O_2956,N_22036,N_19789);
nand UO_2957 (O_2957,N_20035,N_19559);
and UO_2958 (O_2958,N_20422,N_23914);
or UO_2959 (O_2959,N_20924,N_24194);
and UO_2960 (O_2960,N_20691,N_22397);
nor UO_2961 (O_2961,N_20404,N_20968);
and UO_2962 (O_2962,N_23008,N_20425);
and UO_2963 (O_2963,N_22609,N_21601);
xnor UO_2964 (O_2964,N_20251,N_22171);
nor UO_2965 (O_2965,N_21397,N_22804);
nand UO_2966 (O_2966,N_20757,N_22588);
and UO_2967 (O_2967,N_21953,N_22214);
nor UO_2968 (O_2968,N_23160,N_23764);
and UO_2969 (O_2969,N_19728,N_20625);
or UO_2970 (O_2970,N_21715,N_24278);
xor UO_2971 (O_2971,N_19299,N_21803);
nor UO_2972 (O_2972,N_21711,N_21163);
nor UO_2973 (O_2973,N_20967,N_19353);
or UO_2974 (O_2974,N_20482,N_22302);
and UO_2975 (O_2975,N_19968,N_22474);
nand UO_2976 (O_2976,N_22068,N_21171);
nor UO_2977 (O_2977,N_24843,N_24067);
nand UO_2978 (O_2978,N_24512,N_19179);
nand UO_2979 (O_2979,N_21881,N_22347);
nand UO_2980 (O_2980,N_18963,N_24384);
and UO_2981 (O_2981,N_23651,N_22791);
xor UO_2982 (O_2982,N_22787,N_21118);
xor UO_2983 (O_2983,N_24105,N_24182);
or UO_2984 (O_2984,N_21257,N_24617);
xor UO_2985 (O_2985,N_22201,N_23697);
or UO_2986 (O_2986,N_18772,N_19407);
or UO_2987 (O_2987,N_24374,N_24348);
nand UO_2988 (O_2988,N_23773,N_19230);
xor UO_2989 (O_2989,N_22754,N_23027);
or UO_2990 (O_2990,N_24428,N_21012);
or UO_2991 (O_2991,N_23789,N_23959);
or UO_2992 (O_2992,N_20962,N_24060);
nor UO_2993 (O_2993,N_24517,N_22112);
xor UO_2994 (O_2994,N_23390,N_22459);
xnor UO_2995 (O_2995,N_22583,N_24948);
and UO_2996 (O_2996,N_21880,N_24104);
nor UO_2997 (O_2997,N_23050,N_20599);
and UO_2998 (O_2998,N_24163,N_21831);
or UO_2999 (O_2999,N_19500,N_21620);
endmodule