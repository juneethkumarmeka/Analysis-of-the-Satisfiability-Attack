module basic_1000_10000_1500_4_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_758,In_192);
nor U1 (N_1,In_68,In_984);
xnor U2 (N_2,In_342,In_165);
nor U3 (N_3,In_975,In_627);
xor U4 (N_4,In_249,In_147);
xor U5 (N_5,In_177,In_209);
xor U6 (N_6,In_44,In_136);
or U7 (N_7,In_576,In_22);
or U8 (N_8,In_74,In_294);
nand U9 (N_9,In_2,In_940);
or U10 (N_10,In_614,In_795);
nand U11 (N_11,In_461,In_775);
and U12 (N_12,In_547,In_183);
and U13 (N_13,In_536,In_782);
nor U14 (N_14,In_145,In_935);
nand U15 (N_15,In_986,In_685);
or U16 (N_16,In_270,In_252);
nand U17 (N_17,In_699,In_419);
and U18 (N_18,In_691,In_288);
xor U19 (N_19,In_251,In_752);
nand U20 (N_20,In_289,In_222);
and U21 (N_21,In_965,In_428);
nand U22 (N_22,In_989,In_828);
and U23 (N_23,In_676,In_92);
nor U24 (N_24,In_854,In_396);
xnor U25 (N_25,In_861,In_196);
nand U26 (N_26,In_742,In_526);
xor U27 (N_27,In_510,In_487);
and U28 (N_28,In_736,In_615);
nor U29 (N_29,In_149,In_331);
or U30 (N_30,In_114,In_408);
nand U31 (N_31,In_882,In_358);
xor U32 (N_32,In_519,In_592);
and U33 (N_33,In_725,In_416);
nor U34 (N_34,In_640,In_99);
or U35 (N_35,In_637,In_470);
and U36 (N_36,In_52,In_215);
nor U37 (N_37,In_456,In_613);
and U38 (N_38,In_807,In_449);
nor U39 (N_39,In_108,In_537);
and U40 (N_40,In_923,In_697);
nand U41 (N_41,In_818,In_115);
xor U42 (N_42,In_268,In_674);
or U43 (N_43,In_219,In_385);
or U44 (N_44,In_892,In_663);
xnor U45 (N_45,In_822,In_609);
and U46 (N_46,In_857,In_650);
xor U47 (N_47,In_148,In_469);
nor U48 (N_48,In_79,In_798);
xnor U49 (N_49,In_790,In_363);
or U50 (N_50,In_37,In_851);
xnor U51 (N_51,In_178,In_741);
nor U52 (N_52,In_228,In_435);
nor U53 (N_53,In_998,In_506);
nor U54 (N_54,In_937,In_426);
or U55 (N_55,In_922,In_284);
nor U56 (N_56,In_31,In_242);
nor U57 (N_57,In_184,In_625);
or U58 (N_58,In_57,In_719);
or U59 (N_59,In_356,In_459);
and U60 (N_60,In_981,In_554);
or U61 (N_61,In_866,In_71);
and U62 (N_62,In_948,In_66);
nand U63 (N_63,In_722,In_217);
nor U64 (N_64,In_744,In_560);
or U65 (N_65,In_163,In_360);
and U66 (N_66,In_233,In_583);
nor U67 (N_67,In_375,In_6);
nand U68 (N_68,In_75,In_934);
nand U69 (N_69,In_415,In_943);
nand U70 (N_70,In_716,In_496);
or U71 (N_71,In_636,In_684);
and U72 (N_72,In_307,In_82);
xnor U73 (N_73,In_767,In_491);
nor U74 (N_74,In_983,In_831);
nand U75 (N_75,In_900,In_460);
or U76 (N_76,In_9,In_917);
nor U77 (N_77,In_710,In_626);
and U78 (N_78,In_422,In_195);
nand U79 (N_79,In_689,In_484);
nand U80 (N_80,In_25,In_817);
nand U81 (N_81,In_881,In_885);
nor U82 (N_82,In_462,In_988);
xor U83 (N_83,In_81,In_172);
nor U84 (N_84,In_387,In_84);
nor U85 (N_85,In_316,In_11);
nand U86 (N_86,In_494,In_672);
nand U87 (N_87,In_970,In_380);
nor U88 (N_88,In_997,In_378);
and U89 (N_89,In_811,In_906);
and U90 (N_90,In_607,In_117);
or U91 (N_91,In_440,In_389);
xnor U92 (N_92,In_777,In_14);
and U93 (N_93,In_991,In_62);
or U94 (N_94,In_540,In_438);
and U95 (N_95,In_764,In_507);
xnor U96 (N_96,In_442,In_413);
nand U97 (N_97,In_19,In_182);
nor U98 (N_98,In_179,In_221);
or U99 (N_99,In_829,In_443);
or U100 (N_100,In_437,In_271);
nor U101 (N_101,In_224,In_355);
and U102 (N_102,In_478,In_170);
nand U103 (N_103,In_545,In_635);
nand U104 (N_104,In_393,In_314);
or U105 (N_105,In_33,In_175);
xnor U106 (N_106,In_567,In_553);
nand U107 (N_107,In_214,In_717);
xor U108 (N_108,In_283,In_971);
nand U109 (N_109,In_60,In_620);
and U110 (N_110,In_898,In_928);
or U111 (N_111,In_420,In_573);
nand U112 (N_112,In_237,In_511);
and U113 (N_113,In_152,In_612);
nand U114 (N_114,In_543,In_471);
nor U115 (N_115,In_611,In_504);
nor U116 (N_116,In_598,In_982);
nor U117 (N_117,In_464,In_911);
nand U118 (N_118,In_712,In_977);
nand U119 (N_119,In_80,In_968);
nor U120 (N_120,In_141,In_391);
or U121 (N_121,In_439,In_869);
and U122 (N_122,In_867,In_606);
nand U123 (N_123,In_958,In_649);
nand U124 (N_124,In_772,In_601);
or U125 (N_125,In_913,In_564);
or U126 (N_126,In_246,In_571);
nand U127 (N_127,In_30,In_563);
and U128 (N_128,In_847,In_3);
and U129 (N_129,In_18,In_253);
or U130 (N_130,In_97,In_293);
and U131 (N_131,In_967,In_580);
nor U132 (N_132,In_814,In_201);
and U133 (N_133,In_93,In_453);
or U134 (N_134,In_131,In_198);
or U135 (N_135,In_445,In_599);
or U136 (N_136,In_944,In_28);
or U137 (N_137,In_993,In_315);
nor U138 (N_138,In_244,In_529);
or U139 (N_139,In_96,In_879);
nor U140 (N_140,In_451,In_204);
or U141 (N_141,In_846,In_575);
nor U142 (N_142,In_341,In_357);
nand U143 (N_143,In_952,In_208);
and U144 (N_144,In_207,In_29);
nand U145 (N_145,In_538,In_946);
or U146 (N_146,In_267,In_234);
or U147 (N_147,In_150,In_568);
or U148 (N_148,In_347,In_77);
xor U149 (N_149,In_698,In_433);
nand U150 (N_150,In_844,In_258);
and U151 (N_151,In_833,In_572);
nor U152 (N_152,In_754,In_48);
nand U153 (N_153,In_38,In_274);
or U154 (N_154,In_43,In_738);
xor U155 (N_155,In_476,In_327);
nand U156 (N_156,In_513,In_457);
or U157 (N_157,In_305,In_12);
nor U158 (N_158,In_371,In_779);
nor U159 (N_159,In_739,In_299);
and U160 (N_160,In_951,In_978);
or U161 (N_161,In_671,In_144);
and U162 (N_162,In_735,In_254);
nor U163 (N_163,In_713,In_47);
nand U164 (N_164,In_969,In_718);
or U165 (N_165,In_59,In_585);
and U166 (N_166,In_154,In_746);
nand U167 (N_167,In_843,In_326);
and U168 (N_168,In_776,In_231);
or U169 (N_169,In_696,In_365);
nor U170 (N_170,In_499,In_990);
and U171 (N_171,In_191,In_781);
and U172 (N_172,In_412,In_463);
and U173 (N_173,In_105,In_905);
and U174 (N_174,In_54,In_518);
or U175 (N_175,In_311,In_185);
nand U176 (N_176,In_939,In_799);
and U177 (N_177,In_107,In_87);
or U178 (N_178,In_683,In_303);
or U179 (N_179,In_794,In_109);
nand U180 (N_180,In_864,In_956);
nand U181 (N_181,In_600,In_964);
and U182 (N_182,In_474,In_199);
nor U183 (N_183,In_455,In_862);
and U184 (N_184,In_999,In_651);
nor U185 (N_185,In_353,In_382);
xnor U186 (N_186,In_830,In_160);
and U187 (N_187,In_995,In_0);
or U188 (N_188,In_797,In_664);
nor U189 (N_189,In_628,In_826);
and U190 (N_190,In_394,In_584);
nand U191 (N_191,In_174,In_840);
nand U192 (N_192,In_525,In_473);
and U193 (N_193,In_921,In_229);
nand U194 (N_194,In_367,In_240);
nand U195 (N_195,In_912,In_677);
or U196 (N_196,In_961,In_836);
or U197 (N_197,In_317,In_669);
or U198 (N_198,In_559,In_83);
xor U199 (N_199,In_421,In_594);
or U200 (N_200,In_446,In_813);
nor U201 (N_201,In_69,In_51);
and U202 (N_202,In_791,In_390);
nand U203 (N_203,In_424,In_101);
nand U204 (N_204,In_726,In_119);
and U205 (N_205,In_523,In_304);
nand U206 (N_206,In_757,In_220);
or U207 (N_207,In_42,In_629);
nor U208 (N_208,In_528,In_414);
or U209 (N_209,In_659,In_550);
or U210 (N_210,In_116,In_743);
or U211 (N_211,In_227,In_643);
nor U212 (N_212,In_835,In_269);
nor U213 (N_213,In_399,In_361);
or U214 (N_214,In_732,In_740);
xor U215 (N_215,In_280,In_359);
nor U216 (N_216,In_548,In_23);
nand U217 (N_217,In_78,In_909);
nand U218 (N_218,In_624,In_168);
or U219 (N_219,In_789,In_665);
or U220 (N_220,In_296,In_134);
and U221 (N_221,In_448,In_91);
and U222 (N_222,In_475,In_276);
and U223 (N_223,In_401,In_26);
nand U224 (N_224,In_994,In_318);
or U225 (N_225,In_860,In_747);
or U226 (N_226,In_953,In_329);
or U227 (N_227,In_434,In_723);
xor U228 (N_228,In_950,In_886);
xor U229 (N_229,In_495,In_655);
and U230 (N_230,In_549,In_656);
nand U231 (N_231,In_404,In_157);
nand U232 (N_232,In_260,In_652);
nand U233 (N_233,In_588,In_281);
nand U234 (N_234,In_825,In_200);
nand U235 (N_235,In_527,In_121);
nor U236 (N_236,In_302,In_662);
nor U237 (N_237,In_515,In_870);
nor U238 (N_238,In_95,In_631);
and U239 (N_239,In_187,In_858);
xnor U240 (N_240,In_570,In_633);
or U241 (N_241,In_605,In_126);
or U242 (N_242,In_880,In_45);
xnor U243 (N_243,In_481,In_241);
or U244 (N_244,In_945,In_444);
and U245 (N_245,In_376,In_647);
xor U246 (N_246,In_773,In_748);
nor U247 (N_247,In_872,In_16);
xor U248 (N_248,In_369,In_153);
nor U249 (N_249,In_402,In_771);
nand U250 (N_250,In_122,In_286);
or U251 (N_251,In_729,In_661);
and U252 (N_252,In_522,In_930);
nor U253 (N_253,In_158,In_705);
and U254 (N_254,In_841,In_151);
nand U255 (N_255,In_32,In_236);
or U256 (N_256,In_323,In_714);
or U257 (N_257,In_340,In_730);
xor U258 (N_258,In_203,In_348);
or U259 (N_259,In_766,In_125);
and U260 (N_260,In_50,In_164);
and U261 (N_261,In_245,In_534);
and U262 (N_262,In_63,In_188);
nand U263 (N_263,In_155,In_731);
nand U264 (N_264,In_64,In_780);
nand U265 (N_265,In_194,In_992);
and U266 (N_266,In_432,In_763);
nand U267 (N_267,In_985,In_56);
and U268 (N_268,In_497,In_889);
or U269 (N_269,In_875,In_143);
nand U270 (N_270,In_602,In_384);
and U271 (N_271,In_819,In_654);
and U272 (N_272,In_679,In_784);
xor U273 (N_273,In_374,In_239);
and U274 (N_274,In_887,In_816);
or U275 (N_275,In_692,In_914);
xor U276 (N_276,In_319,In_933);
nand U277 (N_277,In_73,In_135);
and U278 (N_278,In_225,In_544);
or U279 (N_279,In_768,In_910);
and U280 (N_280,In_711,In_787);
or U281 (N_281,In_874,In_648);
nor U282 (N_282,In_737,In_397);
or U283 (N_283,In_785,In_346);
nand U284 (N_284,In_166,In_98);
and U285 (N_285,In_388,In_876);
xor U286 (N_286,In_687,In_409);
nor U287 (N_287,In_255,In_339);
and U288 (N_288,In_39,In_34);
nor U289 (N_289,In_610,In_608);
nor U290 (N_290,In_146,In_895);
xor U291 (N_291,In_13,In_514);
or U292 (N_292,In_256,In_520);
or U293 (N_293,In_581,In_411);
nand U294 (N_294,In_290,In_734);
or U295 (N_295,In_796,In_169);
nor U296 (N_296,In_619,In_120);
or U297 (N_297,In_173,In_916);
nor U298 (N_298,In_223,In_800);
nand U299 (N_299,In_405,In_891);
or U300 (N_300,In_332,In_35);
nor U301 (N_301,In_477,In_277);
nand U302 (N_302,In_300,In_959);
or U303 (N_303,In_508,In_960);
nand U304 (N_304,In_878,In_962);
and U305 (N_305,In_377,In_354);
xnor U306 (N_306,In_20,In_102);
nor U307 (N_307,In_366,In_546);
nor U308 (N_308,In_853,In_632);
and U309 (N_309,In_824,In_337);
and U310 (N_310,In_313,In_137);
nor U311 (N_311,In_351,In_657);
nand U312 (N_312,In_618,In_334);
nor U313 (N_313,In_700,In_162);
nor U314 (N_314,In_176,In_901);
nor U315 (N_315,In_352,In_987);
or U316 (N_316,In_46,In_759);
xnor U317 (N_317,In_837,In_61);
and U318 (N_318,In_873,In_658);
nand U319 (N_319,In_535,In_865);
and U320 (N_320,In_480,In_27);
or U321 (N_321,In_349,In_809);
nand U322 (N_322,In_966,In_106);
nor U323 (N_323,In_863,In_450);
nand U324 (N_324,In_498,In_264);
nand U325 (N_325,In_325,In_501);
nor U326 (N_326,In_638,In_769);
nand U327 (N_327,In_820,In_774);
and U328 (N_328,In_915,In_604);
nand U329 (N_329,In_261,In_171);
nor U330 (N_330,In_211,In_938);
nand U331 (N_331,In_750,In_639);
nand U332 (N_332,In_587,In_848);
xor U333 (N_333,In_479,In_262);
nand U334 (N_334,In_15,In_896);
or U335 (N_335,In_193,In_400);
or U336 (N_336,In_695,In_431);
nand U337 (N_337,In_89,In_883);
nor U338 (N_338,In_111,In_423);
nor U339 (N_339,In_980,In_159);
nor U340 (N_340,In_67,In_275);
and U341 (N_341,In_335,In_949);
nand U342 (N_342,In_903,In_941);
nor U343 (N_343,In_715,In_395);
nand U344 (N_344,In_21,In_947);
nand U345 (N_345,In_285,In_556);
nand U346 (N_346,In_466,In_641);
nor U347 (N_347,In_778,In_247);
nor U348 (N_348,In_926,In_180);
or U349 (N_349,In_555,In_517);
or U350 (N_350,In_569,In_336);
and U351 (N_351,In_417,In_623);
and U352 (N_352,In_266,In_113);
and U353 (N_353,In_919,In_877);
and U354 (N_354,In_578,In_642);
nand U355 (N_355,In_668,In_297);
xnor U356 (N_356,In_855,In_675);
and U357 (N_357,In_489,In_407);
or U358 (N_358,In_834,In_871);
nand U359 (N_359,In_680,In_929);
xnor U360 (N_360,In_500,In_706);
and U361 (N_361,In_936,In_441);
nand U362 (N_362,In_644,In_10);
nor U363 (N_363,In_927,In_751);
and U364 (N_364,In_808,In_287);
and U365 (N_365,In_216,In_282);
and U366 (N_366,In_190,In_55);
xnor U367 (N_367,In_894,In_330);
and U368 (N_368,In_907,In_301);
xnor U369 (N_369,In_761,In_823);
nand U370 (N_370,In_156,In_596);
xnor U371 (N_371,In_130,In_686);
nand U372 (N_372,In_379,In_94);
nand U373 (N_373,In_383,In_468);
and U374 (N_374,In_250,In_890);
and U375 (N_375,In_562,In_235);
nor U376 (N_376,In_590,In_272);
nand U377 (N_377,In_322,In_957);
and U378 (N_378,In_565,In_138);
nand U379 (N_379,In_532,In_338);
xor U380 (N_380,In_343,In_802);
or U381 (N_381,In_127,In_492);
nor U382 (N_382,In_447,In_749);
or U383 (N_383,In_257,In_436);
nor U384 (N_384,In_197,In_852);
nor U385 (N_385,In_770,In_972);
nand U386 (N_386,In_653,In_350);
or U387 (N_387,In_503,In_645);
or U388 (N_388,In_308,In_622);
and U389 (N_389,In_5,In_582);
nand U390 (N_390,In_493,In_721);
or U391 (N_391,In_707,In_324);
nor U392 (N_392,In_452,In_189);
and U393 (N_393,In_321,In_310);
nand U394 (N_394,In_41,In_904);
nand U395 (N_395,In_801,In_100);
or U396 (N_396,In_646,In_132);
and U397 (N_397,In_681,In_86);
xor U398 (N_398,In_70,In_124);
or U399 (N_399,In_693,In_278);
nand U400 (N_400,In_372,In_595);
and U401 (N_401,In_557,In_65);
nand U402 (N_402,In_856,In_704);
and U403 (N_403,In_839,In_577);
and U404 (N_404,In_617,In_238);
nor U405 (N_405,In_783,In_815);
or U406 (N_406,In_483,In_205);
nor U407 (N_407,In_850,In_902);
or U408 (N_408,In_454,In_899);
or U409 (N_409,In_678,In_539);
or U410 (N_410,In_821,In_727);
nor U411 (N_411,In_488,In_465);
or U412 (N_412,In_512,In_574);
or U413 (N_413,In_368,In_259);
nor U414 (N_414,In_392,In_974);
or U415 (N_415,In_4,In_243);
and U416 (N_416,In_427,In_248);
and U417 (N_417,In_753,In_973);
nor U418 (N_418,In_118,In_832);
nand U419 (N_419,In_295,In_213);
and U420 (N_420,In_531,In_406);
nor U421 (N_421,In_333,In_104);
and U422 (N_422,In_603,In_806);
nor U423 (N_423,In_803,In_884);
or U424 (N_424,In_103,In_230);
and U425 (N_425,In_425,In_309);
nor U426 (N_426,In_17,In_490);
nor U427 (N_427,In_760,In_673);
nor U428 (N_428,In_58,In_810);
or U429 (N_429,In_931,In_670);
and U430 (N_430,In_85,In_541);
nor U431 (N_431,In_579,In_49);
xor U432 (N_432,In_963,In_1);
nand U433 (N_433,In_942,In_976);
and U434 (N_434,In_667,In_167);
nand U435 (N_435,In_918,In_373);
nand U436 (N_436,In_36,In_467);
or U437 (N_437,In_292,In_7);
and U438 (N_438,In_530,In_868);
and U439 (N_439,In_370,In_897);
and U440 (N_440,In_552,In_932);
nand U441 (N_441,In_634,In_123);
or U442 (N_442,In_908,In_128);
nand U443 (N_443,In_521,In_621);
or U444 (N_444,In_40,In_139);
or U445 (N_445,In_701,In_344);
nand U446 (N_446,In_88,In_226);
nand U447 (N_447,In_566,In_682);
and U448 (N_448,In_842,In_8);
or U449 (N_449,In_129,In_381);
nand U450 (N_450,In_186,In_482);
nor U451 (N_451,In_486,In_690);
nor U452 (N_452,In_765,In_561);
nor U453 (N_453,In_593,In_430);
or U454 (N_454,In_320,In_533);
or U455 (N_455,In_53,In_591);
and U456 (N_456,In_206,In_756);
and U457 (N_457,In_429,In_630);
nand U458 (N_458,In_849,In_812);
or U459 (N_459,In_616,In_306);
and U460 (N_460,In_666,In_328);
xnor U461 (N_461,In_920,In_161);
and U462 (N_462,In_724,In_298);
and U463 (N_463,In_793,In_996);
nor U464 (N_464,In_505,In_133);
or U465 (N_465,In_755,In_733);
or U466 (N_466,In_403,In_597);
nand U467 (N_467,In_142,In_110);
nand U468 (N_468,In_112,In_509);
and U469 (N_469,In_589,In_788);
nand U470 (N_470,In_524,In_586);
or U471 (N_471,In_979,In_859);
xor U472 (N_472,In_212,In_273);
nand U473 (N_473,In_458,In_551);
nand U474 (N_474,In_279,In_516);
nor U475 (N_475,In_924,In_72);
and U476 (N_476,In_398,In_702);
nor U477 (N_477,In_210,In_720);
or U478 (N_478,In_265,In_472);
or U479 (N_479,In_762,In_362);
nor U480 (N_480,In_312,In_703);
or U481 (N_481,In_845,In_140);
or U482 (N_482,In_745,In_345);
and U483 (N_483,In_263,In_893);
nand U484 (N_484,In_708,In_232);
nand U485 (N_485,In_386,In_804);
nand U486 (N_486,In_954,In_485);
or U487 (N_487,In_558,In_410);
nand U488 (N_488,In_888,In_418);
nand U489 (N_489,In_364,In_925);
or U490 (N_490,In_218,In_805);
and U491 (N_491,In_542,In_792);
nand U492 (N_492,In_694,In_202);
nand U493 (N_493,In_955,In_181);
xor U494 (N_494,In_688,In_838);
nor U495 (N_495,In_24,In_728);
nand U496 (N_496,In_709,In_660);
nor U497 (N_497,In_502,In_786);
nor U498 (N_498,In_291,In_76);
nand U499 (N_499,In_827,In_90);
or U500 (N_500,In_985,In_981);
and U501 (N_501,In_158,In_744);
or U502 (N_502,In_533,In_209);
nand U503 (N_503,In_611,In_94);
nor U504 (N_504,In_961,In_914);
and U505 (N_505,In_594,In_942);
and U506 (N_506,In_508,In_590);
nor U507 (N_507,In_199,In_988);
nor U508 (N_508,In_379,In_360);
or U509 (N_509,In_763,In_291);
nand U510 (N_510,In_889,In_965);
and U511 (N_511,In_823,In_715);
nor U512 (N_512,In_164,In_506);
nand U513 (N_513,In_928,In_341);
xor U514 (N_514,In_259,In_318);
nand U515 (N_515,In_195,In_752);
nor U516 (N_516,In_782,In_607);
or U517 (N_517,In_141,In_393);
nor U518 (N_518,In_238,In_515);
nor U519 (N_519,In_489,In_509);
nand U520 (N_520,In_344,In_590);
xnor U521 (N_521,In_364,In_416);
or U522 (N_522,In_610,In_810);
nand U523 (N_523,In_540,In_326);
or U524 (N_524,In_742,In_832);
nor U525 (N_525,In_243,In_646);
nor U526 (N_526,In_17,In_253);
and U527 (N_527,In_677,In_307);
or U528 (N_528,In_519,In_808);
xnor U529 (N_529,In_911,In_761);
or U530 (N_530,In_749,In_97);
and U531 (N_531,In_202,In_604);
nor U532 (N_532,In_743,In_140);
nand U533 (N_533,In_249,In_790);
or U534 (N_534,In_621,In_852);
nor U535 (N_535,In_518,In_688);
nand U536 (N_536,In_275,In_587);
and U537 (N_537,In_631,In_249);
or U538 (N_538,In_66,In_177);
nand U539 (N_539,In_76,In_643);
nor U540 (N_540,In_111,In_354);
and U541 (N_541,In_438,In_709);
nor U542 (N_542,In_109,In_653);
and U543 (N_543,In_991,In_443);
nor U544 (N_544,In_579,In_240);
nand U545 (N_545,In_89,In_206);
nand U546 (N_546,In_119,In_292);
nor U547 (N_547,In_733,In_134);
nand U548 (N_548,In_45,In_631);
nand U549 (N_549,In_755,In_467);
nor U550 (N_550,In_303,In_123);
or U551 (N_551,In_442,In_910);
and U552 (N_552,In_654,In_401);
or U553 (N_553,In_527,In_796);
nand U554 (N_554,In_972,In_239);
or U555 (N_555,In_223,In_286);
nor U556 (N_556,In_567,In_904);
or U557 (N_557,In_68,In_834);
and U558 (N_558,In_711,In_76);
nand U559 (N_559,In_70,In_97);
nor U560 (N_560,In_544,In_564);
nor U561 (N_561,In_223,In_590);
and U562 (N_562,In_968,In_729);
or U563 (N_563,In_250,In_92);
or U564 (N_564,In_506,In_889);
nor U565 (N_565,In_311,In_197);
nor U566 (N_566,In_382,In_653);
nand U567 (N_567,In_820,In_471);
nor U568 (N_568,In_445,In_849);
or U569 (N_569,In_248,In_429);
nand U570 (N_570,In_805,In_56);
nand U571 (N_571,In_286,In_569);
nand U572 (N_572,In_715,In_475);
or U573 (N_573,In_627,In_209);
nor U574 (N_574,In_354,In_385);
and U575 (N_575,In_918,In_767);
and U576 (N_576,In_395,In_308);
or U577 (N_577,In_148,In_866);
or U578 (N_578,In_961,In_815);
nand U579 (N_579,In_909,In_912);
and U580 (N_580,In_90,In_897);
or U581 (N_581,In_392,In_883);
nand U582 (N_582,In_717,In_756);
or U583 (N_583,In_867,In_883);
xor U584 (N_584,In_778,In_96);
nor U585 (N_585,In_350,In_113);
nor U586 (N_586,In_555,In_879);
and U587 (N_587,In_593,In_785);
nor U588 (N_588,In_223,In_787);
nor U589 (N_589,In_17,In_85);
nor U590 (N_590,In_844,In_137);
or U591 (N_591,In_148,In_694);
nand U592 (N_592,In_966,In_162);
xnor U593 (N_593,In_853,In_588);
nor U594 (N_594,In_241,In_343);
xnor U595 (N_595,In_43,In_733);
nor U596 (N_596,In_443,In_340);
nand U597 (N_597,In_903,In_7);
and U598 (N_598,In_152,In_523);
nor U599 (N_599,In_624,In_946);
xnor U600 (N_600,In_703,In_994);
nand U601 (N_601,In_450,In_504);
nand U602 (N_602,In_398,In_37);
and U603 (N_603,In_69,In_497);
nor U604 (N_604,In_999,In_82);
nor U605 (N_605,In_92,In_468);
or U606 (N_606,In_976,In_195);
or U607 (N_607,In_530,In_543);
nand U608 (N_608,In_896,In_707);
nor U609 (N_609,In_392,In_94);
and U610 (N_610,In_309,In_175);
nand U611 (N_611,In_965,In_278);
nand U612 (N_612,In_920,In_866);
xnor U613 (N_613,In_838,In_522);
xor U614 (N_614,In_219,In_81);
nand U615 (N_615,In_325,In_209);
or U616 (N_616,In_187,In_52);
and U617 (N_617,In_47,In_394);
nor U618 (N_618,In_115,In_45);
nand U619 (N_619,In_296,In_818);
and U620 (N_620,In_160,In_321);
and U621 (N_621,In_977,In_779);
nor U622 (N_622,In_499,In_881);
nor U623 (N_623,In_528,In_857);
and U624 (N_624,In_624,In_144);
or U625 (N_625,In_670,In_676);
and U626 (N_626,In_540,In_636);
nand U627 (N_627,In_906,In_44);
nand U628 (N_628,In_136,In_665);
nand U629 (N_629,In_16,In_314);
nand U630 (N_630,In_58,In_740);
nor U631 (N_631,In_803,In_174);
or U632 (N_632,In_234,In_969);
nor U633 (N_633,In_334,In_143);
nor U634 (N_634,In_352,In_529);
or U635 (N_635,In_28,In_184);
nand U636 (N_636,In_494,In_933);
xnor U637 (N_637,In_912,In_178);
nand U638 (N_638,In_999,In_606);
or U639 (N_639,In_668,In_262);
nor U640 (N_640,In_32,In_169);
nand U641 (N_641,In_563,In_841);
and U642 (N_642,In_793,In_92);
nand U643 (N_643,In_306,In_964);
nand U644 (N_644,In_102,In_983);
and U645 (N_645,In_930,In_411);
and U646 (N_646,In_206,In_773);
or U647 (N_647,In_728,In_527);
or U648 (N_648,In_52,In_519);
nor U649 (N_649,In_481,In_302);
nand U650 (N_650,In_722,In_33);
nand U651 (N_651,In_967,In_781);
nor U652 (N_652,In_916,In_532);
or U653 (N_653,In_560,In_659);
nand U654 (N_654,In_625,In_67);
nand U655 (N_655,In_960,In_911);
nor U656 (N_656,In_29,In_948);
and U657 (N_657,In_38,In_199);
xnor U658 (N_658,In_520,In_635);
and U659 (N_659,In_36,In_568);
xnor U660 (N_660,In_831,In_561);
nand U661 (N_661,In_874,In_748);
and U662 (N_662,In_726,In_956);
or U663 (N_663,In_933,In_555);
nand U664 (N_664,In_114,In_886);
nor U665 (N_665,In_950,In_594);
and U666 (N_666,In_870,In_171);
and U667 (N_667,In_480,In_233);
or U668 (N_668,In_325,In_181);
or U669 (N_669,In_355,In_702);
nor U670 (N_670,In_574,In_721);
nand U671 (N_671,In_176,In_30);
or U672 (N_672,In_209,In_777);
xnor U673 (N_673,In_923,In_537);
and U674 (N_674,In_380,In_713);
nor U675 (N_675,In_703,In_78);
nand U676 (N_676,In_312,In_918);
nand U677 (N_677,In_408,In_413);
or U678 (N_678,In_248,In_955);
or U679 (N_679,In_19,In_830);
and U680 (N_680,In_117,In_703);
nand U681 (N_681,In_784,In_552);
and U682 (N_682,In_892,In_460);
nor U683 (N_683,In_328,In_972);
nor U684 (N_684,In_600,In_917);
and U685 (N_685,In_866,In_179);
xnor U686 (N_686,In_608,In_365);
or U687 (N_687,In_426,In_168);
and U688 (N_688,In_275,In_776);
or U689 (N_689,In_98,In_594);
nor U690 (N_690,In_326,In_906);
or U691 (N_691,In_233,In_529);
xor U692 (N_692,In_151,In_711);
nand U693 (N_693,In_181,In_4);
nor U694 (N_694,In_506,In_466);
nor U695 (N_695,In_283,In_161);
and U696 (N_696,In_990,In_459);
and U697 (N_697,In_87,In_601);
xnor U698 (N_698,In_873,In_359);
nand U699 (N_699,In_712,In_914);
and U700 (N_700,In_207,In_19);
nand U701 (N_701,In_853,In_487);
xor U702 (N_702,In_374,In_926);
nor U703 (N_703,In_449,In_879);
nor U704 (N_704,In_831,In_181);
xor U705 (N_705,In_783,In_759);
and U706 (N_706,In_786,In_377);
nand U707 (N_707,In_187,In_656);
or U708 (N_708,In_392,In_704);
xor U709 (N_709,In_198,In_910);
nand U710 (N_710,In_488,In_544);
nor U711 (N_711,In_660,In_15);
nand U712 (N_712,In_280,In_804);
nor U713 (N_713,In_413,In_338);
xor U714 (N_714,In_1,In_483);
and U715 (N_715,In_42,In_594);
nor U716 (N_716,In_178,In_948);
nor U717 (N_717,In_705,In_147);
nand U718 (N_718,In_340,In_163);
nand U719 (N_719,In_989,In_27);
or U720 (N_720,In_271,In_801);
or U721 (N_721,In_735,In_827);
nor U722 (N_722,In_80,In_911);
or U723 (N_723,In_171,In_119);
nor U724 (N_724,In_572,In_337);
and U725 (N_725,In_965,In_654);
nand U726 (N_726,In_731,In_792);
nand U727 (N_727,In_924,In_487);
nand U728 (N_728,In_771,In_584);
nand U729 (N_729,In_182,In_441);
and U730 (N_730,In_289,In_582);
nor U731 (N_731,In_841,In_500);
and U732 (N_732,In_164,In_71);
or U733 (N_733,In_276,In_841);
and U734 (N_734,In_86,In_96);
nor U735 (N_735,In_497,In_495);
and U736 (N_736,In_406,In_501);
and U737 (N_737,In_26,In_90);
nand U738 (N_738,In_698,In_308);
xor U739 (N_739,In_188,In_525);
or U740 (N_740,In_617,In_33);
or U741 (N_741,In_35,In_258);
nand U742 (N_742,In_119,In_597);
and U743 (N_743,In_944,In_138);
and U744 (N_744,In_900,In_671);
or U745 (N_745,In_315,In_191);
or U746 (N_746,In_356,In_289);
nor U747 (N_747,In_214,In_0);
or U748 (N_748,In_249,In_217);
nor U749 (N_749,In_628,In_266);
or U750 (N_750,In_583,In_936);
nand U751 (N_751,In_61,In_461);
and U752 (N_752,In_583,In_238);
nand U753 (N_753,In_726,In_677);
and U754 (N_754,In_300,In_824);
nor U755 (N_755,In_167,In_848);
and U756 (N_756,In_588,In_666);
xnor U757 (N_757,In_286,In_881);
and U758 (N_758,In_924,In_27);
xnor U759 (N_759,In_764,In_582);
or U760 (N_760,In_408,In_777);
or U761 (N_761,In_287,In_252);
and U762 (N_762,In_195,In_627);
xor U763 (N_763,In_936,In_227);
xor U764 (N_764,In_142,In_800);
nand U765 (N_765,In_992,In_443);
nor U766 (N_766,In_815,In_740);
or U767 (N_767,In_833,In_324);
nor U768 (N_768,In_893,In_963);
nand U769 (N_769,In_520,In_174);
xnor U770 (N_770,In_365,In_211);
nor U771 (N_771,In_518,In_854);
or U772 (N_772,In_36,In_721);
nor U773 (N_773,In_108,In_536);
nand U774 (N_774,In_425,In_429);
or U775 (N_775,In_505,In_242);
nand U776 (N_776,In_939,In_26);
xnor U777 (N_777,In_511,In_750);
and U778 (N_778,In_41,In_185);
nor U779 (N_779,In_49,In_149);
or U780 (N_780,In_324,In_542);
nor U781 (N_781,In_168,In_795);
or U782 (N_782,In_388,In_71);
nor U783 (N_783,In_696,In_466);
nor U784 (N_784,In_339,In_128);
and U785 (N_785,In_684,In_901);
and U786 (N_786,In_22,In_396);
and U787 (N_787,In_355,In_724);
and U788 (N_788,In_755,In_6);
nor U789 (N_789,In_574,In_464);
nor U790 (N_790,In_607,In_90);
nor U791 (N_791,In_539,In_544);
and U792 (N_792,In_737,In_245);
or U793 (N_793,In_493,In_570);
xnor U794 (N_794,In_847,In_189);
and U795 (N_795,In_968,In_441);
nor U796 (N_796,In_179,In_367);
nor U797 (N_797,In_269,In_2);
or U798 (N_798,In_546,In_494);
or U799 (N_799,In_304,In_95);
nand U800 (N_800,In_321,In_786);
nand U801 (N_801,In_233,In_387);
and U802 (N_802,In_420,In_729);
nand U803 (N_803,In_780,In_630);
nand U804 (N_804,In_568,In_518);
or U805 (N_805,In_866,In_916);
or U806 (N_806,In_241,In_540);
nor U807 (N_807,In_452,In_637);
or U808 (N_808,In_94,In_626);
nand U809 (N_809,In_987,In_821);
nor U810 (N_810,In_379,In_529);
or U811 (N_811,In_479,In_137);
nand U812 (N_812,In_130,In_7);
nor U813 (N_813,In_71,In_170);
nand U814 (N_814,In_71,In_271);
nor U815 (N_815,In_961,In_96);
nand U816 (N_816,In_356,In_772);
and U817 (N_817,In_275,In_538);
or U818 (N_818,In_785,In_267);
nand U819 (N_819,In_274,In_184);
nor U820 (N_820,In_410,In_168);
and U821 (N_821,In_8,In_96);
nor U822 (N_822,In_556,In_806);
nand U823 (N_823,In_288,In_183);
nand U824 (N_824,In_464,In_786);
nor U825 (N_825,In_461,In_725);
nor U826 (N_826,In_544,In_908);
and U827 (N_827,In_767,In_430);
xnor U828 (N_828,In_73,In_271);
nand U829 (N_829,In_767,In_133);
xnor U830 (N_830,In_725,In_421);
nor U831 (N_831,In_165,In_985);
nor U832 (N_832,In_473,In_11);
xor U833 (N_833,In_305,In_714);
and U834 (N_834,In_736,In_299);
and U835 (N_835,In_333,In_324);
nand U836 (N_836,In_306,In_222);
nand U837 (N_837,In_809,In_940);
and U838 (N_838,In_152,In_576);
or U839 (N_839,In_414,In_259);
nand U840 (N_840,In_658,In_750);
and U841 (N_841,In_309,In_756);
or U842 (N_842,In_630,In_180);
or U843 (N_843,In_30,In_137);
or U844 (N_844,In_848,In_295);
nor U845 (N_845,In_110,In_808);
nand U846 (N_846,In_666,In_950);
nor U847 (N_847,In_238,In_114);
nand U848 (N_848,In_362,In_176);
and U849 (N_849,In_336,In_958);
nor U850 (N_850,In_690,In_501);
or U851 (N_851,In_945,In_841);
or U852 (N_852,In_390,In_942);
and U853 (N_853,In_952,In_866);
nor U854 (N_854,In_994,In_768);
nand U855 (N_855,In_267,In_610);
nand U856 (N_856,In_690,In_612);
nor U857 (N_857,In_909,In_155);
xor U858 (N_858,In_825,In_831);
and U859 (N_859,In_337,In_529);
and U860 (N_860,In_312,In_182);
nor U861 (N_861,In_102,In_490);
xnor U862 (N_862,In_183,In_393);
nand U863 (N_863,In_59,In_893);
nand U864 (N_864,In_502,In_96);
or U865 (N_865,In_441,In_494);
nor U866 (N_866,In_912,In_514);
and U867 (N_867,In_84,In_906);
and U868 (N_868,In_311,In_573);
nor U869 (N_869,In_937,In_526);
nand U870 (N_870,In_956,In_635);
and U871 (N_871,In_59,In_806);
nand U872 (N_872,In_87,In_694);
nor U873 (N_873,In_534,In_400);
or U874 (N_874,In_781,In_146);
or U875 (N_875,In_501,In_881);
or U876 (N_876,In_778,In_576);
or U877 (N_877,In_386,In_237);
nor U878 (N_878,In_813,In_641);
nand U879 (N_879,In_366,In_559);
or U880 (N_880,In_182,In_285);
and U881 (N_881,In_538,In_457);
nand U882 (N_882,In_673,In_44);
xor U883 (N_883,In_762,In_728);
nor U884 (N_884,In_59,In_762);
nor U885 (N_885,In_7,In_316);
and U886 (N_886,In_157,In_79);
xor U887 (N_887,In_879,In_848);
and U888 (N_888,In_697,In_84);
nand U889 (N_889,In_967,In_426);
and U890 (N_890,In_553,In_980);
nand U891 (N_891,In_151,In_651);
nor U892 (N_892,In_722,In_9);
nor U893 (N_893,In_506,In_826);
or U894 (N_894,In_812,In_434);
or U895 (N_895,In_361,In_287);
nand U896 (N_896,In_732,In_945);
or U897 (N_897,In_599,In_360);
nor U898 (N_898,In_120,In_718);
and U899 (N_899,In_93,In_639);
and U900 (N_900,In_238,In_251);
and U901 (N_901,In_149,In_8);
nor U902 (N_902,In_560,In_73);
nor U903 (N_903,In_549,In_714);
nor U904 (N_904,In_780,In_808);
nand U905 (N_905,In_221,In_810);
and U906 (N_906,In_470,In_339);
or U907 (N_907,In_620,In_58);
nor U908 (N_908,In_701,In_242);
nor U909 (N_909,In_139,In_697);
nor U910 (N_910,In_895,In_52);
nor U911 (N_911,In_943,In_998);
xor U912 (N_912,In_614,In_839);
and U913 (N_913,In_473,In_577);
or U914 (N_914,In_856,In_440);
nand U915 (N_915,In_585,In_411);
nand U916 (N_916,In_69,In_805);
or U917 (N_917,In_248,In_23);
nand U918 (N_918,In_991,In_193);
and U919 (N_919,In_610,In_72);
nand U920 (N_920,In_638,In_332);
nand U921 (N_921,In_730,In_621);
nand U922 (N_922,In_990,In_852);
or U923 (N_923,In_768,In_728);
and U924 (N_924,In_996,In_844);
nand U925 (N_925,In_250,In_920);
nor U926 (N_926,In_216,In_757);
and U927 (N_927,In_811,In_537);
nor U928 (N_928,In_697,In_503);
and U929 (N_929,In_520,In_339);
nor U930 (N_930,In_27,In_579);
xnor U931 (N_931,In_815,In_347);
nor U932 (N_932,In_831,In_551);
nor U933 (N_933,In_249,In_336);
nand U934 (N_934,In_295,In_311);
nand U935 (N_935,In_967,In_329);
nand U936 (N_936,In_378,In_356);
nor U937 (N_937,In_869,In_935);
nor U938 (N_938,In_226,In_423);
and U939 (N_939,In_231,In_957);
xnor U940 (N_940,In_286,In_116);
or U941 (N_941,In_528,In_401);
and U942 (N_942,In_629,In_389);
nor U943 (N_943,In_905,In_385);
or U944 (N_944,In_297,In_92);
or U945 (N_945,In_424,In_423);
or U946 (N_946,In_329,In_640);
or U947 (N_947,In_116,In_571);
or U948 (N_948,In_125,In_210);
or U949 (N_949,In_757,In_409);
nor U950 (N_950,In_977,In_591);
xor U951 (N_951,In_519,In_816);
nand U952 (N_952,In_494,In_412);
or U953 (N_953,In_459,In_618);
and U954 (N_954,In_471,In_603);
nor U955 (N_955,In_540,In_188);
xnor U956 (N_956,In_240,In_386);
nand U957 (N_957,In_123,In_850);
nor U958 (N_958,In_114,In_82);
xnor U959 (N_959,In_352,In_516);
nor U960 (N_960,In_422,In_812);
or U961 (N_961,In_328,In_945);
nand U962 (N_962,In_123,In_388);
nor U963 (N_963,In_494,In_153);
nand U964 (N_964,In_334,In_384);
and U965 (N_965,In_17,In_197);
and U966 (N_966,In_423,In_859);
nand U967 (N_967,In_257,In_690);
and U968 (N_968,In_376,In_916);
nor U969 (N_969,In_986,In_961);
and U970 (N_970,In_719,In_309);
nor U971 (N_971,In_144,In_684);
xor U972 (N_972,In_680,In_47);
nor U973 (N_973,In_821,In_175);
xnor U974 (N_974,In_198,In_494);
or U975 (N_975,In_812,In_403);
or U976 (N_976,In_212,In_895);
and U977 (N_977,In_753,In_11);
or U978 (N_978,In_504,In_918);
nor U979 (N_979,In_879,In_680);
and U980 (N_980,In_35,In_828);
and U981 (N_981,In_116,In_371);
or U982 (N_982,In_218,In_704);
xnor U983 (N_983,In_696,In_935);
and U984 (N_984,In_120,In_497);
nor U985 (N_985,In_842,In_136);
nand U986 (N_986,In_512,In_26);
and U987 (N_987,In_342,In_986);
and U988 (N_988,In_60,In_279);
and U989 (N_989,In_974,In_870);
nor U990 (N_990,In_905,In_789);
nor U991 (N_991,In_398,In_443);
nor U992 (N_992,In_795,In_574);
and U993 (N_993,In_756,In_956);
nand U994 (N_994,In_966,In_900);
nor U995 (N_995,In_128,In_510);
and U996 (N_996,In_233,In_902);
and U997 (N_997,In_117,In_490);
or U998 (N_998,In_62,In_471);
or U999 (N_999,In_730,In_450);
nand U1000 (N_1000,In_98,In_187);
or U1001 (N_1001,In_92,In_57);
or U1002 (N_1002,In_585,In_15);
or U1003 (N_1003,In_963,In_457);
nand U1004 (N_1004,In_303,In_83);
and U1005 (N_1005,In_877,In_500);
nor U1006 (N_1006,In_4,In_542);
or U1007 (N_1007,In_57,In_650);
and U1008 (N_1008,In_576,In_889);
and U1009 (N_1009,In_596,In_644);
nand U1010 (N_1010,In_15,In_659);
nand U1011 (N_1011,In_654,In_251);
or U1012 (N_1012,In_818,In_721);
or U1013 (N_1013,In_452,In_339);
nand U1014 (N_1014,In_950,In_849);
and U1015 (N_1015,In_54,In_392);
xnor U1016 (N_1016,In_444,In_626);
or U1017 (N_1017,In_756,In_964);
nand U1018 (N_1018,In_877,In_580);
or U1019 (N_1019,In_433,In_458);
nor U1020 (N_1020,In_866,In_788);
and U1021 (N_1021,In_458,In_239);
nor U1022 (N_1022,In_243,In_215);
and U1023 (N_1023,In_166,In_390);
or U1024 (N_1024,In_222,In_811);
nor U1025 (N_1025,In_410,In_871);
nand U1026 (N_1026,In_613,In_144);
nor U1027 (N_1027,In_876,In_702);
or U1028 (N_1028,In_914,In_542);
nand U1029 (N_1029,In_713,In_874);
nor U1030 (N_1030,In_199,In_350);
and U1031 (N_1031,In_249,In_899);
nand U1032 (N_1032,In_99,In_514);
or U1033 (N_1033,In_502,In_157);
nor U1034 (N_1034,In_328,In_620);
nor U1035 (N_1035,In_494,In_525);
or U1036 (N_1036,In_606,In_471);
nand U1037 (N_1037,In_366,In_631);
nand U1038 (N_1038,In_340,In_31);
nor U1039 (N_1039,In_911,In_465);
xor U1040 (N_1040,In_653,In_694);
xnor U1041 (N_1041,In_310,In_283);
and U1042 (N_1042,In_940,In_843);
and U1043 (N_1043,In_587,In_855);
nand U1044 (N_1044,In_433,In_723);
nand U1045 (N_1045,In_262,In_104);
or U1046 (N_1046,In_308,In_654);
or U1047 (N_1047,In_959,In_673);
or U1048 (N_1048,In_386,In_24);
nor U1049 (N_1049,In_193,In_522);
nand U1050 (N_1050,In_636,In_218);
nand U1051 (N_1051,In_413,In_89);
or U1052 (N_1052,In_893,In_702);
nor U1053 (N_1053,In_961,In_413);
nor U1054 (N_1054,In_818,In_189);
nor U1055 (N_1055,In_733,In_178);
nor U1056 (N_1056,In_720,In_305);
nand U1057 (N_1057,In_663,In_442);
nor U1058 (N_1058,In_457,In_546);
nor U1059 (N_1059,In_433,In_21);
or U1060 (N_1060,In_177,In_348);
and U1061 (N_1061,In_616,In_788);
and U1062 (N_1062,In_214,In_867);
nor U1063 (N_1063,In_269,In_561);
nand U1064 (N_1064,In_228,In_461);
or U1065 (N_1065,In_649,In_550);
nand U1066 (N_1066,In_895,In_43);
nor U1067 (N_1067,In_638,In_496);
nand U1068 (N_1068,In_866,In_618);
and U1069 (N_1069,In_304,In_320);
and U1070 (N_1070,In_117,In_364);
nor U1071 (N_1071,In_178,In_949);
and U1072 (N_1072,In_728,In_784);
nand U1073 (N_1073,In_963,In_173);
nand U1074 (N_1074,In_338,In_600);
and U1075 (N_1075,In_842,In_342);
or U1076 (N_1076,In_148,In_338);
and U1077 (N_1077,In_528,In_31);
nor U1078 (N_1078,In_373,In_438);
nor U1079 (N_1079,In_781,In_306);
nand U1080 (N_1080,In_148,In_929);
and U1081 (N_1081,In_659,In_744);
xor U1082 (N_1082,In_743,In_543);
or U1083 (N_1083,In_887,In_368);
nand U1084 (N_1084,In_73,In_395);
nor U1085 (N_1085,In_125,In_121);
and U1086 (N_1086,In_259,In_936);
and U1087 (N_1087,In_202,In_594);
or U1088 (N_1088,In_109,In_285);
nand U1089 (N_1089,In_242,In_945);
nand U1090 (N_1090,In_229,In_247);
nand U1091 (N_1091,In_563,In_923);
and U1092 (N_1092,In_306,In_280);
and U1093 (N_1093,In_445,In_465);
nor U1094 (N_1094,In_702,In_109);
xor U1095 (N_1095,In_594,In_826);
or U1096 (N_1096,In_206,In_704);
and U1097 (N_1097,In_161,In_857);
xnor U1098 (N_1098,In_599,In_208);
or U1099 (N_1099,In_963,In_879);
or U1100 (N_1100,In_146,In_105);
nor U1101 (N_1101,In_915,In_930);
or U1102 (N_1102,In_644,In_931);
or U1103 (N_1103,In_686,In_962);
or U1104 (N_1104,In_847,In_783);
and U1105 (N_1105,In_39,In_481);
or U1106 (N_1106,In_427,In_266);
and U1107 (N_1107,In_746,In_875);
and U1108 (N_1108,In_337,In_848);
and U1109 (N_1109,In_593,In_140);
or U1110 (N_1110,In_847,In_33);
or U1111 (N_1111,In_682,In_42);
nand U1112 (N_1112,In_871,In_234);
and U1113 (N_1113,In_259,In_731);
xnor U1114 (N_1114,In_731,In_176);
xnor U1115 (N_1115,In_324,In_810);
xor U1116 (N_1116,In_250,In_80);
or U1117 (N_1117,In_5,In_611);
xnor U1118 (N_1118,In_3,In_80);
nor U1119 (N_1119,In_965,In_400);
nand U1120 (N_1120,In_242,In_194);
or U1121 (N_1121,In_352,In_565);
or U1122 (N_1122,In_331,In_247);
nor U1123 (N_1123,In_275,In_884);
or U1124 (N_1124,In_660,In_501);
and U1125 (N_1125,In_886,In_974);
or U1126 (N_1126,In_901,In_786);
nor U1127 (N_1127,In_766,In_496);
nor U1128 (N_1128,In_38,In_486);
or U1129 (N_1129,In_545,In_76);
nand U1130 (N_1130,In_483,In_919);
nor U1131 (N_1131,In_130,In_432);
nor U1132 (N_1132,In_59,In_973);
nand U1133 (N_1133,In_916,In_231);
and U1134 (N_1134,In_929,In_492);
or U1135 (N_1135,In_29,In_976);
and U1136 (N_1136,In_115,In_539);
and U1137 (N_1137,In_610,In_153);
nand U1138 (N_1138,In_168,In_236);
and U1139 (N_1139,In_291,In_188);
nor U1140 (N_1140,In_911,In_539);
and U1141 (N_1141,In_806,In_493);
nor U1142 (N_1142,In_135,In_229);
or U1143 (N_1143,In_265,In_701);
and U1144 (N_1144,In_747,In_278);
nand U1145 (N_1145,In_644,In_593);
nand U1146 (N_1146,In_26,In_568);
nor U1147 (N_1147,In_757,In_545);
and U1148 (N_1148,In_565,In_597);
nand U1149 (N_1149,In_246,In_4);
nor U1150 (N_1150,In_746,In_841);
or U1151 (N_1151,In_307,In_760);
nand U1152 (N_1152,In_517,In_278);
nand U1153 (N_1153,In_340,In_223);
or U1154 (N_1154,In_627,In_689);
xor U1155 (N_1155,In_394,In_610);
and U1156 (N_1156,In_808,In_370);
and U1157 (N_1157,In_981,In_597);
nand U1158 (N_1158,In_905,In_717);
nor U1159 (N_1159,In_940,In_597);
nand U1160 (N_1160,In_433,In_783);
nand U1161 (N_1161,In_792,In_831);
or U1162 (N_1162,In_3,In_649);
xnor U1163 (N_1163,In_287,In_347);
and U1164 (N_1164,In_382,In_237);
and U1165 (N_1165,In_649,In_173);
and U1166 (N_1166,In_211,In_410);
nor U1167 (N_1167,In_243,In_941);
or U1168 (N_1168,In_153,In_177);
or U1169 (N_1169,In_963,In_491);
xor U1170 (N_1170,In_283,In_601);
or U1171 (N_1171,In_446,In_521);
and U1172 (N_1172,In_508,In_874);
nand U1173 (N_1173,In_466,In_918);
nand U1174 (N_1174,In_48,In_822);
xnor U1175 (N_1175,In_592,In_247);
nand U1176 (N_1176,In_873,In_549);
nand U1177 (N_1177,In_35,In_132);
nor U1178 (N_1178,In_274,In_866);
and U1179 (N_1179,In_160,In_884);
nor U1180 (N_1180,In_17,In_105);
nand U1181 (N_1181,In_513,In_32);
xnor U1182 (N_1182,In_374,In_59);
nand U1183 (N_1183,In_109,In_708);
and U1184 (N_1184,In_919,In_69);
xnor U1185 (N_1185,In_885,In_706);
nor U1186 (N_1186,In_220,In_253);
or U1187 (N_1187,In_689,In_39);
or U1188 (N_1188,In_419,In_684);
or U1189 (N_1189,In_762,In_187);
nand U1190 (N_1190,In_516,In_119);
nor U1191 (N_1191,In_93,In_980);
nand U1192 (N_1192,In_879,In_990);
xor U1193 (N_1193,In_589,In_74);
or U1194 (N_1194,In_213,In_928);
nand U1195 (N_1195,In_326,In_44);
nand U1196 (N_1196,In_669,In_681);
nor U1197 (N_1197,In_191,In_489);
nand U1198 (N_1198,In_770,In_896);
nor U1199 (N_1199,In_692,In_904);
and U1200 (N_1200,In_77,In_792);
or U1201 (N_1201,In_702,In_196);
nor U1202 (N_1202,In_176,In_225);
and U1203 (N_1203,In_943,In_188);
or U1204 (N_1204,In_625,In_788);
and U1205 (N_1205,In_347,In_820);
nand U1206 (N_1206,In_414,In_538);
and U1207 (N_1207,In_981,In_382);
or U1208 (N_1208,In_878,In_141);
or U1209 (N_1209,In_444,In_436);
xor U1210 (N_1210,In_440,In_952);
nor U1211 (N_1211,In_213,In_116);
nor U1212 (N_1212,In_966,In_787);
and U1213 (N_1213,In_49,In_153);
and U1214 (N_1214,In_958,In_112);
and U1215 (N_1215,In_439,In_666);
nor U1216 (N_1216,In_881,In_588);
and U1217 (N_1217,In_510,In_623);
or U1218 (N_1218,In_988,In_44);
nor U1219 (N_1219,In_826,In_161);
nor U1220 (N_1220,In_328,In_494);
nor U1221 (N_1221,In_672,In_93);
and U1222 (N_1222,In_262,In_85);
nor U1223 (N_1223,In_139,In_68);
nand U1224 (N_1224,In_645,In_527);
nand U1225 (N_1225,In_20,In_901);
and U1226 (N_1226,In_794,In_898);
nand U1227 (N_1227,In_289,In_448);
xnor U1228 (N_1228,In_234,In_305);
and U1229 (N_1229,In_122,In_521);
and U1230 (N_1230,In_892,In_531);
or U1231 (N_1231,In_307,In_992);
or U1232 (N_1232,In_509,In_118);
nor U1233 (N_1233,In_461,In_37);
and U1234 (N_1234,In_321,In_897);
or U1235 (N_1235,In_22,In_298);
xnor U1236 (N_1236,In_484,In_662);
and U1237 (N_1237,In_491,In_595);
or U1238 (N_1238,In_461,In_58);
and U1239 (N_1239,In_627,In_169);
and U1240 (N_1240,In_894,In_280);
nor U1241 (N_1241,In_128,In_62);
or U1242 (N_1242,In_209,In_817);
nand U1243 (N_1243,In_838,In_334);
xor U1244 (N_1244,In_180,In_143);
xnor U1245 (N_1245,In_716,In_761);
nand U1246 (N_1246,In_638,In_714);
nor U1247 (N_1247,In_803,In_30);
nor U1248 (N_1248,In_152,In_936);
and U1249 (N_1249,In_398,In_828);
and U1250 (N_1250,In_141,In_833);
nor U1251 (N_1251,In_35,In_782);
nor U1252 (N_1252,In_205,In_170);
xor U1253 (N_1253,In_806,In_731);
or U1254 (N_1254,In_229,In_619);
nand U1255 (N_1255,In_300,In_623);
nor U1256 (N_1256,In_505,In_636);
nor U1257 (N_1257,In_798,In_382);
and U1258 (N_1258,In_85,In_728);
nor U1259 (N_1259,In_305,In_41);
nor U1260 (N_1260,In_908,In_347);
or U1261 (N_1261,In_767,In_932);
nand U1262 (N_1262,In_63,In_273);
nor U1263 (N_1263,In_400,In_352);
xnor U1264 (N_1264,In_386,In_783);
nor U1265 (N_1265,In_143,In_475);
and U1266 (N_1266,In_577,In_308);
and U1267 (N_1267,In_647,In_346);
or U1268 (N_1268,In_317,In_540);
and U1269 (N_1269,In_800,In_217);
xor U1270 (N_1270,In_868,In_215);
and U1271 (N_1271,In_916,In_775);
and U1272 (N_1272,In_631,In_890);
nor U1273 (N_1273,In_454,In_978);
nand U1274 (N_1274,In_288,In_520);
nand U1275 (N_1275,In_680,In_586);
nor U1276 (N_1276,In_502,In_305);
nand U1277 (N_1277,In_920,In_56);
and U1278 (N_1278,In_502,In_890);
nor U1279 (N_1279,In_398,In_181);
xnor U1280 (N_1280,In_226,In_112);
nor U1281 (N_1281,In_949,In_944);
nand U1282 (N_1282,In_663,In_686);
or U1283 (N_1283,In_583,In_456);
and U1284 (N_1284,In_589,In_165);
nor U1285 (N_1285,In_692,In_42);
nand U1286 (N_1286,In_373,In_148);
xnor U1287 (N_1287,In_788,In_320);
and U1288 (N_1288,In_949,In_488);
or U1289 (N_1289,In_764,In_643);
xnor U1290 (N_1290,In_868,In_359);
nand U1291 (N_1291,In_305,In_358);
and U1292 (N_1292,In_647,In_183);
and U1293 (N_1293,In_534,In_719);
nor U1294 (N_1294,In_468,In_754);
nand U1295 (N_1295,In_707,In_753);
xnor U1296 (N_1296,In_125,In_434);
nand U1297 (N_1297,In_331,In_189);
or U1298 (N_1298,In_709,In_596);
nand U1299 (N_1299,In_786,In_469);
nand U1300 (N_1300,In_6,In_248);
or U1301 (N_1301,In_847,In_180);
nor U1302 (N_1302,In_629,In_224);
or U1303 (N_1303,In_975,In_822);
or U1304 (N_1304,In_431,In_755);
nand U1305 (N_1305,In_832,In_878);
nand U1306 (N_1306,In_35,In_547);
or U1307 (N_1307,In_754,In_466);
nor U1308 (N_1308,In_958,In_762);
or U1309 (N_1309,In_531,In_899);
nand U1310 (N_1310,In_288,In_287);
nand U1311 (N_1311,In_307,In_71);
and U1312 (N_1312,In_68,In_349);
or U1313 (N_1313,In_363,In_339);
xor U1314 (N_1314,In_979,In_662);
or U1315 (N_1315,In_694,In_140);
or U1316 (N_1316,In_182,In_491);
or U1317 (N_1317,In_363,In_971);
or U1318 (N_1318,In_745,In_993);
or U1319 (N_1319,In_269,In_863);
nand U1320 (N_1320,In_985,In_653);
or U1321 (N_1321,In_120,In_292);
nand U1322 (N_1322,In_18,In_282);
xnor U1323 (N_1323,In_442,In_262);
nand U1324 (N_1324,In_875,In_775);
and U1325 (N_1325,In_155,In_347);
nor U1326 (N_1326,In_717,In_325);
nand U1327 (N_1327,In_102,In_340);
and U1328 (N_1328,In_841,In_357);
nor U1329 (N_1329,In_291,In_707);
and U1330 (N_1330,In_952,In_407);
xnor U1331 (N_1331,In_301,In_322);
nand U1332 (N_1332,In_841,In_950);
nand U1333 (N_1333,In_982,In_153);
nor U1334 (N_1334,In_634,In_803);
or U1335 (N_1335,In_614,In_315);
and U1336 (N_1336,In_325,In_909);
or U1337 (N_1337,In_846,In_867);
or U1338 (N_1338,In_218,In_141);
or U1339 (N_1339,In_609,In_541);
and U1340 (N_1340,In_680,In_73);
or U1341 (N_1341,In_669,In_668);
or U1342 (N_1342,In_492,In_307);
nand U1343 (N_1343,In_624,In_984);
xor U1344 (N_1344,In_521,In_913);
and U1345 (N_1345,In_545,In_672);
nand U1346 (N_1346,In_225,In_604);
and U1347 (N_1347,In_97,In_610);
and U1348 (N_1348,In_433,In_428);
or U1349 (N_1349,In_58,In_523);
or U1350 (N_1350,In_461,In_763);
nand U1351 (N_1351,In_770,In_189);
nand U1352 (N_1352,In_939,In_649);
nand U1353 (N_1353,In_801,In_861);
xnor U1354 (N_1354,In_235,In_205);
nand U1355 (N_1355,In_772,In_86);
or U1356 (N_1356,In_263,In_577);
or U1357 (N_1357,In_193,In_473);
nor U1358 (N_1358,In_104,In_871);
nand U1359 (N_1359,In_356,In_833);
nand U1360 (N_1360,In_474,In_100);
nand U1361 (N_1361,In_61,In_905);
nand U1362 (N_1362,In_850,In_921);
nand U1363 (N_1363,In_701,In_812);
xnor U1364 (N_1364,In_873,In_330);
and U1365 (N_1365,In_594,In_790);
nor U1366 (N_1366,In_198,In_622);
nand U1367 (N_1367,In_281,In_778);
and U1368 (N_1368,In_871,In_596);
nand U1369 (N_1369,In_19,In_235);
xor U1370 (N_1370,In_762,In_404);
nand U1371 (N_1371,In_410,In_231);
or U1372 (N_1372,In_789,In_145);
nor U1373 (N_1373,In_758,In_193);
nand U1374 (N_1374,In_847,In_319);
xor U1375 (N_1375,In_489,In_216);
nor U1376 (N_1376,In_109,In_811);
or U1377 (N_1377,In_998,In_308);
xnor U1378 (N_1378,In_747,In_550);
or U1379 (N_1379,In_687,In_65);
or U1380 (N_1380,In_845,In_819);
nand U1381 (N_1381,In_442,In_425);
and U1382 (N_1382,In_610,In_1);
nor U1383 (N_1383,In_888,In_112);
or U1384 (N_1384,In_346,In_839);
and U1385 (N_1385,In_249,In_76);
and U1386 (N_1386,In_376,In_798);
nor U1387 (N_1387,In_447,In_804);
nor U1388 (N_1388,In_619,In_843);
xor U1389 (N_1389,In_424,In_791);
and U1390 (N_1390,In_331,In_553);
nand U1391 (N_1391,In_118,In_284);
nand U1392 (N_1392,In_569,In_256);
and U1393 (N_1393,In_127,In_91);
xor U1394 (N_1394,In_492,In_448);
or U1395 (N_1395,In_629,In_500);
and U1396 (N_1396,In_207,In_599);
or U1397 (N_1397,In_218,In_558);
and U1398 (N_1398,In_796,In_41);
or U1399 (N_1399,In_186,In_943);
nor U1400 (N_1400,In_197,In_919);
nor U1401 (N_1401,In_432,In_668);
or U1402 (N_1402,In_595,In_188);
and U1403 (N_1403,In_371,In_924);
nand U1404 (N_1404,In_880,In_370);
and U1405 (N_1405,In_344,In_826);
nor U1406 (N_1406,In_306,In_241);
xnor U1407 (N_1407,In_883,In_884);
nor U1408 (N_1408,In_574,In_270);
nor U1409 (N_1409,In_249,In_841);
and U1410 (N_1410,In_889,In_759);
or U1411 (N_1411,In_286,In_75);
or U1412 (N_1412,In_685,In_62);
and U1413 (N_1413,In_890,In_543);
or U1414 (N_1414,In_108,In_653);
and U1415 (N_1415,In_183,In_497);
nand U1416 (N_1416,In_313,In_779);
and U1417 (N_1417,In_150,In_487);
or U1418 (N_1418,In_99,In_616);
nand U1419 (N_1419,In_697,In_338);
nor U1420 (N_1420,In_374,In_164);
and U1421 (N_1421,In_532,In_756);
xor U1422 (N_1422,In_510,In_817);
or U1423 (N_1423,In_107,In_442);
and U1424 (N_1424,In_722,In_539);
xor U1425 (N_1425,In_482,In_910);
or U1426 (N_1426,In_883,In_5);
xnor U1427 (N_1427,In_703,In_329);
nand U1428 (N_1428,In_442,In_132);
nand U1429 (N_1429,In_406,In_108);
or U1430 (N_1430,In_936,In_913);
nand U1431 (N_1431,In_434,In_379);
and U1432 (N_1432,In_924,In_578);
or U1433 (N_1433,In_837,In_37);
or U1434 (N_1434,In_941,In_555);
nand U1435 (N_1435,In_214,In_468);
or U1436 (N_1436,In_360,In_453);
nor U1437 (N_1437,In_869,In_904);
or U1438 (N_1438,In_454,In_617);
nor U1439 (N_1439,In_747,In_84);
nor U1440 (N_1440,In_738,In_16);
or U1441 (N_1441,In_492,In_21);
nor U1442 (N_1442,In_216,In_124);
nand U1443 (N_1443,In_932,In_85);
nand U1444 (N_1444,In_534,In_404);
or U1445 (N_1445,In_909,In_151);
and U1446 (N_1446,In_846,In_621);
and U1447 (N_1447,In_384,In_775);
and U1448 (N_1448,In_166,In_95);
and U1449 (N_1449,In_815,In_257);
xor U1450 (N_1450,In_29,In_199);
or U1451 (N_1451,In_661,In_225);
nor U1452 (N_1452,In_188,In_218);
and U1453 (N_1453,In_618,In_2);
nor U1454 (N_1454,In_546,In_444);
nand U1455 (N_1455,In_601,In_993);
or U1456 (N_1456,In_702,In_957);
nand U1457 (N_1457,In_646,In_102);
and U1458 (N_1458,In_732,In_919);
nor U1459 (N_1459,In_5,In_100);
nor U1460 (N_1460,In_316,In_994);
or U1461 (N_1461,In_167,In_477);
nand U1462 (N_1462,In_969,In_369);
nor U1463 (N_1463,In_839,In_136);
or U1464 (N_1464,In_813,In_298);
or U1465 (N_1465,In_95,In_596);
nand U1466 (N_1466,In_297,In_187);
nor U1467 (N_1467,In_114,In_383);
nand U1468 (N_1468,In_811,In_615);
nand U1469 (N_1469,In_37,In_138);
nor U1470 (N_1470,In_106,In_645);
xor U1471 (N_1471,In_187,In_426);
and U1472 (N_1472,In_507,In_944);
and U1473 (N_1473,In_82,In_396);
and U1474 (N_1474,In_836,In_228);
nor U1475 (N_1475,In_933,In_384);
or U1476 (N_1476,In_878,In_467);
nor U1477 (N_1477,In_972,In_941);
xor U1478 (N_1478,In_344,In_960);
nand U1479 (N_1479,In_32,In_958);
xor U1480 (N_1480,In_448,In_377);
xor U1481 (N_1481,In_145,In_239);
nand U1482 (N_1482,In_123,In_406);
nor U1483 (N_1483,In_157,In_59);
and U1484 (N_1484,In_439,In_120);
nand U1485 (N_1485,In_286,In_748);
nand U1486 (N_1486,In_252,In_654);
or U1487 (N_1487,In_239,In_579);
or U1488 (N_1488,In_1,In_769);
nor U1489 (N_1489,In_8,In_312);
nor U1490 (N_1490,In_339,In_909);
nand U1491 (N_1491,In_876,In_779);
xor U1492 (N_1492,In_867,In_987);
xnor U1493 (N_1493,In_184,In_176);
xor U1494 (N_1494,In_929,In_791);
or U1495 (N_1495,In_283,In_915);
or U1496 (N_1496,In_340,In_399);
nand U1497 (N_1497,In_915,In_724);
nor U1498 (N_1498,In_367,In_204);
nor U1499 (N_1499,In_916,In_968);
or U1500 (N_1500,In_942,In_878);
or U1501 (N_1501,In_989,In_380);
or U1502 (N_1502,In_633,In_876);
and U1503 (N_1503,In_198,In_806);
xor U1504 (N_1504,In_382,In_316);
or U1505 (N_1505,In_760,In_276);
and U1506 (N_1506,In_345,In_405);
or U1507 (N_1507,In_380,In_766);
nand U1508 (N_1508,In_107,In_114);
nor U1509 (N_1509,In_428,In_576);
nand U1510 (N_1510,In_870,In_516);
or U1511 (N_1511,In_770,In_367);
nor U1512 (N_1512,In_85,In_90);
and U1513 (N_1513,In_202,In_153);
xnor U1514 (N_1514,In_660,In_191);
nand U1515 (N_1515,In_336,In_819);
and U1516 (N_1516,In_369,In_514);
nand U1517 (N_1517,In_243,In_305);
nand U1518 (N_1518,In_947,In_285);
nor U1519 (N_1519,In_461,In_539);
and U1520 (N_1520,In_579,In_84);
nand U1521 (N_1521,In_508,In_629);
and U1522 (N_1522,In_789,In_312);
nor U1523 (N_1523,In_352,In_381);
and U1524 (N_1524,In_983,In_272);
and U1525 (N_1525,In_298,In_539);
xnor U1526 (N_1526,In_772,In_774);
or U1527 (N_1527,In_554,In_338);
or U1528 (N_1528,In_664,In_66);
or U1529 (N_1529,In_455,In_861);
and U1530 (N_1530,In_201,In_487);
and U1531 (N_1531,In_538,In_92);
nand U1532 (N_1532,In_418,In_444);
xor U1533 (N_1533,In_825,In_448);
nor U1534 (N_1534,In_214,In_519);
nand U1535 (N_1535,In_193,In_946);
and U1536 (N_1536,In_13,In_910);
xnor U1537 (N_1537,In_30,In_861);
and U1538 (N_1538,In_289,In_692);
or U1539 (N_1539,In_940,In_537);
or U1540 (N_1540,In_661,In_391);
xnor U1541 (N_1541,In_891,In_258);
xnor U1542 (N_1542,In_865,In_16);
or U1543 (N_1543,In_663,In_726);
and U1544 (N_1544,In_521,In_825);
nor U1545 (N_1545,In_237,In_663);
or U1546 (N_1546,In_402,In_902);
nand U1547 (N_1547,In_631,In_280);
and U1548 (N_1548,In_135,In_298);
nand U1549 (N_1549,In_434,In_364);
or U1550 (N_1550,In_155,In_867);
xor U1551 (N_1551,In_724,In_806);
and U1552 (N_1552,In_515,In_881);
nor U1553 (N_1553,In_262,In_268);
or U1554 (N_1554,In_71,In_313);
nand U1555 (N_1555,In_643,In_517);
and U1556 (N_1556,In_260,In_23);
or U1557 (N_1557,In_729,In_536);
and U1558 (N_1558,In_740,In_486);
and U1559 (N_1559,In_930,In_757);
nand U1560 (N_1560,In_658,In_424);
nor U1561 (N_1561,In_749,In_38);
xor U1562 (N_1562,In_443,In_647);
or U1563 (N_1563,In_56,In_835);
nand U1564 (N_1564,In_650,In_381);
and U1565 (N_1565,In_845,In_349);
nor U1566 (N_1566,In_567,In_458);
xor U1567 (N_1567,In_247,In_495);
xnor U1568 (N_1568,In_242,In_167);
and U1569 (N_1569,In_36,In_903);
nor U1570 (N_1570,In_74,In_909);
or U1571 (N_1571,In_650,In_107);
xor U1572 (N_1572,In_963,In_572);
or U1573 (N_1573,In_804,In_833);
or U1574 (N_1574,In_768,In_401);
or U1575 (N_1575,In_944,In_840);
and U1576 (N_1576,In_131,In_329);
xor U1577 (N_1577,In_446,In_644);
or U1578 (N_1578,In_761,In_638);
and U1579 (N_1579,In_538,In_563);
nor U1580 (N_1580,In_320,In_166);
or U1581 (N_1581,In_817,In_600);
or U1582 (N_1582,In_378,In_929);
and U1583 (N_1583,In_200,In_917);
nor U1584 (N_1584,In_403,In_773);
and U1585 (N_1585,In_350,In_808);
xor U1586 (N_1586,In_830,In_133);
nand U1587 (N_1587,In_412,In_303);
or U1588 (N_1588,In_250,In_497);
and U1589 (N_1589,In_462,In_963);
nand U1590 (N_1590,In_223,In_778);
or U1591 (N_1591,In_27,In_742);
nand U1592 (N_1592,In_105,In_259);
or U1593 (N_1593,In_317,In_409);
nand U1594 (N_1594,In_556,In_244);
and U1595 (N_1595,In_997,In_873);
nand U1596 (N_1596,In_413,In_990);
nor U1597 (N_1597,In_28,In_471);
or U1598 (N_1598,In_796,In_206);
or U1599 (N_1599,In_94,In_269);
or U1600 (N_1600,In_221,In_917);
nor U1601 (N_1601,In_861,In_682);
nor U1602 (N_1602,In_285,In_560);
nand U1603 (N_1603,In_105,In_641);
nor U1604 (N_1604,In_763,In_585);
nand U1605 (N_1605,In_267,In_47);
and U1606 (N_1606,In_537,In_231);
nor U1607 (N_1607,In_491,In_667);
nand U1608 (N_1608,In_672,In_376);
nor U1609 (N_1609,In_226,In_956);
xor U1610 (N_1610,In_927,In_28);
nand U1611 (N_1611,In_450,In_55);
nor U1612 (N_1612,In_375,In_129);
and U1613 (N_1613,In_418,In_810);
nand U1614 (N_1614,In_933,In_735);
nand U1615 (N_1615,In_733,In_373);
or U1616 (N_1616,In_11,In_384);
nand U1617 (N_1617,In_223,In_102);
xor U1618 (N_1618,In_96,In_457);
nor U1619 (N_1619,In_898,In_583);
nor U1620 (N_1620,In_223,In_137);
or U1621 (N_1621,In_409,In_670);
xnor U1622 (N_1622,In_459,In_122);
nand U1623 (N_1623,In_310,In_271);
or U1624 (N_1624,In_477,In_198);
nor U1625 (N_1625,In_191,In_87);
xor U1626 (N_1626,In_758,In_85);
nor U1627 (N_1627,In_9,In_156);
nor U1628 (N_1628,In_325,In_678);
xnor U1629 (N_1629,In_276,In_460);
nand U1630 (N_1630,In_760,In_358);
or U1631 (N_1631,In_370,In_900);
or U1632 (N_1632,In_791,In_471);
nand U1633 (N_1633,In_947,In_328);
xnor U1634 (N_1634,In_812,In_93);
xor U1635 (N_1635,In_397,In_0);
and U1636 (N_1636,In_899,In_176);
nor U1637 (N_1637,In_292,In_741);
and U1638 (N_1638,In_247,In_858);
nand U1639 (N_1639,In_858,In_56);
nor U1640 (N_1640,In_132,In_116);
and U1641 (N_1641,In_474,In_743);
or U1642 (N_1642,In_694,In_909);
and U1643 (N_1643,In_384,In_284);
nor U1644 (N_1644,In_584,In_479);
and U1645 (N_1645,In_547,In_411);
nand U1646 (N_1646,In_158,In_62);
or U1647 (N_1647,In_868,In_944);
or U1648 (N_1648,In_672,In_817);
nor U1649 (N_1649,In_701,In_439);
and U1650 (N_1650,In_444,In_134);
and U1651 (N_1651,In_852,In_920);
nor U1652 (N_1652,In_250,In_470);
and U1653 (N_1653,In_932,In_565);
or U1654 (N_1654,In_684,In_654);
and U1655 (N_1655,In_614,In_24);
nand U1656 (N_1656,In_367,In_134);
or U1657 (N_1657,In_43,In_161);
xnor U1658 (N_1658,In_949,In_694);
nor U1659 (N_1659,In_496,In_127);
nand U1660 (N_1660,In_327,In_774);
nand U1661 (N_1661,In_959,In_238);
and U1662 (N_1662,In_561,In_746);
or U1663 (N_1663,In_478,In_135);
nor U1664 (N_1664,In_563,In_152);
nor U1665 (N_1665,In_130,In_909);
nor U1666 (N_1666,In_411,In_850);
and U1667 (N_1667,In_812,In_106);
and U1668 (N_1668,In_436,In_300);
nand U1669 (N_1669,In_835,In_760);
nor U1670 (N_1670,In_3,In_905);
and U1671 (N_1671,In_931,In_712);
nor U1672 (N_1672,In_884,In_621);
or U1673 (N_1673,In_578,In_284);
xor U1674 (N_1674,In_799,In_292);
nand U1675 (N_1675,In_668,In_772);
or U1676 (N_1676,In_584,In_337);
or U1677 (N_1677,In_801,In_86);
or U1678 (N_1678,In_88,In_664);
nand U1679 (N_1679,In_974,In_372);
and U1680 (N_1680,In_785,In_682);
nand U1681 (N_1681,In_83,In_343);
or U1682 (N_1682,In_818,In_70);
nand U1683 (N_1683,In_327,In_312);
xor U1684 (N_1684,In_824,In_564);
nand U1685 (N_1685,In_647,In_554);
or U1686 (N_1686,In_906,In_547);
nor U1687 (N_1687,In_963,In_653);
and U1688 (N_1688,In_725,In_508);
or U1689 (N_1689,In_824,In_568);
and U1690 (N_1690,In_676,In_684);
nand U1691 (N_1691,In_932,In_84);
xor U1692 (N_1692,In_511,In_700);
and U1693 (N_1693,In_995,In_756);
and U1694 (N_1694,In_522,In_296);
nor U1695 (N_1695,In_899,In_318);
nor U1696 (N_1696,In_78,In_631);
and U1697 (N_1697,In_893,In_280);
and U1698 (N_1698,In_648,In_517);
nor U1699 (N_1699,In_579,In_397);
xor U1700 (N_1700,In_979,In_97);
or U1701 (N_1701,In_130,In_373);
or U1702 (N_1702,In_450,In_756);
or U1703 (N_1703,In_16,In_216);
nand U1704 (N_1704,In_30,In_669);
or U1705 (N_1705,In_718,In_164);
nand U1706 (N_1706,In_549,In_950);
nor U1707 (N_1707,In_960,In_422);
nand U1708 (N_1708,In_918,In_150);
or U1709 (N_1709,In_765,In_329);
and U1710 (N_1710,In_574,In_719);
nor U1711 (N_1711,In_776,In_380);
xnor U1712 (N_1712,In_39,In_608);
or U1713 (N_1713,In_638,In_322);
xor U1714 (N_1714,In_665,In_461);
and U1715 (N_1715,In_159,In_619);
or U1716 (N_1716,In_932,In_731);
and U1717 (N_1717,In_465,In_664);
and U1718 (N_1718,In_327,In_944);
and U1719 (N_1719,In_161,In_664);
and U1720 (N_1720,In_96,In_94);
and U1721 (N_1721,In_356,In_993);
and U1722 (N_1722,In_374,In_628);
nor U1723 (N_1723,In_203,In_738);
and U1724 (N_1724,In_787,In_978);
or U1725 (N_1725,In_195,In_749);
nand U1726 (N_1726,In_796,In_114);
nor U1727 (N_1727,In_373,In_695);
and U1728 (N_1728,In_127,In_908);
nand U1729 (N_1729,In_739,In_913);
xor U1730 (N_1730,In_27,In_87);
nand U1731 (N_1731,In_990,In_154);
or U1732 (N_1732,In_314,In_863);
xor U1733 (N_1733,In_475,In_980);
nor U1734 (N_1734,In_783,In_534);
and U1735 (N_1735,In_37,In_843);
nand U1736 (N_1736,In_378,In_439);
nor U1737 (N_1737,In_161,In_556);
or U1738 (N_1738,In_641,In_688);
nand U1739 (N_1739,In_189,In_103);
or U1740 (N_1740,In_469,In_237);
or U1741 (N_1741,In_735,In_276);
and U1742 (N_1742,In_373,In_722);
or U1743 (N_1743,In_498,In_52);
nand U1744 (N_1744,In_55,In_830);
or U1745 (N_1745,In_618,In_205);
nor U1746 (N_1746,In_47,In_340);
xnor U1747 (N_1747,In_222,In_683);
or U1748 (N_1748,In_967,In_315);
nand U1749 (N_1749,In_421,In_907);
and U1750 (N_1750,In_106,In_383);
nor U1751 (N_1751,In_17,In_194);
and U1752 (N_1752,In_28,In_30);
or U1753 (N_1753,In_648,In_929);
nor U1754 (N_1754,In_951,In_120);
and U1755 (N_1755,In_107,In_689);
or U1756 (N_1756,In_969,In_855);
nor U1757 (N_1757,In_456,In_981);
nand U1758 (N_1758,In_779,In_260);
xnor U1759 (N_1759,In_175,In_732);
or U1760 (N_1760,In_912,In_765);
and U1761 (N_1761,In_438,In_368);
nor U1762 (N_1762,In_494,In_934);
and U1763 (N_1763,In_503,In_135);
xnor U1764 (N_1764,In_923,In_173);
nand U1765 (N_1765,In_73,In_635);
nand U1766 (N_1766,In_520,In_643);
nand U1767 (N_1767,In_470,In_606);
nor U1768 (N_1768,In_705,In_243);
or U1769 (N_1769,In_677,In_327);
nor U1770 (N_1770,In_957,In_582);
nor U1771 (N_1771,In_734,In_550);
and U1772 (N_1772,In_773,In_194);
nor U1773 (N_1773,In_623,In_279);
nor U1774 (N_1774,In_429,In_564);
nor U1775 (N_1775,In_906,In_355);
nand U1776 (N_1776,In_809,In_755);
and U1777 (N_1777,In_602,In_428);
nor U1778 (N_1778,In_838,In_947);
or U1779 (N_1779,In_422,In_922);
nor U1780 (N_1780,In_346,In_956);
or U1781 (N_1781,In_139,In_489);
or U1782 (N_1782,In_243,In_890);
nand U1783 (N_1783,In_986,In_551);
nand U1784 (N_1784,In_133,In_949);
and U1785 (N_1785,In_152,In_656);
and U1786 (N_1786,In_139,In_15);
or U1787 (N_1787,In_557,In_50);
or U1788 (N_1788,In_460,In_734);
nand U1789 (N_1789,In_59,In_855);
and U1790 (N_1790,In_810,In_492);
nand U1791 (N_1791,In_189,In_326);
nor U1792 (N_1792,In_244,In_168);
or U1793 (N_1793,In_548,In_492);
xor U1794 (N_1794,In_646,In_429);
nand U1795 (N_1795,In_707,In_28);
and U1796 (N_1796,In_912,In_984);
nor U1797 (N_1797,In_60,In_662);
nand U1798 (N_1798,In_675,In_278);
and U1799 (N_1799,In_434,In_419);
or U1800 (N_1800,In_726,In_835);
and U1801 (N_1801,In_124,In_894);
xor U1802 (N_1802,In_316,In_85);
or U1803 (N_1803,In_36,In_569);
nand U1804 (N_1804,In_601,In_934);
or U1805 (N_1805,In_963,In_582);
nor U1806 (N_1806,In_981,In_240);
nor U1807 (N_1807,In_746,In_192);
nor U1808 (N_1808,In_520,In_660);
nor U1809 (N_1809,In_152,In_125);
nand U1810 (N_1810,In_26,In_686);
and U1811 (N_1811,In_594,In_740);
or U1812 (N_1812,In_791,In_441);
or U1813 (N_1813,In_910,In_439);
and U1814 (N_1814,In_467,In_152);
nor U1815 (N_1815,In_19,In_874);
nor U1816 (N_1816,In_398,In_966);
xor U1817 (N_1817,In_364,In_35);
nor U1818 (N_1818,In_446,In_954);
nor U1819 (N_1819,In_489,In_14);
or U1820 (N_1820,In_390,In_91);
nor U1821 (N_1821,In_51,In_434);
and U1822 (N_1822,In_464,In_530);
or U1823 (N_1823,In_530,In_432);
or U1824 (N_1824,In_482,In_596);
nor U1825 (N_1825,In_868,In_218);
nand U1826 (N_1826,In_769,In_873);
nor U1827 (N_1827,In_398,In_940);
or U1828 (N_1828,In_524,In_781);
and U1829 (N_1829,In_857,In_369);
nor U1830 (N_1830,In_820,In_254);
nor U1831 (N_1831,In_104,In_544);
and U1832 (N_1832,In_66,In_927);
or U1833 (N_1833,In_885,In_279);
xor U1834 (N_1834,In_982,In_116);
nand U1835 (N_1835,In_259,In_660);
and U1836 (N_1836,In_429,In_839);
nor U1837 (N_1837,In_442,In_876);
nand U1838 (N_1838,In_458,In_739);
and U1839 (N_1839,In_138,In_246);
and U1840 (N_1840,In_842,In_316);
nand U1841 (N_1841,In_94,In_629);
and U1842 (N_1842,In_846,In_627);
and U1843 (N_1843,In_786,In_357);
nor U1844 (N_1844,In_101,In_681);
xnor U1845 (N_1845,In_836,In_598);
nand U1846 (N_1846,In_215,In_82);
nand U1847 (N_1847,In_183,In_900);
or U1848 (N_1848,In_74,In_499);
nand U1849 (N_1849,In_442,In_561);
or U1850 (N_1850,In_823,In_810);
xnor U1851 (N_1851,In_717,In_274);
and U1852 (N_1852,In_333,In_206);
nor U1853 (N_1853,In_139,In_991);
nor U1854 (N_1854,In_106,In_210);
and U1855 (N_1855,In_933,In_812);
or U1856 (N_1856,In_604,In_412);
or U1857 (N_1857,In_852,In_220);
xor U1858 (N_1858,In_893,In_197);
or U1859 (N_1859,In_677,In_850);
nand U1860 (N_1860,In_665,In_901);
or U1861 (N_1861,In_421,In_446);
or U1862 (N_1862,In_291,In_621);
and U1863 (N_1863,In_766,In_315);
and U1864 (N_1864,In_623,In_368);
and U1865 (N_1865,In_852,In_123);
or U1866 (N_1866,In_10,In_826);
or U1867 (N_1867,In_64,In_130);
nand U1868 (N_1868,In_495,In_759);
nand U1869 (N_1869,In_196,In_337);
xor U1870 (N_1870,In_697,In_129);
xor U1871 (N_1871,In_263,In_174);
or U1872 (N_1872,In_289,In_577);
and U1873 (N_1873,In_667,In_255);
and U1874 (N_1874,In_792,In_409);
and U1875 (N_1875,In_50,In_488);
and U1876 (N_1876,In_403,In_268);
nand U1877 (N_1877,In_234,In_144);
and U1878 (N_1878,In_72,In_277);
nor U1879 (N_1879,In_442,In_785);
nor U1880 (N_1880,In_382,In_396);
nand U1881 (N_1881,In_941,In_225);
and U1882 (N_1882,In_581,In_853);
nor U1883 (N_1883,In_909,In_802);
and U1884 (N_1884,In_518,In_863);
nand U1885 (N_1885,In_958,In_355);
and U1886 (N_1886,In_194,In_201);
nand U1887 (N_1887,In_909,In_507);
and U1888 (N_1888,In_224,In_281);
nor U1889 (N_1889,In_315,In_928);
nor U1890 (N_1890,In_140,In_656);
and U1891 (N_1891,In_142,In_752);
and U1892 (N_1892,In_958,In_609);
nor U1893 (N_1893,In_895,In_248);
and U1894 (N_1894,In_247,In_877);
or U1895 (N_1895,In_356,In_644);
nand U1896 (N_1896,In_719,In_925);
nor U1897 (N_1897,In_78,In_594);
xor U1898 (N_1898,In_522,In_750);
nand U1899 (N_1899,In_311,In_182);
nor U1900 (N_1900,In_703,In_277);
and U1901 (N_1901,In_519,In_143);
nor U1902 (N_1902,In_494,In_465);
nand U1903 (N_1903,In_767,In_986);
nand U1904 (N_1904,In_683,In_441);
nand U1905 (N_1905,In_845,In_75);
nor U1906 (N_1906,In_978,In_139);
and U1907 (N_1907,In_602,In_219);
and U1908 (N_1908,In_199,In_572);
nand U1909 (N_1909,In_674,In_925);
nand U1910 (N_1910,In_466,In_345);
or U1911 (N_1911,In_272,In_382);
nand U1912 (N_1912,In_868,In_605);
and U1913 (N_1913,In_783,In_519);
nor U1914 (N_1914,In_972,In_253);
and U1915 (N_1915,In_412,In_471);
xnor U1916 (N_1916,In_736,In_908);
or U1917 (N_1917,In_427,In_47);
nand U1918 (N_1918,In_427,In_472);
nand U1919 (N_1919,In_798,In_541);
nor U1920 (N_1920,In_459,In_918);
and U1921 (N_1921,In_91,In_412);
nor U1922 (N_1922,In_470,In_872);
nand U1923 (N_1923,In_507,In_174);
or U1924 (N_1924,In_420,In_872);
and U1925 (N_1925,In_274,In_713);
and U1926 (N_1926,In_410,In_130);
and U1927 (N_1927,In_69,In_46);
nand U1928 (N_1928,In_282,In_517);
and U1929 (N_1929,In_85,In_557);
nand U1930 (N_1930,In_140,In_274);
and U1931 (N_1931,In_905,In_507);
xnor U1932 (N_1932,In_917,In_656);
or U1933 (N_1933,In_394,In_152);
nor U1934 (N_1934,In_508,In_550);
xnor U1935 (N_1935,In_990,In_901);
nor U1936 (N_1936,In_467,In_30);
or U1937 (N_1937,In_683,In_44);
nand U1938 (N_1938,In_795,In_872);
or U1939 (N_1939,In_410,In_101);
nand U1940 (N_1940,In_357,In_172);
nand U1941 (N_1941,In_479,In_845);
nand U1942 (N_1942,In_451,In_540);
or U1943 (N_1943,In_591,In_283);
nand U1944 (N_1944,In_360,In_418);
nand U1945 (N_1945,In_169,In_923);
or U1946 (N_1946,In_808,In_460);
or U1947 (N_1947,In_940,In_300);
nor U1948 (N_1948,In_82,In_69);
nor U1949 (N_1949,In_571,In_362);
or U1950 (N_1950,In_796,In_57);
nor U1951 (N_1951,In_735,In_69);
nor U1952 (N_1952,In_135,In_515);
or U1953 (N_1953,In_622,In_370);
or U1954 (N_1954,In_867,In_928);
nor U1955 (N_1955,In_362,In_146);
nor U1956 (N_1956,In_33,In_988);
or U1957 (N_1957,In_196,In_919);
or U1958 (N_1958,In_708,In_776);
and U1959 (N_1959,In_498,In_871);
or U1960 (N_1960,In_124,In_356);
and U1961 (N_1961,In_686,In_535);
or U1962 (N_1962,In_180,In_774);
nor U1963 (N_1963,In_343,In_437);
nand U1964 (N_1964,In_815,In_879);
nand U1965 (N_1965,In_404,In_183);
nand U1966 (N_1966,In_591,In_979);
xnor U1967 (N_1967,In_804,In_491);
and U1968 (N_1968,In_938,In_172);
or U1969 (N_1969,In_544,In_70);
xnor U1970 (N_1970,In_666,In_924);
nor U1971 (N_1971,In_305,In_556);
nor U1972 (N_1972,In_46,In_714);
nand U1973 (N_1973,In_624,In_777);
nand U1974 (N_1974,In_348,In_361);
xnor U1975 (N_1975,In_866,In_545);
and U1976 (N_1976,In_550,In_525);
or U1977 (N_1977,In_900,In_92);
and U1978 (N_1978,In_742,In_970);
nand U1979 (N_1979,In_922,In_475);
or U1980 (N_1980,In_776,In_325);
nor U1981 (N_1981,In_364,In_716);
and U1982 (N_1982,In_682,In_520);
nor U1983 (N_1983,In_262,In_336);
nor U1984 (N_1984,In_29,In_401);
nor U1985 (N_1985,In_642,In_931);
or U1986 (N_1986,In_229,In_868);
xor U1987 (N_1987,In_503,In_241);
and U1988 (N_1988,In_654,In_3);
xnor U1989 (N_1989,In_738,In_960);
xor U1990 (N_1990,In_563,In_625);
and U1991 (N_1991,In_856,In_658);
or U1992 (N_1992,In_326,In_137);
and U1993 (N_1993,In_70,In_972);
nor U1994 (N_1994,In_748,In_205);
nor U1995 (N_1995,In_334,In_574);
or U1996 (N_1996,In_763,In_177);
xor U1997 (N_1997,In_215,In_65);
and U1998 (N_1998,In_664,In_242);
nand U1999 (N_1999,In_934,In_716);
and U2000 (N_2000,In_331,In_754);
and U2001 (N_2001,In_73,In_838);
xor U2002 (N_2002,In_611,In_937);
nand U2003 (N_2003,In_652,In_341);
or U2004 (N_2004,In_409,In_451);
or U2005 (N_2005,In_564,In_137);
nor U2006 (N_2006,In_400,In_376);
or U2007 (N_2007,In_527,In_8);
or U2008 (N_2008,In_453,In_25);
xnor U2009 (N_2009,In_6,In_714);
nand U2010 (N_2010,In_886,In_923);
and U2011 (N_2011,In_301,In_116);
and U2012 (N_2012,In_241,In_152);
nand U2013 (N_2013,In_832,In_381);
nand U2014 (N_2014,In_27,In_393);
xnor U2015 (N_2015,In_709,In_265);
and U2016 (N_2016,In_106,In_762);
and U2017 (N_2017,In_507,In_928);
nor U2018 (N_2018,In_576,In_408);
nor U2019 (N_2019,In_889,In_864);
xor U2020 (N_2020,In_948,In_706);
nand U2021 (N_2021,In_797,In_248);
nand U2022 (N_2022,In_501,In_410);
xor U2023 (N_2023,In_472,In_398);
xor U2024 (N_2024,In_336,In_842);
and U2025 (N_2025,In_950,In_739);
nand U2026 (N_2026,In_485,In_472);
and U2027 (N_2027,In_477,In_341);
xor U2028 (N_2028,In_422,In_631);
or U2029 (N_2029,In_326,In_494);
or U2030 (N_2030,In_188,In_356);
nand U2031 (N_2031,In_682,In_292);
nor U2032 (N_2032,In_681,In_396);
and U2033 (N_2033,In_796,In_631);
xor U2034 (N_2034,In_149,In_639);
nand U2035 (N_2035,In_17,In_914);
nand U2036 (N_2036,In_360,In_963);
and U2037 (N_2037,In_565,In_289);
or U2038 (N_2038,In_893,In_602);
nand U2039 (N_2039,In_971,In_955);
or U2040 (N_2040,In_850,In_795);
nor U2041 (N_2041,In_120,In_362);
or U2042 (N_2042,In_616,In_770);
nand U2043 (N_2043,In_682,In_851);
nor U2044 (N_2044,In_397,In_862);
nor U2045 (N_2045,In_496,In_275);
nand U2046 (N_2046,In_534,In_412);
nor U2047 (N_2047,In_291,In_28);
and U2048 (N_2048,In_554,In_42);
and U2049 (N_2049,In_53,In_539);
nand U2050 (N_2050,In_399,In_837);
and U2051 (N_2051,In_423,In_229);
and U2052 (N_2052,In_309,In_94);
nand U2053 (N_2053,In_157,In_953);
xor U2054 (N_2054,In_848,In_572);
nand U2055 (N_2055,In_761,In_760);
nand U2056 (N_2056,In_810,In_956);
or U2057 (N_2057,In_587,In_964);
or U2058 (N_2058,In_853,In_172);
nand U2059 (N_2059,In_957,In_414);
xnor U2060 (N_2060,In_340,In_158);
or U2061 (N_2061,In_25,In_904);
xor U2062 (N_2062,In_698,In_427);
and U2063 (N_2063,In_244,In_129);
nor U2064 (N_2064,In_498,In_547);
and U2065 (N_2065,In_100,In_713);
or U2066 (N_2066,In_463,In_285);
nor U2067 (N_2067,In_411,In_133);
and U2068 (N_2068,In_698,In_943);
or U2069 (N_2069,In_206,In_518);
or U2070 (N_2070,In_278,In_411);
or U2071 (N_2071,In_640,In_683);
or U2072 (N_2072,In_380,In_895);
or U2073 (N_2073,In_802,In_610);
nand U2074 (N_2074,In_630,In_101);
and U2075 (N_2075,In_224,In_676);
or U2076 (N_2076,In_792,In_757);
xor U2077 (N_2077,In_223,In_499);
and U2078 (N_2078,In_814,In_878);
or U2079 (N_2079,In_193,In_241);
nor U2080 (N_2080,In_801,In_906);
nand U2081 (N_2081,In_985,In_622);
or U2082 (N_2082,In_894,In_77);
or U2083 (N_2083,In_836,In_129);
or U2084 (N_2084,In_252,In_303);
and U2085 (N_2085,In_943,In_402);
or U2086 (N_2086,In_262,In_181);
nor U2087 (N_2087,In_57,In_186);
or U2088 (N_2088,In_885,In_662);
nor U2089 (N_2089,In_875,In_236);
or U2090 (N_2090,In_549,In_976);
nand U2091 (N_2091,In_262,In_353);
nor U2092 (N_2092,In_318,In_372);
and U2093 (N_2093,In_706,In_220);
nor U2094 (N_2094,In_383,In_422);
nor U2095 (N_2095,In_216,In_206);
xor U2096 (N_2096,In_635,In_602);
nand U2097 (N_2097,In_520,In_248);
and U2098 (N_2098,In_595,In_782);
xnor U2099 (N_2099,In_119,In_439);
nor U2100 (N_2100,In_376,In_831);
or U2101 (N_2101,In_15,In_614);
nor U2102 (N_2102,In_282,In_939);
nor U2103 (N_2103,In_375,In_383);
and U2104 (N_2104,In_750,In_712);
nand U2105 (N_2105,In_423,In_848);
or U2106 (N_2106,In_256,In_984);
nand U2107 (N_2107,In_629,In_931);
nor U2108 (N_2108,In_24,In_83);
and U2109 (N_2109,In_600,In_689);
or U2110 (N_2110,In_536,In_927);
or U2111 (N_2111,In_496,In_670);
or U2112 (N_2112,In_12,In_795);
or U2113 (N_2113,In_897,In_607);
xnor U2114 (N_2114,In_134,In_55);
or U2115 (N_2115,In_823,In_764);
or U2116 (N_2116,In_884,In_999);
and U2117 (N_2117,In_846,In_357);
xor U2118 (N_2118,In_787,In_88);
nand U2119 (N_2119,In_981,In_630);
and U2120 (N_2120,In_362,In_714);
and U2121 (N_2121,In_965,In_704);
nor U2122 (N_2122,In_217,In_991);
xor U2123 (N_2123,In_750,In_626);
nor U2124 (N_2124,In_723,In_913);
or U2125 (N_2125,In_478,In_991);
or U2126 (N_2126,In_384,In_669);
and U2127 (N_2127,In_837,In_635);
nor U2128 (N_2128,In_8,In_408);
nor U2129 (N_2129,In_437,In_17);
nor U2130 (N_2130,In_468,In_212);
and U2131 (N_2131,In_435,In_323);
nand U2132 (N_2132,In_863,In_291);
nor U2133 (N_2133,In_718,In_898);
nor U2134 (N_2134,In_243,In_801);
nor U2135 (N_2135,In_803,In_182);
and U2136 (N_2136,In_981,In_336);
nand U2137 (N_2137,In_637,In_285);
or U2138 (N_2138,In_760,In_872);
and U2139 (N_2139,In_437,In_687);
nor U2140 (N_2140,In_328,In_532);
nand U2141 (N_2141,In_916,In_949);
xor U2142 (N_2142,In_862,In_147);
or U2143 (N_2143,In_819,In_897);
nand U2144 (N_2144,In_615,In_862);
nor U2145 (N_2145,In_839,In_657);
nand U2146 (N_2146,In_67,In_36);
xnor U2147 (N_2147,In_123,In_359);
nor U2148 (N_2148,In_967,In_346);
nor U2149 (N_2149,In_740,In_140);
nand U2150 (N_2150,In_898,In_815);
and U2151 (N_2151,In_21,In_173);
nand U2152 (N_2152,In_487,In_776);
and U2153 (N_2153,In_799,In_883);
nand U2154 (N_2154,In_535,In_423);
and U2155 (N_2155,In_538,In_979);
and U2156 (N_2156,In_939,In_180);
or U2157 (N_2157,In_479,In_236);
nand U2158 (N_2158,In_137,In_629);
nor U2159 (N_2159,In_224,In_985);
nor U2160 (N_2160,In_136,In_542);
nor U2161 (N_2161,In_834,In_700);
nand U2162 (N_2162,In_387,In_879);
nor U2163 (N_2163,In_680,In_761);
and U2164 (N_2164,In_16,In_64);
or U2165 (N_2165,In_670,In_328);
nand U2166 (N_2166,In_398,In_213);
xnor U2167 (N_2167,In_556,In_290);
nand U2168 (N_2168,In_560,In_413);
and U2169 (N_2169,In_481,In_188);
nand U2170 (N_2170,In_919,In_152);
nand U2171 (N_2171,In_352,In_656);
nand U2172 (N_2172,In_794,In_2);
or U2173 (N_2173,In_416,In_540);
or U2174 (N_2174,In_997,In_234);
or U2175 (N_2175,In_923,In_900);
nor U2176 (N_2176,In_68,In_48);
or U2177 (N_2177,In_694,In_36);
and U2178 (N_2178,In_355,In_307);
nand U2179 (N_2179,In_637,In_179);
and U2180 (N_2180,In_973,In_126);
nand U2181 (N_2181,In_620,In_984);
nor U2182 (N_2182,In_671,In_140);
and U2183 (N_2183,In_911,In_306);
and U2184 (N_2184,In_345,In_436);
nand U2185 (N_2185,In_629,In_680);
nor U2186 (N_2186,In_675,In_628);
nand U2187 (N_2187,In_162,In_533);
and U2188 (N_2188,In_174,In_35);
and U2189 (N_2189,In_82,In_858);
and U2190 (N_2190,In_587,In_808);
nand U2191 (N_2191,In_411,In_69);
and U2192 (N_2192,In_831,In_769);
nor U2193 (N_2193,In_149,In_624);
or U2194 (N_2194,In_454,In_623);
or U2195 (N_2195,In_906,In_183);
and U2196 (N_2196,In_11,In_158);
and U2197 (N_2197,In_9,In_457);
or U2198 (N_2198,In_41,In_642);
or U2199 (N_2199,In_624,In_5);
xor U2200 (N_2200,In_667,In_329);
nand U2201 (N_2201,In_157,In_687);
and U2202 (N_2202,In_232,In_201);
and U2203 (N_2203,In_438,In_151);
nor U2204 (N_2204,In_681,In_93);
nor U2205 (N_2205,In_775,In_836);
nand U2206 (N_2206,In_903,In_481);
or U2207 (N_2207,In_441,In_620);
xor U2208 (N_2208,In_237,In_529);
and U2209 (N_2209,In_808,In_312);
and U2210 (N_2210,In_798,In_247);
and U2211 (N_2211,In_582,In_585);
or U2212 (N_2212,In_675,In_827);
nor U2213 (N_2213,In_301,In_287);
nor U2214 (N_2214,In_544,In_220);
xor U2215 (N_2215,In_947,In_275);
nor U2216 (N_2216,In_202,In_457);
nand U2217 (N_2217,In_527,In_164);
nor U2218 (N_2218,In_319,In_133);
or U2219 (N_2219,In_411,In_615);
and U2220 (N_2220,In_60,In_733);
or U2221 (N_2221,In_937,In_52);
or U2222 (N_2222,In_304,In_332);
and U2223 (N_2223,In_913,In_71);
and U2224 (N_2224,In_718,In_322);
and U2225 (N_2225,In_993,In_288);
nor U2226 (N_2226,In_396,In_919);
nor U2227 (N_2227,In_273,In_834);
nor U2228 (N_2228,In_951,In_359);
nand U2229 (N_2229,In_295,In_53);
nand U2230 (N_2230,In_545,In_21);
nor U2231 (N_2231,In_639,In_690);
nand U2232 (N_2232,In_886,In_704);
nor U2233 (N_2233,In_122,In_733);
nand U2234 (N_2234,In_729,In_448);
nor U2235 (N_2235,In_375,In_781);
or U2236 (N_2236,In_901,In_378);
nor U2237 (N_2237,In_193,In_636);
nor U2238 (N_2238,In_736,In_590);
or U2239 (N_2239,In_34,In_678);
nor U2240 (N_2240,In_605,In_785);
and U2241 (N_2241,In_12,In_246);
and U2242 (N_2242,In_953,In_107);
or U2243 (N_2243,In_177,In_10);
nor U2244 (N_2244,In_778,In_528);
nor U2245 (N_2245,In_925,In_882);
or U2246 (N_2246,In_420,In_637);
and U2247 (N_2247,In_790,In_949);
xor U2248 (N_2248,In_820,In_196);
nor U2249 (N_2249,In_905,In_520);
and U2250 (N_2250,In_54,In_811);
nand U2251 (N_2251,In_383,In_600);
nand U2252 (N_2252,In_561,In_574);
nand U2253 (N_2253,In_709,In_801);
nor U2254 (N_2254,In_414,In_396);
nand U2255 (N_2255,In_217,In_400);
xor U2256 (N_2256,In_650,In_407);
and U2257 (N_2257,In_106,In_147);
nand U2258 (N_2258,In_437,In_730);
and U2259 (N_2259,In_651,In_570);
nand U2260 (N_2260,In_920,In_168);
nor U2261 (N_2261,In_422,In_835);
xnor U2262 (N_2262,In_285,In_640);
and U2263 (N_2263,In_73,In_177);
nor U2264 (N_2264,In_665,In_799);
nand U2265 (N_2265,In_229,In_59);
or U2266 (N_2266,In_255,In_981);
nor U2267 (N_2267,In_776,In_142);
nor U2268 (N_2268,In_23,In_665);
nor U2269 (N_2269,In_403,In_285);
and U2270 (N_2270,In_14,In_787);
nand U2271 (N_2271,In_359,In_277);
or U2272 (N_2272,In_739,In_777);
nand U2273 (N_2273,In_967,In_158);
nand U2274 (N_2274,In_795,In_333);
and U2275 (N_2275,In_805,In_235);
and U2276 (N_2276,In_843,In_324);
nor U2277 (N_2277,In_19,In_241);
or U2278 (N_2278,In_482,In_220);
nand U2279 (N_2279,In_703,In_196);
nand U2280 (N_2280,In_992,In_641);
or U2281 (N_2281,In_570,In_761);
and U2282 (N_2282,In_912,In_808);
or U2283 (N_2283,In_895,In_827);
or U2284 (N_2284,In_986,In_867);
or U2285 (N_2285,In_595,In_41);
and U2286 (N_2286,In_830,In_480);
nor U2287 (N_2287,In_337,In_731);
nand U2288 (N_2288,In_117,In_41);
or U2289 (N_2289,In_779,In_619);
or U2290 (N_2290,In_751,In_381);
and U2291 (N_2291,In_220,In_258);
xor U2292 (N_2292,In_387,In_793);
and U2293 (N_2293,In_508,In_67);
and U2294 (N_2294,In_904,In_466);
nor U2295 (N_2295,In_533,In_666);
nand U2296 (N_2296,In_855,In_348);
xor U2297 (N_2297,In_694,In_565);
and U2298 (N_2298,In_894,In_186);
and U2299 (N_2299,In_875,In_861);
or U2300 (N_2300,In_880,In_438);
or U2301 (N_2301,In_394,In_629);
xnor U2302 (N_2302,In_625,In_889);
nor U2303 (N_2303,In_243,In_393);
and U2304 (N_2304,In_349,In_140);
and U2305 (N_2305,In_743,In_538);
xnor U2306 (N_2306,In_109,In_779);
nor U2307 (N_2307,In_886,In_697);
and U2308 (N_2308,In_970,In_217);
or U2309 (N_2309,In_116,In_776);
and U2310 (N_2310,In_850,In_85);
nor U2311 (N_2311,In_800,In_610);
nor U2312 (N_2312,In_562,In_64);
xnor U2313 (N_2313,In_150,In_491);
xnor U2314 (N_2314,In_387,In_171);
or U2315 (N_2315,In_552,In_446);
nand U2316 (N_2316,In_682,In_603);
or U2317 (N_2317,In_614,In_37);
nor U2318 (N_2318,In_885,In_307);
xor U2319 (N_2319,In_722,In_523);
and U2320 (N_2320,In_904,In_358);
xor U2321 (N_2321,In_908,In_450);
and U2322 (N_2322,In_893,In_443);
nor U2323 (N_2323,In_136,In_267);
nand U2324 (N_2324,In_421,In_305);
xnor U2325 (N_2325,In_314,In_490);
nand U2326 (N_2326,In_91,In_715);
and U2327 (N_2327,In_75,In_914);
nor U2328 (N_2328,In_976,In_23);
nor U2329 (N_2329,In_313,In_83);
nand U2330 (N_2330,In_929,In_207);
nand U2331 (N_2331,In_832,In_988);
and U2332 (N_2332,In_520,In_98);
nor U2333 (N_2333,In_451,In_300);
nand U2334 (N_2334,In_971,In_230);
nand U2335 (N_2335,In_345,In_517);
and U2336 (N_2336,In_89,In_754);
and U2337 (N_2337,In_20,In_162);
nor U2338 (N_2338,In_134,In_953);
xnor U2339 (N_2339,In_554,In_137);
and U2340 (N_2340,In_359,In_264);
nand U2341 (N_2341,In_175,In_487);
nand U2342 (N_2342,In_863,In_945);
or U2343 (N_2343,In_447,In_727);
nand U2344 (N_2344,In_225,In_266);
or U2345 (N_2345,In_681,In_671);
nand U2346 (N_2346,In_233,In_545);
and U2347 (N_2347,In_53,In_290);
and U2348 (N_2348,In_467,In_620);
and U2349 (N_2349,In_361,In_989);
nor U2350 (N_2350,In_121,In_115);
nor U2351 (N_2351,In_319,In_107);
and U2352 (N_2352,In_315,In_406);
nand U2353 (N_2353,In_264,In_20);
xnor U2354 (N_2354,In_69,In_184);
and U2355 (N_2355,In_933,In_205);
nand U2356 (N_2356,In_501,In_25);
and U2357 (N_2357,In_674,In_788);
xnor U2358 (N_2358,In_505,In_25);
nand U2359 (N_2359,In_331,In_938);
nand U2360 (N_2360,In_531,In_783);
and U2361 (N_2361,In_139,In_983);
nor U2362 (N_2362,In_258,In_744);
xor U2363 (N_2363,In_777,In_422);
nor U2364 (N_2364,In_694,In_956);
nor U2365 (N_2365,In_877,In_981);
nor U2366 (N_2366,In_343,In_118);
xnor U2367 (N_2367,In_971,In_672);
nand U2368 (N_2368,In_827,In_789);
nor U2369 (N_2369,In_631,In_591);
and U2370 (N_2370,In_241,In_290);
nor U2371 (N_2371,In_451,In_722);
and U2372 (N_2372,In_402,In_945);
or U2373 (N_2373,In_818,In_252);
and U2374 (N_2374,In_616,In_787);
nor U2375 (N_2375,In_289,In_8);
nor U2376 (N_2376,In_458,In_816);
nor U2377 (N_2377,In_902,In_71);
nor U2378 (N_2378,In_16,In_717);
nor U2379 (N_2379,In_592,In_52);
or U2380 (N_2380,In_693,In_875);
nor U2381 (N_2381,In_787,In_296);
or U2382 (N_2382,In_955,In_619);
and U2383 (N_2383,In_430,In_623);
nor U2384 (N_2384,In_368,In_360);
or U2385 (N_2385,In_720,In_419);
or U2386 (N_2386,In_78,In_445);
and U2387 (N_2387,In_192,In_844);
xnor U2388 (N_2388,In_724,In_362);
or U2389 (N_2389,In_490,In_183);
nand U2390 (N_2390,In_321,In_538);
or U2391 (N_2391,In_382,In_262);
or U2392 (N_2392,In_404,In_485);
and U2393 (N_2393,In_199,In_590);
or U2394 (N_2394,In_536,In_129);
nor U2395 (N_2395,In_568,In_468);
xnor U2396 (N_2396,In_682,In_413);
xor U2397 (N_2397,In_790,In_818);
and U2398 (N_2398,In_191,In_760);
nor U2399 (N_2399,In_94,In_870);
and U2400 (N_2400,In_993,In_50);
and U2401 (N_2401,In_903,In_77);
nand U2402 (N_2402,In_43,In_63);
nor U2403 (N_2403,In_220,In_21);
nand U2404 (N_2404,In_989,In_321);
or U2405 (N_2405,In_104,In_256);
nor U2406 (N_2406,In_987,In_123);
nor U2407 (N_2407,In_324,In_949);
nand U2408 (N_2408,In_807,In_81);
nor U2409 (N_2409,In_398,In_651);
nand U2410 (N_2410,In_95,In_913);
xnor U2411 (N_2411,In_553,In_749);
and U2412 (N_2412,In_402,In_583);
xnor U2413 (N_2413,In_15,In_432);
and U2414 (N_2414,In_87,In_510);
nor U2415 (N_2415,In_863,In_464);
xor U2416 (N_2416,In_498,In_708);
and U2417 (N_2417,In_3,In_166);
nor U2418 (N_2418,In_435,In_576);
and U2419 (N_2419,In_808,In_60);
nor U2420 (N_2420,In_452,In_670);
nor U2421 (N_2421,In_943,In_795);
nor U2422 (N_2422,In_79,In_934);
or U2423 (N_2423,In_925,In_148);
and U2424 (N_2424,In_596,In_118);
or U2425 (N_2425,In_446,In_895);
or U2426 (N_2426,In_604,In_386);
or U2427 (N_2427,In_951,In_796);
and U2428 (N_2428,In_23,In_718);
or U2429 (N_2429,In_961,In_555);
nand U2430 (N_2430,In_745,In_308);
and U2431 (N_2431,In_104,In_165);
and U2432 (N_2432,In_398,In_777);
nand U2433 (N_2433,In_438,In_493);
nor U2434 (N_2434,In_696,In_590);
nand U2435 (N_2435,In_698,In_176);
and U2436 (N_2436,In_756,In_981);
or U2437 (N_2437,In_853,In_537);
and U2438 (N_2438,In_192,In_149);
or U2439 (N_2439,In_154,In_240);
or U2440 (N_2440,In_550,In_625);
nand U2441 (N_2441,In_706,In_508);
nor U2442 (N_2442,In_567,In_320);
and U2443 (N_2443,In_724,In_620);
xnor U2444 (N_2444,In_928,In_684);
and U2445 (N_2445,In_975,In_21);
nor U2446 (N_2446,In_159,In_737);
or U2447 (N_2447,In_102,In_830);
nor U2448 (N_2448,In_497,In_662);
or U2449 (N_2449,In_741,In_423);
nor U2450 (N_2450,In_84,In_875);
nand U2451 (N_2451,In_649,In_578);
nand U2452 (N_2452,In_54,In_491);
nor U2453 (N_2453,In_117,In_707);
nand U2454 (N_2454,In_135,In_820);
or U2455 (N_2455,In_625,In_295);
nand U2456 (N_2456,In_608,In_958);
nand U2457 (N_2457,In_628,In_188);
and U2458 (N_2458,In_484,In_168);
nand U2459 (N_2459,In_939,In_875);
nand U2460 (N_2460,In_337,In_294);
or U2461 (N_2461,In_822,In_756);
or U2462 (N_2462,In_972,In_763);
or U2463 (N_2463,In_995,In_757);
or U2464 (N_2464,In_815,In_430);
and U2465 (N_2465,In_776,In_717);
nor U2466 (N_2466,In_490,In_614);
or U2467 (N_2467,In_661,In_513);
nand U2468 (N_2468,In_567,In_128);
nor U2469 (N_2469,In_202,In_485);
xnor U2470 (N_2470,In_425,In_392);
and U2471 (N_2471,In_126,In_948);
or U2472 (N_2472,In_529,In_466);
and U2473 (N_2473,In_533,In_992);
and U2474 (N_2474,In_955,In_307);
nand U2475 (N_2475,In_333,In_535);
or U2476 (N_2476,In_530,In_96);
nor U2477 (N_2477,In_677,In_757);
and U2478 (N_2478,In_712,In_439);
nand U2479 (N_2479,In_92,In_48);
nor U2480 (N_2480,In_602,In_439);
xor U2481 (N_2481,In_662,In_535);
nand U2482 (N_2482,In_251,In_509);
or U2483 (N_2483,In_274,In_242);
nor U2484 (N_2484,In_416,In_706);
nor U2485 (N_2485,In_699,In_867);
or U2486 (N_2486,In_298,In_823);
nand U2487 (N_2487,In_345,In_379);
xor U2488 (N_2488,In_202,In_148);
and U2489 (N_2489,In_311,In_275);
xor U2490 (N_2490,In_635,In_153);
and U2491 (N_2491,In_110,In_958);
and U2492 (N_2492,In_806,In_254);
nor U2493 (N_2493,In_874,In_795);
nor U2494 (N_2494,In_896,In_852);
and U2495 (N_2495,In_344,In_413);
or U2496 (N_2496,In_713,In_233);
or U2497 (N_2497,In_70,In_748);
nand U2498 (N_2498,In_617,In_479);
nand U2499 (N_2499,In_890,In_339);
nand U2500 (N_2500,N_3,N_91);
nand U2501 (N_2501,N_1954,N_1311);
or U2502 (N_2502,N_1785,N_2103);
nor U2503 (N_2503,N_1395,N_1449);
and U2504 (N_2504,N_1869,N_446);
nor U2505 (N_2505,N_2001,N_1400);
nor U2506 (N_2506,N_771,N_1905);
or U2507 (N_2507,N_974,N_424);
nand U2508 (N_2508,N_85,N_648);
xnor U2509 (N_2509,N_978,N_1857);
xor U2510 (N_2510,N_2336,N_975);
xnor U2511 (N_2511,N_2016,N_854);
nand U2512 (N_2512,N_62,N_514);
or U2513 (N_2513,N_2012,N_1994);
or U2514 (N_2514,N_1758,N_1223);
and U2515 (N_2515,N_1889,N_618);
or U2516 (N_2516,N_1258,N_905);
nor U2517 (N_2517,N_2000,N_1689);
and U2518 (N_2518,N_1038,N_574);
nor U2519 (N_2519,N_2047,N_311);
nand U2520 (N_2520,N_1229,N_1313);
nand U2521 (N_2521,N_960,N_100);
and U2522 (N_2522,N_2044,N_48);
and U2523 (N_2523,N_1517,N_1530);
or U2524 (N_2524,N_2295,N_2228);
nand U2525 (N_2525,N_1903,N_470);
nor U2526 (N_2526,N_1690,N_713);
xor U2527 (N_2527,N_669,N_1061);
nor U2528 (N_2528,N_1507,N_235);
nor U2529 (N_2529,N_1686,N_888);
nor U2530 (N_2530,N_177,N_855);
and U2531 (N_2531,N_1640,N_1763);
nand U2532 (N_2532,N_993,N_1430);
and U2533 (N_2533,N_682,N_1001);
or U2534 (N_2534,N_2102,N_1329);
and U2535 (N_2535,N_355,N_109);
nand U2536 (N_2536,N_461,N_112);
nand U2537 (N_2537,N_373,N_1124);
or U2538 (N_2538,N_1121,N_237);
and U2539 (N_2539,N_788,N_943);
xnor U2540 (N_2540,N_1823,N_687);
and U2541 (N_2541,N_2219,N_2490);
nor U2542 (N_2542,N_360,N_1221);
nor U2543 (N_2543,N_2128,N_1284);
nor U2544 (N_2544,N_1660,N_500);
nand U2545 (N_2545,N_1842,N_1594);
nor U2546 (N_2546,N_558,N_2360);
nand U2547 (N_2547,N_376,N_1318);
nand U2548 (N_2548,N_396,N_665);
nor U2549 (N_2549,N_738,N_2056);
nor U2550 (N_2550,N_583,N_1032);
nor U2551 (N_2551,N_220,N_1780);
nand U2552 (N_2552,N_904,N_371);
and U2553 (N_2553,N_1563,N_1157);
nor U2554 (N_2554,N_1973,N_908);
or U2555 (N_2555,N_1685,N_757);
xnor U2556 (N_2556,N_43,N_1183);
nand U2557 (N_2557,N_348,N_1465);
xnor U2558 (N_2558,N_1002,N_831);
nand U2559 (N_2559,N_404,N_1150);
xor U2560 (N_2560,N_1564,N_1567);
and U2561 (N_2561,N_924,N_268);
nor U2562 (N_2562,N_764,N_2062);
or U2563 (N_2563,N_929,N_2401);
and U2564 (N_2564,N_1845,N_245);
xnor U2565 (N_2565,N_1621,N_578);
and U2566 (N_2566,N_292,N_2278);
xor U2567 (N_2567,N_473,N_659);
nor U2568 (N_2568,N_796,N_1543);
or U2569 (N_2569,N_1969,N_2028);
or U2570 (N_2570,N_737,N_415);
nand U2571 (N_2571,N_466,N_1021);
or U2572 (N_2572,N_663,N_156);
or U2573 (N_2573,N_9,N_2216);
nor U2574 (N_2574,N_381,N_1541);
and U2575 (N_2575,N_2106,N_1631);
or U2576 (N_2576,N_1531,N_1244);
nand U2577 (N_2577,N_2158,N_2305);
nand U2578 (N_2578,N_107,N_1379);
nor U2579 (N_2579,N_2151,N_2112);
nor U2580 (N_2580,N_399,N_1585);
and U2581 (N_2581,N_793,N_1704);
nand U2582 (N_2582,N_2324,N_1017);
and U2583 (N_2583,N_1866,N_389);
or U2584 (N_2584,N_654,N_482);
nand U2585 (N_2585,N_2380,N_295);
and U2586 (N_2586,N_1321,N_1848);
nand U2587 (N_2587,N_1746,N_800);
nor U2588 (N_2588,N_1418,N_2017);
xor U2589 (N_2589,N_1119,N_834);
or U2590 (N_2590,N_159,N_170);
and U2591 (N_2591,N_288,N_693);
and U2592 (N_2592,N_1436,N_1282);
nand U2593 (N_2593,N_860,N_1941);
or U2594 (N_2594,N_1601,N_1495);
or U2595 (N_2595,N_2250,N_780);
nor U2596 (N_2596,N_762,N_1518);
xor U2597 (N_2597,N_1250,N_2002);
nand U2598 (N_2598,N_602,N_1225);
and U2599 (N_2599,N_24,N_1407);
or U2600 (N_2600,N_787,N_1374);
nand U2601 (N_2601,N_1359,N_178);
nand U2602 (N_2602,N_1478,N_306);
or U2603 (N_2603,N_1044,N_1814);
nand U2604 (N_2604,N_2217,N_1565);
and U2605 (N_2605,N_845,N_952);
nand U2606 (N_2606,N_572,N_329);
nor U2607 (N_2607,N_703,N_606);
or U2608 (N_2608,N_312,N_1298);
nand U2609 (N_2609,N_1700,N_2284);
and U2610 (N_2610,N_950,N_2111);
and U2611 (N_2611,N_2184,N_430);
nand U2612 (N_2612,N_1308,N_1280);
and U2613 (N_2613,N_129,N_2197);
or U2614 (N_2614,N_973,N_1514);
and U2615 (N_2615,N_1090,N_2456);
and U2616 (N_2616,N_681,N_401);
nand U2617 (N_2617,N_1634,N_2432);
nand U2618 (N_2618,N_621,N_1067);
and U2619 (N_2619,N_1656,N_941);
nand U2620 (N_2620,N_808,N_2472);
nor U2621 (N_2621,N_1492,N_105);
and U2622 (N_2622,N_42,N_1429);
and U2623 (N_2623,N_633,N_1205);
or U2624 (N_2624,N_2408,N_22);
and U2625 (N_2625,N_289,N_2413);
and U2626 (N_2626,N_885,N_1019);
nor U2627 (N_2627,N_1932,N_1421);
nor U2628 (N_2628,N_1187,N_586);
or U2629 (N_2629,N_164,N_365);
or U2630 (N_2630,N_1415,N_439);
and U2631 (N_2631,N_1115,N_2267);
and U2632 (N_2632,N_321,N_436);
nand U2633 (N_2633,N_632,N_1159);
or U2634 (N_2634,N_2188,N_990);
nand U2635 (N_2635,N_1336,N_1428);
or U2636 (N_2636,N_1508,N_2160);
nor U2637 (N_2637,N_2109,N_864);
and U2638 (N_2638,N_706,N_1772);
or U2639 (N_2639,N_95,N_607);
nand U2640 (N_2640,N_2174,N_464);
or U2641 (N_2641,N_479,N_1828);
nand U2642 (N_2642,N_2351,N_1123);
xor U2643 (N_2643,N_1341,N_1007);
nand U2644 (N_2644,N_1859,N_769);
and U2645 (N_2645,N_1087,N_2434);
nand U2646 (N_2646,N_1940,N_622);
or U2647 (N_2647,N_684,N_1697);
nand U2648 (N_2648,N_2343,N_387);
nor U2649 (N_2649,N_284,N_2390);
nand U2650 (N_2650,N_1650,N_2213);
or U2651 (N_2651,N_1511,N_1695);
and U2652 (N_2652,N_2076,N_1745);
nor U2653 (N_2653,N_1176,N_1060);
nor U2654 (N_2654,N_1461,N_71);
or U2655 (N_2655,N_58,N_1910);
or U2656 (N_2656,N_1880,N_1611);
nand U2657 (N_2657,N_2280,N_688);
or U2658 (N_2658,N_856,N_133);
or U2659 (N_2659,N_1748,N_1977);
nor U2660 (N_2660,N_2354,N_2320);
or U2661 (N_2661,N_379,N_502);
nor U2662 (N_2662,N_1575,N_729);
or U2663 (N_2663,N_2149,N_816);
nand U2664 (N_2664,N_1481,N_2207);
and U2665 (N_2665,N_417,N_1014);
nor U2666 (N_2666,N_1579,N_1292);
nand U2667 (N_2667,N_2078,N_1606);
and U2668 (N_2668,N_140,N_1155);
and U2669 (N_2669,N_799,N_677);
nor U2670 (N_2670,N_82,N_900);
nand U2671 (N_2671,N_314,N_1965);
nor U2672 (N_2672,N_1996,N_2362);
nand U2673 (N_2673,N_2210,N_413);
nor U2674 (N_2674,N_127,N_2033);
nor U2675 (N_2675,N_1295,N_539);
nand U2676 (N_2676,N_751,N_2127);
xor U2677 (N_2677,N_1818,N_165);
nand U2678 (N_2678,N_1271,N_1143);
xnor U2679 (N_2679,N_1358,N_1993);
nor U2680 (N_2680,N_1939,N_720);
nor U2681 (N_2681,N_748,N_471);
nor U2682 (N_2682,N_614,N_1571);
and U2683 (N_2683,N_2435,N_942);
and U2684 (N_2684,N_180,N_1058);
or U2685 (N_2685,N_2371,N_1004);
or U2686 (N_2686,N_1300,N_1312);
xnor U2687 (N_2687,N_2161,N_1424);
and U2688 (N_2688,N_1317,N_694);
and U2689 (N_2689,N_255,N_779);
or U2690 (N_2690,N_1749,N_2482);
nor U2691 (N_2691,N_2347,N_917);
or U2692 (N_2692,N_2148,N_2124);
or U2693 (N_2693,N_1082,N_1947);
nor U2694 (N_2694,N_867,N_625);
and U2695 (N_2695,N_216,N_655);
or U2696 (N_2696,N_316,N_512);
nor U2697 (N_2697,N_927,N_711);
and U2698 (N_2698,N_1608,N_610);
nor U2699 (N_2699,N_2259,N_1171);
xnor U2700 (N_2700,N_505,N_1139);
nor U2701 (N_2701,N_1375,N_1405);
nand U2702 (N_2702,N_397,N_1274);
nand U2703 (N_2703,N_1373,N_346);
nand U2704 (N_2704,N_1109,N_1735);
nand U2705 (N_2705,N_304,N_2166);
or U2706 (N_2706,N_2176,N_670);
and U2707 (N_2707,N_712,N_422);
xnor U2708 (N_2708,N_1990,N_901);
nand U2709 (N_2709,N_281,N_2282);
or U2710 (N_2710,N_1684,N_1979);
nor U2711 (N_2711,N_273,N_293);
xnor U2712 (N_2712,N_962,N_822);
nand U2713 (N_2713,N_996,N_650);
nand U2714 (N_2714,N_2476,N_1417);
nor U2715 (N_2715,N_752,N_675);
or U2716 (N_2716,N_1453,N_1211);
or U2717 (N_2717,N_274,N_1587);
xor U2718 (N_2718,N_278,N_2455);
nor U2719 (N_2719,N_1811,N_1085);
nor U2720 (N_2720,N_2052,N_1533);
or U2721 (N_2721,N_1288,N_238);
or U2722 (N_2722,N_1501,N_28);
and U2723 (N_2723,N_242,N_361);
or U2724 (N_2724,N_1141,N_2199);
or U2725 (N_2725,N_560,N_679);
nor U2726 (N_2726,N_233,N_549);
or U2727 (N_2727,N_1149,N_2234);
nor U2728 (N_2728,N_1265,N_1129);
nor U2729 (N_2729,N_398,N_297);
and U2730 (N_2730,N_438,N_1125);
or U2731 (N_2731,N_478,N_1668);
nand U2732 (N_2732,N_1948,N_2429);
or U2733 (N_2733,N_1978,N_1437);
nand U2734 (N_2734,N_7,N_102);
nand U2735 (N_2735,N_652,N_1907);
nor U2736 (N_2736,N_2157,N_637);
and U2737 (N_2737,N_857,N_1548);
or U2738 (N_2738,N_582,N_349);
or U2739 (N_2739,N_2359,N_948);
nand U2740 (N_2740,N_685,N_132);
nand U2741 (N_2741,N_1051,N_1204);
nand U2742 (N_2742,N_605,N_364);
nand U2743 (N_2743,N_1868,N_1664);
and U2744 (N_2744,N_511,N_411);
and U2745 (N_2745,N_267,N_761);
or U2746 (N_2746,N_967,N_148);
or U2747 (N_2747,N_2181,N_567);
nand U2748 (N_2748,N_897,N_2412);
or U2749 (N_2749,N_2192,N_1739);
and U2750 (N_2750,N_1703,N_1368);
nor U2751 (N_2751,N_280,N_2437);
nor U2752 (N_2752,N_2085,N_15);
or U2753 (N_2753,N_1266,N_118);
nand U2754 (N_2754,N_2431,N_1456);
or U2755 (N_2755,N_2236,N_214);
or U2756 (N_2756,N_353,N_1070);
xnor U2757 (N_2757,N_1706,N_1542);
and U2758 (N_2758,N_589,N_807);
nor U2759 (N_2759,N_671,N_2366);
and U2760 (N_2760,N_696,N_219);
nand U2761 (N_2761,N_963,N_1738);
and U2762 (N_2762,N_1655,N_997);
nand U2763 (N_2763,N_1184,N_2226);
nand U2764 (N_2764,N_468,N_254);
and U2765 (N_2765,N_1851,N_898);
or U2766 (N_2766,N_2154,N_664);
and U2767 (N_2767,N_1452,N_958);
or U2768 (N_2768,N_2196,N_344);
nor U2769 (N_2769,N_2008,N_1815);
and U2770 (N_2770,N_1853,N_1997);
nand U2771 (N_2771,N_172,N_1161);
nand U2772 (N_2772,N_1008,N_1263);
and U2773 (N_2773,N_2096,N_225);
or U2774 (N_2774,N_1186,N_395);
nor U2775 (N_2775,N_585,N_1247);
or U2776 (N_2776,N_809,N_2398);
nand U2777 (N_2777,N_667,N_1914);
and U2778 (N_2778,N_1830,N_1849);
xor U2779 (N_2779,N_619,N_440);
or U2780 (N_2780,N_535,N_1888);
and U2781 (N_2781,N_592,N_453);
and U2782 (N_2782,N_1722,N_1612);
and U2783 (N_2783,N_1307,N_676);
or U2784 (N_2784,N_2443,N_2302);
or U2785 (N_2785,N_609,N_2095);
and U2786 (N_2786,N_678,N_647);
nor U2787 (N_2787,N_561,N_634);
nor U2788 (N_2788,N_86,N_335);
and U2789 (N_2789,N_2406,N_881);
nand U2790 (N_2790,N_1647,N_1215);
and U2791 (N_2791,N_1470,N_200);
xor U2792 (N_2792,N_162,N_207);
nand U2793 (N_2793,N_1100,N_81);
and U2794 (N_2794,N_240,N_1576);
nor U2795 (N_2795,N_1281,N_2043);
or U2796 (N_2796,N_1991,N_1391);
or U2797 (N_2797,N_1596,N_735);
nor U2798 (N_2798,N_253,N_1434);
xor U2799 (N_2799,N_358,N_1714);
and U2800 (N_2800,N_2121,N_1515);
nor U2801 (N_2801,N_269,N_2377);
or U2802 (N_2802,N_340,N_1315);
nand U2803 (N_2803,N_756,N_1503);
nor U2804 (N_2804,N_137,N_1682);
nand U2805 (N_2805,N_1457,N_26);
nand U2806 (N_2806,N_1455,N_1393);
nor U2807 (N_2807,N_2481,N_1654);
nand U2808 (N_2808,N_1534,N_2457);
nor U2809 (N_2809,N_1097,N_155);
nor U2810 (N_2810,N_940,N_1408);
or U2811 (N_2811,N_698,N_244);
and U2812 (N_2812,N_1702,N_1108);
nand U2813 (N_2813,N_403,N_893);
nand U2814 (N_2814,N_965,N_914);
nand U2815 (N_2815,N_343,N_111);
or U2816 (N_2816,N_227,N_1724);
or U2817 (N_2817,N_2469,N_463);
nor U2818 (N_2818,N_188,N_2187);
nor U2819 (N_2819,N_1794,N_1102);
xnor U2820 (N_2820,N_1716,N_640);
or U2821 (N_2821,N_2290,N_1071);
nand U2822 (N_2822,N_772,N_460);
and U2823 (N_2823,N_717,N_1648);
and U2824 (N_2824,N_1080,N_931);
and U2825 (N_2825,N_122,N_1768);
nor U2826 (N_2826,N_103,N_2089);
and U2827 (N_2827,N_31,N_319);
nor U2828 (N_2828,N_2485,N_1766);
xor U2829 (N_2829,N_2271,N_1111);
nand U2830 (N_2830,N_425,N_1825);
or U2831 (N_2831,N_275,N_1251);
xor U2832 (N_2832,N_530,N_547);
or U2833 (N_2833,N_1767,N_230);
xor U2834 (N_2834,N_1504,N_1202);
nand U2835 (N_2835,N_84,N_2009);
and U2836 (N_2836,N_1052,N_489);
nand U2837 (N_2837,N_811,N_983);
nor U2838 (N_2838,N_2275,N_2376);
or U2839 (N_2839,N_1175,N_879);
and U2840 (N_2840,N_345,N_1091);
or U2841 (N_2841,N_2143,N_570);
xnor U2842 (N_2842,N_176,N_442);
nor U2843 (N_2843,N_972,N_2385);
nand U2844 (N_2844,N_1595,N_2306);
or U2845 (N_2845,N_884,N_1834);
nor U2846 (N_2846,N_926,N_141);
nand U2847 (N_2847,N_1839,N_1908);
and U2848 (N_2848,N_486,N_2316);
and U2849 (N_2849,N_458,N_1870);
and U2850 (N_2850,N_2365,N_2262);
nor U2851 (N_2851,N_1927,N_179);
nor U2852 (N_2852,N_2198,N_1591);
nand U2853 (N_2853,N_265,N_827);
nand U2854 (N_2854,N_2387,N_722);
nand U2855 (N_2855,N_596,N_2243);
and U2856 (N_2856,N_1566,N_2036);
xor U2857 (N_2857,N_1035,N_1444);
or U2858 (N_2858,N_638,N_1387);
nor U2859 (N_2859,N_2314,N_742);
and U2860 (N_2860,N_2086,N_2200);
xnor U2861 (N_2861,N_1832,N_862);
xnor U2862 (N_2862,N_217,N_870);
and U2863 (N_2863,N_2007,N_2222);
or U2864 (N_2864,N_2375,N_1633);
and U2865 (N_2865,N_2446,N_333);
nand U2866 (N_2866,N_1054,N_382);
and U2867 (N_2867,N_765,N_1305);
and U2868 (N_2868,N_1104,N_1289);
xor U2869 (N_2869,N_1382,N_98);
nand U2870 (N_2870,N_2214,N_1872);
or U2871 (N_2871,N_1077,N_153);
or U2872 (N_2872,N_2020,N_90);
and U2873 (N_2873,N_1414,N_192);
nor U2874 (N_2874,N_2242,N_1302);
nand U2875 (N_2875,N_185,N_1902);
or U2876 (N_2876,N_557,N_88);
and U2877 (N_2877,N_1602,N_515);
nor U2878 (N_2878,N_2318,N_823);
nand U2879 (N_2879,N_2268,N_2497);
nand U2880 (N_2880,N_690,N_970);
and U2881 (N_2881,N_0,N_1193);
or U2882 (N_2882,N_1380,N_104);
nand U2883 (N_2883,N_1063,N_1147);
nand U2884 (N_2884,N_1637,N_794);
and U2885 (N_2885,N_858,N_2323);
nand U2886 (N_2886,N_380,N_69);
or U2887 (N_2887,N_2063,N_2313);
nor U2888 (N_2888,N_1411,N_1933);
and U2889 (N_2889,N_2110,N_56);
nor U2890 (N_2890,N_418,N_1412);
xnor U2891 (N_2891,N_1360,N_2114);
nor U2892 (N_2892,N_2042,N_2321);
xor U2893 (N_2893,N_408,N_1256);
nor U2894 (N_2894,N_1526,N_2133);
nor U2895 (N_2895,N_1181,N_296);
nor U2896 (N_2896,N_736,N_951);
and U2897 (N_2897,N_2358,N_1747);
nor U2898 (N_2898,N_1086,N_1831);
nor U2899 (N_2899,N_1337,N_2066);
nor U2900 (N_2900,N_459,N_612);
or U2901 (N_2901,N_171,N_981);
and U2902 (N_2902,N_2247,N_2150);
or U2903 (N_2903,N_1756,N_1334);
and U2904 (N_2904,N_2051,N_1093);
nor U2905 (N_2905,N_469,N_1871);
or U2906 (N_2906,N_302,N_1043);
nand U2907 (N_2907,N_1460,N_39);
and U2908 (N_2908,N_328,N_394);
nor U2909 (N_2909,N_841,N_215);
xor U2910 (N_2910,N_64,N_1210);
and U2911 (N_2911,N_339,N_1917);
and U2912 (N_2912,N_1134,N_1527);
or U2913 (N_2913,N_2131,N_641);
or U2914 (N_2914,N_32,N_878);
xor U2915 (N_2915,N_1055,N_2445);
nor U2916 (N_2916,N_270,N_1169);
or U2917 (N_2917,N_1588,N_1369);
or U2918 (N_2918,N_1192,N_1667);
nand U2919 (N_2919,N_1764,N_1687);
nand U2920 (N_2920,N_542,N_427);
and U2921 (N_2921,N_1810,N_1034);
nor U2922 (N_2922,N_2010,N_492);
or U2923 (N_2923,N_1180,N_501);
nor U2924 (N_2924,N_384,N_2125);
nand U2925 (N_2925,N_20,N_301);
nor U2926 (N_2926,N_2378,N_1715);
and U2927 (N_2927,N_1774,N_1583);
nor U2928 (N_2928,N_2264,N_1665);
xor U2929 (N_2929,N_2239,N_1796);
nor U2930 (N_2930,N_54,N_1326);
xor U2931 (N_2931,N_2088,N_126);
nand U2932 (N_2932,N_1487,N_523);
xnor U2933 (N_2933,N_1370,N_1220);
nand U2934 (N_2934,N_2025,N_2240);
and U2935 (N_2935,N_1826,N_2183);
or U2936 (N_2936,N_475,N_1502);
nor U2937 (N_2937,N_571,N_1688);
or U2938 (N_2938,N_1846,N_1935);
xor U2939 (N_2939,N_147,N_462);
or U2940 (N_2940,N_2297,N_1419);
nand U2941 (N_2941,N_806,N_476);
and U2942 (N_2942,N_80,N_77);
or U2943 (N_2943,N_1628,N_1805);
nand U2944 (N_2944,N_1584,N_1658);
and U2945 (N_2945,N_65,N_1362);
and U2946 (N_2946,N_636,N_1867);
and U2947 (N_2947,N_2159,N_1620);
nor U2948 (N_2948,N_2209,N_323);
nor U2949 (N_2949,N_1381,N_1365);
and U2950 (N_2950,N_1781,N_1775);
nand U2951 (N_2951,N_1743,N_1555);
nand U2952 (N_2952,N_1203,N_27);
and U2953 (N_2953,N_101,N_2484);
nand U2954 (N_2954,N_957,N_2458);
or U2955 (N_2955,N_2251,N_2249);
nor U2956 (N_2956,N_932,N_55);
nand U2957 (N_2957,N_1904,N_35);
and U2958 (N_2958,N_218,N_844);
and U2959 (N_2959,N_1913,N_1962);
nand U2960 (N_2960,N_1331,N_852);
and U2961 (N_2961,N_1551,N_849);
and U2962 (N_2962,N_541,N_1041);
or U2963 (N_2963,N_1968,N_1011);
nor U2964 (N_2964,N_2163,N_290);
nand U2965 (N_2965,N_2393,N_828);
xnor U2966 (N_2966,N_142,N_1540);
or U2967 (N_2967,N_631,N_1301);
and U2968 (N_2968,N_1122,N_1653);
nor U2969 (N_2969,N_193,N_1286);
nor U2970 (N_2970,N_1674,N_2130);
or U2971 (N_2971,N_838,N_1338);
or U2972 (N_2972,N_1178,N_1046);
nor U2973 (N_2973,N_1581,N_2334);
nor U2974 (N_2974,N_843,N_493);
or U2975 (N_2975,N_1158,N_2263);
or U2976 (N_2976,N_1110,N_1844);
nor U2977 (N_2977,N_2330,N_2077);
and U2978 (N_2978,N_2361,N_2097);
or U2979 (N_2979,N_282,N_2064);
nand U2980 (N_2980,N_123,N_1999);
xnor U2981 (N_2981,N_93,N_1590);
nand U2982 (N_2982,N_1092,N_666);
xnor U2983 (N_2983,N_37,N_2221);
nand U2984 (N_2984,N_2193,N_947);
nand U2985 (N_2985,N_774,N_2231);
nand U2986 (N_2986,N_2005,N_2092);
nand U2987 (N_2987,N_1835,N_1522);
and U2988 (N_2988,N_710,N_1222);
and U2989 (N_2989,N_2289,N_2255);
or U2990 (N_2990,N_423,N_1445);
and U2991 (N_2991,N_1882,N_2105);
nor U2992 (N_2992,N_1652,N_1242);
and U2993 (N_2993,N_1883,N_1212);
and U2994 (N_2994,N_2203,N_1026);
nor U2995 (N_2995,N_1335,N_1603);
nand U2996 (N_2996,N_151,N_1829);
or U2997 (N_2997,N_789,N_1974);
nand U2998 (N_2998,N_47,N_1539);
or U2999 (N_2999,N_1279,N_1226);
nand U3000 (N_3000,N_2332,N_763);
and U3001 (N_3001,N_236,N_1864);
and U3002 (N_3002,N_1490,N_1493);
or U3003 (N_3003,N_672,N_1744);
xor U3004 (N_3004,N_555,N_1050);
and U3005 (N_3005,N_1448,N_1692);
xnor U3006 (N_3006,N_1995,N_2147);
nand U3007 (N_3007,N_930,N_548);
or U3008 (N_3008,N_998,N_994);
nand U3009 (N_3009,N_1779,N_1736);
or U3010 (N_3010,N_702,N_144);
nand U3011 (N_3011,N_601,N_2495);
or U3012 (N_3012,N_1909,N_414);
nor U3013 (N_3013,N_1466,N_726);
nor U3014 (N_3014,N_2450,N_851);
nor U3015 (N_3015,N_1390,N_1033);
nand U3016 (N_3016,N_2060,N_1693);
nand U3017 (N_3017,N_1151,N_1270);
or U3018 (N_3018,N_830,N_1167);
nor U3019 (N_3019,N_1484,N_2451);
nand U3020 (N_3020,N_1980,N_241);
nor U3021 (N_3021,N_1626,N_1246);
and U3022 (N_3022,N_1398,N_1394);
and U3023 (N_3023,N_1958,N_1750);
nand U3024 (N_3024,N_1770,N_1072);
or U3025 (N_3025,N_1728,N_1410);
or U3026 (N_3026,N_2177,N_2101);
and U3027 (N_3027,N_368,N_2244);
nor U3028 (N_3028,N_1521,N_1740);
nor U3029 (N_3029,N_1544,N_441);
nand U3030 (N_3030,N_456,N_2107);
nand U3031 (N_3031,N_2442,N_317);
or U3032 (N_3032,N_2357,N_2459);
nor U3033 (N_3033,N_1855,N_2462);
nand U3034 (N_3034,N_1788,N_758);
nor U3035 (N_3035,N_1000,N_431);
xor U3036 (N_3036,N_680,N_2340);
nand U3037 (N_3037,N_1837,N_1510);
or U3038 (N_3038,N_206,N_829);
or U3039 (N_3039,N_260,N_291);
xnor U3040 (N_3040,N_2003,N_2322);
or U3041 (N_3041,N_1079,N_161);
nor U3042 (N_3042,N_991,N_1152);
and U3043 (N_3043,N_2307,N_2254);
xor U3044 (N_3044,N_375,N_2232);
nand U3045 (N_3045,N_83,N_33);
nor U3046 (N_3046,N_277,N_2355);
nor U3047 (N_3047,N_322,N_921);
nor U3048 (N_3048,N_2394,N_2169);
xor U3049 (N_3049,N_1873,N_2396);
or U3050 (N_3050,N_11,N_125);
xnor U3051 (N_3051,N_1349,N_143);
nand U3052 (N_3052,N_2212,N_805);
or U3053 (N_3053,N_434,N_577);
nand U3054 (N_3054,N_2379,N_1801);
or U3055 (N_3055,N_2152,N_1918);
nand U3056 (N_3056,N_2488,N_1309);
nor U3057 (N_3057,N_797,N_2304);
nand U3058 (N_3058,N_1949,N_1045);
and U3059 (N_3059,N_134,N_923);
nor U3060 (N_3060,N_1627,N_94);
and U3061 (N_3061,N_1934,N_2329);
xor U3062 (N_3062,N_1480,N_1031);
or U3063 (N_3063,N_108,N_2137);
xnor U3064 (N_3064,N_1875,N_1887);
nor U3065 (N_3065,N_2015,N_795);
and U3066 (N_3066,N_1189,N_1707);
or U3067 (N_3067,N_964,N_1401);
nand U3068 (N_3068,N_259,N_2486);
and U3069 (N_3069,N_2333,N_533);
and U3070 (N_3070,N_692,N_1694);
nand U3071 (N_3071,N_727,N_1946);
xnor U3072 (N_3072,N_846,N_2027);
or U3073 (N_3073,N_2397,N_212);
and U3074 (N_3074,N_2168,N_629);
nand U3075 (N_3075,N_714,N_400);
nand U3076 (N_3076,N_725,N_980);
and U3077 (N_3077,N_2464,N_1821);
nor U3078 (N_3078,N_1921,N_1708);
and U3079 (N_3079,N_1732,N_2410);
or U3080 (N_3080,N_2024,N_877);
nor U3081 (N_3081,N_1196,N_697);
nand U3082 (N_3082,N_2053,N_2447);
or U3083 (N_3083,N_1224,N_956);
or U3084 (N_3084,N_810,N_2208);
or U3085 (N_3085,N_1885,N_1377);
or U3086 (N_3086,N_704,N_1617);
or U3087 (N_3087,N_1959,N_1190);
nand U3088 (N_3088,N_1012,N_1353);
nand U3089 (N_3089,N_517,N_859);
nand U3090 (N_3090,N_1886,N_581);
and U3091 (N_3091,N_1162,N_324);
or U3092 (N_3092,N_372,N_2248);
or U3093 (N_3093,N_1784,N_231);
or U3094 (N_3094,N_2019,N_1130);
nand U3095 (N_3095,N_2134,N_2489);
nand U3096 (N_3096,N_821,N_166);
or U3097 (N_3097,N_773,N_915);
xor U3098 (N_3098,N_889,N_1267);
nand U3099 (N_3099,N_250,N_1236);
nor U3100 (N_3100,N_283,N_2310);
nor U3101 (N_3101,N_1138,N_1881);
or U3102 (N_3102,N_1354,N_536);
nand U3103 (N_3103,N_2083,N_2480);
or U3104 (N_3104,N_1351,N_2145);
nor U3105 (N_3105,N_136,N_1389);
or U3106 (N_3106,N_745,N_2465);
nor U3107 (N_3107,N_540,N_1472);
or U3108 (N_3108,N_2073,N_521);
nand U3109 (N_3109,N_41,N_1876);
or U3110 (N_3110,N_1852,N_124);
nor U3111 (N_3111,N_2004,N_1643);
nand U3112 (N_3112,N_1915,N_429);
nand U3113 (N_3113,N_971,N_2068);
and U3114 (N_3114,N_485,N_1435);
and U3115 (N_3115,N_1485,N_92);
nor U3116 (N_3116,N_1489,N_2466);
and U3117 (N_3117,N_1614,N_1854);
and U3118 (N_3118,N_1062,N_2285);
or U3119 (N_3119,N_1113,N_472);
or U3120 (N_3120,N_2475,N_1464);
or U3121 (N_3121,N_2233,N_2238);
xnor U3122 (N_3122,N_565,N_2082);
xnor U3123 (N_3123,N_272,N_791);
nand U3124 (N_3124,N_1524,N_496);
and U3125 (N_3125,N_1005,N_1207);
and U3126 (N_3126,N_2468,N_1096);
and U3127 (N_3127,N_2090,N_2421);
xor U3128 (N_3128,N_695,N_1233);
xor U3129 (N_3129,N_228,N_167);
and U3130 (N_3130,N_986,N_853);
nand U3131 (N_3131,N_1642,N_1230);
or U3132 (N_3132,N_1433,N_370);
nor U3133 (N_3133,N_1535,N_2138);
and U3134 (N_3134,N_933,N_305);
or U3135 (N_3135,N_1597,N_2402);
and U3136 (N_3136,N_1078,N_604);
nor U3137 (N_3137,N_2294,N_2315);
nand U3138 (N_3138,N_2218,N_1164);
or U3139 (N_3139,N_1296,N_1850);
or U3140 (N_3140,N_25,N_2279);
nand U3141 (N_3141,N_562,N_1127);
and U3142 (N_3142,N_537,N_1593);
or U3143 (N_3143,N_875,N_263);
and U3144 (N_3144,N_1237,N_44);
nor U3145 (N_3145,N_1348,N_1833);
and U3146 (N_3146,N_17,N_1901);
or U3147 (N_3147,N_989,N_1355);
or U3148 (N_3148,N_691,N_1483);
and U3149 (N_3149,N_783,N_815);
and U3150 (N_3150,N_686,N_2287);
nor U3151 (N_3151,N_545,N_1425);
or U3152 (N_3152,N_1500,N_2140);
xnor U3153 (N_3153,N_1812,N_2414);
or U3154 (N_3154,N_2374,N_1672);
nand U3155 (N_3155,N_559,N_1496);
and U3156 (N_3156,N_320,N_1179);
or U3157 (N_3157,N_1559,N_739);
or U3158 (N_3158,N_2129,N_1094);
nand U3159 (N_3159,N_2352,N_222);
or U3160 (N_3160,N_546,N_1275);
and U3161 (N_3161,N_1926,N_1509);
nand U3162 (N_3162,N_210,N_833);
or U3163 (N_3163,N_2417,N_174);
or U3164 (N_3164,N_910,N_519);
and U3165 (N_3165,N_1976,N_733);
nand U3166 (N_3166,N_1762,N_405);
and U3167 (N_3167,N_920,N_1937);
and U3168 (N_3168,N_1499,N_2339);
xnor U3169 (N_3169,N_525,N_919);
nand U3170 (N_3170,N_45,N_936);
xor U3171 (N_3171,N_2449,N_1966);
nor U3172 (N_3172,N_868,N_117);
and U3173 (N_3173,N_630,N_2191);
and U3174 (N_3174,N_1804,N_508);
or U3175 (N_3175,N_1806,N_1101);
xor U3176 (N_3176,N_247,N_2026);
nor U3177 (N_3177,N_2049,N_871);
nor U3178 (N_3178,N_1659,N_1911);
nand U3179 (N_3179,N_2126,N_728);
nand U3180 (N_3180,N_649,N_1897);
or U3181 (N_3181,N_705,N_208);
nor U3182 (N_3182,N_911,N_310);
or U3183 (N_3183,N_2418,N_781);
and U3184 (N_3184,N_1984,N_116);
xnor U3185 (N_3185,N_2415,N_2453);
nor U3186 (N_3186,N_2054,N_550);
or U3187 (N_3187,N_2266,N_131);
and U3188 (N_3188,N_448,N_1609);
xor U3189 (N_3189,N_1952,N_2368);
and U3190 (N_3190,N_1793,N_2309);
and U3191 (N_3191,N_378,N_988);
or U3192 (N_3192,N_1105,N_1142);
nand U3193 (N_3193,N_1049,N_1053);
and U3194 (N_3194,N_2496,N_976);
or U3195 (N_3195,N_266,N_2006);
nand U3196 (N_3196,N_1771,N_1757);
nand U3197 (N_3197,N_1971,N_67);
xor U3198 (N_3198,N_366,N_1200);
and U3199 (N_3199,N_490,N_700);
nor U3200 (N_3200,N_1332,N_1396);
nand U3201 (N_3201,N_138,N_1622);
nor U3202 (N_3202,N_1022,N_1549);
nand U3203 (N_3203,N_68,N_568);
and U3204 (N_3204,N_205,N_1371);
and U3205 (N_3205,N_616,N_1476);
nor U3206 (N_3206,N_556,N_2498);
nor U3207 (N_3207,N_1231,N_2428);
or U3208 (N_3208,N_38,N_1325);
and U3209 (N_3209,N_1333,N_61);
nor U3210 (N_3210,N_286,N_1938);
or U3211 (N_3211,N_644,N_1303);
or U3212 (N_3212,N_257,N_985);
nor U3213 (N_3213,N_603,N_30);
nand U3214 (N_3214,N_2093,N_1208);
nor U3215 (N_3215,N_2331,N_2115);
xnor U3216 (N_3216,N_2031,N_928);
or U3217 (N_3217,N_1083,N_1255);
and U3218 (N_3218,N_1813,N_1213);
nand U3219 (N_3219,N_1386,N_110);
or U3220 (N_3220,N_1891,N_564);
and U3221 (N_3221,N_309,N_1107);
or U3222 (N_3222,N_1198,N_1894);
nand U3223 (N_3223,N_1592,N_279);
nand U3224 (N_3224,N_873,N_21);
or U3225 (N_3225,N_1450,N_175);
xnor U3226 (N_3226,N_1777,N_307);
or U3227 (N_3227,N_850,N_895);
or U3228 (N_3228,N_2035,N_2416);
nand U3229 (N_3229,N_1754,N_600);
or U3230 (N_3230,N_599,N_2389);
and U3231 (N_3231,N_992,N_2438);
nor U3232 (N_3232,N_552,N_1737);
nand U3233 (N_3233,N_465,N_674);
xnor U3234 (N_3234,N_454,N_2439);
nand U3235 (N_3235,N_1285,N_1725);
nor U3236 (N_3236,N_861,N_1018);
nand U3237 (N_3237,N_2225,N_451);
or U3238 (N_3238,N_198,N_1800);
or U3239 (N_3239,N_2272,N_1961);
nor U3240 (N_3240,N_1195,N_2312);
or U3241 (N_3241,N_1955,N_1136);
nand U3242 (N_3242,N_1103,N_2286);
nor U3243 (N_3243,N_2386,N_1709);
xor U3244 (N_3244,N_1214,N_1273);
nand U3245 (N_3245,N_1992,N_1761);
nor U3246 (N_3246,N_1020,N_2202);
nand U3247 (N_3247,N_836,N_1987);
or U3248 (N_3248,N_1858,N_551);
and U3249 (N_3249,N_1406,N_1028);
or U3250 (N_3250,N_1168,N_6);
or U3251 (N_3251,N_1137,N_1272);
nor U3252 (N_3252,N_2296,N_2229);
or U3253 (N_3253,N_352,N_457);
nor U3254 (N_3254,N_213,N_78);
and U3255 (N_3255,N_1657,N_1459);
or U3256 (N_3256,N_1118,N_318);
and U3257 (N_3257,N_907,N_1206);
nor U3258 (N_3258,N_2440,N_1194);
nor U3259 (N_3259,N_2023,N_1884);
nor U3260 (N_3260,N_1350,N_1420);
and U3261 (N_3261,N_1865,N_2261);
and U3262 (N_3262,N_2189,N_443);
or U3263 (N_3263,N_747,N_145);
and U3264 (N_3264,N_2132,N_643);
or U3265 (N_3265,N_2194,N_2349);
or U3266 (N_3266,N_2204,N_1191);
nand U3267 (N_3267,N_264,N_2317);
nor U3268 (N_3268,N_2460,N_1816);
nor U3269 (N_3269,N_1343,N_494);
and U3270 (N_3270,N_2098,N_1975);
and U3271 (N_3271,N_1441,N_2409);
and U3272 (N_3272,N_2483,N_2084);
nand U3273 (N_3273,N_1967,N_801);
nand U3274 (N_3274,N_128,N_2473);
or U3275 (N_3275,N_730,N_1890);
nand U3276 (N_3276,N_863,N_70);
nor U3277 (N_3277,N_1342,N_628);
and U3278 (N_3278,N_392,N_913);
nand U3279 (N_3279,N_369,N_1068);
nand U3280 (N_3280,N_657,N_719);
and U3281 (N_3281,N_518,N_2383);
and U3282 (N_3282,N_1919,N_1730);
xor U3283 (N_3283,N_1619,N_1177);
xnor U3284 (N_3284,N_969,N_906);
nor U3285 (N_3285,N_1545,N_918);
xor U3286 (N_3286,N_1426,N_966);
nand U3287 (N_3287,N_2190,N_1573);
nand U3288 (N_3288,N_1719,N_1943);
nand U3289 (N_3289,N_474,N_1027);
and U3290 (N_3290,N_10,N_946);
or U3291 (N_3291,N_491,N_481);
and U3292 (N_3292,N_14,N_635);
or U3293 (N_3293,N_554,N_1416);
and U3294 (N_3294,N_553,N_89);
nand U3295 (N_3295,N_1023,N_2117);
or U3296 (N_3296,N_755,N_2059);
and U3297 (N_3297,N_1742,N_412);
nor U3298 (N_3298,N_2433,N_1261);
nor U3299 (N_3299,N_1277,N_334);
or U3300 (N_3300,N_934,N_977);
and U3301 (N_3301,N_1625,N_590);
or U3302 (N_3302,N_114,N_203);
and U3303 (N_3303,N_734,N_1712);
nor U3304 (N_3304,N_778,N_1646);
and U3305 (N_3305,N_683,N_1451);
nand U3306 (N_3306,N_1446,N_2364);
nand U3307 (N_3307,N_1537,N_385);
nand U3308 (N_3308,N_1232,N_1799);
nor U3309 (N_3309,N_357,N_2032);
nand U3310 (N_3310,N_1755,N_1165);
and U3311 (N_3311,N_1892,N_1384);
nand U3312 (N_3312,N_1600,N_2441);
and U3313 (N_3313,N_1488,N_699);
nand U3314 (N_3314,N_2463,N_1661);
and U3315 (N_3315,N_2499,N_945);
and U3316 (N_3316,N_199,N_909);
nand U3317 (N_3317,N_731,N_416);
and U3318 (N_3318,N_49,N_189);
or U3319 (N_3319,N_2345,N_374);
nand U3320 (N_3320,N_1820,N_1432);
or U3321 (N_3321,N_1344,N_709);
nand U3322 (N_3322,N_2029,N_79);
nor U3323 (N_3323,N_1057,N_2420);
or U3324 (N_3324,N_1069,N_354);
or U3325 (N_3325,N_341,N_421);
nor U3326 (N_3326,N_1388,N_195);
or U3327 (N_3327,N_1615,N_1328);
and U3328 (N_3328,N_1638,N_1402);
or U3329 (N_3329,N_1951,N_1721);
and U3330 (N_3330,N_1928,N_1988);
or U3331 (N_3331,N_2372,N_1803);
and U3332 (N_3332,N_1582,N_2070);
nand U3333 (N_3333,N_209,N_315);
nand U3334 (N_3334,N_584,N_507);
nor U3335 (N_3335,N_1970,N_1632);
or U3336 (N_3336,N_2477,N_2100);
nor U3337 (N_3337,N_1316,N_1486);
nand U3338 (N_3338,N_1916,N_239);
and U3339 (N_3339,N_1676,N_2072);
and U3340 (N_3340,N_2094,N_1442);
nand U3341 (N_3341,N_313,N_1753);
or U3342 (N_3342,N_529,N_2099);
and U3343 (N_3343,N_2153,N_1982);
and U3344 (N_3344,N_782,N_534);
or U3345 (N_3345,N_1003,N_1572);
and U3346 (N_3346,N_723,N_2079);
or U3347 (N_3347,N_226,N_2356);
nor U3348 (N_3348,N_1607,N_76);
and U3349 (N_3349,N_721,N_46);
and U3350 (N_3350,N_120,N_1084);
and U3351 (N_3351,N_150,N_1324);
and U3352 (N_3352,N_2171,N_2311);
nand U3353 (N_3353,N_347,N_569);
xnor U3354 (N_3354,N_812,N_1729);
nor U3355 (N_3355,N_2452,N_820);
or U3356 (N_3356,N_880,N_617);
nor U3357 (N_3357,N_1216,N_2328);
nand U3358 (N_3358,N_1536,N_984);
nor U3359 (N_3359,N_2424,N_1929);
nand U3360 (N_3360,N_938,N_1473);
or U3361 (N_3361,N_1899,N_2426);
or U3362 (N_3362,N_350,N_1577);
and U3363 (N_3363,N_2392,N_211);
nand U3364 (N_3364,N_2206,N_1505);
and U3365 (N_3365,N_2388,N_1128);
xnor U3366 (N_3366,N_1320,N_767);
nor U3367 (N_3367,N_2113,N_2080);
nand U3368 (N_3368,N_1252,N_1731);
xnor U3369 (N_3369,N_527,N_194);
xnor U3370 (N_3370,N_949,N_1817);
xor U3371 (N_3371,N_819,N_1454);
nand U3372 (N_3372,N_1557,N_2201);
nor U3373 (N_3373,N_169,N_1025);
nand U3374 (N_3374,N_563,N_2081);
or U3375 (N_3375,N_1802,N_2303);
nand U3376 (N_3376,N_708,N_202);
or U3377 (N_3377,N_2430,N_503);
or U3378 (N_3378,N_444,N_367);
nor U3379 (N_3379,N_1713,N_1059);
xor U3380 (N_3380,N_1669,N_447);
or U3381 (N_3381,N_1269,N_326);
or U3382 (N_3382,N_1024,N_407);
nor U3383 (N_3383,N_1895,N_1680);
and U3384 (N_3384,N_2422,N_1808);
and U3385 (N_3385,N_509,N_1116);
and U3386 (N_3386,N_1691,N_477);
xor U3387 (N_3387,N_435,N_1720);
or U3388 (N_3388,N_1726,N_2419);
nor U3389 (N_3389,N_848,N_2014);
nor U3390 (N_3390,N_912,N_1791);
or U3391 (N_3391,N_876,N_701);
or U3392 (N_3392,N_256,N_2155);
and U3393 (N_3393,N_2467,N_1786);
and U3394 (N_3394,N_303,N_1030);
xnor U3395 (N_3395,N_1898,N_1241);
nand U3396 (N_3396,N_2346,N_2173);
xnor U3397 (N_3397,N_840,N_19);
nand U3398 (N_3398,N_2227,N_1048);
nor U3399 (N_3399,N_2353,N_2011);
nor U3400 (N_3400,N_1245,N_1874);
nor U3401 (N_3401,N_246,N_595);
or U3402 (N_3402,N_1945,N_1010);
nor U3403 (N_3403,N_1383,N_2348);
or U3404 (N_3404,N_1219,N_1639);
or U3405 (N_3405,N_1561,N_2436);
xor U3406 (N_3406,N_1843,N_1963);
and U3407 (N_3407,N_624,N_1291);
nor U3408 (N_3408,N_342,N_620);
nand U3409 (N_3409,N_598,N_299);
or U3410 (N_3410,N_2136,N_1462);
nor U3411 (N_3411,N_1532,N_363);
or U3412 (N_3412,N_2425,N_2382);
and U3413 (N_3413,N_869,N_2404);
or U3414 (N_3414,N_954,N_1227);
or U3415 (N_3415,N_1340,N_935);
and U3416 (N_3416,N_409,N_1399);
and U3417 (N_3417,N_1751,N_2492);
xnor U3418 (N_3418,N_660,N_2048);
xnor U3419 (N_3419,N_1173,N_2277);
or U3420 (N_3420,N_13,N_2120);
or U3421 (N_3421,N_432,N_1560);
and U3422 (N_3422,N_29,N_1930);
and U3423 (N_3423,N_1960,N_2108);
or U3424 (N_3424,N_1064,N_1586);
nand U3425 (N_3425,N_2224,N_1076);
nand U3426 (N_3426,N_1723,N_1956);
nor U3427 (N_3427,N_377,N_645);
nor U3428 (N_3428,N_770,N_8);
nand U3429 (N_3429,N_627,N_2162);
nand U3430 (N_3430,N_2400,N_1578);
nand U3431 (N_3431,N_2065,N_2230);
xnor U3432 (N_3432,N_959,N_2179);
nor U3433 (N_3433,N_1790,N_2075);
nand U3434 (N_3434,N_168,N_1782);
nand U3435 (N_3435,N_1427,N_1131);
or U3436 (N_3436,N_835,N_1797);
nand U3437 (N_3437,N_1185,N_1479);
and U3438 (N_3438,N_201,N_825);
and U3439 (N_3439,N_1931,N_847);
nand U3440 (N_3440,N_716,N_2061);
or U3441 (N_3441,N_445,N_1132);
and U3442 (N_3442,N_1009,N_1356);
or U3443 (N_3443,N_87,N_115);
and U3444 (N_3444,N_2,N_2369);
nand U3445 (N_3445,N_1896,N_594);
or U3446 (N_3446,N_1678,N_1322);
or U3447 (N_3447,N_1964,N_522);
nand U3448 (N_3448,N_1644,N_4);
and U3449 (N_3449,N_149,N_813);
nand U3450 (N_3450,N_99,N_2350);
xor U3451 (N_3451,N_146,N_1120);
nand U3452 (N_3452,N_646,N_73);
and U3453 (N_3453,N_2205,N_154);
and U3454 (N_3454,N_597,N_1188);
nand U3455 (N_3455,N_2270,N_2291);
nor U3456 (N_3456,N_651,N_759);
or U3457 (N_3457,N_1618,N_1361);
nand U3458 (N_3458,N_248,N_1081);
or U3459 (N_3459,N_1015,N_1314);
and U3460 (N_3460,N_75,N_1819);
or U3461 (N_3461,N_1297,N_2370);
nor U3462 (N_3462,N_1809,N_1569);
or U3463 (N_3463,N_1413,N_2327);
nor U3464 (N_3464,N_1243,N_2269);
xor U3465 (N_3465,N_1163,N_1604);
or U3466 (N_3466,N_261,N_1209);
nor U3467 (N_3467,N_1073,N_2427);
xnor U3468 (N_3468,N_2344,N_1822);
xor U3469 (N_3469,N_891,N_1795);
xnor U3470 (N_3470,N_642,N_2235);
nor U3471 (N_3471,N_2299,N_1013);
nor U3472 (N_3472,N_1662,N_187);
and U3473 (N_3473,N_1841,N_1174);
nand U3474 (N_3474,N_338,N_1364);
nor U3475 (N_3475,N_1506,N_513);
nand U3476 (N_3476,N_955,N_1431);
and U3477 (N_3477,N_784,N_573);
nor U3478 (N_3478,N_776,N_1438);
nand U3479 (N_3479,N_1519,N_662);
and U3480 (N_3480,N_426,N_1513);
and U3481 (N_3481,N_1346,N_1673);
and U3482 (N_3482,N_433,N_2067);
and U3483 (N_3483,N_1998,N_1112);
nand U3484 (N_3484,N_1469,N_135);
xnor U3485 (N_3485,N_882,N_1893);
nand U3486 (N_3486,N_243,N_1260);
nor U3487 (N_3487,N_325,N_2087);
or U3488 (N_3488,N_287,N_689);
nor U3489 (N_3489,N_899,N_995);
and U3490 (N_3490,N_1262,N_190);
nand U3491 (N_3491,N_818,N_184);
or U3492 (N_3492,N_1924,N_1906);
nand U3493 (N_3493,N_1006,N_152);
or U3494 (N_3494,N_1516,N_1240);
or U3495 (N_3495,N_768,N_1523);
nand U3496 (N_3496,N_1773,N_524);
and U3497 (N_3497,N_1789,N_1616);
or U3498 (N_3498,N_839,N_1630);
and U3499 (N_3499,N_97,N_386);
nand U3500 (N_3500,N_987,N_2491);
or U3501 (N_3501,N_1037,N_1319);
nor U3502 (N_3502,N_1985,N_2338);
xnor U3503 (N_3503,N_191,N_1016);
nand U3504 (N_3504,N_1144,N_2487);
and U3505 (N_3505,N_1259,N_2252);
nor U3506 (N_3506,N_232,N_1290);
and U3507 (N_3507,N_1404,N_12);
and U3508 (N_3508,N_1649,N_57);
nand U3509 (N_3509,N_1294,N_872);
nor U3510 (N_3510,N_1040,N_1681);
nor U3511 (N_3511,N_2265,N_276);
or U3512 (N_3512,N_2045,N_52);
and U3513 (N_3513,N_1683,N_1923);
and U3514 (N_3514,N_1953,N_1172);
or U3515 (N_3515,N_362,N_2246);
or U3516 (N_3516,N_181,N_1409);
xnor U3517 (N_3517,N_1423,N_1599);
nor U3518 (N_3518,N_1234,N_300);
and U3519 (N_3519,N_51,N_2104);
and U3520 (N_3520,N_1264,N_483);
nand U3521 (N_3521,N_1133,N_2381);
nor U3522 (N_3522,N_746,N_894);
or U3523 (N_3523,N_2164,N_1912);
nor U3524 (N_3524,N_2215,N_1525);
and U3525 (N_3525,N_1878,N_1352);
or U3526 (N_3526,N_1787,N_1114);
or U3527 (N_3527,N_2384,N_532);
nor U3528 (N_3528,N_1357,N_2185);
or U3529 (N_3529,N_1268,N_1166);
nor U3530 (N_3530,N_2123,N_163);
nand U3531 (N_3531,N_626,N_2258);
nand U3532 (N_3532,N_1863,N_1199);
xnor U3533 (N_3533,N_258,N_2411);
and U3534 (N_3534,N_495,N_224);
and U3535 (N_3535,N_1553,N_2395);
and U3536 (N_3536,N_1836,N_182);
xnor U3537 (N_3537,N_1718,N_890);
and U3538 (N_3538,N_2170,N_467);
nand U3539 (N_3539,N_824,N_2363);
nor U3540 (N_3540,N_2301,N_390);
nor U3541 (N_3541,N_2274,N_1847);
and U3542 (N_3542,N_2038,N_1666);
or U3543 (N_3543,N_802,N_18);
or U3544 (N_3544,N_1253,N_2405);
or U3545 (N_3545,N_16,N_1636);
and U3546 (N_3546,N_1463,N_249);
or U3547 (N_3547,N_1679,N_96);
and U3548 (N_3548,N_2135,N_121);
nand U3549 (N_3549,N_1546,N_50);
nor U3550 (N_3550,N_1705,N_1276);
nand U3551 (N_3551,N_2037,N_754);
or U3552 (N_3552,N_1972,N_204);
nand U3553 (N_3553,N_2142,N_1474);
or U3554 (N_3554,N_1042,N_1778);
and U3555 (N_3555,N_526,N_673);
nand U3556 (N_3556,N_866,N_1776);
nor U3557 (N_3557,N_1156,N_883);
nor U3558 (N_3558,N_661,N_2167);
or U3559 (N_3559,N_1944,N_1293);
nand U3560 (N_3560,N_450,N_798);
and U3561 (N_3561,N_2407,N_2139);
or U3562 (N_3562,N_750,N_615);
xor U3563 (N_3563,N_1623,N_2165);
nand U3564 (N_3564,N_1957,N_2319);
nor U3565 (N_3565,N_785,N_944);
or U3566 (N_3566,N_388,N_575);
or U3567 (N_3567,N_1089,N_1986);
nand U3568 (N_3568,N_2175,N_113);
nand U3569 (N_3569,N_865,N_1367);
nor U3570 (N_3570,N_1512,N_40);
nor U3571 (N_3571,N_1447,N_1477);
xor U3572 (N_3572,N_2373,N_903);
or U3573 (N_3573,N_1624,N_234);
or U3574 (N_3574,N_308,N_2257);
nor U3575 (N_3575,N_66,N_1827);
xor U3576 (N_3576,N_1363,N_1248);
nand U3577 (N_3577,N_1182,N_1306);
and U3578 (N_3578,N_623,N_1397);
or U3579 (N_3579,N_1556,N_2245);
and U3580 (N_3580,N_2118,N_1);
xnor U3581 (N_3581,N_1752,N_2057);
nand U3582 (N_3582,N_2342,N_999);
nand U3583 (N_3583,N_1099,N_2367);
and U3584 (N_3584,N_2276,N_766);
and U3585 (N_3585,N_2335,N_1547);
or U3586 (N_3586,N_1323,N_1378);
nor U3587 (N_3587,N_2069,N_1824);
or U3588 (N_3588,N_2186,N_939);
or U3589 (N_3589,N_1135,N_1862);
or U3590 (N_3590,N_1936,N_1698);
nand U3591 (N_3591,N_488,N_1140);
nor U3592 (N_3592,N_916,N_1498);
nor U3593 (N_3593,N_1088,N_1339);
xor U3594 (N_3594,N_1385,N_1562);
xnor U3595 (N_3595,N_327,N_351);
nand U3596 (N_3596,N_229,N_498);
nor U3597 (N_3597,N_1218,N_1580);
nand U3598 (N_3598,N_1925,N_2055);
nand U3599 (N_3599,N_2293,N_1983);
nand U3600 (N_3600,N_2058,N_516);
nor U3601 (N_3601,N_106,N_1475);
and U3602 (N_3602,N_1677,N_1651);
nor U3603 (N_3603,N_196,N_2013);
or U3604 (N_3604,N_886,N_1098);
or U3605 (N_3605,N_922,N_925);
or U3606 (N_3606,N_803,N_1574);
nand U3607 (N_3607,N_1497,N_2391);
or U3608 (N_3608,N_1491,N_2471);
nand U3609 (N_3609,N_1670,N_2292);
nand U3610 (N_3610,N_1458,N_1257);
nand U3611 (N_3611,N_953,N_1170);
and U3612 (N_3612,N_1235,N_1074);
nand U3613 (N_3613,N_504,N_1154);
and U3614 (N_3614,N_1699,N_593);
nor U3615 (N_3615,N_59,N_1900);
nand U3616 (N_3616,N_2308,N_74);
and U3617 (N_3617,N_1467,N_588);
or U3618 (N_3618,N_2146,N_1733);
nor U3619 (N_3619,N_2423,N_826);
and U3620 (N_3620,N_449,N_2474);
or U3621 (N_3621,N_1671,N_1552);
nand U3622 (N_3622,N_1613,N_544);
nor U3623 (N_3623,N_1372,N_63);
or U3624 (N_3624,N_2256,N_1570);
and U3625 (N_3625,N_2341,N_1403);
or U3626 (N_3626,N_1126,N_1310);
or U3627 (N_3627,N_937,N_1482);
xor U3628 (N_3628,N_1734,N_1065);
or U3629 (N_3629,N_2220,N_1529);
xnor U3630 (N_3630,N_543,N_1066);
nand U3631 (N_3631,N_510,N_968);
or U3632 (N_3632,N_804,N_391);
and U3633 (N_3633,N_452,N_832);
nor U3634 (N_3634,N_1117,N_1075);
nor U3635 (N_3635,N_1717,N_157);
nand U3636 (N_3636,N_2493,N_1920);
nor U3637 (N_3637,N_656,N_1922);
and U3638 (N_3638,N_1807,N_887);
and U3639 (N_3639,N_2040,N_2470);
or U3640 (N_3640,N_2260,N_1605);
and U3641 (N_3641,N_715,N_1520);
xnor U3642 (N_3642,N_1347,N_2074);
nand U3643 (N_3643,N_2461,N_580);
or U3644 (N_3644,N_2211,N_2180);
xnor U3645 (N_3645,N_892,N_1840);
nand U3646 (N_3646,N_1710,N_1422);
nor U3647 (N_3647,N_1727,N_743);
nor U3648 (N_3648,N_2119,N_1783);
xor U3649 (N_3649,N_2071,N_2454);
or U3650 (N_3650,N_528,N_2326);
and U3651 (N_3651,N_1330,N_2241);
or U3652 (N_3652,N_1981,N_591);
or U3653 (N_3653,N_2091,N_139);
xor U3654 (N_3654,N_1769,N_1238);
or U3655 (N_3655,N_740,N_5);
or U3656 (N_3656,N_896,N_1641);
nor U3657 (N_3657,N_566,N_786);
xnor U3658 (N_3658,N_1696,N_1760);
and U3659 (N_3659,N_579,N_1392);
or U3660 (N_3660,N_1197,N_428);
nand U3661 (N_3661,N_1145,N_2195);
nor U3662 (N_3662,N_639,N_53);
nand U3663 (N_3663,N_1217,N_1345);
and U3664 (N_3664,N_1039,N_1798);
xnor U3665 (N_3665,N_1598,N_1439);
nand U3666 (N_3666,N_744,N_480);
nor U3667 (N_3667,N_359,N_2399);
nand U3668 (N_3668,N_332,N_1471);
nor U3669 (N_3669,N_2298,N_197);
and U3670 (N_3670,N_837,N_1254);
nor U3671 (N_3671,N_2237,N_1879);
and U3672 (N_3672,N_2403,N_1239);
or U3673 (N_3673,N_2122,N_1568);
nor U3674 (N_3674,N_1759,N_1249);
nand U3675 (N_3675,N_760,N_2144);
xor U3676 (N_3676,N_2325,N_383);
nor U3677 (N_3677,N_1856,N_1538);
nand U3678 (N_3678,N_2034,N_2022);
xnor U3679 (N_3679,N_499,N_1029);
nand U3680 (N_3680,N_2182,N_1304);
or U3681 (N_3681,N_72,N_1146);
and U3682 (N_3682,N_753,N_1153);
xnor U3683 (N_3683,N_531,N_2448);
and U3684 (N_3684,N_1228,N_2288);
nand U3685 (N_3685,N_790,N_707);
nor U3686 (N_3686,N_356,N_576);
and U3687 (N_3687,N_34,N_252);
or U3688 (N_3688,N_60,N_2141);
or U3689 (N_3689,N_1663,N_1675);
nor U3690 (N_3690,N_1106,N_1201);
and U3691 (N_3691,N_2300,N_337);
and U3692 (N_3692,N_1494,N_1366);
nor U3693 (N_3693,N_1838,N_1942);
nor U3694 (N_3694,N_1860,N_1468);
nand U3695 (N_3695,N_1528,N_1148);
nand U3696 (N_3696,N_1741,N_874);
nor U3697 (N_3697,N_842,N_420);
nand U3698 (N_3698,N_221,N_2478);
and U3699 (N_3699,N_587,N_814);
and U3700 (N_3700,N_961,N_538);
or U3701 (N_3701,N_130,N_262);
or U3702 (N_3702,N_2253,N_2444);
nand U3703 (N_3703,N_2273,N_455);
xnor U3704 (N_3704,N_1589,N_653);
nand U3705 (N_3705,N_119,N_1989);
and U3706 (N_3706,N_2337,N_1440);
or U3707 (N_3707,N_1283,N_173);
nor U3708 (N_3708,N_724,N_298);
nor U3709 (N_3709,N_186,N_658);
nor U3710 (N_3710,N_23,N_2039);
nand U3711 (N_3711,N_1950,N_223);
nand U3712 (N_3712,N_741,N_1160);
or U3713 (N_3713,N_2116,N_668);
nand U3714 (N_3714,N_160,N_2283);
nor U3715 (N_3715,N_402,N_1635);
or U3716 (N_3716,N_2021,N_2281);
nand U3717 (N_3717,N_775,N_1877);
nand U3718 (N_3718,N_419,N_183);
and U3719 (N_3719,N_2223,N_718);
nor U3720 (N_3720,N_1550,N_613);
and U3721 (N_3721,N_2050,N_817);
nor U3722 (N_3722,N_2041,N_979);
nor U3723 (N_3723,N_1376,N_437);
nor U3724 (N_3724,N_1056,N_1278);
or U3725 (N_3725,N_1036,N_1645);
or U3726 (N_3726,N_2046,N_1095);
or U3727 (N_3727,N_336,N_251);
nand U3728 (N_3728,N_2172,N_294);
and U3729 (N_3729,N_520,N_732);
nand U3730 (N_3730,N_497,N_1765);
or U3731 (N_3731,N_1554,N_1861);
or U3732 (N_3732,N_1711,N_36);
and U3733 (N_3733,N_1610,N_2479);
nor U3734 (N_3734,N_608,N_1287);
nor U3735 (N_3735,N_792,N_1327);
or U3736 (N_3736,N_902,N_2018);
or U3737 (N_3737,N_285,N_1047);
or U3738 (N_3738,N_1629,N_1701);
and U3739 (N_3739,N_1443,N_1792);
or U3740 (N_3740,N_271,N_777);
nand U3741 (N_3741,N_158,N_2156);
and U3742 (N_3742,N_2494,N_1558);
nor U3743 (N_3743,N_982,N_749);
and U3744 (N_3744,N_410,N_331);
nor U3745 (N_3745,N_611,N_2030);
nand U3746 (N_3746,N_506,N_406);
and U3747 (N_3747,N_487,N_484);
nor U3748 (N_3748,N_330,N_393);
nor U3749 (N_3749,N_1299,N_2178);
xnor U3750 (N_3750,N_1505,N_1091);
and U3751 (N_3751,N_239,N_1384);
nand U3752 (N_3752,N_359,N_508);
and U3753 (N_3753,N_2021,N_444);
nand U3754 (N_3754,N_969,N_1810);
or U3755 (N_3755,N_95,N_510);
nand U3756 (N_3756,N_1625,N_2343);
nor U3757 (N_3757,N_1373,N_751);
xor U3758 (N_3758,N_1383,N_2273);
nor U3759 (N_3759,N_2372,N_641);
or U3760 (N_3760,N_2385,N_2052);
and U3761 (N_3761,N_834,N_1639);
xor U3762 (N_3762,N_1102,N_1660);
nand U3763 (N_3763,N_1703,N_139);
xnor U3764 (N_3764,N_1090,N_1397);
nand U3765 (N_3765,N_753,N_1776);
nand U3766 (N_3766,N_2215,N_299);
nand U3767 (N_3767,N_2249,N_1678);
or U3768 (N_3768,N_1683,N_2458);
and U3769 (N_3769,N_1141,N_1362);
and U3770 (N_3770,N_2428,N_722);
nor U3771 (N_3771,N_172,N_1440);
xor U3772 (N_3772,N_1807,N_861);
or U3773 (N_3773,N_328,N_1702);
nor U3774 (N_3774,N_2145,N_2415);
nand U3775 (N_3775,N_1528,N_1888);
and U3776 (N_3776,N_602,N_2459);
or U3777 (N_3777,N_1942,N_2310);
and U3778 (N_3778,N_97,N_1183);
nand U3779 (N_3779,N_76,N_1827);
nand U3780 (N_3780,N_149,N_302);
or U3781 (N_3781,N_2280,N_2345);
nand U3782 (N_3782,N_1446,N_1215);
nor U3783 (N_3783,N_77,N_1145);
and U3784 (N_3784,N_1599,N_576);
or U3785 (N_3785,N_2111,N_37);
nand U3786 (N_3786,N_1923,N_2379);
nor U3787 (N_3787,N_227,N_1831);
nor U3788 (N_3788,N_1304,N_701);
xor U3789 (N_3789,N_2130,N_2200);
or U3790 (N_3790,N_984,N_567);
nor U3791 (N_3791,N_1839,N_749);
or U3792 (N_3792,N_1235,N_1084);
or U3793 (N_3793,N_131,N_806);
nor U3794 (N_3794,N_427,N_2161);
and U3795 (N_3795,N_125,N_2253);
nand U3796 (N_3796,N_1850,N_447);
or U3797 (N_3797,N_1296,N_1833);
and U3798 (N_3798,N_2348,N_2009);
xnor U3799 (N_3799,N_1156,N_2211);
nor U3800 (N_3800,N_1620,N_1144);
and U3801 (N_3801,N_978,N_1348);
xnor U3802 (N_3802,N_860,N_2424);
nor U3803 (N_3803,N_633,N_875);
and U3804 (N_3804,N_2492,N_1643);
nand U3805 (N_3805,N_1730,N_2217);
nand U3806 (N_3806,N_4,N_1431);
nand U3807 (N_3807,N_2281,N_2166);
and U3808 (N_3808,N_1864,N_2318);
and U3809 (N_3809,N_1469,N_1108);
nor U3810 (N_3810,N_1924,N_971);
and U3811 (N_3811,N_978,N_1180);
or U3812 (N_3812,N_1050,N_988);
nand U3813 (N_3813,N_1571,N_937);
xnor U3814 (N_3814,N_1064,N_608);
or U3815 (N_3815,N_1761,N_1083);
xor U3816 (N_3816,N_1233,N_404);
or U3817 (N_3817,N_389,N_216);
xnor U3818 (N_3818,N_1081,N_661);
and U3819 (N_3819,N_439,N_2012);
nor U3820 (N_3820,N_1592,N_1139);
or U3821 (N_3821,N_1699,N_909);
nand U3822 (N_3822,N_971,N_1492);
or U3823 (N_3823,N_892,N_356);
or U3824 (N_3824,N_807,N_2160);
or U3825 (N_3825,N_323,N_1590);
or U3826 (N_3826,N_1654,N_1545);
nor U3827 (N_3827,N_789,N_2172);
nor U3828 (N_3828,N_2168,N_1610);
nand U3829 (N_3829,N_2436,N_608);
nand U3830 (N_3830,N_1588,N_2162);
and U3831 (N_3831,N_658,N_1100);
or U3832 (N_3832,N_1874,N_732);
or U3833 (N_3833,N_1225,N_881);
nor U3834 (N_3834,N_1573,N_219);
xnor U3835 (N_3835,N_2458,N_1957);
nand U3836 (N_3836,N_2355,N_2429);
nand U3837 (N_3837,N_1890,N_340);
xnor U3838 (N_3838,N_2351,N_2461);
nor U3839 (N_3839,N_1823,N_1193);
nand U3840 (N_3840,N_332,N_2168);
and U3841 (N_3841,N_2230,N_906);
or U3842 (N_3842,N_1647,N_1387);
nand U3843 (N_3843,N_1699,N_886);
nand U3844 (N_3844,N_1279,N_1089);
nor U3845 (N_3845,N_659,N_1502);
nor U3846 (N_3846,N_1054,N_1851);
or U3847 (N_3847,N_2322,N_1103);
or U3848 (N_3848,N_2210,N_208);
nor U3849 (N_3849,N_1328,N_1234);
nand U3850 (N_3850,N_500,N_63);
or U3851 (N_3851,N_489,N_1240);
nor U3852 (N_3852,N_2086,N_382);
and U3853 (N_3853,N_1960,N_428);
and U3854 (N_3854,N_1720,N_1053);
or U3855 (N_3855,N_104,N_2231);
nor U3856 (N_3856,N_208,N_1747);
and U3857 (N_3857,N_358,N_1149);
xnor U3858 (N_3858,N_1117,N_1132);
or U3859 (N_3859,N_73,N_2031);
nand U3860 (N_3860,N_286,N_452);
nand U3861 (N_3861,N_1494,N_654);
and U3862 (N_3862,N_1152,N_2261);
or U3863 (N_3863,N_2185,N_2493);
nand U3864 (N_3864,N_1502,N_2002);
xor U3865 (N_3865,N_763,N_162);
nand U3866 (N_3866,N_1089,N_932);
nor U3867 (N_3867,N_2337,N_1919);
or U3868 (N_3868,N_34,N_1068);
nor U3869 (N_3869,N_592,N_440);
nand U3870 (N_3870,N_1709,N_1864);
or U3871 (N_3871,N_82,N_1674);
and U3872 (N_3872,N_205,N_797);
nand U3873 (N_3873,N_2498,N_1153);
xnor U3874 (N_3874,N_2361,N_1412);
and U3875 (N_3875,N_442,N_1918);
or U3876 (N_3876,N_1044,N_2122);
and U3877 (N_3877,N_1355,N_1833);
nor U3878 (N_3878,N_138,N_1071);
nand U3879 (N_3879,N_662,N_1990);
or U3880 (N_3880,N_1609,N_1876);
nor U3881 (N_3881,N_1168,N_1121);
nor U3882 (N_3882,N_480,N_1947);
nand U3883 (N_3883,N_345,N_2140);
xor U3884 (N_3884,N_1931,N_1638);
or U3885 (N_3885,N_1714,N_430);
nor U3886 (N_3886,N_1281,N_1726);
or U3887 (N_3887,N_856,N_232);
nand U3888 (N_3888,N_2351,N_1477);
or U3889 (N_3889,N_1458,N_586);
and U3890 (N_3890,N_1118,N_976);
nand U3891 (N_3891,N_2087,N_834);
nor U3892 (N_3892,N_269,N_1484);
and U3893 (N_3893,N_576,N_1724);
and U3894 (N_3894,N_2415,N_2142);
nand U3895 (N_3895,N_1041,N_2277);
xnor U3896 (N_3896,N_1606,N_6);
and U3897 (N_3897,N_1785,N_2198);
nor U3898 (N_3898,N_742,N_346);
or U3899 (N_3899,N_140,N_911);
nor U3900 (N_3900,N_74,N_787);
nor U3901 (N_3901,N_1369,N_111);
and U3902 (N_3902,N_570,N_1055);
nand U3903 (N_3903,N_842,N_2232);
nor U3904 (N_3904,N_989,N_1346);
nand U3905 (N_3905,N_1226,N_1790);
nand U3906 (N_3906,N_540,N_1203);
nand U3907 (N_3907,N_1046,N_1963);
or U3908 (N_3908,N_503,N_1969);
nand U3909 (N_3909,N_2094,N_237);
or U3910 (N_3910,N_2325,N_2488);
nand U3911 (N_3911,N_1128,N_1628);
xnor U3912 (N_3912,N_2379,N_1031);
nand U3913 (N_3913,N_1033,N_542);
nor U3914 (N_3914,N_677,N_888);
and U3915 (N_3915,N_884,N_1473);
xnor U3916 (N_3916,N_2418,N_1115);
or U3917 (N_3917,N_1937,N_15);
or U3918 (N_3918,N_848,N_865);
nand U3919 (N_3919,N_836,N_1699);
or U3920 (N_3920,N_1684,N_245);
and U3921 (N_3921,N_334,N_677);
or U3922 (N_3922,N_305,N_1857);
nand U3923 (N_3923,N_1186,N_1432);
and U3924 (N_3924,N_296,N_1996);
xnor U3925 (N_3925,N_2399,N_1534);
and U3926 (N_3926,N_1713,N_2076);
and U3927 (N_3927,N_2414,N_1860);
nor U3928 (N_3928,N_101,N_44);
nand U3929 (N_3929,N_1905,N_704);
and U3930 (N_3930,N_851,N_1976);
nand U3931 (N_3931,N_2158,N_1716);
or U3932 (N_3932,N_2102,N_1992);
nand U3933 (N_3933,N_96,N_89);
or U3934 (N_3934,N_464,N_1778);
xor U3935 (N_3935,N_2174,N_2271);
nand U3936 (N_3936,N_1967,N_883);
and U3937 (N_3937,N_1588,N_2368);
nand U3938 (N_3938,N_21,N_712);
xor U3939 (N_3939,N_1695,N_694);
nand U3940 (N_3940,N_460,N_752);
nor U3941 (N_3941,N_27,N_1018);
or U3942 (N_3942,N_1523,N_2253);
nand U3943 (N_3943,N_1270,N_2145);
nor U3944 (N_3944,N_1440,N_1301);
nor U3945 (N_3945,N_1000,N_566);
nor U3946 (N_3946,N_647,N_513);
and U3947 (N_3947,N_950,N_1702);
and U3948 (N_3948,N_482,N_127);
nor U3949 (N_3949,N_1131,N_1339);
nand U3950 (N_3950,N_1470,N_1763);
nand U3951 (N_3951,N_2407,N_962);
nor U3952 (N_3952,N_1959,N_1021);
or U3953 (N_3953,N_993,N_1233);
or U3954 (N_3954,N_799,N_1692);
nor U3955 (N_3955,N_564,N_466);
nand U3956 (N_3956,N_1552,N_783);
and U3957 (N_3957,N_2210,N_1530);
nand U3958 (N_3958,N_1935,N_178);
nor U3959 (N_3959,N_690,N_567);
and U3960 (N_3960,N_1368,N_1743);
nand U3961 (N_3961,N_95,N_28);
or U3962 (N_3962,N_641,N_248);
xor U3963 (N_3963,N_12,N_840);
nand U3964 (N_3964,N_1940,N_2168);
nand U3965 (N_3965,N_396,N_271);
and U3966 (N_3966,N_1945,N_488);
or U3967 (N_3967,N_2096,N_1838);
nand U3968 (N_3968,N_2211,N_1489);
or U3969 (N_3969,N_2388,N_1093);
nor U3970 (N_3970,N_1813,N_971);
or U3971 (N_3971,N_1588,N_764);
or U3972 (N_3972,N_241,N_85);
and U3973 (N_3973,N_1470,N_1);
and U3974 (N_3974,N_1770,N_2456);
nor U3975 (N_3975,N_194,N_2322);
or U3976 (N_3976,N_2403,N_973);
and U3977 (N_3977,N_2291,N_1114);
nand U3978 (N_3978,N_2199,N_1854);
or U3979 (N_3979,N_1333,N_1140);
xnor U3980 (N_3980,N_1248,N_966);
and U3981 (N_3981,N_261,N_1012);
or U3982 (N_3982,N_1095,N_2437);
and U3983 (N_3983,N_1753,N_2272);
or U3984 (N_3984,N_768,N_1660);
and U3985 (N_3985,N_1528,N_523);
nand U3986 (N_3986,N_1247,N_1483);
nand U3987 (N_3987,N_202,N_423);
nand U3988 (N_3988,N_1188,N_203);
or U3989 (N_3989,N_249,N_1319);
xnor U3990 (N_3990,N_513,N_1604);
or U3991 (N_3991,N_1121,N_196);
or U3992 (N_3992,N_2238,N_2001);
nand U3993 (N_3993,N_929,N_608);
nand U3994 (N_3994,N_297,N_1943);
nand U3995 (N_3995,N_978,N_1231);
nand U3996 (N_3996,N_1545,N_1130);
or U3997 (N_3997,N_1066,N_2205);
or U3998 (N_3998,N_1607,N_183);
nor U3999 (N_3999,N_815,N_2280);
or U4000 (N_4000,N_1044,N_431);
nor U4001 (N_4001,N_629,N_1708);
nand U4002 (N_4002,N_2299,N_150);
and U4003 (N_4003,N_2066,N_1827);
or U4004 (N_4004,N_1701,N_1914);
and U4005 (N_4005,N_1244,N_803);
nand U4006 (N_4006,N_817,N_882);
and U4007 (N_4007,N_2184,N_2312);
and U4008 (N_4008,N_2382,N_1053);
and U4009 (N_4009,N_757,N_1941);
or U4010 (N_4010,N_1942,N_1300);
or U4011 (N_4011,N_2371,N_273);
nor U4012 (N_4012,N_687,N_27);
xnor U4013 (N_4013,N_410,N_1574);
nor U4014 (N_4014,N_804,N_1809);
nor U4015 (N_4015,N_578,N_1096);
and U4016 (N_4016,N_1105,N_409);
or U4017 (N_4017,N_1694,N_1783);
or U4018 (N_4018,N_1254,N_1773);
or U4019 (N_4019,N_1277,N_1024);
or U4020 (N_4020,N_211,N_1567);
nor U4021 (N_4021,N_899,N_1691);
nor U4022 (N_4022,N_997,N_2021);
or U4023 (N_4023,N_1868,N_1711);
or U4024 (N_4024,N_899,N_667);
nand U4025 (N_4025,N_1917,N_618);
or U4026 (N_4026,N_594,N_278);
xnor U4027 (N_4027,N_398,N_1182);
xor U4028 (N_4028,N_2183,N_1203);
and U4029 (N_4029,N_1322,N_2396);
or U4030 (N_4030,N_1690,N_1846);
xnor U4031 (N_4031,N_790,N_2057);
or U4032 (N_4032,N_1549,N_36);
nand U4033 (N_4033,N_724,N_1527);
nor U4034 (N_4034,N_2115,N_1936);
and U4035 (N_4035,N_2183,N_33);
and U4036 (N_4036,N_231,N_873);
xor U4037 (N_4037,N_2009,N_1419);
or U4038 (N_4038,N_528,N_2105);
nor U4039 (N_4039,N_1221,N_406);
and U4040 (N_4040,N_2160,N_1667);
or U4041 (N_4041,N_1784,N_351);
nand U4042 (N_4042,N_994,N_1045);
nor U4043 (N_4043,N_1382,N_1368);
nand U4044 (N_4044,N_2419,N_1394);
nor U4045 (N_4045,N_134,N_2089);
xor U4046 (N_4046,N_1299,N_906);
or U4047 (N_4047,N_1178,N_2094);
nand U4048 (N_4048,N_1678,N_1102);
nor U4049 (N_4049,N_310,N_1881);
nor U4050 (N_4050,N_1795,N_1867);
nand U4051 (N_4051,N_1706,N_145);
nor U4052 (N_4052,N_1058,N_1528);
or U4053 (N_4053,N_596,N_2071);
nand U4054 (N_4054,N_155,N_2307);
nor U4055 (N_4055,N_114,N_1934);
nand U4056 (N_4056,N_2260,N_2042);
nor U4057 (N_4057,N_481,N_1498);
nor U4058 (N_4058,N_134,N_1894);
nor U4059 (N_4059,N_1486,N_101);
and U4060 (N_4060,N_3,N_2272);
nor U4061 (N_4061,N_1167,N_1719);
or U4062 (N_4062,N_1418,N_611);
nor U4063 (N_4063,N_22,N_2026);
and U4064 (N_4064,N_2033,N_667);
nand U4065 (N_4065,N_1581,N_733);
nand U4066 (N_4066,N_1754,N_2130);
nor U4067 (N_4067,N_2084,N_883);
nor U4068 (N_4068,N_1902,N_538);
nand U4069 (N_4069,N_2498,N_1078);
and U4070 (N_4070,N_226,N_2068);
nand U4071 (N_4071,N_1175,N_458);
nor U4072 (N_4072,N_70,N_108);
xnor U4073 (N_4073,N_145,N_983);
and U4074 (N_4074,N_1108,N_2364);
nor U4075 (N_4075,N_1205,N_379);
and U4076 (N_4076,N_1970,N_506);
nor U4077 (N_4077,N_1976,N_568);
and U4078 (N_4078,N_1861,N_1742);
and U4079 (N_4079,N_1042,N_431);
and U4080 (N_4080,N_1021,N_420);
or U4081 (N_4081,N_469,N_1594);
and U4082 (N_4082,N_1665,N_483);
and U4083 (N_4083,N_2179,N_1864);
and U4084 (N_4084,N_1995,N_2031);
and U4085 (N_4085,N_183,N_1896);
nand U4086 (N_4086,N_361,N_1495);
nor U4087 (N_4087,N_1316,N_541);
nand U4088 (N_4088,N_397,N_1523);
nand U4089 (N_4089,N_2163,N_1092);
or U4090 (N_4090,N_1909,N_1141);
nor U4091 (N_4091,N_2348,N_1657);
or U4092 (N_4092,N_480,N_1210);
nor U4093 (N_4093,N_1205,N_1438);
or U4094 (N_4094,N_942,N_1178);
nand U4095 (N_4095,N_633,N_1566);
or U4096 (N_4096,N_1807,N_1137);
nand U4097 (N_4097,N_335,N_753);
and U4098 (N_4098,N_859,N_1617);
and U4099 (N_4099,N_2093,N_2277);
and U4100 (N_4100,N_1020,N_1041);
nand U4101 (N_4101,N_1894,N_2367);
or U4102 (N_4102,N_2281,N_2171);
nor U4103 (N_4103,N_1934,N_462);
nand U4104 (N_4104,N_1218,N_1093);
nor U4105 (N_4105,N_1229,N_1671);
nor U4106 (N_4106,N_890,N_1601);
or U4107 (N_4107,N_610,N_1448);
and U4108 (N_4108,N_2122,N_325);
nor U4109 (N_4109,N_1159,N_2007);
nand U4110 (N_4110,N_878,N_64);
nor U4111 (N_4111,N_47,N_2482);
nand U4112 (N_4112,N_801,N_158);
or U4113 (N_4113,N_1516,N_2116);
and U4114 (N_4114,N_267,N_1423);
nand U4115 (N_4115,N_1121,N_918);
and U4116 (N_4116,N_89,N_2275);
nor U4117 (N_4117,N_206,N_91);
and U4118 (N_4118,N_1281,N_1398);
nand U4119 (N_4119,N_483,N_1781);
nand U4120 (N_4120,N_1066,N_99);
nand U4121 (N_4121,N_785,N_495);
or U4122 (N_4122,N_2400,N_1141);
xor U4123 (N_4123,N_1377,N_856);
xor U4124 (N_4124,N_507,N_782);
nand U4125 (N_4125,N_2102,N_1725);
nand U4126 (N_4126,N_1969,N_719);
nor U4127 (N_4127,N_113,N_2015);
and U4128 (N_4128,N_748,N_1261);
and U4129 (N_4129,N_1029,N_104);
nor U4130 (N_4130,N_2122,N_738);
nand U4131 (N_4131,N_279,N_1771);
and U4132 (N_4132,N_1882,N_198);
nor U4133 (N_4133,N_1407,N_2350);
nand U4134 (N_4134,N_510,N_1746);
nor U4135 (N_4135,N_218,N_344);
and U4136 (N_4136,N_1693,N_565);
nor U4137 (N_4137,N_1477,N_369);
nand U4138 (N_4138,N_843,N_2216);
and U4139 (N_4139,N_1454,N_1513);
and U4140 (N_4140,N_522,N_2367);
or U4141 (N_4141,N_1626,N_2299);
nand U4142 (N_4142,N_1197,N_88);
and U4143 (N_4143,N_420,N_1510);
and U4144 (N_4144,N_107,N_220);
or U4145 (N_4145,N_1093,N_62);
and U4146 (N_4146,N_404,N_772);
or U4147 (N_4147,N_2049,N_796);
nor U4148 (N_4148,N_1742,N_1643);
or U4149 (N_4149,N_1610,N_1828);
and U4150 (N_4150,N_1920,N_2413);
or U4151 (N_4151,N_204,N_1306);
nor U4152 (N_4152,N_990,N_2297);
or U4153 (N_4153,N_2275,N_1434);
or U4154 (N_4154,N_797,N_590);
nand U4155 (N_4155,N_361,N_584);
nor U4156 (N_4156,N_224,N_871);
nand U4157 (N_4157,N_2174,N_876);
xnor U4158 (N_4158,N_591,N_2186);
and U4159 (N_4159,N_1523,N_2495);
nand U4160 (N_4160,N_615,N_1944);
and U4161 (N_4161,N_2120,N_488);
nor U4162 (N_4162,N_986,N_1975);
and U4163 (N_4163,N_300,N_591);
nor U4164 (N_4164,N_935,N_668);
or U4165 (N_4165,N_711,N_2462);
and U4166 (N_4166,N_1355,N_2236);
nand U4167 (N_4167,N_1044,N_439);
or U4168 (N_4168,N_2062,N_470);
nand U4169 (N_4169,N_1767,N_2477);
and U4170 (N_4170,N_781,N_1025);
or U4171 (N_4171,N_2245,N_1187);
nand U4172 (N_4172,N_1615,N_1849);
nand U4173 (N_4173,N_847,N_212);
or U4174 (N_4174,N_1888,N_970);
nand U4175 (N_4175,N_635,N_2358);
xor U4176 (N_4176,N_1496,N_1208);
nor U4177 (N_4177,N_2155,N_529);
nor U4178 (N_4178,N_2000,N_236);
and U4179 (N_4179,N_679,N_1535);
nand U4180 (N_4180,N_1007,N_1987);
and U4181 (N_4181,N_2324,N_1173);
or U4182 (N_4182,N_22,N_1837);
xnor U4183 (N_4183,N_2166,N_468);
xnor U4184 (N_4184,N_2173,N_367);
xnor U4185 (N_4185,N_1140,N_116);
and U4186 (N_4186,N_1931,N_948);
and U4187 (N_4187,N_1280,N_1628);
nand U4188 (N_4188,N_1057,N_1969);
nor U4189 (N_4189,N_2292,N_249);
and U4190 (N_4190,N_1770,N_1904);
or U4191 (N_4191,N_1263,N_1102);
and U4192 (N_4192,N_544,N_1479);
and U4193 (N_4193,N_1974,N_646);
and U4194 (N_4194,N_46,N_1041);
nor U4195 (N_4195,N_1324,N_1737);
nand U4196 (N_4196,N_629,N_1102);
and U4197 (N_4197,N_117,N_143);
nand U4198 (N_4198,N_2460,N_466);
and U4199 (N_4199,N_1601,N_874);
and U4200 (N_4200,N_2345,N_2489);
and U4201 (N_4201,N_1660,N_2470);
nand U4202 (N_4202,N_1338,N_1380);
nor U4203 (N_4203,N_1835,N_2242);
and U4204 (N_4204,N_1306,N_1508);
xnor U4205 (N_4205,N_136,N_2084);
or U4206 (N_4206,N_452,N_2053);
or U4207 (N_4207,N_2252,N_138);
and U4208 (N_4208,N_895,N_2221);
or U4209 (N_4209,N_500,N_1950);
nor U4210 (N_4210,N_1359,N_680);
nand U4211 (N_4211,N_1202,N_1854);
nand U4212 (N_4212,N_412,N_1312);
or U4213 (N_4213,N_178,N_2309);
and U4214 (N_4214,N_1653,N_430);
nand U4215 (N_4215,N_296,N_2119);
nor U4216 (N_4216,N_291,N_2216);
and U4217 (N_4217,N_807,N_816);
nand U4218 (N_4218,N_1219,N_641);
or U4219 (N_4219,N_657,N_1977);
nor U4220 (N_4220,N_1810,N_1556);
nand U4221 (N_4221,N_2463,N_1318);
nand U4222 (N_4222,N_2340,N_1408);
nand U4223 (N_4223,N_1264,N_349);
and U4224 (N_4224,N_1570,N_1397);
nor U4225 (N_4225,N_991,N_1747);
or U4226 (N_4226,N_157,N_1674);
or U4227 (N_4227,N_2480,N_117);
or U4228 (N_4228,N_35,N_1937);
and U4229 (N_4229,N_550,N_2458);
and U4230 (N_4230,N_171,N_32);
nand U4231 (N_4231,N_1244,N_1663);
nor U4232 (N_4232,N_999,N_499);
nor U4233 (N_4233,N_810,N_566);
or U4234 (N_4234,N_31,N_1826);
and U4235 (N_4235,N_886,N_2337);
nand U4236 (N_4236,N_2015,N_1332);
or U4237 (N_4237,N_387,N_637);
nand U4238 (N_4238,N_831,N_2272);
or U4239 (N_4239,N_682,N_1546);
nor U4240 (N_4240,N_1373,N_86);
nor U4241 (N_4241,N_1360,N_31);
or U4242 (N_4242,N_313,N_928);
or U4243 (N_4243,N_996,N_623);
or U4244 (N_4244,N_1449,N_541);
or U4245 (N_4245,N_2395,N_115);
nor U4246 (N_4246,N_2335,N_2316);
nor U4247 (N_4247,N_2211,N_327);
or U4248 (N_4248,N_1416,N_656);
and U4249 (N_4249,N_1634,N_517);
nand U4250 (N_4250,N_1715,N_1064);
nand U4251 (N_4251,N_232,N_1024);
nand U4252 (N_4252,N_540,N_1785);
xor U4253 (N_4253,N_935,N_1028);
or U4254 (N_4254,N_485,N_992);
nand U4255 (N_4255,N_418,N_658);
nand U4256 (N_4256,N_707,N_1313);
or U4257 (N_4257,N_1668,N_28);
and U4258 (N_4258,N_696,N_1035);
or U4259 (N_4259,N_2430,N_1572);
nand U4260 (N_4260,N_346,N_448);
nand U4261 (N_4261,N_1009,N_1878);
nand U4262 (N_4262,N_1895,N_1174);
or U4263 (N_4263,N_534,N_1922);
or U4264 (N_4264,N_2218,N_1785);
and U4265 (N_4265,N_906,N_879);
nand U4266 (N_4266,N_153,N_946);
or U4267 (N_4267,N_1481,N_1222);
nor U4268 (N_4268,N_1748,N_1345);
nor U4269 (N_4269,N_1221,N_1623);
nand U4270 (N_4270,N_755,N_2431);
or U4271 (N_4271,N_1056,N_2145);
nand U4272 (N_4272,N_158,N_395);
and U4273 (N_4273,N_415,N_2412);
nor U4274 (N_4274,N_1528,N_1893);
xor U4275 (N_4275,N_853,N_2259);
nor U4276 (N_4276,N_2343,N_881);
or U4277 (N_4277,N_1360,N_1329);
or U4278 (N_4278,N_1221,N_660);
xnor U4279 (N_4279,N_141,N_47);
and U4280 (N_4280,N_1507,N_1383);
and U4281 (N_4281,N_2375,N_1565);
and U4282 (N_4282,N_952,N_1405);
or U4283 (N_4283,N_1957,N_511);
xnor U4284 (N_4284,N_1184,N_1236);
or U4285 (N_4285,N_2462,N_1476);
nand U4286 (N_4286,N_2088,N_1785);
or U4287 (N_4287,N_736,N_1394);
or U4288 (N_4288,N_1743,N_1038);
and U4289 (N_4289,N_2084,N_1380);
and U4290 (N_4290,N_1731,N_1638);
and U4291 (N_4291,N_123,N_2310);
nor U4292 (N_4292,N_1278,N_2475);
nand U4293 (N_4293,N_2396,N_1213);
xnor U4294 (N_4294,N_1518,N_639);
nor U4295 (N_4295,N_493,N_1591);
nand U4296 (N_4296,N_546,N_898);
and U4297 (N_4297,N_1234,N_1531);
or U4298 (N_4298,N_593,N_898);
xnor U4299 (N_4299,N_2136,N_1063);
or U4300 (N_4300,N_861,N_1853);
xnor U4301 (N_4301,N_467,N_732);
and U4302 (N_4302,N_2230,N_2330);
and U4303 (N_4303,N_1586,N_150);
nor U4304 (N_4304,N_26,N_1522);
nand U4305 (N_4305,N_1729,N_1837);
xnor U4306 (N_4306,N_390,N_733);
nor U4307 (N_4307,N_394,N_1555);
and U4308 (N_4308,N_1616,N_2340);
nor U4309 (N_4309,N_1706,N_2055);
and U4310 (N_4310,N_344,N_2337);
or U4311 (N_4311,N_58,N_1519);
and U4312 (N_4312,N_184,N_2156);
nand U4313 (N_4313,N_1411,N_927);
and U4314 (N_4314,N_1761,N_383);
or U4315 (N_4315,N_1651,N_2225);
nor U4316 (N_4316,N_1272,N_1362);
nor U4317 (N_4317,N_50,N_1517);
xor U4318 (N_4318,N_439,N_2031);
nor U4319 (N_4319,N_821,N_1958);
nor U4320 (N_4320,N_62,N_1863);
xnor U4321 (N_4321,N_1151,N_1354);
and U4322 (N_4322,N_13,N_1387);
or U4323 (N_4323,N_2229,N_209);
nand U4324 (N_4324,N_2145,N_2469);
or U4325 (N_4325,N_623,N_496);
xnor U4326 (N_4326,N_381,N_1212);
nor U4327 (N_4327,N_1996,N_1351);
and U4328 (N_4328,N_2268,N_370);
xnor U4329 (N_4329,N_908,N_12);
and U4330 (N_4330,N_1155,N_1460);
nor U4331 (N_4331,N_1996,N_955);
or U4332 (N_4332,N_1282,N_1413);
nand U4333 (N_4333,N_983,N_2020);
xnor U4334 (N_4334,N_1091,N_1301);
nor U4335 (N_4335,N_2485,N_2446);
nand U4336 (N_4336,N_11,N_2220);
or U4337 (N_4337,N_891,N_2239);
xor U4338 (N_4338,N_18,N_2111);
and U4339 (N_4339,N_2110,N_76);
nor U4340 (N_4340,N_686,N_268);
or U4341 (N_4341,N_1475,N_2246);
and U4342 (N_4342,N_115,N_1536);
nand U4343 (N_4343,N_460,N_1445);
and U4344 (N_4344,N_1090,N_1389);
and U4345 (N_4345,N_118,N_2113);
nand U4346 (N_4346,N_329,N_540);
or U4347 (N_4347,N_1146,N_640);
or U4348 (N_4348,N_2032,N_972);
nand U4349 (N_4349,N_638,N_2415);
nand U4350 (N_4350,N_2369,N_994);
nand U4351 (N_4351,N_474,N_101);
or U4352 (N_4352,N_974,N_656);
nor U4353 (N_4353,N_1279,N_407);
or U4354 (N_4354,N_1493,N_1688);
or U4355 (N_4355,N_1294,N_788);
and U4356 (N_4356,N_574,N_1167);
nand U4357 (N_4357,N_1546,N_2453);
nor U4358 (N_4358,N_1219,N_685);
and U4359 (N_4359,N_1041,N_75);
or U4360 (N_4360,N_229,N_602);
nor U4361 (N_4361,N_2144,N_1329);
or U4362 (N_4362,N_14,N_297);
nand U4363 (N_4363,N_1606,N_513);
nor U4364 (N_4364,N_918,N_752);
nand U4365 (N_4365,N_1448,N_1450);
or U4366 (N_4366,N_557,N_1470);
and U4367 (N_4367,N_1592,N_310);
nor U4368 (N_4368,N_875,N_652);
and U4369 (N_4369,N_2150,N_566);
xnor U4370 (N_4370,N_1058,N_2172);
and U4371 (N_4371,N_1440,N_1860);
and U4372 (N_4372,N_514,N_277);
nor U4373 (N_4373,N_2492,N_1665);
and U4374 (N_4374,N_303,N_836);
nor U4375 (N_4375,N_1556,N_1677);
nor U4376 (N_4376,N_985,N_886);
nand U4377 (N_4377,N_2407,N_2343);
xnor U4378 (N_4378,N_1064,N_521);
nor U4379 (N_4379,N_2252,N_2025);
nor U4380 (N_4380,N_1494,N_37);
nand U4381 (N_4381,N_1554,N_1266);
nor U4382 (N_4382,N_1578,N_2101);
and U4383 (N_4383,N_780,N_2260);
xor U4384 (N_4384,N_1406,N_1799);
nand U4385 (N_4385,N_362,N_1926);
or U4386 (N_4386,N_2105,N_1875);
or U4387 (N_4387,N_116,N_847);
xor U4388 (N_4388,N_2001,N_2054);
and U4389 (N_4389,N_2316,N_771);
or U4390 (N_4390,N_1034,N_1414);
and U4391 (N_4391,N_352,N_1011);
or U4392 (N_4392,N_749,N_1725);
or U4393 (N_4393,N_626,N_1242);
nand U4394 (N_4394,N_20,N_545);
and U4395 (N_4395,N_1017,N_1780);
xnor U4396 (N_4396,N_1481,N_1153);
nor U4397 (N_4397,N_387,N_2336);
nand U4398 (N_4398,N_1808,N_1996);
or U4399 (N_4399,N_1879,N_608);
and U4400 (N_4400,N_1060,N_2463);
or U4401 (N_4401,N_71,N_2029);
or U4402 (N_4402,N_2365,N_643);
or U4403 (N_4403,N_1049,N_2387);
or U4404 (N_4404,N_1371,N_796);
nand U4405 (N_4405,N_32,N_192);
and U4406 (N_4406,N_610,N_1562);
and U4407 (N_4407,N_1590,N_189);
nor U4408 (N_4408,N_1885,N_614);
nand U4409 (N_4409,N_961,N_798);
and U4410 (N_4410,N_2032,N_255);
xnor U4411 (N_4411,N_2203,N_1974);
and U4412 (N_4412,N_2020,N_448);
xor U4413 (N_4413,N_1007,N_2494);
nand U4414 (N_4414,N_327,N_1476);
xor U4415 (N_4415,N_276,N_591);
nand U4416 (N_4416,N_1958,N_1333);
nor U4417 (N_4417,N_1364,N_370);
or U4418 (N_4418,N_1767,N_848);
nand U4419 (N_4419,N_720,N_1813);
and U4420 (N_4420,N_981,N_1686);
or U4421 (N_4421,N_2429,N_1628);
xor U4422 (N_4422,N_1745,N_1451);
and U4423 (N_4423,N_655,N_960);
nor U4424 (N_4424,N_420,N_2056);
and U4425 (N_4425,N_2316,N_1156);
nand U4426 (N_4426,N_936,N_1947);
nand U4427 (N_4427,N_38,N_1);
or U4428 (N_4428,N_1380,N_1130);
xnor U4429 (N_4429,N_299,N_1942);
or U4430 (N_4430,N_1793,N_1464);
and U4431 (N_4431,N_1503,N_291);
or U4432 (N_4432,N_2397,N_967);
and U4433 (N_4433,N_2069,N_229);
nand U4434 (N_4434,N_150,N_240);
xor U4435 (N_4435,N_1508,N_2385);
and U4436 (N_4436,N_2160,N_1048);
nand U4437 (N_4437,N_1614,N_667);
xor U4438 (N_4438,N_1650,N_1533);
or U4439 (N_4439,N_2331,N_949);
nand U4440 (N_4440,N_1623,N_164);
nand U4441 (N_4441,N_1759,N_1933);
nand U4442 (N_4442,N_556,N_1991);
nor U4443 (N_4443,N_817,N_1113);
and U4444 (N_4444,N_771,N_159);
or U4445 (N_4445,N_1633,N_1605);
nand U4446 (N_4446,N_2496,N_2275);
and U4447 (N_4447,N_2475,N_708);
or U4448 (N_4448,N_1946,N_1218);
and U4449 (N_4449,N_451,N_949);
or U4450 (N_4450,N_564,N_1958);
xor U4451 (N_4451,N_1219,N_1733);
nor U4452 (N_4452,N_209,N_698);
nor U4453 (N_4453,N_1939,N_1026);
and U4454 (N_4454,N_1334,N_1409);
and U4455 (N_4455,N_2401,N_1774);
nand U4456 (N_4456,N_1218,N_2357);
and U4457 (N_4457,N_1646,N_245);
nand U4458 (N_4458,N_271,N_2294);
nand U4459 (N_4459,N_223,N_151);
nand U4460 (N_4460,N_1222,N_667);
nand U4461 (N_4461,N_276,N_1950);
nor U4462 (N_4462,N_1942,N_286);
nor U4463 (N_4463,N_1742,N_2190);
and U4464 (N_4464,N_2492,N_704);
and U4465 (N_4465,N_782,N_1209);
and U4466 (N_4466,N_212,N_2216);
nor U4467 (N_4467,N_1389,N_1483);
and U4468 (N_4468,N_1209,N_2468);
or U4469 (N_4469,N_558,N_1383);
nand U4470 (N_4470,N_1204,N_955);
and U4471 (N_4471,N_1244,N_710);
or U4472 (N_4472,N_418,N_1506);
nor U4473 (N_4473,N_47,N_1802);
nor U4474 (N_4474,N_105,N_2310);
or U4475 (N_4475,N_53,N_2146);
or U4476 (N_4476,N_1073,N_1094);
nand U4477 (N_4477,N_1665,N_2406);
nand U4478 (N_4478,N_347,N_1218);
and U4479 (N_4479,N_1298,N_1703);
nor U4480 (N_4480,N_627,N_1556);
nor U4481 (N_4481,N_610,N_1985);
and U4482 (N_4482,N_553,N_692);
or U4483 (N_4483,N_2245,N_1892);
xnor U4484 (N_4484,N_982,N_1824);
xor U4485 (N_4485,N_1795,N_761);
nor U4486 (N_4486,N_230,N_569);
or U4487 (N_4487,N_752,N_2336);
or U4488 (N_4488,N_517,N_1131);
or U4489 (N_4489,N_2078,N_2497);
nand U4490 (N_4490,N_1491,N_2428);
and U4491 (N_4491,N_1267,N_1738);
nand U4492 (N_4492,N_825,N_2319);
or U4493 (N_4493,N_1989,N_1842);
nor U4494 (N_4494,N_1542,N_350);
and U4495 (N_4495,N_1911,N_119);
nand U4496 (N_4496,N_639,N_1317);
and U4497 (N_4497,N_1522,N_1342);
nor U4498 (N_4498,N_918,N_1043);
nand U4499 (N_4499,N_1807,N_1419);
nand U4500 (N_4500,N_166,N_900);
or U4501 (N_4501,N_1851,N_2411);
nand U4502 (N_4502,N_2488,N_2444);
xnor U4503 (N_4503,N_1049,N_1974);
nand U4504 (N_4504,N_1468,N_544);
nor U4505 (N_4505,N_1952,N_1187);
nor U4506 (N_4506,N_1102,N_301);
nand U4507 (N_4507,N_388,N_459);
and U4508 (N_4508,N_1329,N_1770);
and U4509 (N_4509,N_2122,N_1372);
or U4510 (N_4510,N_914,N_1119);
or U4511 (N_4511,N_218,N_1071);
or U4512 (N_4512,N_1561,N_1178);
or U4513 (N_4513,N_1991,N_2256);
and U4514 (N_4514,N_2086,N_1451);
nand U4515 (N_4515,N_25,N_1998);
or U4516 (N_4516,N_2191,N_178);
nand U4517 (N_4517,N_1237,N_539);
nor U4518 (N_4518,N_2319,N_603);
nand U4519 (N_4519,N_108,N_2324);
nor U4520 (N_4520,N_67,N_2010);
nor U4521 (N_4521,N_1374,N_288);
and U4522 (N_4522,N_1337,N_858);
nor U4523 (N_4523,N_2461,N_1406);
nand U4524 (N_4524,N_27,N_1827);
nand U4525 (N_4525,N_1586,N_2455);
nand U4526 (N_4526,N_1255,N_152);
or U4527 (N_4527,N_849,N_528);
or U4528 (N_4528,N_2360,N_1373);
nand U4529 (N_4529,N_1301,N_562);
or U4530 (N_4530,N_1973,N_2403);
and U4531 (N_4531,N_759,N_670);
nor U4532 (N_4532,N_1087,N_653);
or U4533 (N_4533,N_684,N_1847);
and U4534 (N_4534,N_2246,N_623);
nand U4535 (N_4535,N_1071,N_282);
nor U4536 (N_4536,N_874,N_264);
nand U4537 (N_4537,N_510,N_1966);
nand U4538 (N_4538,N_253,N_7);
xor U4539 (N_4539,N_1577,N_1554);
nor U4540 (N_4540,N_1818,N_2037);
nand U4541 (N_4541,N_633,N_1902);
or U4542 (N_4542,N_211,N_609);
and U4543 (N_4543,N_2459,N_1990);
nand U4544 (N_4544,N_1706,N_2276);
or U4545 (N_4545,N_14,N_2327);
or U4546 (N_4546,N_345,N_2249);
nand U4547 (N_4547,N_183,N_2476);
xor U4548 (N_4548,N_1716,N_1241);
or U4549 (N_4549,N_1185,N_1135);
xnor U4550 (N_4550,N_963,N_1538);
xor U4551 (N_4551,N_522,N_2462);
nand U4552 (N_4552,N_1330,N_1046);
and U4553 (N_4553,N_1102,N_2451);
xor U4554 (N_4554,N_2471,N_1039);
and U4555 (N_4555,N_177,N_1239);
and U4556 (N_4556,N_1861,N_1557);
and U4557 (N_4557,N_331,N_1340);
or U4558 (N_4558,N_1044,N_941);
nand U4559 (N_4559,N_323,N_1987);
and U4560 (N_4560,N_582,N_1447);
nor U4561 (N_4561,N_2401,N_1623);
nor U4562 (N_4562,N_1462,N_529);
nor U4563 (N_4563,N_1019,N_2093);
nor U4564 (N_4564,N_790,N_1586);
nor U4565 (N_4565,N_1394,N_81);
and U4566 (N_4566,N_1932,N_751);
or U4567 (N_4567,N_869,N_851);
or U4568 (N_4568,N_1974,N_755);
nand U4569 (N_4569,N_2080,N_2276);
nor U4570 (N_4570,N_423,N_1398);
or U4571 (N_4571,N_2426,N_1340);
xor U4572 (N_4572,N_1682,N_2004);
or U4573 (N_4573,N_2084,N_246);
and U4574 (N_4574,N_831,N_2172);
nand U4575 (N_4575,N_444,N_2464);
nand U4576 (N_4576,N_1542,N_224);
or U4577 (N_4577,N_113,N_2434);
nand U4578 (N_4578,N_623,N_2170);
nor U4579 (N_4579,N_506,N_882);
xor U4580 (N_4580,N_2044,N_1633);
and U4581 (N_4581,N_75,N_298);
and U4582 (N_4582,N_30,N_1193);
nor U4583 (N_4583,N_1985,N_2103);
nor U4584 (N_4584,N_408,N_1124);
or U4585 (N_4585,N_1816,N_1310);
nand U4586 (N_4586,N_732,N_365);
xor U4587 (N_4587,N_1606,N_2310);
or U4588 (N_4588,N_1521,N_170);
nand U4589 (N_4589,N_321,N_1213);
nand U4590 (N_4590,N_35,N_2350);
and U4591 (N_4591,N_1853,N_241);
and U4592 (N_4592,N_650,N_249);
or U4593 (N_4593,N_371,N_534);
or U4594 (N_4594,N_1015,N_169);
and U4595 (N_4595,N_2350,N_1332);
and U4596 (N_4596,N_1842,N_337);
or U4597 (N_4597,N_2133,N_1950);
xor U4598 (N_4598,N_1841,N_407);
nand U4599 (N_4599,N_68,N_83);
or U4600 (N_4600,N_385,N_921);
nand U4601 (N_4601,N_1656,N_1807);
and U4602 (N_4602,N_1019,N_2246);
nand U4603 (N_4603,N_2134,N_873);
nor U4604 (N_4604,N_585,N_725);
or U4605 (N_4605,N_59,N_424);
or U4606 (N_4606,N_1623,N_947);
nor U4607 (N_4607,N_1616,N_631);
nor U4608 (N_4608,N_1783,N_1717);
and U4609 (N_4609,N_2025,N_1080);
nand U4610 (N_4610,N_788,N_1370);
nor U4611 (N_4611,N_2321,N_855);
xor U4612 (N_4612,N_791,N_1442);
nor U4613 (N_4613,N_1652,N_1850);
xnor U4614 (N_4614,N_1767,N_1023);
and U4615 (N_4615,N_2409,N_1291);
or U4616 (N_4616,N_31,N_2023);
or U4617 (N_4617,N_672,N_276);
xnor U4618 (N_4618,N_2298,N_1258);
or U4619 (N_4619,N_739,N_486);
and U4620 (N_4620,N_1,N_1961);
nand U4621 (N_4621,N_1070,N_1410);
nand U4622 (N_4622,N_873,N_2012);
xor U4623 (N_4623,N_1929,N_1873);
nand U4624 (N_4624,N_414,N_1949);
nand U4625 (N_4625,N_2358,N_1537);
nand U4626 (N_4626,N_425,N_2214);
or U4627 (N_4627,N_1575,N_796);
and U4628 (N_4628,N_2031,N_200);
or U4629 (N_4629,N_637,N_525);
xnor U4630 (N_4630,N_1233,N_1177);
nor U4631 (N_4631,N_2264,N_1114);
or U4632 (N_4632,N_2090,N_191);
xor U4633 (N_4633,N_1418,N_536);
xnor U4634 (N_4634,N_1821,N_1450);
nor U4635 (N_4635,N_1746,N_2031);
nand U4636 (N_4636,N_61,N_1891);
and U4637 (N_4637,N_1302,N_2439);
nand U4638 (N_4638,N_1644,N_2188);
xor U4639 (N_4639,N_1901,N_1064);
and U4640 (N_4640,N_609,N_2312);
nor U4641 (N_4641,N_2352,N_2274);
nor U4642 (N_4642,N_2182,N_1455);
nor U4643 (N_4643,N_16,N_2383);
nor U4644 (N_4644,N_1747,N_1715);
xnor U4645 (N_4645,N_319,N_256);
nor U4646 (N_4646,N_348,N_1112);
and U4647 (N_4647,N_246,N_1921);
or U4648 (N_4648,N_519,N_1546);
nor U4649 (N_4649,N_432,N_846);
nand U4650 (N_4650,N_1024,N_792);
or U4651 (N_4651,N_382,N_1228);
nand U4652 (N_4652,N_2006,N_1231);
nor U4653 (N_4653,N_1035,N_2052);
nor U4654 (N_4654,N_489,N_2283);
nand U4655 (N_4655,N_707,N_356);
or U4656 (N_4656,N_1127,N_602);
nand U4657 (N_4657,N_1100,N_2224);
and U4658 (N_4658,N_2346,N_1049);
nor U4659 (N_4659,N_903,N_2068);
nor U4660 (N_4660,N_2087,N_1924);
nand U4661 (N_4661,N_479,N_2161);
or U4662 (N_4662,N_986,N_2137);
nand U4663 (N_4663,N_1618,N_1347);
nand U4664 (N_4664,N_540,N_874);
nor U4665 (N_4665,N_1368,N_732);
nor U4666 (N_4666,N_1404,N_1054);
nand U4667 (N_4667,N_2177,N_127);
nand U4668 (N_4668,N_920,N_2369);
nor U4669 (N_4669,N_1530,N_1205);
or U4670 (N_4670,N_90,N_1318);
xnor U4671 (N_4671,N_737,N_2233);
or U4672 (N_4672,N_445,N_1797);
nor U4673 (N_4673,N_1905,N_467);
nor U4674 (N_4674,N_2410,N_753);
and U4675 (N_4675,N_968,N_383);
and U4676 (N_4676,N_2064,N_1441);
and U4677 (N_4677,N_750,N_1936);
nand U4678 (N_4678,N_886,N_698);
nor U4679 (N_4679,N_2457,N_2124);
nand U4680 (N_4680,N_1598,N_1726);
or U4681 (N_4681,N_2320,N_1810);
nor U4682 (N_4682,N_571,N_580);
xnor U4683 (N_4683,N_2450,N_219);
or U4684 (N_4684,N_637,N_104);
and U4685 (N_4685,N_632,N_1308);
nand U4686 (N_4686,N_2286,N_803);
or U4687 (N_4687,N_264,N_2188);
nor U4688 (N_4688,N_1989,N_1925);
nand U4689 (N_4689,N_91,N_471);
or U4690 (N_4690,N_45,N_813);
or U4691 (N_4691,N_1424,N_629);
or U4692 (N_4692,N_955,N_1608);
or U4693 (N_4693,N_242,N_345);
or U4694 (N_4694,N_790,N_702);
or U4695 (N_4695,N_1866,N_854);
and U4696 (N_4696,N_80,N_1576);
nor U4697 (N_4697,N_2277,N_157);
nand U4698 (N_4698,N_2189,N_405);
nor U4699 (N_4699,N_1317,N_1665);
nor U4700 (N_4700,N_1846,N_896);
xor U4701 (N_4701,N_1180,N_1030);
nand U4702 (N_4702,N_1604,N_672);
and U4703 (N_4703,N_2267,N_1850);
nor U4704 (N_4704,N_213,N_430);
or U4705 (N_4705,N_2324,N_1267);
and U4706 (N_4706,N_2102,N_41);
and U4707 (N_4707,N_2394,N_580);
or U4708 (N_4708,N_117,N_235);
xnor U4709 (N_4709,N_1974,N_1802);
nand U4710 (N_4710,N_1321,N_51);
nor U4711 (N_4711,N_1276,N_2461);
nor U4712 (N_4712,N_570,N_1013);
and U4713 (N_4713,N_345,N_347);
xor U4714 (N_4714,N_432,N_2329);
and U4715 (N_4715,N_1789,N_622);
nor U4716 (N_4716,N_1203,N_177);
nor U4717 (N_4717,N_152,N_1749);
or U4718 (N_4718,N_630,N_977);
or U4719 (N_4719,N_1656,N_515);
nor U4720 (N_4720,N_915,N_2150);
or U4721 (N_4721,N_1638,N_958);
and U4722 (N_4722,N_1580,N_604);
nor U4723 (N_4723,N_54,N_2420);
nor U4724 (N_4724,N_1831,N_1561);
and U4725 (N_4725,N_527,N_534);
nor U4726 (N_4726,N_1081,N_1791);
and U4727 (N_4727,N_1701,N_1361);
or U4728 (N_4728,N_484,N_397);
nor U4729 (N_4729,N_682,N_1907);
and U4730 (N_4730,N_2378,N_1709);
nand U4731 (N_4731,N_1174,N_1336);
and U4732 (N_4732,N_954,N_1318);
nand U4733 (N_4733,N_1308,N_1549);
nand U4734 (N_4734,N_2114,N_1626);
nor U4735 (N_4735,N_823,N_916);
nor U4736 (N_4736,N_1586,N_1230);
xnor U4737 (N_4737,N_762,N_1003);
nor U4738 (N_4738,N_49,N_1742);
or U4739 (N_4739,N_1230,N_733);
and U4740 (N_4740,N_567,N_1140);
nand U4741 (N_4741,N_434,N_2452);
xor U4742 (N_4742,N_943,N_1910);
xnor U4743 (N_4743,N_1099,N_1800);
and U4744 (N_4744,N_2489,N_1555);
or U4745 (N_4745,N_41,N_1899);
or U4746 (N_4746,N_2499,N_2296);
or U4747 (N_4747,N_2391,N_1138);
xnor U4748 (N_4748,N_348,N_1637);
nor U4749 (N_4749,N_1592,N_2380);
and U4750 (N_4750,N_481,N_1185);
nor U4751 (N_4751,N_1398,N_2176);
nand U4752 (N_4752,N_852,N_348);
nand U4753 (N_4753,N_2231,N_911);
and U4754 (N_4754,N_1622,N_435);
and U4755 (N_4755,N_570,N_2315);
or U4756 (N_4756,N_1676,N_663);
xnor U4757 (N_4757,N_572,N_996);
nand U4758 (N_4758,N_2429,N_2418);
nand U4759 (N_4759,N_1835,N_541);
and U4760 (N_4760,N_340,N_2335);
or U4761 (N_4761,N_1939,N_1997);
or U4762 (N_4762,N_1609,N_2194);
nor U4763 (N_4763,N_2146,N_1326);
or U4764 (N_4764,N_7,N_756);
nor U4765 (N_4765,N_2280,N_2259);
or U4766 (N_4766,N_1195,N_1356);
xor U4767 (N_4767,N_1893,N_66);
nor U4768 (N_4768,N_1346,N_336);
nand U4769 (N_4769,N_1825,N_1212);
nand U4770 (N_4770,N_1927,N_909);
or U4771 (N_4771,N_1298,N_1216);
nor U4772 (N_4772,N_963,N_1541);
xnor U4773 (N_4773,N_2132,N_567);
and U4774 (N_4774,N_212,N_2458);
nand U4775 (N_4775,N_1125,N_2225);
or U4776 (N_4776,N_1877,N_1625);
or U4777 (N_4777,N_524,N_856);
or U4778 (N_4778,N_1327,N_1291);
or U4779 (N_4779,N_525,N_1312);
and U4780 (N_4780,N_1662,N_80);
and U4781 (N_4781,N_852,N_646);
nand U4782 (N_4782,N_1643,N_1826);
nand U4783 (N_4783,N_1533,N_1517);
nand U4784 (N_4784,N_115,N_1530);
nand U4785 (N_4785,N_377,N_990);
nor U4786 (N_4786,N_1327,N_1585);
or U4787 (N_4787,N_1064,N_1558);
and U4788 (N_4788,N_2448,N_828);
nor U4789 (N_4789,N_856,N_2361);
and U4790 (N_4790,N_1266,N_1514);
nand U4791 (N_4791,N_1097,N_1434);
and U4792 (N_4792,N_1733,N_124);
nand U4793 (N_4793,N_234,N_1690);
nor U4794 (N_4794,N_1846,N_1112);
nor U4795 (N_4795,N_930,N_2446);
nand U4796 (N_4796,N_1031,N_2301);
nor U4797 (N_4797,N_1666,N_411);
or U4798 (N_4798,N_288,N_1488);
nand U4799 (N_4799,N_532,N_270);
nor U4800 (N_4800,N_848,N_887);
nor U4801 (N_4801,N_1562,N_1982);
nor U4802 (N_4802,N_1018,N_1117);
or U4803 (N_4803,N_2321,N_2072);
or U4804 (N_4804,N_2107,N_372);
nand U4805 (N_4805,N_2425,N_426);
nor U4806 (N_4806,N_2029,N_1940);
xnor U4807 (N_4807,N_531,N_212);
nor U4808 (N_4808,N_2038,N_1314);
or U4809 (N_4809,N_1691,N_1365);
nand U4810 (N_4810,N_1056,N_1121);
nor U4811 (N_4811,N_1819,N_406);
nor U4812 (N_4812,N_1539,N_1092);
nor U4813 (N_4813,N_1102,N_1023);
and U4814 (N_4814,N_2027,N_1618);
nand U4815 (N_4815,N_1853,N_2428);
nor U4816 (N_4816,N_2377,N_2322);
nand U4817 (N_4817,N_506,N_117);
or U4818 (N_4818,N_391,N_163);
nand U4819 (N_4819,N_1957,N_1472);
or U4820 (N_4820,N_64,N_1767);
or U4821 (N_4821,N_1475,N_2439);
nor U4822 (N_4822,N_615,N_1631);
nor U4823 (N_4823,N_597,N_966);
nand U4824 (N_4824,N_1331,N_2342);
or U4825 (N_4825,N_1096,N_1274);
or U4826 (N_4826,N_1013,N_1022);
or U4827 (N_4827,N_2214,N_1209);
nor U4828 (N_4828,N_722,N_1255);
nor U4829 (N_4829,N_1892,N_1424);
or U4830 (N_4830,N_425,N_323);
and U4831 (N_4831,N_1190,N_167);
nand U4832 (N_4832,N_44,N_1304);
nor U4833 (N_4833,N_2010,N_183);
or U4834 (N_4834,N_454,N_1225);
or U4835 (N_4835,N_1911,N_957);
nand U4836 (N_4836,N_2497,N_847);
nand U4837 (N_4837,N_47,N_1583);
xnor U4838 (N_4838,N_1003,N_138);
nor U4839 (N_4839,N_1077,N_1931);
or U4840 (N_4840,N_1182,N_244);
nand U4841 (N_4841,N_1733,N_1777);
nor U4842 (N_4842,N_445,N_1019);
and U4843 (N_4843,N_1448,N_2197);
nand U4844 (N_4844,N_323,N_684);
xnor U4845 (N_4845,N_1428,N_2495);
nand U4846 (N_4846,N_339,N_1397);
xnor U4847 (N_4847,N_1222,N_1037);
nand U4848 (N_4848,N_1286,N_1507);
or U4849 (N_4849,N_1101,N_1248);
nand U4850 (N_4850,N_1974,N_843);
nor U4851 (N_4851,N_454,N_1299);
nand U4852 (N_4852,N_1031,N_334);
and U4853 (N_4853,N_1193,N_2141);
nand U4854 (N_4854,N_1075,N_330);
nand U4855 (N_4855,N_2279,N_1866);
nor U4856 (N_4856,N_728,N_1355);
and U4857 (N_4857,N_989,N_490);
nand U4858 (N_4858,N_1948,N_1255);
nor U4859 (N_4859,N_2310,N_1190);
or U4860 (N_4860,N_2492,N_1917);
nand U4861 (N_4861,N_904,N_658);
nand U4862 (N_4862,N_1983,N_1252);
nor U4863 (N_4863,N_119,N_2396);
nand U4864 (N_4864,N_231,N_1517);
or U4865 (N_4865,N_1327,N_1442);
nand U4866 (N_4866,N_2312,N_190);
nor U4867 (N_4867,N_2499,N_959);
nand U4868 (N_4868,N_2063,N_810);
or U4869 (N_4869,N_163,N_1362);
and U4870 (N_4870,N_209,N_1054);
and U4871 (N_4871,N_276,N_30);
nand U4872 (N_4872,N_2051,N_1623);
xnor U4873 (N_4873,N_1918,N_1909);
nand U4874 (N_4874,N_90,N_506);
and U4875 (N_4875,N_2090,N_1585);
nand U4876 (N_4876,N_1831,N_667);
and U4877 (N_4877,N_1142,N_2373);
and U4878 (N_4878,N_1305,N_2245);
or U4879 (N_4879,N_1155,N_974);
nor U4880 (N_4880,N_146,N_1995);
xnor U4881 (N_4881,N_1562,N_2353);
nand U4882 (N_4882,N_2250,N_1041);
and U4883 (N_4883,N_264,N_114);
nand U4884 (N_4884,N_180,N_495);
xor U4885 (N_4885,N_2028,N_2045);
nor U4886 (N_4886,N_1021,N_1587);
or U4887 (N_4887,N_1478,N_1115);
nor U4888 (N_4888,N_1766,N_392);
nor U4889 (N_4889,N_89,N_2252);
nor U4890 (N_4890,N_1662,N_1461);
nor U4891 (N_4891,N_1995,N_646);
nand U4892 (N_4892,N_35,N_883);
nor U4893 (N_4893,N_918,N_2101);
nand U4894 (N_4894,N_165,N_1744);
nand U4895 (N_4895,N_2386,N_1708);
nor U4896 (N_4896,N_941,N_2299);
nor U4897 (N_4897,N_1533,N_551);
nor U4898 (N_4898,N_193,N_1516);
or U4899 (N_4899,N_2408,N_705);
and U4900 (N_4900,N_749,N_1459);
or U4901 (N_4901,N_998,N_432);
and U4902 (N_4902,N_304,N_19);
nand U4903 (N_4903,N_784,N_1613);
nor U4904 (N_4904,N_655,N_1968);
or U4905 (N_4905,N_608,N_406);
or U4906 (N_4906,N_378,N_1889);
or U4907 (N_4907,N_1263,N_1474);
or U4908 (N_4908,N_1025,N_65);
nor U4909 (N_4909,N_2220,N_600);
nand U4910 (N_4910,N_1093,N_947);
nor U4911 (N_4911,N_362,N_1437);
nand U4912 (N_4912,N_2274,N_1578);
nor U4913 (N_4913,N_116,N_1420);
nand U4914 (N_4914,N_1062,N_2426);
nor U4915 (N_4915,N_1860,N_1628);
nand U4916 (N_4916,N_368,N_2283);
or U4917 (N_4917,N_1519,N_54);
and U4918 (N_4918,N_1526,N_549);
and U4919 (N_4919,N_2412,N_2446);
xnor U4920 (N_4920,N_839,N_740);
or U4921 (N_4921,N_196,N_2365);
nor U4922 (N_4922,N_1774,N_1992);
or U4923 (N_4923,N_168,N_1300);
nor U4924 (N_4924,N_1105,N_336);
nor U4925 (N_4925,N_1366,N_1426);
or U4926 (N_4926,N_639,N_961);
and U4927 (N_4927,N_2155,N_993);
and U4928 (N_4928,N_2392,N_1855);
nor U4929 (N_4929,N_1286,N_941);
or U4930 (N_4930,N_2177,N_2351);
or U4931 (N_4931,N_406,N_679);
or U4932 (N_4932,N_1028,N_1509);
nor U4933 (N_4933,N_758,N_987);
nand U4934 (N_4934,N_2129,N_1562);
or U4935 (N_4935,N_1715,N_1935);
nor U4936 (N_4936,N_128,N_1731);
xor U4937 (N_4937,N_261,N_1558);
nor U4938 (N_4938,N_527,N_2408);
xor U4939 (N_4939,N_1995,N_1667);
nor U4940 (N_4940,N_412,N_1612);
nand U4941 (N_4941,N_2328,N_645);
nor U4942 (N_4942,N_1744,N_2254);
nor U4943 (N_4943,N_1570,N_107);
nor U4944 (N_4944,N_2257,N_671);
or U4945 (N_4945,N_8,N_1889);
nand U4946 (N_4946,N_699,N_1416);
nand U4947 (N_4947,N_1928,N_1073);
or U4948 (N_4948,N_729,N_2286);
or U4949 (N_4949,N_18,N_841);
or U4950 (N_4950,N_2012,N_1815);
nor U4951 (N_4951,N_224,N_1413);
and U4952 (N_4952,N_1418,N_1682);
xor U4953 (N_4953,N_1512,N_1564);
nor U4954 (N_4954,N_2183,N_2294);
nand U4955 (N_4955,N_1323,N_1214);
and U4956 (N_4956,N_180,N_110);
and U4957 (N_4957,N_2315,N_2313);
or U4958 (N_4958,N_242,N_130);
nor U4959 (N_4959,N_2250,N_2106);
nand U4960 (N_4960,N_1055,N_9);
and U4961 (N_4961,N_269,N_1529);
xnor U4962 (N_4962,N_1176,N_1992);
nand U4963 (N_4963,N_911,N_2412);
and U4964 (N_4964,N_1906,N_735);
or U4965 (N_4965,N_933,N_255);
nand U4966 (N_4966,N_446,N_740);
xnor U4967 (N_4967,N_2284,N_1473);
xnor U4968 (N_4968,N_1211,N_400);
nor U4969 (N_4969,N_1749,N_1131);
xnor U4970 (N_4970,N_277,N_925);
nand U4971 (N_4971,N_2009,N_1592);
and U4972 (N_4972,N_2150,N_1142);
or U4973 (N_4973,N_929,N_999);
and U4974 (N_4974,N_558,N_2080);
and U4975 (N_4975,N_57,N_209);
and U4976 (N_4976,N_325,N_1674);
or U4977 (N_4977,N_265,N_1041);
and U4978 (N_4978,N_875,N_1742);
nor U4979 (N_4979,N_986,N_340);
nand U4980 (N_4980,N_1059,N_163);
nor U4981 (N_4981,N_180,N_255);
or U4982 (N_4982,N_610,N_930);
nand U4983 (N_4983,N_1520,N_1466);
and U4984 (N_4984,N_1282,N_1907);
xnor U4985 (N_4985,N_2047,N_280);
or U4986 (N_4986,N_2179,N_1761);
and U4987 (N_4987,N_1306,N_1075);
nor U4988 (N_4988,N_1914,N_2230);
nand U4989 (N_4989,N_2152,N_2312);
or U4990 (N_4990,N_1138,N_2096);
nand U4991 (N_4991,N_1499,N_1711);
nand U4992 (N_4992,N_457,N_1343);
or U4993 (N_4993,N_1913,N_1664);
and U4994 (N_4994,N_2300,N_1515);
xor U4995 (N_4995,N_115,N_1193);
nor U4996 (N_4996,N_433,N_1542);
and U4997 (N_4997,N_71,N_2193);
nor U4998 (N_4998,N_354,N_1102);
and U4999 (N_4999,N_1943,N_2215);
nor U5000 (N_5000,N_4404,N_3840);
nand U5001 (N_5001,N_4302,N_2762);
or U5002 (N_5002,N_3397,N_3565);
nand U5003 (N_5003,N_3601,N_3387);
xor U5004 (N_5004,N_3544,N_4028);
or U5005 (N_5005,N_4792,N_3677);
or U5006 (N_5006,N_4517,N_3663);
and U5007 (N_5007,N_4694,N_2855);
nand U5008 (N_5008,N_2773,N_4596);
nor U5009 (N_5009,N_2723,N_4498);
or U5010 (N_5010,N_4865,N_3498);
xor U5011 (N_5011,N_3585,N_2508);
or U5012 (N_5012,N_3484,N_4668);
and U5013 (N_5013,N_4593,N_3288);
or U5014 (N_5014,N_3383,N_3562);
nand U5015 (N_5015,N_2738,N_3316);
or U5016 (N_5016,N_2629,N_3633);
and U5017 (N_5017,N_4120,N_3309);
nor U5018 (N_5018,N_4351,N_4034);
nand U5019 (N_5019,N_3742,N_4383);
or U5020 (N_5020,N_2826,N_3209);
nand U5021 (N_5021,N_2842,N_2811);
or U5022 (N_5022,N_3375,N_3963);
and U5023 (N_5023,N_3342,N_3481);
nand U5024 (N_5024,N_3207,N_4598);
or U5025 (N_5025,N_2816,N_3875);
and U5026 (N_5026,N_4967,N_3867);
or U5027 (N_5027,N_4512,N_2505);
and U5028 (N_5028,N_4379,N_2840);
and U5029 (N_5029,N_3907,N_2654);
xor U5030 (N_5030,N_3324,N_4176);
nor U5031 (N_5031,N_3512,N_4925);
xor U5032 (N_5032,N_3317,N_4943);
nand U5033 (N_5033,N_4180,N_3169);
nor U5034 (N_5034,N_2831,N_4101);
nor U5035 (N_5035,N_4049,N_4775);
nor U5036 (N_5036,N_2748,N_3529);
nor U5037 (N_5037,N_2830,N_3142);
and U5038 (N_5038,N_3129,N_4990);
nand U5039 (N_5039,N_4684,N_4154);
nor U5040 (N_5040,N_3398,N_2512);
or U5041 (N_5041,N_2917,N_3403);
xnor U5042 (N_5042,N_3208,N_4195);
nor U5043 (N_5043,N_3351,N_4393);
or U5044 (N_5044,N_3872,N_2945);
nand U5045 (N_5045,N_4421,N_3639);
xor U5046 (N_5046,N_4810,N_3292);
xor U5047 (N_5047,N_2670,N_4892);
nor U5048 (N_5048,N_2506,N_3311);
xor U5049 (N_5049,N_4224,N_3011);
or U5050 (N_5050,N_3115,N_4485);
nor U5051 (N_5051,N_3451,N_3181);
or U5052 (N_5052,N_2550,N_4141);
and U5053 (N_5053,N_3100,N_4181);
or U5054 (N_5054,N_4402,N_4928);
nand U5055 (N_5055,N_4249,N_3096);
xor U5056 (N_5056,N_3640,N_3732);
or U5057 (N_5057,N_4396,N_3791);
nand U5058 (N_5058,N_2535,N_4375);
nor U5059 (N_5059,N_4853,N_3438);
nor U5060 (N_5060,N_2839,N_3273);
nor U5061 (N_5061,N_4663,N_2967);
nor U5062 (N_5062,N_4132,N_2931);
nand U5063 (N_5063,N_3097,N_4709);
xnor U5064 (N_5064,N_3727,N_4585);
nand U5065 (N_5065,N_3682,N_3658);
or U5066 (N_5066,N_4378,N_3087);
or U5067 (N_5067,N_2521,N_4069);
xnor U5068 (N_5068,N_2824,N_2782);
or U5069 (N_5069,N_4236,N_4398);
nor U5070 (N_5070,N_4414,N_3153);
nand U5071 (N_5071,N_4183,N_3814);
and U5072 (N_5072,N_2769,N_4146);
or U5073 (N_5073,N_4873,N_4160);
and U5074 (N_5074,N_3084,N_3884);
or U5075 (N_5075,N_4059,N_4995);
nand U5076 (N_5076,N_4969,N_3635);
nand U5077 (N_5077,N_3491,N_2780);
and U5078 (N_5078,N_4891,N_3604);
or U5079 (N_5079,N_3740,N_4215);
xor U5080 (N_5080,N_2717,N_3574);
nor U5081 (N_5081,N_4561,N_3165);
xnor U5082 (N_5082,N_4425,N_4122);
nand U5083 (N_5083,N_3137,N_3701);
nand U5084 (N_5084,N_3305,N_4908);
and U5085 (N_5085,N_4608,N_3012);
nand U5086 (N_5086,N_4446,N_4764);
and U5087 (N_5087,N_3001,N_4948);
nand U5088 (N_5088,N_2631,N_4364);
and U5089 (N_5089,N_3920,N_3401);
xor U5090 (N_5090,N_3217,N_3507);
nand U5091 (N_5091,N_4964,N_2609);
and U5092 (N_5092,N_3098,N_3124);
nand U5093 (N_5093,N_3447,N_4455);
and U5094 (N_5094,N_4124,N_3193);
nand U5095 (N_5095,N_3693,N_3159);
or U5096 (N_5096,N_2792,N_3712);
or U5097 (N_5097,N_4554,N_4348);
xor U5098 (N_5098,N_3670,N_2563);
or U5099 (N_5099,N_3690,N_3263);
nor U5100 (N_5100,N_3487,N_4475);
and U5101 (N_5101,N_4650,N_4788);
nor U5102 (N_5102,N_4898,N_2763);
nor U5103 (N_5103,N_3276,N_3478);
and U5104 (N_5104,N_4316,N_3952);
nand U5105 (N_5105,N_4340,N_4603);
nand U5106 (N_5106,N_3282,N_2971);
and U5107 (N_5107,N_2895,N_3702);
nor U5108 (N_5108,N_4202,N_2600);
or U5109 (N_5109,N_4574,N_3514);
nand U5110 (N_5110,N_4060,N_4695);
or U5111 (N_5111,N_2972,N_4371);
or U5112 (N_5112,N_2926,N_2531);
and U5113 (N_5113,N_3573,N_3081);
nor U5114 (N_5114,N_2869,N_3564);
and U5115 (N_5115,N_4386,N_4391);
nor U5116 (N_5116,N_4291,N_4743);
nand U5117 (N_5117,N_4263,N_3474);
nor U5118 (N_5118,N_4165,N_3789);
or U5119 (N_5119,N_4271,N_3848);
or U5120 (N_5120,N_4790,N_3272);
nor U5121 (N_5121,N_2779,N_4392);
nand U5122 (N_5122,N_4061,N_4468);
or U5123 (N_5123,N_3518,N_3265);
and U5124 (N_5124,N_4056,N_3306);
xor U5125 (N_5125,N_4685,N_2844);
nand U5126 (N_5126,N_2676,N_2529);
or U5127 (N_5127,N_4084,N_2975);
nand U5128 (N_5128,N_4712,N_4701);
or U5129 (N_5129,N_4870,N_4965);
nor U5130 (N_5130,N_4228,N_4765);
xor U5131 (N_5131,N_3349,N_4845);
and U5132 (N_5132,N_4368,N_2851);
nor U5133 (N_5133,N_4354,N_2599);
xnor U5134 (N_5134,N_3899,N_3915);
nor U5135 (N_5135,N_2700,N_2680);
nor U5136 (N_5136,N_4630,N_3245);
or U5137 (N_5137,N_4867,N_3123);
nand U5138 (N_5138,N_3620,N_3869);
nand U5139 (N_5139,N_3384,N_2897);
xor U5140 (N_5140,N_3061,N_2865);
and U5141 (N_5141,N_2705,N_3569);
nor U5142 (N_5142,N_3331,N_4921);
nand U5143 (N_5143,N_3535,N_2520);
nand U5144 (N_5144,N_4131,N_4234);
or U5145 (N_5145,N_4331,N_2827);
or U5146 (N_5146,N_4460,N_3589);
and U5147 (N_5147,N_3737,N_4589);
nor U5148 (N_5148,N_3505,N_4530);
and U5149 (N_5149,N_3857,N_2577);
or U5150 (N_5150,N_4725,N_3798);
or U5151 (N_5151,N_4282,N_2746);
nor U5152 (N_5152,N_3261,N_4547);
and U5153 (N_5153,N_3592,N_2591);
and U5154 (N_5154,N_4086,N_4038);
and U5155 (N_5155,N_3628,N_2857);
and U5156 (N_5156,N_4994,N_3025);
nand U5157 (N_5157,N_4535,N_3266);
or U5158 (N_5158,N_4706,N_4168);
and U5159 (N_5159,N_4940,N_4631);
nand U5160 (N_5160,N_4436,N_4923);
nand U5161 (N_5161,N_2704,N_4044);
nor U5162 (N_5162,N_3860,N_4403);
or U5163 (N_5163,N_4828,N_3005);
xnor U5164 (N_5164,N_4434,N_4611);
or U5165 (N_5165,N_4273,N_3902);
nand U5166 (N_5166,N_2904,N_2775);
xor U5167 (N_5167,N_2836,N_4666);
and U5168 (N_5168,N_3988,N_3026);
and U5169 (N_5169,N_3216,N_4824);
nand U5170 (N_5170,N_3195,N_4255);
nor U5171 (N_5171,N_2856,N_4619);
and U5172 (N_5172,N_4689,N_3104);
nand U5173 (N_5173,N_4629,N_3392);
nand U5174 (N_5174,N_2527,N_4014);
nor U5175 (N_5175,N_4313,N_4651);
nor U5176 (N_5176,N_4047,N_3768);
or U5177 (N_5177,N_3364,N_4099);
or U5178 (N_5178,N_4238,N_4641);
nand U5179 (N_5179,N_4926,N_3625);
or U5180 (N_5180,N_3386,N_2502);
or U5181 (N_5181,N_4791,N_3782);
and U5182 (N_5182,N_4886,N_4872);
nor U5183 (N_5183,N_4051,N_4301);
nand U5184 (N_5184,N_3239,N_3551);
xor U5185 (N_5185,N_2879,N_4411);
xnor U5186 (N_5186,N_4516,N_4799);
nand U5187 (N_5187,N_4907,N_3004);
nand U5188 (N_5188,N_3360,N_3843);
nor U5189 (N_5189,N_4423,N_3959);
nor U5190 (N_5190,N_4841,N_3232);
and U5191 (N_5191,N_3321,N_3906);
or U5192 (N_5192,N_3422,N_2913);
nand U5193 (N_5193,N_2647,N_4570);
or U5194 (N_5194,N_2530,N_3739);
or U5195 (N_5195,N_3876,N_2691);
nand U5196 (N_5196,N_2803,N_4521);
or U5197 (N_5197,N_4072,N_3699);
nor U5198 (N_5198,N_3885,N_4197);
or U5199 (N_5199,N_4532,N_3796);
nand U5200 (N_5200,N_3287,N_2832);
or U5201 (N_5201,N_3520,N_4473);
and U5202 (N_5202,N_3548,N_4357);
xor U5203 (N_5203,N_4728,N_3431);
nand U5204 (N_5204,N_3488,N_3674);
nand U5205 (N_5205,N_3524,N_3400);
and U5206 (N_5206,N_4092,N_3199);
or U5207 (N_5207,N_2988,N_4537);
and U5208 (N_5208,N_3652,N_2616);
nand U5209 (N_5209,N_3378,N_4678);
nor U5210 (N_5210,N_4062,N_3079);
nor U5211 (N_5211,N_3347,N_3729);
nor U5212 (N_5212,N_2656,N_2932);
or U5213 (N_5213,N_2923,N_3746);
and U5214 (N_5214,N_4345,N_3893);
nor U5215 (N_5215,N_3469,N_2852);
or U5216 (N_5216,N_3913,N_2545);
nand U5217 (N_5217,N_4671,N_4178);
nor U5218 (N_5218,N_3215,N_3174);
and U5219 (N_5219,N_3615,N_3271);
and U5220 (N_5220,N_4729,N_4250);
nor U5221 (N_5221,N_3458,N_2644);
and U5222 (N_5222,N_4174,N_4735);
and U5223 (N_5223,N_2947,N_4707);
or U5224 (N_5224,N_3500,N_3108);
and U5225 (N_5225,N_3171,N_3968);
nand U5226 (N_5226,N_4491,N_4214);
and U5227 (N_5227,N_3979,N_2959);
or U5228 (N_5228,N_4595,N_4858);
nand U5229 (N_5229,N_2754,N_4232);
or U5230 (N_5230,N_3489,N_4219);
nand U5231 (N_5231,N_4594,N_3462);
xnor U5232 (N_5232,N_2513,N_4989);
and U5233 (N_5233,N_4638,N_2804);
nor U5234 (N_5234,N_3611,N_3736);
or U5235 (N_5235,N_3058,N_3894);
and U5236 (N_5236,N_4055,N_2871);
nand U5237 (N_5237,N_3095,N_4453);
or U5238 (N_5238,N_2651,N_4677);
xor U5239 (N_5239,N_2685,N_3040);
xor U5240 (N_5240,N_3371,N_4551);
nor U5241 (N_5241,N_3766,N_4657);
nor U5242 (N_5242,N_3803,N_4006);
nand U5243 (N_5243,N_4447,N_2737);
nor U5244 (N_5244,N_4022,N_3643);
or U5245 (N_5245,N_4519,N_4557);
nor U5246 (N_5246,N_4693,N_3607);
nor U5247 (N_5247,N_4114,N_4785);
nand U5248 (N_5248,N_4067,N_3441);
nand U5249 (N_5249,N_3577,N_3036);
and U5250 (N_5250,N_4253,N_4427);
nor U5251 (N_5251,N_2756,N_3301);
or U5252 (N_5252,N_4767,N_4040);
nor U5253 (N_5253,N_3747,N_2949);
and U5254 (N_5254,N_2618,N_4157);
and U5255 (N_5255,N_3424,N_2874);
and U5256 (N_5256,N_4991,N_2678);
and U5257 (N_5257,N_4981,N_3890);
nor U5258 (N_5258,N_2747,N_2817);
or U5259 (N_5259,N_3667,N_4642);
xnor U5260 (N_5260,N_4544,N_4935);
and U5261 (N_5261,N_2781,N_3163);
xor U5262 (N_5262,N_4441,N_2681);
nand U5263 (N_5263,N_3328,N_4199);
or U5264 (N_5264,N_4772,N_3303);
and U5265 (N_5265,N_2559,N_3408);
xnor U5266 (N_5266,N_3878,N_4279);
and U5267 (N_5267,N_4992,N_3405);
or U5268 (N_5268,N_4390,N_3109);
or U5269 (N_5269,N_3918,N_4419);
nand U5270 (N_5270,N_2937,N_3626);
nand U5271 (N_5271,N_4106,N_2673);
xnor U5272 (N_5272,N_2999,N_4352);
nor U5273 (N_5273,N_4996,N_3764);
and U5274 (N_5274,N_3089,N_4801);
or U5275 (N_5275,N_4459,N_2507);
nand U5276 (N_5276,N_3781,N_3343);
nand U5277 (N_5277,N_2946,N_4098);
nand U5278 (N_5278,N_4346,N_3322);
nand U5279 (N_5279,N_2511,N_4334);
nor U5280 (N_5280,N_4325,N_2594);
and U5281 (N_5281,N_4959,N_3989);
xor U5282 (N_5282,N_3563,N_4080);
and U5283 (N_5283,N_4456,N_3657);
nand U5284 (N_5284,N_4829,N_3866);
xor U5285 (N_5285,N_3049,N_2846);
and U5286 (N_5286,N_4280,N_3641);
nor U5287 (N_5287,N_3310,N_4531);
and U5288 (N_5288,N_4887,N_4927);
and U5289 (N_5289,N_3943,N_2900);
xnor U5290 (N_5290,N_3332,N_3119);
nor U5291 (N_5291,N_4087,N_2720);
or U5292 (N_5292,N_4874,N_2605);
nor U5293 (N_5293,N_3183,N_4888);
and U5294 (N_5294,N_3511,N_2572);
xor U5295 (N_5295,N_3919,N_4477);
and U5296 (N_5296,N_4756,N_2884);
nor U5297 (N_5297,N_3121,N_4920);
nand U5298 (N_5298,N_3996,N_4033);
nand U5299 (N_5299,N_4633,N_4504);
nand U5300 (N_5300,N_3226,N_3809);
nand U5301 (N_5301,N_3300,N_3912);
and U5302 (N_5302,N_4781,N_2902);
nor U5303 (N_5303,N_4711,N_3825);
nor U5304 (N_5304,N_2861,N_3391);
nand U5305 (N_5305,N_2794,N_2663);
or U5306 (N_5306,N_4451,N_4111);
or U5307 (N_5307,N_2984,N_2761);
and U5308 (N_5308,N_2974,N_4645);
nand U5309 (N_5309,N_3683,N_2981);
xnor U5310 (N_5310,N_4283,N_3720);
nor U5311 (N_5311,N_3991,N_4448);
or U5312 (N_5312,N_4803,N_2948);
xnor U5313 (N_5313,N_2751,N_2944);
nor U5314 (N_5314,N_3140,N_2930);
xnor U5315 (N_5315,N_4945,N_4140);
and U5316 (N_5316,N_4230,N_2658);
or U5317 (N_5317,N_2684,N_3584);
nand U5318 (N_5318,N_3721,N_4076);
xor U5319 (N_5319,N_4546,N_3760);
nand U5320 (N_5320,N_3889,N_4982);
or U5321 (N_5321,N_4564,N_4635);
xnor U5322 (N_5322,N_4272,N_3964);
or U5323 (N_5323,N_3823,N_4761);
or U5324 (N_5324,N_3992,N_4085);
nand U5325 (N_5325,N_4961,N_4401);
nor U5326 (N_5326,N_4513,N_3075);
or U5327 (N_5327,N_2584,N_4245);
nor U5328 (N_5328,N_4248,N_3839);
nor U5329 (N_5329,N_4039,N_4387);
or U5330 (N_5330,N_2634,N_4605);
nor U5331 (N_5331,N_4221,N_4186);
or U5332 (N_5332,N_4856,N_3538);
and U5333 (N_5333,N_4822,N_3810);
nand U5334 (N_5334,N_3466,N_4899);
and U5335 (N_5335,N_4933,N_4295);
or U5336 (N_5336,N_4924,N_3554);
or U5337 (N_5337,N_4138,N_3182);
and U5338 (N_5338,N_3185,N_3304);
and U5339 (N_5339,N_4013,N_4161);
or U5340 (N_5340,N_4628,N_3880);
nor U5341 (N_5341,N_3837,N_4147);
nor U5342 (N_5342,N_4363,N_4911);
nand U5343 (N_5343,N_4335,N_4237);
and U5344 (N_5344,N_3196,N_3528);
nor U5345 (N_5345,N_3495,N_3204);
and U5346 (N_5346,N_3981,N_2834);
xor U5347 (N_5347,N_2885,N_3479);
nor U5348 (N_5348,N_4164,N_2850);
nor U5349 (N_5349,N_2553,N_2696);
and U5350 (N_5350,N_3399,N_3990);
xor U5351 (N_5351,N_3619,N_4063);
or U5352 (N_5352,N_4377,N_3138);
nand U5353 (N_5353,N_2568,N_3064);
nor U5354 (N_5354,N_3561,N_4835);
nand U5355 (N_5355,N_4052,N_3853);
xor U5356 (N_5356,N_4023,N_4590);
or U5357 (N_5357,N_4261,N_2725);
or U5358 (N_5358,N_3955,N_3082);
nor U5359 (N_5359,N_2822,N_4332);
nor U5360 (N_5360,N_3013,N_3960);
nor U5361 (N_5361,N_3033,N_4601);
and U5362 (N_5362,N_4958,N_3694);
or U5363 (N_5363,N_4620,N_4481);
nand U5364 (N_5364,N_3523,N_4714);
and U5365 (N_5365,N_3556,N_3937);
or U5366 (N_5366,N_3243,N_2873);
nand U5367 (N_5367,N_4222,N_4568);
and U5368 (N_5368,N_4486,N_4418);
nand U5369 (N_5369,N_3223,N_4552);
nor U5370 (N_5370,N_4526,N_2886);
and U5371 (N_5371,N_3010,N_3629);
and U5372 (N_5372,N_4527,N_4819);
and U5373 (N_5373,N_4470,N_4339);
xnor U5374 (N_5374,N_2783,N_4242);
nor U5375 (N_5375,N_2745,N_3923);
xnor U5376 (N_5376,N_4278,N_3380);
nand U5377 (N_5377,N_3756,N_4464);
nor U5378 (N_5378,N_3419,N_4614);
nand U5379 (N_5379,N_3056,N_4407);
nand U5380 (N_5380,N_2878,N_3672);
and U5381 (N_5381,N_2743,N_4478);
nor U5382 (N_5382,N_4745,N_3503);
or U5383 (N_5383,N_2922,N_4832);
and U5384 (N_5384,N_3800,N_2966);
or U5385 (N_5385,N_4094,N_3143);
or U5386 (N_5386,N_3319,N_2820);
or U5387 (N_5387,N_4751,N_2706);
or U5388 (N_5388,N_3833,N_3352);
or U5389 (N_5389,N_3785,N_2955);
nand U5390 (N_5390,N_3314,N_4749);
and U5391 (N_5391,N_3131,N_4244);
nor U5392 (N_5392,N_4980,N_3726);
or U5393 (N_5393,N_3647,N_4754);
and U5394 (N_5394,N_4844,N_2564);
nor U5395 (N_5395,N_4548,N_2710);
nand U5396 (N_5396,N_4833,N_3016);
and U5397 (N_5397,N_2613,N_3339);
nand U5398 (N_5398,N_3333,N_4905);
and U5399 (N_5399,N_4871,N_4962);
nor U5400 (N_5400,N_2801,N_3454);
or U5401 (N_5401,N_3394,N_4815);
or U5402 (N_5402,N_3407,N_4988);
or U5403 (N_5403,N_2582,N_2735);
nand U5404 (N_5404,N_3444,N_3390);
and U5405 (N_5405,N_4576,N_3817);
xnor U5406 (N_5406,N_2938,N_4834);
xnor U5407 (N_5407,N_4704,N_4660);
nand U5408 (N_5408,N_3020,N_2894);
nand U5409 (N_5409,N_4042,N_4308);
or U5410 (N_5410,N_4875,N_3425);
nand U5411 (N_5411,N_4944,N_4826);
nor U5412 (N_5412,N_3455,N_3376);
nand U5413 (N_5413,N_3961,N_4682);
xor U5414 (N_5414,N_2750,N_3490);
and U5415 (N_5415,N_3771,N_2731);
nand U5416 (N_5416,N_4912,N_4732);
xor U5417 (N_5417,N_3815,N_3480);
nor U5418 (N_5418,N_2730,N_2632);
or U5419 (N_5419,N_3030,N_2573);
or U5420 (N_5420,N_3231,N_3997);
or U5421 (N_5421,N_3887,N_2669);
xnor U5422 (N_5422,N_3521,N_2538);
or U5423 (N_5423,N_2786,N_4632);
or U5424 (N_5424,N_3173,N_3218);
nor U5425 (N_5425,N_3168,N_4771);
nor U5426 (N_5426,N_3356,N_4342);
and U5427 (N_5427,N_3687,N_3935);
and U5428 (N_5428,N_3982,N_4951);
and U5429 (N_5429,N_2662,N_2778);
nand U5430 (N_5430,N_3734,N_3200);
nand U5431 (N_5431,N_4960,N_4720);
nand U5432 (N_5432,N_2790,N_4229);
and U5433 (N_5433,N_3679,N_2619);
or U5434 (N_5434,N_4410,N_4285);
and U5435 (N_5435,N_2934,N_4538);
or U5436 (N_5436,N_4173,N_4264);
nand U5437 (N_5437,N_4857,N_2526);
nor U5438 (N_5438,N_2668,N_3717);
and U5439 (N_5439,N_2627,N_4191);
nand U5440 (N_5440,N_4484,N_3227);
nor U5441 (N_5441,N_3286,N_2636);
nand U5442 (N_5442,N_3616,N_4035);
and U5443 (N_5443,N_3229,N_3427);
or U5444 (N_5444,N_2915,N_4012);
nor U5445 (N_5445,N_4747,N_4742);
or U5446 (N_5446,N_3618,N_3113);
nand U5447 (N_5447,N_4766,N_4697);
and U5448 (N_5448,N_4104,N_4373);
nand U5449 (N_5449,N_2648,N_3938);
nand U5450 (N_5450,N_4814,N_4939);
or U5451 (N_5451,N_3127,N_4068);
xnor U5452 (N_5452,N_4399,N_2522);
nor U5453 (N_5453,N_3801,N_2875);
and U5454 (N_5454,N_2893,N_2909);
and U5455 (N_5455,N_3206,N_2569);
nand U5456 (N_5456,N_3336,N_4643);
nand U5457 (N_5457,N_3829,N_4490);
and U5458 (N_5458,N_3692,N_3522);
nor U5459 (N_5459,N_4949,N_2712);
xnor U5460 (N_5460,N_3656,N_4209);
nand U5461 (N_5461,N_2500,N_4139);
nand U5462 (N_5462,N_4226,N_4942);
nor U5463 (N_5463,N_2918,N_3579);
and U5464 (N_5464,N_4362,N_3192);
or U5465 (N_5465,N_3086,N_3358);
and U5466 (N_5466,N_4208,N_2694);
nor U5467 (N_5467,N_4626,N_3002);
nor U5468 (N_5468,N_2766,N_3450);
and U5469 (N_5469,N_2808,N_3307);
nor U5470 (N_5470,N_3877,N_4699);
nand U5471 (N_5471,N_3006,N_3983);
or U5472 (N_5472,N_2642,N_4883);
nand U5473 (N_5473,N_4247,N_4567);
or U5474 (N_5474,N_2742,N_4880);
nand U5475 (N_5475,N_4324,N_3492);
or U5476 (N_5476,N_3105,N_3854);
and U5477 (N_5477,N_3892,N_4471);
and U5478 (N_5478,N_4003,N_2760);
nor U5479 (N_5479,N_4240,N_4406);
or U5480 (N_5480,N_4480,N_2965);
and U5481 (N_5481,N_4162,N_2727);
or U5482 (N_5482,N_3921,N_4549);
and U5483 (N_5483,N_2798,N_3290);
nor U5484 (N_5484,N_3015,N_2604);
xor U5485 (N_5485,N_3664,N_4838);
xnor U5486 (N_5486,N_2994,N_4338);
nand U5487 (N_5487,N_4037,N_3686);
or U5488 (N_5488,N_2578,N_3707);
nor U5489 (N_5489,N_2825,N_2867);
nor U5490 (N_5490,N_4010,N_4416);
nor U5491 (N_5491,N_3954,N_2576);
or U5492 (N_5492,N_2877,N_2567);
nor U5493 (N_5493,N_3552,N_2608);
or U5494 (N_5494,N_4457,N_3780);
nand U5495 (N_5495,N_3297,N_3439);
or U5496 (N_5496,N_3666,N_3705);
and U5497 (N_5497,N_3270,N_3128);
nand U5498 (N_5498,N_2963,N_4592);
or U5499 (N_5499,N_2718,N_4007);
nor U5500 (N_5500,N_4435,N_3659);
or U5501 (N_5501,N_3112,N_3795);
and U5502 (N_5502,N_4125,N_4509);
or U5503 (N_5503,N_4428,N_4683);
and U5504 (N_5504,N_3068,N_4499);
or U5505 (N_5505,N_4661,N_4506);
nand U5506 (N_5506,N_2837,N_4021);
nand U5507 (N_5507,N_2848,N_3244);
or U5508 (N_5508,N_4654,N_3588);
nor U5509 (N_5509,N_3925,N_3980);
or U5510 (N_5510,N_4947,N_4999);
nor U5511 (N_5511,N_2518,N_2528);
or U5512 (N_5512,N_4467,N_2853);
or U5513 (N_5513,N_3032,N_4836);
nand U5514 (N_5514,N_4800,N_3409);
nor U5515 (N_5515,N_3211,N_3130);
xor U5516 (N_5516,N_4687,N_2517);
and U5517 (N_5517,N_2639,N_4726);
nand U5518 (N_5518,N_4913,N_4482);
and U5519 (N_5519,N_4167,N_2702);
nand U5520 (N_5520,N_3028,N_4864);
xor U5521 (N_5521,N_4586,N_4903);
and U5522 (N_5522,N_3586,N_3753);
or U5523 (N_5523,N_3648,N_3224);
and U5524 (N_5524,N_2806,N_4653);
nor U5525 (N_5525,N_2541,N_3463);
or U5526 (N_5526,N_4625,N_3597);
and U5527 (N_5527,N_3327,N_2667);
xnor U5528 (N_5528,N_3994,N_4545);
nand U5529 (N_5529,N_4050,N_3776);
or U5530 (N_5530,N_2698,N_2734);
xor U5531 (N_5531,N_3818,N_2595);
and U5532 (N_5532,N_2593,N_2996);
and U5533 (N_5533,N_3967,N_3668);
nand U5534 (N_5534,N_2916,N_2849);
or U5535 (N_5535,N_3238,N_4806);
or U5536 (N_5536,N_4266,N_3177);
nand U5537 (N_5537,N_2711,N_4372);
and U5538 (N_5538,N_2561,N_2544);
and U5539 (N_5539,N_4169,N_2688);
nor U5540 (N_5540,N_4137,N_4500);
or U5541 (N_5541,N_3078,N_4667);
xor U5542 (N_5542,N_3471,N_2701);
or U5543 (N_5543,N_2805,N_2795);
or U5544 (N_5544,N_4895,N_4757);
and U5545 (N_5545,N_3379,N_4813);
nand U5546 (N_5546,N_2713,N_3900);
and U5547 (N_5547,N_3141,N_3922);
and U5548 (N_5548,N_4317,N_2733);
nand U5549 (N_5549,N_3186,N_3660);
or U5550 (N_5550,N_3267,N_4979);
nand U5551 (N_5551,N_4438,N_4299);
nor U5552 (N_5552,N_4616,N_3473);
nor U5553 (N_5553,N_4287,N_2920);
nand U5554 (N_5554,N_3019,N_3696);
nor U5555 (N_5555,N_3757,N_4112);
and U5556 (N_5556,N_4175,N_3516);
or U5557 (N_5557,N_4311,N_4105);
or U5558 (N_5558,N_3695,N_3851);
and U5559 (N_5559,N_3236,N_3188);
nor U5560 (N_5560,N_4479,N_4179);
or U5561 (N_5561,N_4569,N_3911);
or U5562 (N_5562,N_3816,N_2606);
and U5563 (N_5563,N_4144,N_3513);
and U5564 (N_5564,N_2579,N_3050);
nor U5565 (N_5565,N_4495,N_3256);
xnor U5566 (N_5566,N_2829,N_3340);
and U5567 (N_5567,N_3031,N_4524);
and U5568 (N_5568,N_3559,N_3651);
or U5569 (N_5569,N_2504,N_4922);
or U5570 (N_5570,N_4001,N_4307);
nor U5571 (N_5571,N_4148,N_2941);
and U5572 (N_5572,N_4349,N_3014);
or U5573 (N_5573,N_3536,N_2635);
nand U5574 (N_5574,N_3067,N_4655);
nor U5575 (N_5575,N_4627,N_3320);
nor U5576 (N_5576,N_3539,N_3710);
nor U5577 (N_5577,N_3752,N_3234);
and U5578 (N_5578,N_4213,N_3842);
or U5579 (N_5579,N_3421,N_4851);
nand U5580 (N_5580,N_2768,N_4776);
nand U5581 (N_5581,N_3350,N_4839);
nand U5582 (N_5582,N_4974,N_3284);
and U5583 (N_5583,N_2814,N_3099);
nor U5584 (N_5584,N_3293,N_3362);
nor U5585 (N_5585,N_3653,N_4797);
and U5586 (N_5586,N_3578,N_2940);
or U5587 (N_5587,N_3461,N_3681);
nor U5588 (N_5588,N_4878,N_4894);
xnor U5589 (N_5589,N_2860,N_2772);
or U5590 (N_5590,N_3060,N_3608);
nand U5591 (N_5591,N_4724,N_4511);
and U5592 (N_5592,N_4768,N_3669);
nor U5593 (N_5593,N_4158,N_4591);
nand U5594 (N_5594,N_3046,N_2728);
xor U5595 (N_5595,N_4290,N_4323);
nor U5596 (N_5596,N_3819,N_3494);
xnor U5597 (N_5597,N_4674,N_2942);
nand U5598 (N_5598,N_4444,N_3735);
and U5599 (N_5599,N_4413,N_3811);
and U5600 (N_5600,N_4600,N_4388);
and U5601 (N_5601,N_4153,N_4095);
nand U5602 (N_5602,N_3945,N_2719);
and U5603 (N_5603,N_3632,N_4750);
and U5604 (N_5604,N_2683,N_4848);
nor U5605 (N_5605,N_4426,N_3323);
nor U5606 (N_5606,N_4077,N_3373);
and U5607 (N_5607,N_3326,N_3631);
and U5608 (N_5608,N_4821,N_4716);
nor U5609 (N_5609,N_4201,N_4816);
or U5610 (N_5610,N_4505,N_2556);
xor U5611 (N_5611,N_4795,N_3600);
and U5612 (N_5612,N_3827,N_3936);
nor U5613 (N_5613,N_3429,N_2630);
and U5614 (N_5614,N_3769,N_3393);
and U5615 (N_5615,N_4910,N_4659);
nor U5616 (N_5616,N_2809,N_4649);
xnor U5617 (N_5617,N_4252,N_4450);
nand U5618 (N_5618,N_2586,N_2689);
or U5619 (N_5619,N_4204,N_4755);
and U5620 (N_5620,N_3225,N_2764);
and U5621 (N_5621,N_2907,N_4970);
and U5622 (N_5622,N_3312,N_3508);
and U5623 (N_5623,N_3804,N_3576);
and U5624 (N_5624,N_4405,N_2665);
nor U5625 (N_5625,N_4454,N_3103);
xnor U5626 (N_5626,N_4070,N_4284);
or U5627 (N_5627,N_4058,N_3684);
nand U5628 (N_5628,N_4030,N_3091);
nor U5629 (N_5629,N_3269,N_3414);
and U5630 (N_5630,N_3570,N_3415);
and U5631 (N_5631,N_3504,N_4431);
nand U5632 (N_5632,N_2810,N_2744);
and U5633 (N_5633,N_2515,N_3714);
nor U5634 (N_5634,N_2858,N_3527);
nand U5635 (N_5635,N_4128,N_4318);
xnor U5636 (N_5636,N_2641,N_3395);
nand U5637 (N_5637,N_4270,N_4936);
nor U5638 (N_5638,N_3434,N_3122);
nand U5639 (N_5639,N_4353,N_3155);
or U5640 (N_5640,N_4127,N_3080);
or U5641 (N_5641,N_3420,N_4937);
nand U5642 (N_5642,N_2876,N_3661);
and U5643 (N_5643,N_3560,N_4329);
and U5644 (N_5644,N_4126,N_3285);
nor U5645 (N_5645,N_2715,N_2666);
nand U5646 (N_5646,N_2539,N_3767);
nor U5647 (N_5647,N_4409,N_4938);
or U5648 (N_5648,N_3178,N_2912);
nor U5649 (N_5649,N_4304,N_2525);
or U5650 (N_5650,N_4846,N_2953);
or U5651 (N_5651,N_3172,N_4376);
and U5652 (N_5652,N_2986,N_4739);
nand U5653 (N_5653,N_4235,N_3606);
or U5654 (N_5654,N_3724,N_3274);
or U5655 (N_5655,N_3042,N_3251);
nand U5656 (N_5656,N_3998,N_4019);
nand U5657 (N_5657,N_3634,N_3744);
nor U5658 (N_5658,N_3410,N_4577);
nor U5659 (N_5659,N_4024,N_3949);
or U5660 (N_5660,N_2952,N_3870);
and U5661 (N_5661,N_4356,N_4177);
nand U5662 (N_5662,N_4367,N_3905);
or U5663 (N_5663,N_4787,N_2721);
or U5664 (N_5664,N_3330,N_3531);
or U5665 (N_5665,N_3987,N_4840);
xor U5666 (N_5666,N_2514,N_4027);
nor U5667 (N_5667,N_3189,N_3416);
nor U5668 (N_5668,N_4066,N_4314);
xor U5669 (N_5669,N_4020,N_3435);
or U5670 (N_5670,N_2960,N_3580);
or U5671 (N_5671,N_3248,N_3709);
nand U5672 (N_5672,N_4090,N_3318);
and U5673 (N_5673,N_4550,N_3749);
or U5674 (N_5674,N_3133,N_4784);
and U5675 (N_5675,N_4676,N_4529);
nand U5676 (N_5676,N_4812,N_4502);
xor U5677 (N_5677,N_3179,N_3368);
nand U5678 (N_5678,N_4171,N_3406);
nor U5679 (N_5679,N_2581,N_4748);
nor U5680 (N_5680,N_2962,N_2716);
or U5681 (N_5681,N_3065,N_4617);
or U5682 (N_5682,N_3916,N_4559);
nor U5683 (N_5683,N_3649,N_4599);
nor U5684 (N_5684,N_4487,N_3557);
xnor U5685 (N_5685,N_4863,N_4831);
and U5686 (N_5686,N_4476,N_2939);
and U5687 (N_5687,N_4474,N_4514);
xnor U5688 (N_5688,N_2924,N_4966);
or U5689 (N_5689,N_4103,N_3745);
or U5690 (N_5690,N_4902,N_4786);
nor U5691 (N_5691,N_2859,N_2571);
xnor U5692 (N_5692,N_4389,N_4262);
or U5693 (N_5693,N_4277,N_4862);
nand U5694 (N_5694,N_2818,N_3228);
and U5695 (N_5695,N_3700,N_4135);
and U5696 (N_5696,N_4953,N_2970);
nor U5697 (N_5697,N_4385,N_3547);
nand U5698 (N_5698,N_4646,N_2976);
nor U5699 (N_5699,N_4461,N_4963);
nor U5700 (N_5700,N_4719,N_3044);
nor U5701 (N_5701,N_2575,N_3161);
nor U5702 (N_5702,N_4759,N_3930);
nand U5703 (N_5703,N_4700,N_4496);
nand U5704 (N_5704,N_3506,N_4956);
nand U5705 (N_5705,N_4736,N_3623);
or U5706 (N_5706,N_4107,N_2776);
nor U5707 (N_5707,N_2724,N_3971);
nor U5708 (N_5708,N_3793,N_3978);
nor U5709 (N_5709,N_2602,N_3039);
nand U5710 (N_5710,N_3382,N_4884);
or U5711 (N_5711,N_4350,N_2969);
or U5712 (N_5712,N_3374,N_3176);
nand U5713 (N_5713,N_3370,N_3775);
nor U5714 (N_5714,N_3969,N_2548);
nand U5715 (N_5715,N_4648,N_4652);
nand U5716 (N_5716,N_4769,N_4777);
nor U5717 (N_5717,N_3928,N_2800);
nand U5718 (N_5718,N_3277,N_4134);
and U5719 (N_5719,N_4877,N_4011);
or U5720 (N_5720,N_4796,N_3457);
or U5721 (N_5721,N_3262,N_4859);
nand U5722 (N_5722,N_3750,N_2793);
nand U5723 (N_5723,N_4805,N_3214);
and U5724 (N_5724,N_3650,N_4246);
xor U5725 (N_5725,N_2828,N_2961);
xnor U5726 (N_5726,N_2767,N_2664);
nor U5727 (N_5727,N_2625,N_3045);
xor U5728 (N_5728,N_4896,N_3071);
xor U5729 (N_5729,N_4225,N_3581);
or U5730 (N_5730,N_3537,N_4117);
and U5731 (N_5731,N_4415,N_3873);
nand U5732 (N_5732,N_3882,N_2695);
or U5733 (N_5733,N_4233,N_4065);
or U5734 (N_5734,N_4097,N_4205);
or U5735 (N_5735,N_2552,N_4566);
and U5736 (N_5736,N_4664,N_2903);
nor U5737 (N_5737,N_3765,N_3533);
nor U5738 (N_5738,N_2753,N_3891);
nand U5739 (N_5739,N_3023,N_4741);
nor U5740 (N_5740,N_3985,N_4489);
xnor U5741 (N_5741,N_4347,N_3367);
and U5742 (N_5742,N_2870,N_4395);
nand U5743 (N_5743,N_3126,N_3160);
nand U5744 (N_5744,N_4281,N_4185);
and U5745 (N_5745,N_2697,N_4762);
nand U5746 (N_5746,N_2612,N_3909);
and U5747 (N_5747,N_3591,N_3365);
and U5748 (N_5748,N_3456,N_4578);
nand U5749 (N_5749,N_3540,N_4916);
or U5750 (N_5750,N_4093,N_3198);
nand U5751 (N_5751,N_4184,N_3895);
or U5752 (N_5752,N_3530,N_3638);
nand U5753 (N_5753,N_4520,N_2882);
xor U5754 (N_5754,N_2864,N_4088);
nor U5755 (N_5755,N_3497,N_2554);
and U5756 (N_5756,N_2570,N_2785);
nor U5757 (N_5757,N_4906,N_3283);
xor U5758 (N_5758,N_3908,N_4503);
and U5759 (N_5759,N_4571,N_3164);
nor U5760 (N_5760,N_3790,N_4430);
or U5761 (N_5761,N_3369,N_3417);
and U5762 (N_5762,N_3107,N_4523);
nor U5763 (N_5763,N_2950,N_3976);
or U5764 (N_5764,N_3502,N_3864);
or U5765 (N_5765,N_2633,N_2919);
nor U5766 (N_5766,N_3610,N_3636);
nor U5767 (N_5767,N_4703,N_2610);
and U5768 (N_5768,N_3812,N_2674);
nor U5769 (N_5769,N_3975,N_3341);
and U5770 (N_5770,N_3759,N_4533);
nand U5771 (N_5771,N_3865,N_3841);
xnor U5772 (N_5772,N_4847,N_4897);
nor U5773 (N_5773,N_3637,N_4931);
nand U5774 (N_5774,N_3838,N_3135);
and U5775 (N_5775,N_3003,N_4289);
nor U5776 (N_5776,N_4934,N_2660);
nand U5777 (N_5777,N_2566,N_3685);
or U5778 (N_5778,N_3595,N_4046);
nor U5779 (N_5779,N_3831,N_4054);
nor U5780 (N_5780,N_3110,N_4692);
and U5781 (N_5781,N_4889,N_3599);
or U5782 (N_5782,N_2546,N_3230);
nor U5783 (N_5783,N_4142,N_3132);
nand U5784 (N_5784,N_4494,N_4579);
nor U5785 (N_5785,N_3871,N_4384);
or U5786 (N_5786,N_4151,N_3213);
nor U5787 (N_5787,N_2843,N_3241);
nand U5788 (N_5788,N_3029,N_4602);
xnor U5789 (N_5789,N_3718,N_4647);
nor U5790 (N_5790,N_2890,N_3706);
and U5791 (N_5791,N_3550,N_2643);
nand U5792 (N_5792,N_3472,N_2555);
nor U5793 (N_5793,N_2929,N_4987);
nor U5794 (N_5794,N_4015,N_4861);
nor U5795 (N_5795,N_4018,N_3073);
nor U5796 (N_5796,N_3296,N_4187);
or U5797 (N_5797,N_4669,N_4048);
nand U5798 (N_5798,N_3069,N_3294);
or U5799 (N_5799,N_3467,N_4918);
or U5800 (N_5800,N_4330,N_3542);
and U5801 (N_5801,N_2819,N_4452);
nor U5802 (N_5802,N_3904,N_3381);
and U5803 (N_5803,N_4621,N_2914);
or U5804 (N_5804,N_2911,N_3334);
nand U5805 (N_5805,N_4227,N_3047);
nor U5806 (N_5806,N_4303,N_3719);
or U5807 (N_5807,N_3972,N_4917);
nand U5808 (N_5808,N_3125,N_3662);
or U5809 (N_5809,N_4424,N_2722);
nand U5810 (N_5810,N_4809,N_3778);
nor U5811 (N_5811,N_3847,N_3784);
nand U5812 (N_5812,N_3673,N_2905);
and U5813 (N_5813,N_3910,N_4256);
xor U5814 (N_5814,N_3541,N_3355);
nor U5815 (N_5815,N_4344,N_4536);
or U5816 (N_5816,N_4294,N_2872);
or U5817 (N_5817,N_4089,N_4705);
nor U5818 (N_5818,N_3807,N_3946);
nand U5819 (N_5819,N_4773,N_4820);
or U5820 (N_5820,N_2935,N_3571);
nor U5821 (N_5821,N_2973,N_2928);
or U5822 (N_5822,N_3802,N_2758);
or U5823 (N_5823,N_2770,N_2791);
xnor U5824 (N_5824,N_2887,N_3594);
or U5825 (N_5825,N_4310,N_4793);
xnor U5826 (N_5826,N_4116,N_3883);
nor U5827 (N_5827,N_3680,N_3501);
or U5828 (N_5828,N_2925,N_2835);
nor U5829 (N_5829,N_3826,N_3037);
nand U5830 (N_5830,N_3144,N_4518);
or U5831 (N_5831,N_3085,N_4522);
or U5832 (N_5832,N_3748,N_2534);
or U5833 (N_5833,N_3934,N_3868);
or U5834 (N_5834,N_2759,N_4562);
nor U5835 (N_5835,N_4016,N_3762);
nand U5836 (N_5836,N_3222,N_3116);
or U5837 (N_5837,N_2789,N_4254);
and U5838 (N_5838,N_3596,N_3197);
nor U5839 (N_5839,N_4971,N_4432);
or U5840 (N_5840,N_4540,N_3313);
nand U5841 (N_5841,N_3275,N_4609);
nand U5842 (N_5842,N_4618,N_4580);
nor U5843 (N_5843,N_4315,N_4539);
nand U5844 (N_5844,N_4328,N_3805);
or U5845 (N_5845,N_4182,N_3281);
or U5846 (N_5846,N_4510,N_2777);
nand U5847 (N_5847,N_3052,N_4890);
or U5848 (N_5848,N_2655,N_4381);
and U5849 (N_5849,N_3062,N_4400);
xor U5850 (N_5850,N_3924,N_4275);
or U5851 (N_5851,N_3957,N_2866);
and U5852 (N_5852,N_4681,N_4818);
and U5853 (N_5853,N_2736,N_2741);
nor U5854 (N_5854,N_4727,N_3973);
nor U5855 (N_5855,N_2901,N_2549);
nor U5856 (N_5856,N_2958,N_3357);
nor U5857 (N_5857,N_4239,N_4558);
xor U5858 (N_5858,N_3947,N_4108);
xor U5859 (N_5859,N_3250,N_3053);
xnor U5860 (N_5860,N_4525,N_3691);
nor U5861 (N_5861,N_3622,N_2841);
nand U5862 (N_5862,N_3773,N_4129);
and U5863 (N_5863,N_4734,N_4972);
nand U5864 (N_5864,N_3092,N_3148);
nand U5865 (N_5865,N_4998,N_3205);
nor U5866 (N_5866,N_4556,N_3555);
and U5867 (N_5867,N_2813,N_4710);
xor U5868 (N_5868,N_4733,N_3830);
and U5869 (N_5869,N_2596,N_2542);
nand U5870 (N_5870,N_3102,N_3411);
nand U5871 (N_5871,N_2765,N_3077);
nand U5872 (N_5872,N_4955,N_4901);
nand U5873 (N_5873,N_4855,N_3428);
xnor U5874 (N_5874,N_3510,N_3496);
or U5875 (N_5875,N_2682,N_4825);
and U5876 (N_5876,N_2615,N_3743);
or U5877 (N_5877,N_3903,N_4983);
nand U5878 (N_5878,N_2657,N_3146);
xor U5879 (N_5879,N_3822,N_3389);
or U5880 (N_5880,N_2752,N_3995);
xor U5881 (N_5881,N_3385,N_4698);
and U5882 (N_5882,N_2621,N_3792);
nor U5883 (N_5883,N_3470,N_2686);
nand U5884 (N_5884,N_4206,N_4783);
xor U5885 (N_5885,N_3820,N_4868);
or U5886 (N_5886,N_3728,N_4365);
or U5887 (N_5887,N_4096,N_3605);
or U5888 (N_5888,N_2880,N_3627);
nor U5889 (N_5889,N_4534,N_2796);
and U5890 (N_5890,N_3448,N_4041);
and U5891 (N_5891,N_3136,N_3219);
or U5892 (N_5892,N_2645,N_3246);
nor U5893 (N_5893,N_3654,N_4573);
nand U5894 (N_5894,N_2990,N_3167);
and U5895 (N_5895,N_3476,N_3445);
and U5896 (N_5896,N_4690,N_3703);
or U5897 (N_5897,N_3888,N_4194);
and U5898 (N_5898,N_4243,N_4560);
nor U5899 (N_5899,N_4722,N_3150);
nor U5900 (N_5900,N_4572,N_3212);
nand U5901 (N_5901,N_4866,N_4193);
or U5902 (N_5902,N_4778,N_4553);
nand U5903 (N_5903,N_2964,N_4823);
and U5904 (N_5904,N_3779,N_3716);
and U5905 (N_5905,N_2951,N_4133);
xor U5906 (N_5906,N_3593,N_4420);
or U5907 (N_5907,N_2927,N_2799);
and U5908 (N_5908,N_3157,N_3532);
nand U5909 (N_5909,N_3233,N_4443);
and U5910 (N_5910,N_4145,N_3074);
or U5911 (N_5911,N_4909,N_2892);
or U5912 (N_5912,N_2652,N_4770);
and U5913 (N_5913,N_4492,N_4429);
and U5914 (N_5914,N_4119,N_4369);
nor U5915 (N_5915,N_3708,N_2891);
and U5916 (N_5916,N_4672,N_2580);
nand U5917 (N_5917,N_3566,N_4223);
nor U5918 (N_5918,N_4497,N_2650);
xor U5919 (N_5919,N_4869,N_3298);
or U5920 (N_5920,N_3147,N_4541);
or U5921 (N_5921,N_4189,N_3242);
and U5922 (N_5922,N_4686,N_4738);
nand U5923 (N_5923,N_4582,N_3220);
nor U5924 (N_5924,N_4408,N_3452);
xnor U5925 (N_5925,N_3509,N_4581);
or U5926 (N_5926,N_4740,N_4082);
and U5927 (N_5927,N_4774,N_4029);
nor U5928 (N_5928,N_4721,N_2896);
nor U5929 (N_5929,N_4118,N_3499);
nand U5930 (N_5930,N_3354,N_4269);
and U5931 (N_5931,N_2523,N_2862);
xor U5932 (N_5932,N_3072,N_3372);
and U5933 (N_5933,N_4673,N_2998);
nor U5934 (N_5934,N_3835,N_4919);
nand U5935 (N_5935,N_3291,N_3898);
nand U5936 (N_5936,N_2692,N_3359);
nor U5937 (N_5937,N_2687,N_3970);
nand U5938 (N_5938,N_3070,N_4110);
nand U5939 (N_5939,N_2707,N_4850);
and U5940 (N_5940,N_3856,N_3783);
nor U5941 (N_5941,N_3896,N_4798);
nand U5942 (N_5942,N_3777,N_2910);
nand U5943 (N_5943,N_2588,N_4071);
xor U5944 (N_5944,N_2598,N_4045);
or U5945 (N_5945,N_4900,N_2649);
xnor U5946 (N_5946,N_3493,N_3879);
and U5947 (N_5947,N_2757,N_4297);
xor U5948 (N_5948,N_2978,N_3966);
nor U5949 (N_5949,N_4296,N_3051);
nand U5950 (N_5950,N_3088,N_2653);
and U5951 (N_5951,N_4433,N_2624);
nor U5952 (N_5952,N_4360,N_2671);
nand U5953 (N_5953,N_4439,N_2985);
and U5954 (N_5954,N_2708,N_4188);
nand U5955 (N_5955,N_3240,N_3035);
nor U5956 (N_5956,N_3845,N_3027);
or U5957 (N_5957,N_3252,N_3139);
or U5958 (N_5958,N_3034,N_4904);
or U5959 (N_5959,N_4437,N_4422);
or U5960 (N_5960,N_2543,N_4984);
xor U5961 (N_5961,N_3237,N_4613);
and U5962 (N_5962,N_2991,N_2821);
or U5963 (N_5963,N_2954,N_3465);
or U5964 (N_5964,N_3254,N_3950);
nor U5965 (N_5965,N_3446,N_3624);
nand U5966 (N_5966,N_2592,N_3007);
nand U5967 (N_5967,N_3738,N_4102);
nand U5968 (N_5968,N_4472,N_3598);
nor U5969 (N_5969,N_2547,N_2638);
nand U5970 (N_5970,N_3449,N_3733);
nor U5971 (N_5971,N_2815,N_2997);
nand U5972 (N_5972,N_3808,N_3436);
nor U5973 (N_5973,N_4292,N_2562);
or U5974 (N_5974,N_4469,N_3711);
or U5975 (N_5975,N_4136,N_3083);
or U5976 (N_5976,N_3402,N_4542);
or U5977 (N_5977,N_4932,N_2620);
and U5978 (N_5978,N_4837,N_3788);
or U5979 (N_5979,N_3418,N_4968);
xor U5980 (N_5980,N_3118,N_3430);
and U5981 (N_5981,N_3396,N_2956);
or U5982 (N_5982,N_2646,N_3345);
and U5983 (N_5983,N_4656,N_4032);
or U5984 (N_5984,N_3302,N_4083);
and U5985 (N_5985,N_3751,N_3862);
or U5986 (N_5986,N_3849,N_3715);
nand U5987 (N_5987,N_3253,N_4753);
and U5988 (N_5988,N_2524,N_3114);
or U5989 (N_5989,N_4708,N_4008);
xnor U5990 (N_5990,N_3268,N_3642);
or U5991 (N_5991,N_4298,N_4337);
nor U5992 (N_5992,N_4217,N_3363);
nand U5993 (N_5993,N_4170,N_3187);
nor U5994 (N_5994,N_3602,N_3093);
xor U5995 (N_5995,N_4043,N_3308);
and U5996 (N_5996,N_4212,N_3993);
nand U5997 (N_5997,N_4081,N_4691);
or U5998 (N_5998,N_3786,N_4808);
nor U5999 (N_5999,N_4612,N_3678);
and U6000 (N_6000,N_2881,N_3413);
or U6001 (N_6001,N_3346,N_4882);
nand U6002 (N_6002,N_3048,N_3247);
or U6003 (N_6003,N_4218,N_4881);
nor U6004 (N_6004,N_3299,N_4543);
and U6005 (N_6005,N_3821,N_4555);
or U6006 (N_6006,N_2802,N_3850);
and U6007 (N_6007,N_2797,N_4361);
or U6008 (N_6008,N_3787,N_3054);
and U6009 (N_6009,N_3958,N_4306);
nor U6010 (N_6010,N_2854,N_3933);
or U6011 (N_6011,N_4241,N_4597);
or U6012 (N_6012,N_4231,N_2863);
nor U6013 (N_6013,N_3858,N_4274);
nand U6014 (N_6014,N_3377,N_3149);
or U6015 (N_6015,N_2532,N_3423);
or U6016 (N_6016,N_2992,N_2628);
nor U6017 (N_6017,N_3799,N_4057);
nand U6018 (N_6018,N_2601,N_4575);
nor U6019 (N_6019,N_3617,N_4779);
or U6020 (N_6020,N_3688,N_3043);
nand U6021 (N_6021,N_4718,N_4879);
nor U6022 (N_6022,N_4073,N_4259);
nor U6023 (N_6023,N_3180,N_4341);
nor U6024 (N_6024,N_3567,N_2537);
and U6025 (N_6025,N_4196,N_4440);
nand U6026 (N_6026,N_3117,N_4370);
xnor U6027 (N_6027,N_3475,N_2607);
or U6028 (N_6028,N_3433,N_3583);
and U6029 (N_6029,N_2787,N_3426);
and U6030 (N_6030,N_2503,N_4326);
and U6031 (N_6031,N_3442,N_3986);
and U6032 (N_6032,N_3453,N_4053);
xnor U6033 (N_6033,N_3412,N_4078);
nand U6034 (N_6034,N_4031,N_4830);
nand U6035 (N_6035,N_3863,N_3194);
and U6036 (N_6036,N_2626,N_4563);
and U6037 (N_6037,N_4152,N_4207);
or U6038 (N_6038,N_3468,N_4293);
nor U6039 (N_6039,N_4528,N_3534);
nor U6040 (N_6040,N_3366,N_4143);
xnor U6041 (N_6041,N_3754,N_4005);
and U6042 (N_6042,N_3017,N_2868);
or U6043 (N_6043,N_4954,N_4565);
and U6044 (N_6044,N_4319,N_2603);
nand U6045 (N_6045,N_3725,N_3755);
nor U6046 (N_6046,N_4679,N_2943);
and U6047 (N_6047,N_4763,N_2995);
nand U6048 (N_6048,N_3644,N_4688);
or U6049 (N_6049,N_2732,N_3582);
xor U6050 (N_6050,N_3901,N_2968);
xor U6051 (N_6051,N_2551,N_2982);
and U6052 (N_6052,N_3443,N_4852);
or U6053 (N_6053,N_4914,N_4794);
nor U6054 (N_6054,N_4463,N_4975);
and U6055 (N_6055,N_3704,N_3834);
nand U6056 (N_6056,N_4488,N_3432);
nor U6057 (N_6057,N_4300,N_3932);
or U6058 (N_6058,N_4758,N_2729);
nand U6059 (N_6059,N_4807,N_3055);
or U6060 (N_6060,N_2533,N_4752);
and U6061 (N_6061,N_3337,N_3645);
or U6062 (N_6062,N_4493,N_2774);
xnor U6063 (N_6063,N_3931,N_2519);
or U6064 (N_6064,N_4604,N_2536);
or U6065 (N_6065,N_3477,N_2560);
nor U6066 (N_6066,N_4017,N_4731);
nor U6067 (N_6067,N_4288,N_3741);
or U6068 (N_6068,N_4382,N_4744);
and U6069 (N_6069,N_3927,N_4715);
xor U6070 (N_6070,N_4946,N_3646);
nor U6071 (N_6071,N_3630,N_3772);
and U6072 (N_6072,N_4680,N_3190);
nor U6073 (N_6073,N_4359,N_3774);
and U6074 (N_6074,N_3941,N_4210);
nand U6075 (N_6075,N_3621,N_3111);
xor U6076 (N_6076,N_4320,N_3329);
or U6077 (N_6077,N_4827,N_4622);
nor U6078 (N_6078,N_4109,N_3344);
nand U6079 (N_6079,N_4941,N_3152);
nor U6080 (N_6080,N_4026,N_4166);
or U6081 (N_6081,N_3460,N_2597);
nand U6082 (N_6082,N_4305,N_2540);
nor U6083 (N_6083,N_4100,N_4746);
or U6084 (N_6084,N_3881,N_3024);
and U6085 (N_6085,N_3038,N_4216);
nor U6086 (N_6086,N_2921,N_3977);
or U6087 (N_6087,N_3485,N_2987);
or U6088 (N_6088,N_3170,N_3101);
or U6089 (N_6089,N_4079,N_4115);
and U6090 (N_6090,N_3525,N_3158);
and U6091 (N_6091,N_4713,N_3761);
and U6092 (N_6092,N_3951,N_3549);
nand U6093 (N_6093,N_3066,N_4321);
and U6094 (N_6094,N_4159,N_4483);
nor U6095 (N_6095,N_3543,N_3090);
or U6096 (N_6096,N_2838,N_4993);
xnor U6097 (N_6097,N_4782,N_4358);
nand U6098 (N_6098,N_2617,N_4615);
or U6099 (N_6099,N_2672,N_4155);
nor U6100 (N_6100,N_2558,N_3175);
and U6101 (N_6101,N_4004,N_4333);
or U6102 (N_6102,N_4121,N_4265);
nor U6103 (N_6103,N_3094,N_4817);
and U6104 (N_6104,N_3713,N_3948);
or U6105 (N_6105,N_3731,N_3763);
nor U6106 (N_6106,N_4929,N_4976);
and U6107 (N_6107,N_3515,N_4412);
or U6108 (N_6108,N_4036,N_4665);
or U6109 (N_6109,N_3572,N_3151);
nand U6110 (N_6110,N_4624,N_2590);
and U6111 (N_6111,N_4515,N_2714);
nand U6112 (N_6112,N_3295,N_3353);
xnor U6113 (N_6113,N_4952,N_3846);
xnor U6114 (N_6114,N_3348,N_2771);
and U6115 (N_6115,N_4997,N_3852);
nor U6116 (N_6116,N_3076,N_3264);
nand U6117 (N_6117,N_4336,N_2587);
and U6118 (N_6118,N_3440,N_3203);
nand U6119 (N_6119,N_3770,N_2661);
nand U6120 (N_6120,N_3553,N_2693);
nor U6121 (N_6121,N_3184,N_4804);
or U6122 (N_6122,N_3824,N_2690);
nor U6123 (N_6123,N_4780,N_3897);
or U6124 (N_6124,N_3939,N_3965);
nor U6125 (N_6125,N_2699,N_3154);
nand U6126 (N_6126,N_3202,N_4366);
and U6127 (N_6127,N_3984,N_2740);
nor U6128 (N_6128,N_2908,N_3162);
nor U6129 (N_6129,N_2675,N_4025);
nor U6130 (N_6130,N_4309,N_3614);
and U6131 (N_6131,N_3797,N_4260);
nor U6132 (N_6132,N_3855,N_3258);
xnor U6133 (N_6133,N_3280,N_4192);
nor U6134 (N_6134,N_3519,N_3612);
and U6135 (N_6135,N_4466,N_3874);
xor U6136 (N_6136,N_3145,N_2833);
nand U6137 (N_6137,N_3018,N_2565);
nand U6138 (N_6138,N_4723,N_3526);
xor U6139 (N_6139,N_4258,N_2888);
or U6140 (N_6140,N_4860,N_2677);
or U6141 (N_6141,N_4172,N_3517);
and U6142 (N_6142,N_4639,N_2933);
nor U6143 (N_6143,N_2784,N_4675);
xnor U6144 (N_6144,N_2845,N_4257);
and U6145 (N_6145,N_3315,N_3260);
and U6146 (N_6146,N_2883,N_2516);
and U6147 (N_6147,N_4075,N_3041);
nand U6148 (N_6148,N_4607,N_4449);
nor U6149 (N_6149,N_3813,N_4445);
nand U6150 (N_6150,N_3655,N_4637);
nor U6151 (N_6151,N_2899,N_4267);
or U6152 (N_6152,N_3255,N_4811);
nand U6153 (N_6153,N_3235,N_2755);
or U6154 (N_6154,N_3483,N_2726);
xor U6155 (N_6155,N_3459,N_3279);
nand U6156 (N_6156,N_3009,N_3388);
nand U6157 (N_6157,N_4950,N_3730);
or U6158 (N_6158,N_4312,N_4696);
nand U6159 (N_6159,N_4286,N_3249);
and U6160 (N_6160,N_2898,N_3999);
nor U6161 (N_6161,N_4442,N_2589);
nor U6162 (N_6162,N_3063,N_2557);
nor U6163 (N_6163,N_2659,N_3166);
nor U6164 (N_6164,N_4760,N_3259);
xnor U6165 (N_6165,N_4583,N_4957);
nor U6166 (N_6166,N_3437,N_4251);
nand U6167 (N_6167,N_2509,N_3059);
nand U6168 (N_6168,N_2989,N_4973);
nor U6169 (N_6169,N_4000,N_4355);
nand U6170 (N_6170,N_3335,N_3794);
or U6171 (N_6171,N_4074,N_4501);
or U6172 (N_6172,N_2936,N_4584);
xor U6173 (N_6173,N_3361,N_3917);
nand U6174 (N_6174,N_3221,N_4717);
nand U6175 (N_6175,N_4374,N_3057);
xnor U6176 (N_6176,N_4802,N_2807);
or U6177 (N_6177,N_2788,N_4002);
nor U6178 (N_6178,N_4276,N_4462);
and U6179 (N_6179,N_3836,N_3953);
and U6180 (N_6180,N_2640,N_2623);
and U6181 (N_6181,N_4064,N_4789);
or U6182 (N_6182,N_2983,N_2812);
xnor U6183 (N_6183,N_2611,N_3926);
nand U6184 (N_6184,N_3120,N_3558);
nand U6185 (N_6185,N_4915,N_3257);
or U6186 (N_6186,N_3278,N_3671);
nand U6187 (N_6187,N_3338,N_4397);
or U6188 (N_6188,N_3000,N_4091);
and U6189 (N_6189,N_4268,N_2847);
or U6190 (N_6190,N_4885,N_2957);
and U6191 (N_6191,N_3486,N_3828);
and U6192 (N_6192,N_4394,N_4610);
and U6193 (N_6193,N_3289,N_3568);
or U6194 (N_6194,N_4203,N_4644);
nor U6195 (N_6195,N_4843,N_4458);
nor U6196 (N_6196,N_3942,N_3940);
xor U6197 (N_6197,N_4327,N_4156);
nand U6198 (N_6198,N_3698,N_2510);
and U6199 (N_6199,N_4198,N_3021);
and U6200 (N_6200,N_3859,N_4636);
and U6201 (N_6201,N_4634,N_2906);
nor U6202 (N_6202,N_3886,N_4113);
nor U6203 (N_6203,N_2709,N_4623);
xnor U6204 (N_6204,N_2703,N_3914);
or U6205 (N_6205,N_4190,N_4702);
or U6206 (N_6206,N_2585,N_3022);
xor U6207 (N_6207,N_4876,N_4849);
nand U6208 (N_6208,N_4465,N_4606);
or U6209 (N_6209,N_4893,N_3832);
nor U6210 (N_6210,N_4211,N_3546);
nand U6211 (N_6211,N_4149,N_3844);
nor U6212 (N_6212,N_3134,N_4123);
nand U6213 (N_6213,N_3722,N_3974);
nand U6214 (N_6214,N_3156,N_4009);
and U6215 (N_6215,N_4930,N_3944);
xor U6216 (N_6216,N_3587,N_4343);
or U6217 (N_6217,N_3325,N_4380);
or U6218 (N_6218,N_4507,N_4986);
nor U6219 (N_6219,N_3482,N_4978);
nand U6220 (N_6220,N_2574,N_2739);
nand U6221 (N_6221,N_3665,N_2749);
or U6222 (N_6222,N_3404,N_2993);
and U6223 (N_6223,N_4662,N_2979);
nor U6224 (N_6224,N_4640,N_2679);
nor U6225 (N_6225,N_4220,N_2622);
or U6226 (N_6226,N_4130,N_3758);
xnor U6227 (N_6227,N_4417,N_3675);
xnor U6228 (N_6228,N_4200,N_4658);
nor U6229 (N_6229,N_2980,N_3106);
nor U6230 (N_6230,N_4730,N_3191);
nor U6231 (N_6231,N_2977,N_3956);
or U6232 (N_6232,N_4977,N_3603);
xnor U6233 (N_6233,N_4163,N_3590);
or U6234 (N_6234,N_4508,N_2583);
and U6235 (N_6235,N_4854,N_3723);
xnor U6236 (N_6236,N_4842,N_3697);
xor U6237 (N_6237,N_3861,N_3201);
or U6238 (N_6238,N_2501,N_4737);
nand U6239 (N_6239,N_3929,N_3545);
nor U6240 (N_6240,N_3613,N_2614);
and U6241 (N_6241,N_3676,N_3575);
or U6242 (N_6242,N_4150,N_3609);
nand U6243 (N_6243,N_4322,N_4587);
or U6244 (N_6244,N_4670,N_3689);
nor U6245 (N_6245,N_3806,N_3962);
and U6246 (N_6246,N_2637,N_4985);
nor U6247 (N_6247,N_3008,N_4588);
and U6248 (N_6248,N_2889,N_3464);
and U6249 (N_6249,N_3210,N_2823);
nand U6250 (N_6250,N_3022,N_3929);
and U6251 (N_6251,N_3946,N_4808);
and U6252 (N_6252,N_4545,N_3739);
and U6253 (N_6253,N_3896,N_4594);
or U6254 (N_6254,N_4947,N_3396);
xor U6255 (N_6255,N_4731,N_3754);
nor U6256 (N_6256,N_3825,N_4120);
xor U6257 (N_6257,N_2864,N_2924);
nand U6258 (N_6258,N_3353,N_3589);
and U6259 (N_6259,N_4761,N_4236);
nor U6260 (N_6260,N_3413,N_2678);
and U6261 (N_6261,N_3023,N_2973);
and U6262 (N_6262,N_4775,N_4291);
and U6263 (N_6263,N_3795,N_3126);
and U6264 (N_6264,N_2835,N_3775);
and U6265 (N_6265,N_4546,N_4046);
or U6266 (N_6266,N_4166,N_3800);
or U6267 (N_6267,N_2749,N_4780);
nand U6268 (N_6268,N_3848,N_3639);
or U6269 (N_6269,N_4673,N_3582);
or U6270 (N_6270,N_4673,N_3789);
and U6271 (N_6271,N_4731,N_4970);
nor U6272 (N_6272,N_3555,N_4329);
nor U6273 (N_6273,N_3313,N_3314);
or U6274 (N_6274,N_2717,N_3317);
and U6275 (N_6275,N_3103,N_3955);
nand U6276 (N_6276,N_2815,N_3523);
or U6277 (N_6277,N_4265,N_4321);
nand U6278 (N_6278,N_4262,N_3263);
or U6279 (N_6279,N_3506,N_4911);
and U6280 (N_6280,N_3384,N_2746);
and U6281 (N_6281,N_2776,N_2639);
nand U6282 (N_6282,N_3004,N_4772);
xor U6283 (N_6283,N_3706,N_2543);
nand U6284 (N_6284,N_3449,N_3609);
nand U6285 (N_6285,N_3511,N_3672);
and U6286 (N_6286,N_4317,N_4685);
and U6287 (N_6287,N_3567,N_3332);
or U6288 (N_6288,N_3778,N_2907);
and U6289 (N_6289,N_4274,N_2998);
or U6290 (N_6290,N_4892,N_4082);
nor U6291 (N_6291,N_3603,N_2949);
and U6292 (N_6292,N_3646,N_4456);
or U6293 (N_6293,N_3923,N_3593);
nor U6294 (N_6294,N_3010,N_4044);
nor U6295 (N_6295,N_3701,N_2580);
or U6296 (N_6296,N_2986,N_4219);
or U6297 (N_6297,N_2642,N_4922);
nand U6298 (N_6298,N_4382,N_3701);
or U6299 (N_6299,N_3310,N_3380);
or U6300 (N_6300,N_3153,N_4685);
or U6301 (N_6301,N_2946,N_4766);
nand U6302 (N_6302,N_4730,N_3557);
xnor U6303 (N_6303,N_4405,N_4128);
nand U6304 (N_6304,N_4464,N_4276);
nor U6305 (N_6305,N_3862,N_4167);
nor U6306 (N_6306,N_4912,N_4781);
xnor U6307 (N_6307,N_2543,N_4706);
and U6308 (N_6308,N_3409,N_4011);
nand U6309 (N_6309,N_3752,N_3691);
nor U6310 (N_6310,N_4240,N_2627);
nand U6311 (N_6311,N_4771,N_4370);
nor U6312 (N_6312,N_3804,N_3614);
xor U6313 (N_6313,N_4643,N_2642);
nor U6314 (N_6314,N_2704,N_3419);
and U6315 (N_6315,N_4017,N_4849);
and U6316 (N_6316,N_4053,N_3494);
nand U6317 (N_6317,N_3749,N_3368);
and U6318 (N_6318,N_3288,N_3629);
nor U6319 (N_6319,N_4850,N_3337);
nand U6320 (N_6320,N_2661,N_2937);
xor U6321 (N_6321,N_4902,N_4839);
nor U6322 (N_6322,N_3106,N_2804);
nor U6323 (N_6323,N_2949,N_4901);
nor U6324 (N_6324,N_3738,N_4519);
nand U6325 (N_6325,N_3238,N_4408);
nand U6326 (N_6326,N_3962,N_4157);
or U6327 (N_6327,N_2896,N_3822);
nor U6328 (N_6328,N_4272,N_4901);
xor U6329 (N_6329,N_3486,N_2995);
and U6330 (N_6330,N_3578,N_4918);
nand U6331 (N_6331,N_4657,N_2675);
nor U6332 (N_6332,N_3578,N_3825);
and U6333 (N_6333,N_2883,N_3467);
or U6334 (N_6334,N_4736,N_4391);
nor U6335 (N_6335,N_2940,N_3693);
xnor U6336 (N_6336,N_4865,N_2707);
or U6337 (N_6337,N_4682,N_3290);
nor U6338 (N_6338,N_2891,N_4349);
nor U6339 (N_6339,N_3917,N_2957);
nor U6340 (N_6340,N_2542,N_2995);
nor U6341 (N_6341,N_2998,N_3213);
and U6342 (N_6342,N_4617,N_3510);
nor U6343 (N_6343,N_4838,N_4325);
and U6344 (N_6344,N_2583,N_2714);
or U6345 (N_6345,N_2545,N_3908);
or U6346 (N_6346,N_3045,N_2799);
nor U6347 (N_6347,N_3932,N_3174);
nand U6348 (N_6348,N_2785,N_4804);
nor U6349 (N_6349,N_3726,N_2962);
or U6350 (N_6350,N_2841,N_4714);
or U6351 (N_6351,N_3038,N_4638);
or U6352 (N_6352,N_4115,N_3530);
xnor U6353 (N_6353,N_2568,N_4436);
and U6354 (N_6354,N_4841,N_2943);
and U6355 (N_6355,N_4269,N_3353);
nand U6356 (N_6356,N_3305,N_4375);
or U6357 (N_6357,N_3314,N_4479);
nor U6358 (N_6358,N_3771,N_4571);
or U6359 (N_6359,N_4081,N_4667);
or U6360 (N_6360,N_4244,N_4027);
nor U6361 (N_6361,N_2686,N_4523);
nor U6362 (N_6362,N_2624,N_4233);
nor U6363 (N_6363,N_3763,N_3724);
and U6364 (N_6364,N_3161,N_4767);
xnor U6365 (N_6365,N_4459,N_4935);
xor U6366 (N_6366,N_4677,N_4752);
or U6367 (N_6367,N_2961,N_2922);
or U6368 (N_6368,N_4714,N_3322);
nor U6369 (N_6369,N_3981,N_2595);
or U6370 (N_6370,N_3128,N_3557);
nor U6371 (N_6371,N_3887,N_4603);
nor U6372 (N_6372,N_3607,N_3798);
or U6373 (N_6373,N_4872,N_3724);
and U6374 (N_6374,N_3224,N_3584);
nor U6375 (N_6375,N_4448,N_3936);
nand U6376 (N_6376,N_3765,N_4069);
nor U6377 (N_6377,N_4516,N_3057);
nand U6378 (N_6378,N_2847,N_3547);
nand U6379 (N_6379,N_3009,N_3442);
and U6380 (N_6380,N_3929,N_4188);
nand U6381 (N_6381,N_3182,N_3896);
and U6382 (N_6382,N_2596,N_2769);
nand U6383 (N_6383,N_4867,N_2861);
or U6384 (N_6384,N_4019,N_4584);
nand U6385 (N_6385,N_2535,N_4266);
and U6386 (N_6386,N_3075,N_2510);
or U6387 (N_6387,N_3160,N_4295);
or U6388 (N_6388,N_3463,N_3609);
and U6389 (N_6389,N_4032,N_3906);
and U6390 (N_6390,N_4318,N_4172);
nand U6391 (N_6391,N_4421,N_2592);
or U6392 (N_6392,N_2766,N_3495);
xor U6393 (N_6393,N_4712,N_2817);
or U6394 (N_6394,N_2955,N_4221);
nand U6395 (N_6395,N_3711,N_4763);
and U6396 (N_6396,N_2651,N_2566);
xor U6397 (N_6397,N_3534,N_4135);
nor U6398 (N_6398,N_2933,N_2757);
nor U6399 (N_6399,N_4627,N_2977);
nand U6400 (N_6400,N_3869,N_2994);
or U6401 (N_6401,N_4389,N_4155);
nor U6402 (N_6402,N_4810,N_3967);
or U6403 (N_6403,N_2769,N_4726);
nand U6404 (N_6404,N_3866,N_4839);
nand U6405 (N_6405,N_3080,N_3621);
nand U6406 (N_6406,N_2971,N_2547);
and U6407 (N_6407,N_4734,N_4301);
or U6408 (N_6408,N_3260,N_4988);
nand U6409 (N_6409,N_2667,N_4552);
or U6410 (N_6410,N_4826,N_2698);
xor U6411 (N_6411,N_2771,N_4696);
nand U6412 (N_6412,N_4789,N_3580);
nor U6413 (N_6413,N_3014,N_3559);
and U6414 (N_6414,N_4121,N_4286);
and U6415 (N_6415,N_4302,N_2876);
or U6416 (N_6416,N_2721,N_4032);
nand U6417 (N_6417,N_3351,N_3850);
or U6418 (N_6418,N_2948,N_4152);
nor U6419 (N_6419,N_3570,N_2776);
and U6420 (N_6420,N_2942,N_4461);
nor U6421 (N_6421,N_4414,N_3457);
or U6422 (N_6422,N_4500,N_3224);
nand U6423 (N_6423,N_3618,N_3342);
nand U6424 (N_6424,N_3058,N_3136);
and U6425 (N_6425,N_2505,N_3795);
and U6426 (N_6426,N_3603,N_3295);
nor U6427 (N_6427,N_3658,N_4578);
or U6428 (N_6428,N_2679,N_4495);
nand U6429 (N_6429,N_4890,N_4619);
nor U6430 (N_6430,N_4900,N_3117);
nand U6431 (N_6431,N_3241,N_3779);
and U6432 (N_6432,N_3279,N_4395);
nor U6433 (N_6433,N_3570,N_4425);
and U6434 (N_6434,N_3459,N_3125);
nand U6435 (N_6435,N_4163,N_4603);
xnor U6436 (N_6436,N_3852,N_2823);
or U6437 (N_6437,N_4066,N_2517);
or U6438 (N_6438,N_3362,N_3739);
nor U6439 (N_6439,N_4308,N_4008);
nor U6440 (N_6440,N_4232,N_4993);
or U6441 (N_6441,N_4778,N_4918);
and U6442 (N_6442,N_2565,N_3727);
or U6443 (N_6443,N_2663,N_2748);
nor U6444 (N_6444,N_2706,N_2833);
nand U6445 (N_6445,N_4792,N_3989);
and U6446 (N_6446,N_3858,N_3392);
and U6447 (N_6447,N_3489,N_4165);
and U6448 (N_6448,N_3492,N_3262);
and U6449 (N_6449,N_2786,N_4864);
and U6450 (N_6450,N_4172,N_4459);
or U6451 (N_6451,N_3179,N_4197);
nand U6452 (N_6452,N_4123,N_2726);
nor U6453 (N_6453,N_3844,N_3644);
and U6454 (N_6454,N_2661,N_2708);
and U6455 (N_6455,N_4101,N_4965);
and U6456 (N_6456,N_2903,N_4135);
or U6457 (N_6457,N_4836,N_2626);
or U6458 (N_6458,N_3328,N_3925);
nor U6459 (N_6459,N_4367,N_4430);
nand U6460 (N_6460,N_4745,N_4895);
and U6461 (N_6461,N_3302,N_4232);
xor U6462 (N_6462,N_3033,N_2586);
nor U6463 (N_6463,N_4043,N_3938);
and U6464 (N_6464,N_3602,N_2931);
or U6465 (N_6465,N_3919,N_4798);
nand U6466 (N_6466,N_2931,N_4267);
nand U6467 (N_6467,N_3760,N_3490);
or U6468 (N_6468,N_2981,N_2755);
or U6469 (N_6469,N_2502,N_4578);
and U6470 (N_6470,N_4225,N_3646);
nand U6471 (N_6471,N_3943,N_3155);
or U6472 (N_6472,N_4456,N_3357);
xor U6473 (N_6473,N_2521,N_3204);
nor U6474 (N_6474,N_3023,N_2597);
nand U6475 (N_6475,N_2588,N_2717);
or U6476 (N_6476,N_4643,N_2675);
nor U6477 (N_6477,N_4864,N_4254);
xnor U6478 (N_6478,N_4411,N_3527);
nor U6479 (N_6479,N_4954,N_2510);
nand U6480 (N_6480,N_3848,N_2775);
xnor U6481 (N_6481,N_4903,N_3171);
nor U6482 (N_6482,N_3174,N_4985);
nor U6483 (N_6483,N_3244,N_3401);
or U6484 (N_6484,N_3634,N_3559);
or U6485 (N_6485,N_2966,N_2542);
or U6486 (N_6486,N_4835,N_3296);
or U6487 (N_6487,N_4616,N_3857);
nand U6488 (N_6488,N_2988,N_2598);
nand U6489 (N_6489,N_3492,N_2992);
nor U6490 (N_6490,N_3542,N_4521);
and U6491 (N_6491,N_3283,N_2888);
xor U6492 (N_6492,N_4636,N_3714);
or U6493 (N_6493,N_4250,N_4461);
xor U6494 (N_6494,N_4011,N_3073);
nand U6495 (N_6495,N_3297,N_3137);
nor U6496 (N_6496,N_4420,N_4727);
nor U6497 (N_6497,N_3735,N_2999);
nand U6498 (N_6498,N_3996,N_3857);
and U6499 (N_6499,N_4531,N_4044);
and U6500 (N_6500,N_3910,N_4925);
nor U6501 (N_6501,N_2739,N_3489);
and U6502 (N_6502,N_3990,N_2879);
nor U6503 (N_6503,N_2634,N_2569);
and U6504 (N_6504,N_4192,N_2879);
nor U6505 (N_6505,N_4887,N_3993);
and U6506 (N_6506,N_2962,N_4339);
nor U6507 (N_6507,N_4613,N_2545);
nand U6508 (N_6508,N_3701,N_3761);
and U6509 (N_6509,N_4343,N_3458);
and U6510 (N_6510,N_2535,N_3070);
and U6511 (N_6511,N_4653,N_4257);
nor U6512 (N_6512,N_4313,N_3061);
xnor U6513 (N_6513,N_3988,N_3735);
nand U6514 (N_6514,N_3088,N_3838);
and U6515 (N_6515,N_4962,N_4523);
nand U6516 (N_6516,N_4108,N_3247);
and U6517 (N_6517,N_3741,N_3831);
and U6518 (N_6518,N_2635,N_3371);
and U6519 (N_6519,N_4838,N_4489);
or U6520 (N_6520,N_4501,N_4992);
nand U6521 (N_6521,N_2527,N_3449);
or U6522 (N_6522,N_4991,N_3937);
nand U6523 (N_6523,N_4078,N_2962);
or U6524 (N_6524,N_3516,N_2737);
or U6525 (N_6525,N_3852,N_3381);
nor U6526 (N_6526,N_3749,N_2592);
nor U6527 (N_6527,N_3809,N_3862);
and U6528 (N_6528,N_3366,N_4874);
or U6529 (N_6529,N_4346,N_3213);
nor U6530 (N_6530,N_4639,N_2728);
or U6531 (N_6531,N_4680,N_2741);
xnor U6532 (N_6532,N_3780,N_4664);
and U6533 (N_6533,N_4963,N_2808);
nor U6534 (N_6534,N_3717,N_3641);
xnor U6535 (N_6535,N_3558,N_3459);
nor U6536 (N_6536,N_3241,N_3011);
nand U6537 (N_6537,N_4782,N_3134);
nor U6538 (N_6538,N_4559,N_2778);
or U6539 (N_6539,N_3696,N_3908);
and U6540 (N_6540,N_2725,N_4828);
nor U6541 (N_6541,N_3486,N_3294);
or U6542 (N_6542,N_2944,N_4869);
or U6543 (N_6543,N_4327,N_3856);
nand U6544 (N_6544,N_4062,N_3379);
nor U6545 (N_6545,N_3194,N_2990);
nor U6546 (N_6546,N_4818,N_2709);
or U6547 (N_6547,N_3963,N_3360);
or U6548 (N_6548,N_2520,N_3442);
nor U6549 (N_6549,N_2952,N_4601);
nor U6550 (N_6550,N_3647,N_3498);
or U6551 (N_6551,N_3563,N_3390);
nor U6552 (N_6552,N_3695,N_2666);
nor U6553 (N_6553,N_2591,N_3370);
nand U6554 (N_6554,N_4831,N_3073);
and U6555 (N_6555,N_3202,N_3950);
nor U6556 (N_6556,N_2582,N_3989);
nand U6557 (N_6557,N_3936,N_3502);
and U6558 (N_6558,N_3223,N_2643);
or U6559 (N_6559,N_4197,N_4134);
nand U6560 (N_6560,N_3281,N_3275);
nand U6561 (N_6561,N_4996,N_3539);
or U6562 (N_6562,N_4847,N_3331);
and U6563 (N_6563,N_3772,N_4950);
or U6564 (N_6564,N_4016,N_3076);
and U6565 (N_6565,N_2844,N_4795);
nor U6566 (N_6566,N_4634,N_4197);
nand U6567 (N_6567,N_3090,N_3490);
and U6568 (N_6568,N_3207,N_4333);
or U6569 (N_6569,N_4433,N_3257);
nor U6570 (N_6570,N_3149,N_2731);
nor U6571 (N_6571,N_3530,N_4850);
and U6572 (N_6572,N_3426,N_4604);
nor U6573 (N_6573,N_3389,N_4522);
nand U6574 (N_6574,N_4841,N_3304);
and U6575 (N_6575,N_2954,N_3027);
and U6576 (N_6576,N_3811,N_4649);
nor U6577 (N_6577,N_3444,N_3522);
nor U6578 (N_6578,N_3188,N_4957);
nand U6579 (N_6579,N_2895,N_3361);
or U6580 (N_6580,N_3753,N_4058);
or U6581 (N_6581,N_4333,N_4639);
xnor U6582 (N_6582,N_3218,N_2974);
or U6583 (N_6583,N_4053,N_3685);
and U6584 (N_6584,N_2583,N_3210);
or U6585 (N_6585,N_4704,N_3363);
nand U6586 (N_6586,N_4997,N_3442);
and U6587 (N_6587,N_4025,N_3258);
nand U6588 (N_6588,N_4957,N_3619);
nor U6589 (N_6589,N_4404,N_3585);
xor U6590 (N_6590,N_4176,N_4813);
nor U6591 (N_6591,N_4042,N_3876);
nand U6592 (N_6592,N_3792,N_3750);
and U6593 (N_6593,N_2568,N_3111);
nor U6594 (N_6594,N_4412,N_3786);
or U6595 (N_6595,N_4291,N_3209);
nand U6596 (N_6596,N_3602,N_2845);
or U6597 (N_6597,N_4972,N_3940);
or U6598 (N_6598,N_2639,N_4180);
nor U6599 (N_6599,N_3787,N_3925);
nand U6600 (N_6600,N_3673,N_3587);
or U6601 (N_6601,N_2708,N_4018);
nand U6602 (N_6602,N_4992,N_3311);
nor U6603 (N_6603,N_4788,N_3007);
xor U6604 (N_6604,N_4624,N_3652);
or U6605 (N_6605,N_3622,N_3954);
or U6606 (N_6606,N_4352,N_2957);
and U6607 (N_6607,N_2924,N_4363);
nand U6608 (N_6608,N_2500,N_3689);
or U6609 (N_6609,N_4439,N_4105);
nor U6610 (N_6610,N_2558,N_4833);
nand U6611 (N_6611,N_3758,N_2596);
xnor U6612 (N_6612,N_3427,N_3831);
xnor U6613 (N_6613,N_2798,N_4667);
xnor U6614 (N_6614,N_4386,N_3958);
or U6615 (N_6615,N_4662,N_4170);
nand U6616 (N_6616,N_4961,N_3214);
nor U6617 (N_6617,N_3095,N_3314);
nand U6618 (N_6618,N_2710,N_3771);
and U6619 (N_6619,N_2901,N_4821);
or U6620 (N_6620,N_3937,N_4919);
nor U6621 (N_6621,N_4377,N_2548);
and U6622 (N_6622,N_2654,N_4324);
nand U6623 (N_6623,N_3884,N_2965);
or U6624 (N_6624,N_4860,N_4622);
and U6625 (N_6625,N_3737,N_3516);
nand U6626 (N_6626,N_3150,N_3358);
or U6627 (N_6627,N_3153,N_2737);
or U6628 (N_6628,N_3900,N_2566);
xor U6629 (N_6629,N_3710,N_3196);
or U6630 (N_6630,N_4094,N_3486);
or U6631 (N_6631,N_3849,N_4152);
nand U6632 (N_6632,N_4492,N_3724);
and U6633 (N_6633,N_2533,N_3969);
and U6634 (N_6634,N_3052,N_4562);
and U6635 (N_6635,N_2870,N_3505);
and U6636 (N_6636,N_3164,N_4317);
and U6637 (N_6637,N_3867,N_4225);
and U6638 (N_6638,N_3147,N_4613);
nor U6639 (N_6639,N_4638,N_2881);
nor U6640 (N_6640,N_3631,N_2810);
and U6641 (N_6641,N_3450,N_4237);
nor U6642 (N_6642,N_2754,N_3402);
nand U6643 (N_6643,N_4992,N_2809);
and U6644 (N_6644,N_3865,N_3611);
and U6645 (N_6645,N_3200,N_3128);
nor U6646 (N_6646,N_2822,N_4419);
or U6647 (N_6647,N_2748,N_2734);
nand U6648 (N_6648,N_3812,N_4300);
nand U6649 (N_6649,N_4759,N_3517);
nand U6650 (N_6650,N_3918,N_4902);
and U6651 (N_6651,N_4775,N_4411);
and U6652 (N_6652,N_4393,N_2662);
and U6653 (N_6653,N_2871,N_3089);
nor U6654 (N_6654,N_2864,N_3161);
and U6655 (N_6655,N_4487,N_4194);
nand U6656 (N_6656,N_3903,N_3749);
xnor U6657 (N_6657,N_4770,N_3155);
and U6658 (N_6658,N_3880,N_2624);
or U6659 (N_6659,N_3693,N_4041);
nand U6660 (N_6660,N_3069,N_3559);
and U6661 (N_6661,N_2787,N_4107);
nor U6662 (N_6662,N_3609,N_4410);
and U6663 (N_6663,N_2825,N_3831);
nor U6664 (N_6664,N_3477,N_4487);
nor U6665 (N_6665,N_3804,N_2714);
and U6666 (N_6666,N_2762,N_3369);
nand U6667 (N_6667,N_3194,N_3437);
and U6668 (N_6668,N_4681,N_3622);
and U6669 (N_6669,N_4494,N_3673);
nand U6670 (N_6670,N_3959,N_4263);
nand U6671 (N_6671,N_3921,N_4666);
or U6672 (N_6672,N_4250,N_4534);
and U6673 (N_6673,N_4838,N_4554);
nor U6674 (N_6674,N_3781,N_3540);
nor U6675 (N_6675,N_3315,N_4570);
nand U6676 (N_6676,N_2996,N_3466);
or U6677 (N_6677,N_2839,N_4341);
xnor U6678 (N_6678,N_3598,N_3825);
nand U6679 (N_6679,N_2942,N_2593);
nand U6680 (N_6680,N_4409,N_4615);
nand U6681 (N_6681,N_4608,N_2510);
or U6682 (N_6682,N_4776,N_4874);
or U6683 (N_6683,N_4373,N_3682);
or U6684 (N_6684,N_3626,N_3711);
nor U6685 (N_6685,N_4726,N_3289);
nand U6686 (N_6686,N_4411,N_2613);
xnor U6687 (N_6687,N_4210,N_3243);
nand U6688 (N_6688,N_4517,N_3535);
xor U6689 (N_6689,N_3504,N_2712);
nand U6690 (N_6690,N_4954,N_3806);
nand U6691 (N_6691,N_4928,N_3493);
nor U6692 (N_6692,N_4897,N_3886);
xnor U6693 (N_6693,N_4082,N_3830);
nand U6694 (N_6694,N_3393,N_2876);
and U6695 (N_6695,N_3842,N_4067);
nor U6696 (N_6696,N_4116,N_3897);
nor U6697 (N_6697,N_2906,N_2896);
and U6698 (N_6698,N_2674,N_2829);
nor U6699 (N_6699,N_3166,N_3728);
or U6700 (N_6700,N_3442,N_4272);
or U6701 (N_6701,N_4394,N_2702);
or U6702 (N_6702,N_2554,N_3425);
nor U6703 (N_6703,N_4814,N_2629);
xnor U6704 (N_6704,N_3550,N_3086);
and U6705 (N_6705,N_3057,N_4890);
nand U6706 (N_6706,N_4800,N_3407);
xor U6707 (N_6707,N_2635,N_4740);
nor U6708 (N_6708,N_3115,N_4801);
or U6709 (N_6709,N_4782,N_2651);
and U6710 (N_6710,N_4437,N_3174);
nor U6711 (N_6711,N_4063,N_4819);
nand U6712 (N_6712,N_3006,N_3568);
nand U6713 (N_6713,N_3037,N_4608);
nor U6714 (N_6714,N_3459,N_3303);
nor U6715 (N_6715,N_4695,N_3000);
and U6716 (N_6716,N_3037,N_3324);
and U6717 (N_6717,N_4158,N_2795);
or U6718 (N_6718,N_4235,N_2597);
nand U6719 (N_6719,N_4868,N_3973);
nor U6720 (N_6720,N_4696,N_4161);
and U6721 (N_6721,N_3886,N_3102);
xor U6722 (N_6722,N_4816,N_4110);
and U6723 (N_6723,N_2947,N_4349);
nand U6724 (N_6724,N_2616,N_3282);
or U6725 (N_6725,N_4241,N_4669);
xnor U6726 (N_6726,N_4476,N_3441);
nor U6727 (N_6727,N_3259,N_2838);
nor U6728 (N_6728,N_3796,N_4718);
and U6729 (N_6729,N_4114,N_4928);
xor U6730 (N_6730,N_4347,N_4316);
or U6731 (N_6731,N_3051,N_4595);
nor U6732 (N_6732,N_4684,N_3535);
nor U6733 (N_6733,N_3191,N_2584);
nand U6734 (N_6734,N_4468,N_4255);
nor U6735 (N_6735,N_4947,N_4501);
xor U6736 (N_6736,N_4612,N_3915);
and U6737 (N_6737,N_3254,N_4697);
xnor U6738 (N_6738,N_3872,N_3467);
or U6739 (N_6739,N_4975,N_4520);
nand U6740 (N_6740,N_4571,N_4881);
or U6741 (N_6741,N_2635,N_4205);
and U6742 (N_6742,N_4462,N_4450);
and U6743 (N_6743,N_4087,N_4973);
nand U6744 (N_6744,N_3030,N_4427);
nand U6745 (N_6745,N_4178,N_4697);
and U6746 (N_6746,N_4066,N_4557);
nor U6747 (N_6747,N_4425,N_3966);
or U6748 (N_6748,N_4407,N_4828);
or U6749 (N_6749,N_4999,N_2863);
nand U6750 (N_6750,N_3498,N_4741);
nand U6751 (N_6751,N_3742,N_2954);
or U6752 (N_6752,N_2570,N_2604);
xor U6753 (N_6753,N_4425,N_3206);
and U6754 (N_6754,N_3504,N_4435);
nor U6755 (N_6755,N_3305,N_2703);
nor U6756 (N_6756,N_3371,N_3647);
nor U6757 (N_6757,N_3388,N_3462);
or U6758 (N_6758,N_3882,N_3749);
nor U6759 (N_6759,N_4581,N_4454);
or U6760 (N_6760,N_3701,N_3130);
nor U6761 (N_6761,N_2591,N_4056);
nand U6762 (N_6762,N_2971,N_2743);
or U6763 (N_6763,N_4613,N_2769);
nor U6764 (N_6764,N_2580,N_4904);
and U6765 (N_6765,N_4011,N_3859);
and U6766 (N_6766,N_4746,N_4311);
nand U6767 (N_6767,N_4959,N_3748);
and U6768 (N_6768,N_4018,N_3391);
nor U6769 (N_6769,N_2921,N_2834);
and U6770 (N_6770,N_4498,N_3189);
nand U6771 (N_6771,N_4566,N_4640);
or U6772 (N_6772,N_2906,N_3452);
xnor U6773 (N_6773,N_2534,N_4689);
nor U6774 (N_6774,N_3105,N_3516);
and U6775 (N_6775,N_3486,N_4234);
nor U6776 (N_6776,N_3528,N_4421);
and U6777 (N_6777,N_4439,N_4277);
xnor U6778 (N_6778,N_3979,N_3606);
nor U6779 (N_6779,N_4888,N_3150);
and U6780 (N_6780,N_3622,N_4426);
nor U6781 (N_6781,N_2779,N_3674);
or U6782 (N_6782,N_4717,N_3153);
or U6783 (N_6783,N_4147,N_3833);
nand U6784 (N_6784,N_2659,N_4386);
nor U6785 (N_6785,N_4582,N_2609);
nand U6786 (N_6786,N_3702,N_3877);
xor U6787 (N_6787,N_2523,N_4056);
or U6788 (N_6788,N_3178,N_4412);
nor U6789 (N_6789,N_4759,N_3104);
nor U6790 (N_6790,N_3579,N_3587);
or U6791 (N_6791,N_4588,N_3911);
nand U6792 (N_6792,N_3518,N_4415);
nand U6793 (N_6793,N_4007,N_3549);
nand U6794 (N_6794,N_3702,N_3613);
nand U6795 (N_6795,N_4547,N_3685);
nor U6796 (N_6796,N_2923,N_2910);
nand U6797 (N_6797,N_3611,N_4811);
or U6798 (N_6798,N_2660,N_3089);
or U6799 (N_6799,N_3706,N_3635);
and U6800 (N_6800,N_3613,N_4697);
nand U6801 (N_6801,N_4728,N_4847);
or U6802 (N_6802,N_4997,N_4481);
nand U6803 (N_6803,N_4227,N_3118);
nor U6804 (N_6804,N_3974,N_3066);
nand U6805 (N_6805,N_2665,N_2780);
and U6806 (N_6806,N_3549,N_4302);
and U6807 (N_6807,N_4864,N_3916);
nor U6808 (N_6808,N_2917,N_2828);
and U6809 (N_6809,N_2930,N_2933);
nand U6810 (N_6810,N_2662,N_4352);
nand U6811 (N_6811,N_2943,N_4000);
or U6812 (N_6812,N_4745,N_2949);
and U6813 (N_6813,N_3327,N_3742);
or U6814 (N_6814,N_4757,N_2860);
nor U6815 (N_6815,N_4401,N_4468);
xor U6816 (N_6816,N_3107,N_4619);
nor U6817 (N_6817,N_3930,N_3256);
nand U6818 (N_6818,N_2793,N_3159);
xor U6819 (N_6819,N_3572,N_3062);
or U6820 (N_6820,N_3785,N_3419);
and U6821 (N_6821,N_4557,N_3823);
nand U6822 (N_6822,N_3559,N_4256);
or U6823 (N_6823,N_2840,N_3118);
nand U6824 (N_6824,N_3638,N_4990);
nand U6825 (N_6825,N_4971,N_3100);
or U6826 (N_6826,N_3727,N_4678);
and U6827 (N_6827,N_4265,N_3493);
or U6828 (N_6828,N_3826,N_4004);
and U6829 (N_6829,N_3230,N_4323);
or U6830 (N_6830,N_2735,N_3041);
and U6831 (N_6831,N_3701,N_4086);
xnor U6832 (N_6832,N_3989,N_2984);
and U6833 (N_6833,N_4530,N_3617);
nor U6834 (N_6834,N_2706,N_4839);
and U6835 (N_6835,N_2664,N_3145);
nor U6836 (N_6836,N_4508,N_4733);
and U6837 (N_6837,N_2923,N_3404);
or U6838 (N_6838,N_3548,N_3064);
xor U6839 (N_6839,N_4961,N_2741);
or U6840 (N_6840,N_3247,N_3474);
or U6841 (N_6841,N_3186,N_3414);
nand U6842 (N_6842,N_2683,N_3759);
or U6843 (N_6843,N_2745,N_2856);
or U6844 (N_6844,N_3124,N_4465);
and U6845 (N_6845,N_3447,N_4493);
nand U6846 (N_6846,N_3050,N_4179);
nand U6847 (N_6847,N_3830,N_2976);
nand U6848 (N_6848,N_4585,N_3749);
nor U6849 (N_6849,N_4950,N_3566);
nor U6850 (N_6850,N_3848,N_4461);
nand U6851 (N_6851,N_4695,N_3652);
and U6852 (N_6852,N_3473,N_3495);
and U6853 (N_6853,N_4732,N_4888);
and U6854 (N_6854,N_4941,N_4305);
or U6855 (N_6855,N_3406,N_2592);
or U6856 (N_6856,N_4590,N_4044);
nor U6857 (N_6857,N_4981,N_2822);
nand U6858 (N_6858,N_4145,N_4712);
nand U6859 (N_6859,N_3897,N_2897);
nand U6860 (N_6860,N_4556,N_3871);
nand U6861 (N_6861,N_3378,N_2604);
and U6862 (N_6862,N_3251,N_4628);
nor U6863 (N_6863,N_4054,N_4690);
or U6864 (N_6864,N_4138,N_3334);
or U6865 (N_6865,N_3360,N_3423);
nor U6866 (N_6866,N_3791,N_3083);
or U6867 (N_6867,N_3597,N_2915);
and U6868 (N_6868,N_4827,N_2667);
or U6869 (N_6869,N_2719,N_3981);
nand U6870 (N_6870,N_3496,N_4132);
and U6871 (N_6871,N_4253,N_3157);
and U6872 (N_6872,N_3415,N_3997);
xnor U6873 (N_6873,N_2672,N_4531);
and U6874 (N_6874,N_3183,N_3424);
nor U6875 (N_6875,N_4480,N_4335);
or U6876 (N_6876,N_4228,N_4873);
or U6877 (N_6877,N_3938,N_2983);
nor U6878 (N_6878,N_4247,N_4383);
or U6879 (N_6879,N_2500,N_3164);
nor U6880 (N_6880,N_4763,N_3811);
and U6881 (N_6881,N_4347,N_4947);
nor U6882 (N_6882,N_3945,N_4076);
and U6883 (N_6883,N_3375,N_3506);
and U6884 (N_6884,N_3707,N_4437);
or U6885 (N_6885,N_4133,N_4679);
and U6886 (N_6886,N_4949,N_4301);
nand U6887 (N_6887,N_4205,N_2903);
xnor U6888 (N_6888,N_3745,N_4700);
or U6889 (N_6889,N_2962,N_3066);
nor U6890 (N_6890,N_4025,N_3297);
and U6891 (N_6891,N_3252,N_4687);
nor U6892 (N_6892,N_3101,N_4267);
or U6893 (N_6893,N_3764,N_3490);
nand U6894 (N_6894,N_3832,N_3111);
and U6895 (N_6895,N_4664,N_4908);
nand U6896 (N_6896,N_4491,N_4843);
nand U6897 (N_6897,N_3168,N_2649);
and U6898 (N_6898,N_4045,N_3068);
nand U6899 (N_6899,N_2813,N_3101);
and U6900 (N_6900,N_4072,N_3179);
or U6901 (N_6901,N_4690,N_4813);
nand U6902 (N_6902,N_2962,N_4053);
nor U6903 (N_6903,N_3879,N_4716);
and U6904 (N_6904,N_2806,N_2864);
xor U6905 (N_6905,N_4127,N_3446);
xnor U6906 (N_6906,N_3466,N_3600);
nor U6907 (N_6907,N_3759,N_3894);
nand U6908 (N_6908,N_3361,N_3500);
xnor U6909 (N_6909,N_4975,N_4095);
nor U6910 (N_6910,N_2644,N_4208);
or U6911 (N_6911,N_4371,N_4598);
nor U6912 (N_6912,N_3281,N_4558);
and U6913 (N_6913,N_2956,N_3056);
nor U6914 (N_6914,N_4688,N_4803);
or U6915 (N_6915,N_4548,N_4167);
nand U6916 (N_6916,N_2878,N_4958);
nor U6917 (N_6917,N_4924,N_4637);
or U6918 (N_6918,N_4907,N_3962);
nand U6919 (N_6919,N_4488,N_4171);
or U6920 (N_6920,N_4967,N_4681);
nand U6921 (N_6921,N_2843,N_4043);
nand U6922 (N_6922,N_3584,N_4285);
or U6923 (N_6923,N_4803,N_2934);
and U6924 (N_6924,N_2868,N_4615);
nor U6925 (N_6925,N_4473,N_4756);
or U6926 (N_6926,N_3126,N_3760);
xnor U6927 (N_6927,N_3361,N_2808);
nand U6928 (N_6928,N_3467,N_3949);
nand U6929 (N_6929,N_2520,N_2992);
and U6930 (N_6930,N_3960,N_4096);
nor U6931 (N_6931,N_4864,N_3741);
or U6932 (N_6932,N_4961,N_4462);
or U6933 (N_6933,N_2517,N_3678);
nor U6934 (N_6934,N_4911,N_4159);
xor U6935 (N_6935,N_4722,N_2977);
nand U6936 (N_6936,N_4757,N_3997);
and U6937 (N_6937,N_3164,N_2508);
nor U6938 (N_6938,N_2713,N_4341);
nand U6939 (N_6939,N_3514,N_4800);
nand U6940 (N_6940,N_4209,N_4443);
or U6941 (N_6941,N_4904,N_4263);
nor U6942 (N_6942,N_4789,N_2625);
and U6943 (N_6943,N_3469,N_3723);
nand U6944 (N_6944,N_2981,N_4225);
nor U6945 (N_6945,N_2829,N_4615);
nand U6946 (N_6946,N_3417,N_3748);
xor U6947 (N_6947,N_4814,N_2647);
nand U6948 (N_6948,N_4489,N_3989);
and U6949 (N_6949,N_4922,N_3268);
nand U6950 (N_6950,N_2671,N_4075);
nand U6951 (N_6951,N_3405,N_2781);
or U6952 (N_6952,N_3757,N_3760);
and U6953 (N_6953,N_4106,N_2522);
nor U6954 (N_6954,N_3319,N_4154);
nand U6955 (N_6955,N_3005,N_4821);
nor U6956 (N_6956,N_3476,N_4801);
and U6957 (N_6957,N_3942,N_3928);
nor U6958 (N_6958,N_3246,N_4998);
nor U6959 (N_6959,N_3822,N_4240);
nor U6960 (N_6960,N_3107,N_2615);
or U6961 (N_6961,N_4038,N_3490);
and U6962 (N_6962,N_2943,N_4886);
or U6963 (N_6963,N_2897,N_3150);
nor U6964 (N_6964,N_4204,N_4827);
nand U6965 (N_6965,N_4339,N_4209);
nand U6966 (N_6966,N_4572,N_4407);
or U6967 (N_6967,N_4459,N_4456);
nand U6968 (N_6968,N_4177,N_3505);
and U6969 (N_6969,N_2663,N_2763);
nand U6970 (N_6970,N_4779,N_4694);
or U6971 (N_6971,N_3735,N_4308);
xnor U6972 (N_6972,N_4282,N_4789);
xnor U6973 (N_6973,N_4814,N_2602);
and U6974 (N_6974,N_3790,N_2839);
and U6975 (N_6975,N_3877,N_2963);
or U6976 (N_6976,N_3915,N_4177);
or U6977 (N_6977,N_4947,N_4136);
or U6978 (N_6978,N_4556,N_3877);
nand U6979 (N_6979,N_2693,N_4953);
nor U6980 (N_6980,N_3813,N_3360);
nor U6981 (N_6981,N_4836,N_2943);
and U6982 (N_6982,N_2520,N_3128);
nor U6983 (N_6983,N_3238,N_2960);
or U6984 (N_6984,N_3902,N_4690);
nor U6985 (N_6985,N_4197,N_2877);
or U6986 (N_6986,N_4983,N_4178);
nor U6987 (N_6987,N_4923,N_3415);
nor U6988 (N_6988,N_3542,N_2650);
nor U6989 (N_6989,N_3707,N_4772);
or U6990 (N_6990,N_4324,N_4301);
xnor U6991 (N_6991,N_3160,N_2976);
and U6992 (N_6992,N_3234,N_4820);
nand U6993 (N_6993,N_4310,N_4421);
nor U6994 (N_6994,N_4056,N_3025);
xor U6995 (N_6995,N_2678,N_4146);
and U6996 (N_6996,N_4049,N_4512);
and U6997 (N_6997,N_2732,N_4825);
or U6998 (N_6998,N_4982,N_2866);
or U6999 (N_6999,N_2638,N_2981);
nand U7000 (N_7000,N_4945,N_4246);
and U7001 (N_7001,N_4745,N_4446);
nor U7002 (N_7002,N_3775,N_4582);
or U7003 (N_7003,N_4642,N_4278);
xor U7004 (N_7004,N_4458,N_4095);
nand U7005 (N_7005,N_2523,N_4326);
nor U7006 (N_7006,N_3598,N_3719);
nor U7007 (N_7007,N_3575,N_3104);
xor U7008 (N_7008,N_4008,N_2759);
and U7009 (N_7009,N_3712,N_3308);
nand U7010 (N_7010,N_2906,N_3743);
nand U7011 (N_7011,N_2905,N_3949);
and U7012 (N_7012,N_4770,N_3615);
nand U7013 (N_7013,N_4734,N_3545);
and U7014 (N_7014,N_4507,N_4702);
and U7015 (N_7015,N_4898,N_4712);
or U7016 (N_7016,N_3714,N_2552);
nand U7017 (N_7017,N_3593,N_4658);
nand U7018 (N_7018,N_4044,N_4660);
nand U7019 (N_7019,N_2556,N_3671);
nor U7020 (N_7020,N_2896,N_3437);
nor U7021 (N_7021,N_3546,N_4802);
or U7022 (N_7022,N_3325,N_4372);
xor U7023 (N_7023,N_4262,N_4376);
nand U7024 (N_7024,N_4124,N_4578);
nand U7025 (N_7025,N_3865,N_4195);
or U7026 (N_7026,N_3134,N_4395);
nand U7027 (N_7027,N_4412,N_4739);
and U7028 (N_7028,N_3102,N_3677);
and U7029 (N_7029,N_3605,N_4110);
or U7030 (N_7030,N_4429,N_4295);
and U7031 (N_7031,N_2953,N_4980);
nor U7032 (N_7032,N_2610,N_3312);
xor U7033 (N_7033,N_3774,N_4954);
or U7034 (N_7034,N_4381,N_3357);
nor U7035 (N_7035,N_4667,N_3982);
or U7036 (N_7036,N_3990,N_4344);
nand U7037 (N_7037,N_3765,N_3101);
nand U7038 (N_7038,N_4914,N_4948);
nor U7039 (N_7039,N_4015,N_3797);
nand U7040 (N_7040,N_2535,N_4531);
or U7041 (N_7041,N_4772,N_3922);
and U7042 (N_7042,N_2659,N_4368);
nand U7043 (N_7043,N_4005,N_2631);
or U7044 (N_7044,N_4497,N_4971);
and U7045 (N_7045,N_3203,N_3597);
or U7046 (N_7046,N_2661,N_3406);
nand U7047 (N_7047,N_2771,N_4596);
and U7048 (N_7048,N_3402,N_3476);
nor U7049 (N_7049,N_2878,N_4078);
and U7050 (N_7050,N_4977,N_3766);
nand U7051 (N_7051,N_4672,N_3815);
xor U7052 (N_7052,N_3566,N_3490);
or U7053 (N_7053,N_3678,N_4806);
xor U7054 (N_7054,N_3130,N_4880);
and U7055 (N_7055,N_2614,N_3106);
nand U7056 (N_7056,N_3701,N_4651);
or U7057 (N_7057,N_3849,N_3427);
nor U7058 (N_7058,N_3203,N_4183);
or U7059 (N_7059,N_4585,N_3767);
and U7060 (N_7060,N_3089,N_4148);
nor U7061 (N_7061,N_4785,N_4631);
or U7062 (N_7062,N_4968,N_3782);
nand U7063 (N_7063,N_2870,N_4025);
xor U7064 (N_7064,N_4660,N_4725);
and U7065 (N_7065,N_4129,N_2888);
or U7066 (N_7066,N_2605,N_4087);
and U7067 (N_7067,N_4308,N_2855);
xor U7068 (N_7068,N_2749,N_2954);
nand U7069 (N_7069,N_4092,N_3527);
or U7070 (N_7070,N_3491,N_2552);
or U7071 (N_7071,N_3647,N_3981);
and U7072 (N_7072,N_4676,N_4037);
nor U7073 (N_7073,N_4745,N_4906);
nor U7074 (N_7074,N_3438,N_4774);
nand U7075 (N_7075,N_4231,N_4147);
or U7076 (N_7076,N_3900,N_3974);
nand U7077 (N_7077,N_2813,N_4888);
or U7078 (N_7078,N_3134,N_4647);
nor U7079 (N_7079,N_2885,N_3849);
nor U7080 (N_7080,N_4629,N_2524);
nor U7081 (N_7081,N_4949,N_3704);
and U7082 (N_7082,N_3243,N_2913);
and U7083 (N_7083,N_3202,N_2580);
nand U7084 (N_7084,N_2745,N_3220);
and U7085 (N_7085,N_3497,N_3861);
and U7086 (N_7086,N_3394,N_2501);
nor U7087 (N_7087,N_4507,N_4660);
nand U7088 (N_7088,N_2752,N_2561);
nor U7089 (N_7089,N_4146,N_4112);
nand U7090 (N_7090,N_2872,N_3492);
xnor U7091 (N_7091,N_3729,N_2669);
and U7092 (N_7092,N_4286,N_3665);
nand U7093 (N_7093,N_2837,N_3222);
or U7094 (N_7094,N_3772,N_3986);
and U7095 (N_7095,N_3914,N_4462);
nor U7096 (N_7096,N_3520,N_3627);
or U7097 (N_7097,N_4939,N_4867);
and U7098 (N_7098,N_4973,N_4004);
nor U7099 (N_7099,N_4624,N_4930);
and U7100 (N_7100,N_3847,N_3581);
or U7101 (N_7101,N_4122,N_2637);
nand U7102 (N_7102,N_4854,N_2772);
and U7103 (N_7103,N_3029,N_4350);
nand U7104 (N_7104,N_3866,N_2552);
or U7105 (N_7105,N_3335,N_2953);
nand U7106 (N_7106,N_2992,N_3078);
xnor U7107 (N_7107,N_2696,N_3572);
nand U7108 (N_7108,N_3273,N_4199);
nand U7109 (N_7109,N_2794,N_3006);
and U7110 (N_7110,N_3161,N_4432);
or U7111 (N_7111,N_4180,N_2822);
or U7112 (N_7112,N_3128,N_4866);
or U7113 (N_7113,N_3226,N_2890);
and U7114 (N_7114,N_3577,N_3813);
nand U7115 (N_7115,N_3553,N_3208);
nor U7116 (N_7116,N_4006,N_4329);
nor U7117 (N_7117,N_4146,N_4955);
nor U7118 (N_7118,N_4927,N_3386);
nor U7119 (N_7119,N_2970,N_3472);
and U7120 (N_7120,N_3750,N_3751);
xnor U7121 (N_7121,N_4964,N_3697);
or U7122 (N_7122,N_3400,N_4446);
nor U7123 (N_7123,N_4969,N_3468);
and U7124 (N_7124,N_3755,N_2973);
and U7125 (N_7125,N_4771,N_4488);
and U7126 (N_7126,N_4087,N_4504);
nor U7127 (N_7127,N_2917,N_3009);
or U7128 (N_7128,N_4307,N_3596);
nor U7129 (N_7129,N_3744,N_3311);
nor U7130 (N_7130,N_3679,N_2912);
and U7131 (N_7131,N_3256,N_4029);
or U7132 (N_7132,N_4362,N_2853);
or U7133 (N_7133,N_3568,N_4141);
and U7134 (N_7134,N_2512,N_3302);
or U7135 (N_7135,N_3042,N_4221);
nor U7136 (N_7136,N_2567,N_3519);
or U7137 (N_7137,N_3940,N_4679);
and U7138 (N_7138,N_4260,N_4250);
nor U7139 (N_7139,N_3471,N_3456);
and U7140 (N_7140,N_3089,N_3634);
or U7141 (N_7141,N_2725,N_3044);
nor U7142 (N_7142,N_3678,N_2708);
or U7143 (N_7143,N_4148,N_3803);
xor U7144 (N_7144,N_4553,N_4006);
nor U7145 (N_7145,N_4139,N_3055);
or U7146 (N_7146,N_3874,N_3000);
and U7147 (N_7147,N_3686,N_2810);
or U7148 (N_7148,N_3824,N_3712);
nand U7149 (N_7149,N_2948,N_2636);
nor U7150 (N_7150,N_4812,N_3792);
and U7151 (N_7151,N_3688,N_3844);
and U7152 (N_7152,N_2696,N_3528);
and U7153 (N_7153,N_4476,N_2531);
nor U7154 (N_7154,N_4350,N_3103);
nor U7155 (N_7155,N_4706,N_2933);
nand U7156 (N_7156,N_4970,N_2947);
or U7157 (N_7157,N_4066,N_3713);
nor U7158 (N_7158,N_3070,N_2533);
nand U7159 (N_7159,N_4991,N_3282);
xor U7160 (N_7160,N_2737,N_2718);
xor U7161 (N_7161,N_4840,N_2834);
nor U7162 (N_7162,N_3931,N_4060);
nand U7163 (N_7163,N_4749,N_4928);
nor U7164 (N_7164,N_3213,N_3934);
and U7165 (N_7165,N_4413,N_3564);
nor U7166 (N_7166,N_4998,N_4820);
nor U7167 (N_7167,N_4310,N_4029);
nand U7168 (N_7168,N_4677,N_4112);
and U7169 (N_7169,N_4748,N_4181);
nor U7170 (N_7170,N_2840,N_2523);
xor U7171 (N_7171,N_4342,N_4146);
or U7172 (N_7172,N_3033,N_2778);
nor U7173 (N_7173,N_3836,N_2996);
xnor U7174 (N_7174,N_2992,N_3910);
or U7175 (N_7175,N_3599,N_2589);
nand U7176 (N_7176,N_3667,N_4770);
and U7177 (N_7177,N_2703,N_2567);
xnor U7178 (N_7178,N_3184,N_4622);
nand U7179 (N_7179,N_3826,N_4852);
or U7180 (N_7180,N_2505,N_4685);
nand U7181 (N_7181,N_4738,N_3635);
nand U7182 (N_7182,N_2828,N_3215);
nand U7183 (N_7183,N_3732,N_4697);
and U7184 (N_7184,N_3088,N_4122);
or U7185 (N_7185,N_3545,N_2710);
or U7186 (N_7186,N_4175,N_3793);
nor U7187 (N_7187,N_4211,N_4681);
xnor U7188 (N_7188,N_4935,N_4150);
and U7189 (N_7189,N_2594,N_3146);
and U7190 (N_7190,N_4114,N_4528);
nor U7191 (N_7191,N_3250,N_2958);
xor U7192 (N_7192,N_3297,N_4230);
and U7193 (N_7193,N_4668,N_4921);
or U7194 (N_7194,N_4957,N_2969);
nor U7195 (N_7195,N_4453,N_4350);
nand U7196 (N_7196,N_3285,N_3284);
nor U7197 (N_7197,N_3415,N_2557);
or U7198 (N_7198,N_4086,N_4197);
and U7199 (N_7199,N_2781,N_3104);
nor U7200 (N_7200,N_3844,N_3739);
and U7201 (N_7201,N_3197,N_3794);
and U7202 (N_7202,N_2739,N_3093);
nor U7203 (N_7203,N_4179,N_4826);
xor U7204 (N_7204,N_3083,N_3254);
nand U7205 (N_7205,N_3375,N_4876);
and U7206 (N_7206,N_3223,N_3810);
or U7207 (N_7207,N_4567,N_4094);
and U7208 (N_7208,N_4866,N_2625);
or U7209 (N_7209,N_3414,N_2987);
nand U7210 (N_7210,N_3495,N_2607);
nand U7211 (N_7211,N_3936,N_3279);
nand U7212 (N_7212,N_4621,N_4367);
or U7213 (N_7213,N_3079,N_3871);
xor U7214 (N_7214,N_4180,N_2517);
nor U7215 (N_7215,N_3298,N_2633);
nand U7216 (N_7216,N_2864,N_4735);
nor U7217 (N_7217,N_3863,N_2682);
or U7218 (N_7218,N_2626,N_2564);
nand U7219 (N_7219,N_3331,N_3757);
or U7220 (N_7220,N_4073,N_4510);
nor U7221 (N_7221,N_2938,N_3340);
nand U7222 (N_7222,N_4901,N_4704);
nand U7223 (N_7223,N_3948,N_3911);
nor U7224 (N_7224,N_4163,N_4066);
nor U7225 (N_7225,N_4532,N_4521);
nand U7226 (N_7226,N_2648,N_4826);
and U7227 (N_7227,N_4244,N_2519);
xor U7228 (N_7228,N_4739,N_4594);
and U7229 (N_7229,N_2890,N_4424);
nand U7230 (N_7230,N_4562,N_3838);
or U7231 (N_7231,N_3659,N_2907);
nand U7232 (N_7232,N_3777,N_3442);
xor U7233 (N_7233,N_4104,N_2983);
or U7234 (N_7234,N_3745,N_3938);
nor U7235 (N_7235,N_3379,N_4228);
or U7236 (N_7236,N_3417,N_4712);
nor U7237 (N_7237,N_3486,N_3195);
or U7238 (N_7238,N_3628,N_3400);
or U7239 (N_7239,N_4804,N_4507);
nor U7240 (N_7240,N_3848,N_4644);
nor U7241 (N_7241,N_3901,N_2625);
nand U7242 (N_7242,N_3249,N_3552);
and U7243 (N_7243,N_4971,N_3928);
and U7244 (N_7244,N_2827,N_3204);
or U7245 (N_7245,N_2699,N_4872);
nand U7246 (N_7246,N_4550,N_2976);
nand U7247 (N_7247,N_4010,N_2528);
nand U7248 (N_7248,N_3096,N_2543);
nand U7249 (N_7249,N_3239,N_3921);
and U7250 (N_7250,N_3784,N_4873);
xor U7251 (N_7251,N_4666,N_3693);
nor U7252 (N_7252,N_4851,N_4272);
or U7253 (N_7253,N_4233,N_2951);
xnor U7254 (N_7254,N_4060,N_4464);
nand U7255 (N_7255,N_3973,N_2883);
and U7256 (N_7256,N_4083,N_3144);
and U7257 (N_7257,N_3153,N_4588);
and U7258 (N_7258,N_4570,N_3591);
and U7259 (N_7259,N_4137,N_4051);
nand U7260 (N_7260,N_2905,N_4265);
nor U7261 (N_7261,N_2882,N_3174);
nor U7262 (N_7262,N_2927,N_4377);
nor U7263 (N_7263,N_3442,N_2558);
nor U7264 (N_7264,N_3426,N_4277);
nor U7265 (N_7265,N_4277,N_3763);
nand U7266 (N_7266,N_3381,N_3041);
and U7267 (N_7267,N_3991,N_2759);
nor U7268 (N_7268,N_3398,N_4617);
xnor U7269 (N_7269,N_2654,N_3965);
or U7270 (N_7270,N_3193,N_4517);
xor U7271 (N_7271,N_4885,N_2624);
nand U7272 (N_7272,N_2920,N_4936);
nor U7273 (N_7273,N_4410,N_4243);
or U7274 (N_7274,N_4530,N_4290);
nand U7275 (N_7275,N_4141,N_4264);
and U7276 (N_7276,N_3653,N_3402);
or U7277 (N_7277,N_2551,N_4373);
nand U7278 (N_7278,N_4290,N_3659);
or U7279 (N_7279,N_3786,N_4828);
and U7280 (N_7280,N_4158,N_4440);
nand U7281 (N_7281,N_3178,N_2715);
nand U7282 (N_7282,N_3036,N_2733);
nor U7283 (N_7283,N_4557,N_3028);
xor U7284 (N_7284,N_4256,N_2910);
nand U7285 (N_7285,N_3440,N_3303);
nand U7286 (N_7286,N_2747,N_4128);
or U7287 (N_7287,N_4350,N_4366);
nand U7288 (N_7288,N_2738,N_3131);
nand U7289 (N_7289,N_3320,N_2627);
and U7290 (N_7290,N_3140,N_3686);
nor U7291 (N_7291,N_4608,N_4854);
or U7292 (N_7292,N_3638,N_4495);
nor U7293 (N_7293,N_2847,N_2619);
xnor U7294 (N_7294,N_3103,N_3884);
or U7295 (N_7295,N_4405,N_4388);
nand U7296 (N_7296,N_2931,N_2911);
and U7297 (N_7297,N_3243,N_2617);
or U7298 (N_7298,N_3319,N_3621);
and U7299 (N_7299,N_2676,N_4305);
and U7300 (N_7300,N_2643,N_2748);
nand U7301 (N_7301,N_3935,N_2653);
nor U7302 (N_7302,N_3185,N_3819);
nor U7303 (N_7303,N_4642,N_4716);
or U7304 (N_7304,N_4552,N_4689);
and U7305 (N_7305,N_2885,N_3638);
and U7306 (N_7306,N_4495,N_3119);
nand U7307 (N_7307,N_4556,N_3991);
and U7308 (N_7308,N_2604,N_3281);
and U7309 (N_7309,N_2802,N_4238);
nor U7310 (N_7310,N_4433,N_4744);
or U7311 (N_7311,N_4921,N_2725);
or U7312 (N_7312,N_3749,N_3057);
or U7313 (N_7313,N_3119,N_3147);
and U7314 (N_7314,N_4409,N_3982);
or U7315 (N_7315,N_4131,N_4302);
nor U7316 (N_7316,N_3785,N_3502);
nand U7317 (N_7317,N_2718,N_4261);
nor U7318 (N_7318,N_2828,N_2808);
and U7319 (N_7319,N_4961,N_3225);
or U7320 (N_7320,N_4785,N_3276);
and U7321 (N_7321,N_3446,N_4388);
nand U7322 (N_7322,N_4898,N_3014);
or U7323 (N_7323,N_2707,N_3423);
and U7324 (N_7324,N_3514,N_4724);
or U7325 (N_7325,N_4375,N_2635);
nand U7326 (N_7326,N_4407,N_3228);
nand U7327 (N_7327,N_2828,N_3905);
nand U7328 (N_7328,N_4408,N_3429);
or U7329 (N_7329,N_3934,N_4758);
nand U7330 (N_7330,N_2628,N_2816);
and U7331 (N_7331,N_2665,N_2639);
nor U7332 (N_7332,N_4651,N_2855);
and U7333 (N_7333,N_4450,N_3874);
nand U7334 (N_7334,N_2825,N_4968);
nand U7335 (N_7335,N_4628,N_2813);
and U7336 (N_7336,N_3544,N_4263);
and U7337 (N_7337,N_4508,N_4202);
and U7338 (N_7338,N_3617,N_3155);
and U7339 (N_7339,N_2826,N_2912);
nor U7340 (N_7340,N_4811,N_3975);
nand U7341 (N_7341,N_4982,N_3121);
and U7342 (N_7342,N_2980,N_4643);
or U7343 (N_7343,N_2682,N_2548);
nor U7344 (N_7344,N_4948,N_3762);
or U7345 (N_7345,N_3014,N_4235);
nand U7346 (N_7346,N_3804,N_3942);
nand U7347 (N_7347,N_2981,N_2935);
and U7348 (N_7348,N_3107,N_4802);
xor U7349 (N_7349,N_2573,N_3459);
nand U7350 (N_7350,N_2561,N_3963);
nor U7351 (N_7351,N_4909,N_4004);
and U7352 (N_7352,N_3971,N_2758);
nor U7353 (N_7353,N_3080,N_4302);
or U7354 (N_7354,N_3884,N_4032);
nor U7355 (N_7355,N_4660,N_4439);
nand U7356 (N_7356,N_2911,N_3308);
or U7357 (N_7357,N_3536,N_4324);
nand U7358 (N_7358,N_4578,N_3618);
or U7359 (N_7359,N_2560,N_3348);
nand U7360 (N_7360,N_2711,N_2529);
or U7361 (N_7361,N_3328,N_3868);
or U7362 (N_7362,N_4805,N_3626);
nand U7363 (N_7363,N_3269,N_3634);
and U7364 (N_7364,N_4454,N_3005);
or U7365 (N_7365,N_2607,N_4570);
nand U7366 (N_7366,N_4492,N_4732);
or U7367 (N_7367,N_4775,N_2621);
nor U7368 (N_7368,N_4375,N_2621);
and U7369 (N_7369,N_3105,N_4037);
xnor U7370 (N_7370,N_4399,N_3040);
xnor U7371 (N_7371,N_2642,N_4483);
nand U7372 (N_7372,N_4285,N_2828);
and U7373 (N_7373,N_4001,N_3277);
and U7374 (N_7374,N_3616,N_4894);
nand U7375 (N_7375,N_3890,N_4104);
and U7376 (N_7376,N_4240,N_4133);
nand U7377 (N_7377,N_3747,N_3943);
or U7378 (N_7378,N_4613,N_4710);
nor U7379 (N_7379,N_2786,N_3128);
nor U7380 (N_7380,N_2678,N_4542);
nor U7381 (N_7381,N_4345,N_3355);
and U7382 (N_7382,N_3843,N_4320);
nor U7383 (N_7383,N_3505,N_2773);
nand U7384 (N_7384,N_4464,N_2625);
and U7385 (N_7385,N_4086,N_4791);
and U7386 (N_7386,N_2786,N_2583);
and U7387 (N_7387,N_3466,N_4885);
nor U7388 (N_7388,N_2981,N_2990);
and U7389 (N_7389,N_2811,N_4345);
or U7390 (N_7390,N_4793,N_4431);
nand U7391 (N_7391,N_4174,N_4342);
and U7392 (N_7392,N_4261,N_3792);
nand U7393 (N_7393,N_2527,N_3373);
or U7394 (N_7394,N_2551,N_4225);
or U7395 (N_7395,N_2908,N_3002);
and U7396 (N_7396,N_2980,N_2787);
or U7397 (N_7397,N_4177,N_4961);
nand U7398 (N_7398,N_3452,N_3513);
nor U7399 (N_7399,N_4712,N_4052);
nand U7400 (N_7400,N_4520,N_4782);
xor U7401 (N_7401,N_4087,N_4004);
nand U7402 (N_7402,N_3386,N_2918);
nor U7403 (N_7403,N_3284,N_3806);
and U7404 (N_7404,N_3337,N_4634);
and U7405 (N_7405,N_4256,N_3086);
xnor U7406 (N_7406,N_4843,N_4465);
and U7407 (N_7407,N_4177,N_3012);
nor U7408 (N_7408,N_2975,N_4095);
or U7409 (N_7409,N_4011,N_4575);
or U7410 (N_7410,N_3662,N_3492);
xnor U7411 (N_7411,N_2682,N_3041);
xor U7412 (N_7412,N_4420,N_2504);
xnor U7413 (N_7413,N_4318,N_4812);
or U7414 (N_7414,N_2584,N_3037);
nor U7415 (N_7415,N_3187,N_4613);
and U7416 (N_7416,N_4835,N_3749);
and U7417 (N_7417,N_2555,N_3834);
nand U7418 (N_7418,N_2974,N_2624);
and U7419 (N_7419,N_3308,N_3261);
nand U7420 (N_7420,N_3595,N_4666);
xnor U7421 (N_7421,N_4331,N_4871);
or U7422 (N_7422,N_3119,N_2761);
and U7423 (N_7423,N_4468,N_3231);
nand U7424 (N_7424,N_3503,N_4123);
xor U7425 (N_7425,N_4168,N_3047);
nor U7426 (N_7426,N_2561,N_4048);
or U7427 (N_7427,N_2580,N_4712);
nor U7428 (N_7428,N_4889,N_4768);
and U7429 (N_7429,N_2515,N_2944);
nand U7430 (N_7430,N_4056,N_3533);
nand U7431 (N_7431,N_4629,N_4268);
nor U7432 (N_7432,N_4928,N_2782);
xor U7433 (N_7433,N_3980,N_3723);
or U7434 (N_7434,N_2748,N_4026);
nor U7435 (N_7435,N_4469,N_4271);
and U7436 (N_7436,N_3530,N_4574);
nand U7437 (N_7437,N_2941,N_3214);
and U7438 (N_7438,N_2900,N_4011);
or U7439 (N_7439,N_3707,N_3524);
nor U7440 (N_7440,N_3280,N_4475);
or U7441 (N_7441,N_3793,N_4898);
xor U7442 (N_7442,N_2511,N_3470);
nor U7443 (N_7443,N_3796,N_4391);
and U7444 (N_7444,N_2943,N_4347);
nand U7445 (N_7445,N_3086,N_2598);
xor U7446 (N_7446,N_4069,N_4075);
or U7447 (N_7447,N_3728,N_3007);
or U7448 (N_7448,N_4562,N_2887);
and U7449 (N_7449,N_3431,N_3819);
or U7450 (N_7450,N_3360,N_3573);
nand U7451 (N_7451,N_3057,N_3539);
or U7452 (N_7452,N_3839,N_2655);
nor U7453 (N_7453,N_3490,N_3352);
or U7454 (N_7454,N_2970,N_4052);
or U7455 (N_7455,N_3686,N_3931);
xnor U7456 (N_7456,N_4669,N_4466);
nand U7457 (N_7457,N_4141,N_2583);
and U7458 (N_7458,N_4495,N_3899);
nor U7459 (N_7459,N_3399,N_3797);
nand U7460 (N_7460,N_3392,N_4095);
or U7461 (N_7461,N_2826,N_3154);
nand U7462 (N_7462,N_3296,N_4234);
xor U7463 (N_7463,N_3043,N_3904);
and U7464 (N_7464,N_4245,N_2647);
nand U7465 (N_7465,N_3194,N_3073);
nand U7466 (N_7466,N_3886,N_3485);
nand U7467 (N_7467,N_4608,N_3736);
nand U7468 (N_7468,N_3811,N_3215);
nor U7469 (N_7469,N_3060,N_4485);
nor U7470 (N_7470,N_3386,N_4631);
or U7471 (N_7471,N_3443,N_4898);
or U7472 (N_7472,N_3815,N_4282);
nor U7473 (N_7473,N_3801,N_4618);
and U7474 (N_7474,N_3435,N_4489);
nand U7475 (N_7475,N_4718,N_4496);
nand U7476 (N_7476,N_2874,N_3041);
or U7477 (N_7477,N_4607,N_3559);
and U7478 (N_7478,N_3201,N_4044);
nor U7479 (N_7479,N_2779,N_2719);
and U7480 (N_7480,N_3930,N_3730);
nor U7481 (N_7481,N_4995,N_4310);
nand U7482 (N_7482,N_4524,N_3048);
or U7483 (N_7483,N_3402,N_4053);
and U7484 (N_7484,N_3492,N_2796);
xor U7485 (N_7485,N_3690,N_2671);
nand U7486 (N_7486,N_3336,N_4439);
nand U7487 (N_7487,N_2805,N_3224);
and U7488 (N_7488,N_4632,N_3318);
and U7489 (N_7489,N_3377,N_4063);
nand U7490 (N_7490,N_3376,N_4531);
or U7491 (N_7491,N_2636,N_4969);
and U7492 (N_7492,N_3400,N_4720);
xnor U7493 (N_7493,N_3377,N_4140);
or U7494 (N_7494,N_4359,N_3883);
nand U7495 (N_7495,N_4515,N_3980);
and U7496 (N_7496,N_3011,N_3570);
nand U7497 (N_7497,N_3491,N_4856);
nor U7498 (N_7498,N_3645,N_4843);
nand U7499 (N_7499,N_2572,N_2964);
and U7500 (N_7500,N_5753,N_6508);
xor U7501 (N_7501,N_6513,N_5217);
nor U7502 (N_7502,N_5768,N_5782);
nor U7503 (N_7503,N_7166,N_5830);
or U7504 (N_7504,N_5426,N_6658);
or U7505 (N_7505,N_5542,N_6523);
nand U7506 (N_7506,N_5271,N_5225);
or U7507 (N_7507,N_5843,N_5256);
or U7508 (N_7508,N_6354,N_7223);
nand U7509 (N_7509,N_5284,N_6649);
or U7510 (N_7510,N_6707,N_7212);
nor U7511 (N_7511,N_6998,N_5053);
nor U7512 (N_7512,N_6047,N_7145);
or U7513 (N_7513,N_6352,N_7332);
and U7514 (N_7514,N_5041,N_6547);
and U7515 (N_7515,N_5896,N_6457);
nand U7516 (N_7516,N_7063,N_7181);
nand U7517 (N_7517,N_5370,N_6371);
or U7518 (N_7518,N_5465,N_6032);
nor U7519 (N_7519,N_7200,N_5481);
xor U7520 (N_7520,N_5847,N_6312);
or U7521 (N_7521,N_7498,N_5093);
and U7522 (N_7522,N_6974,N_5791);
xnor U7523 (N_7523,N_6507,N_7033);
nor U7524 (N_7524,N_7019,N_5937);
nor U7525 (N_7525,N_5566,N_5659);
nand U7526 (N_7526,N_6398,N_6267);
or U7527 (N_7527,N_5196,N_5004);
nand U7528 (N_7528,N_5761,N_5429);
and U7529 (N_7529,N_6820,N_6294);
nand U7530 (N_7530,N_6551,N_6586);
nor U7531 (N_7531,N_6782,N_5805);
nand U7532 (N_7532,N_6151,N_6275);
nand U7533 (N_7533,N_5997,N_6051);
nand U7534 (N_7534,N_5668,N_5605);
nand U7535 (N_7535,N_7132,N_5671);
or U7536 (N_7536,N_7262,N_5441);
nor U7537 (N_7537,N_6688,N_5210);
nor U7538 (N_7538,N_6126,N_6915);
or U7539 (N_7539,N_7221,N_5518);
nand U7540 (N_7540,N_6827,N_6856);
nand U7541 (N_7541,N_6852,N_6105);
or U7542 (N_7542,N_7308,N_6740);
and U7543 (N_7543,N_7403,N_6530);
and U7544 (N_7544,N_5034,N_6988);
and U7545 (N_7545,N_5186,N_5974);
or U7546 (N_7546,N_6799,N_5918);
or U7547 (N_7547,N_5283,N_6565);
xnor U7548 (N_7548,N_6971,N_5374);
or U7549 (N_7549,N_7040,N_6607);
nor U7550 (N_7550,N_5475,N_7390);
nor U7551 (N_7551,N_7198,N_6015);
nor U7552 (N_7552,N_5988,N_5935);
nand U7553 (N_7553,N_5815,N_5721);
and U7554 (N_7554,N_7278,N_6385);
or U7555 (N_7555,N_6448,N_6737);
and U7556 (N_7556,N_5427,N_5823);
and U7557 (N_7557,N_5373,N_5158);
nor U7558 (N_7558,N_5458,N_6125);
and U7559 (N_7559,N_6948,N_6415);
and U7560 (N_7560,N_6578,N_5509);
and U7561 (N_7561,N_5389,N_5541);
nand U7562 (N_7562,N_6980,N_6609);
or U7563 (N_7563,N_5252,N_5015);
nor U7564 (N_7564,N_5218,N_7456);
xor U7565 (N_7565,N_5088,N_5716);
and U7566 (N_7566,N_5706,N_7338);
nor U7567 (N_7567,N_5163,N_7068);
or U7568 (N_7568,N_6640,N_5246);
and U7569 (N_7569,N_6169,N_7232);
and U7570 (N_7570,N_5244,N_7002);
or U7571 (N_7571,N_7071,N_6045);
nand U7572 (N_7572,N_6800,N_6058);
or U7573 (N_7573,N_5369,N_5002);
nor U7574 (N_7574,N_6285,N_5548);
nand U7575 (N_7575,N_6491,N_5870);
nand U7576 (N_7576,N_5075,N_5872);
nand U7577 (N_7577,N_6817,N_6531);
nor U7578 (N_7578,N_5781,N_5946);
and U7579 (N_7579,N_5836,N_6502);
and U7580 (N_7580,N_6109,N_7399);
and U7581 (N_7581,N_7315,N_6227);
nor U7582 (N_7582,N_6435,N_5808);
nor U7583 (N_7583,N_6766,N_6183);
or U7584 (N_7584,N_5590,N_6437);
or U7585 (N_7585,N_5061,N_5645);
or U7586 (N_7586,N_5938,N_6629);
or U7587 (N_7587,N_6121,N_5521);
nor U7588 (N_7588,N_5037,N_6452);
xor U7589 (N_7589,N_5071,N_7154);
nor U7590 (N_7590,N_6024,N_7446);
and U7591 (N_7591,N_6346,N_6391);
nand U7592 (N_7592,N_5251,N_5139);
and U7593 (N_7593,N_5547,N_7072);
and U7594 (N_7594,N_6672,N_7133);
nand U7595 (N_7595,N_6310,N_6886);
and U7596 (N_7596,N_6619,N_5038);
nor U7597 (N_7597,N_6806,N_5729);
or U7598 (N_7598,N_5174,N_6921);
and U7599 (N_7599,N_6914,N_5249);
xor U7600 (N_7600,N_6095,N_6009);
or U7601 (N_7601,N_5105,N_6160);
nand U7602 (N_7602,N_5673,N_5488);
xnor U7603 (N_7603,N_7324,N_6156);
nor U7604 (N_7604,N_6305,N_5470);
nand U7605 (N_7605,N_6651,N_6842);
and U7606 (N_7606,N_6152,N_6959);
xnor U7607 (N_7607,N_5709,N_5885);
nor U7608 (N_7608,N_5670,N_5189);
and U7609 (N_7609,N_5437,N_5422);
nand U7610 (N_7610,N_5893,N_5274);
and U7611 (N_7611,N_6529,N_6796);
or U7612 (N_7612,N_5192,N_7065);
nand U7613 (N_7613,N_5886,N_6725);
nor U7614 (N_7614,N_5773,N_7138);
nand U7615 (N_7615,N_5372,N_6142);
and U7616 (N_7616,N_5308,N_5181);
nor U7617 (N_7617,N_5469,N_5179);
xor U7618 (N_7618,N_6108,N_5471);
and U7619 (N_7619,N_7481,N_6464);
nor U7620 (N_7620,N_5787,N_5309);
nand U7621 (N_7621,N_6489,N_5151);
xnor U7622 (N_7622,N_5046,N_6844);
nand U7623 (N_7623,N_6055,N_6991);
nor U7624 (N_7624,N_6315,N_6159);
and U7625 (N_7625,N_6035,N_7067);
or U7626 (N_7626,N_6996,N_6610);
nor U7627 (N_7627,N_5914,N_5492);
nor U7628 (N_7628,N_7062,N_6481);
nand U7629 (N_7629,N_5124,N_5926);
nor U7630 (N_7630,N_7092,N_6898);
xor U7631 (N_7631,N_5734,N_5934);
nor U7632 (N_7632,N_5193,N_7417);
and U7633 (N_7633,N_6957,N_5042);
nand U7634 (N_7634,N_5097,N_6364);
and U7635 (N_7635,N_5685,N_5056);
nand U7636 (N_7636,N_5126,N_6040);
nor U7637 (N_7637,N_7034,N_5204);
or U7638 (N_7638,N_6247,N_6136);
or U7639 (N_7639,N_5330,N_6734);
or U7640 (N_7640,N_5882,N_6556);
nor U7641 (N_7641,N_7116,N_5695);
xnor U7642 (N_7642,N_5577,N_6116);
or U7643 (N_7643,N_6573,N_7393);
xnor U7644 (N_7644,N_6103,N_5275);
or U7645 (N_7645,N_6910,N_5107);
nand U7646 (N_7646,N_7080,N_6695);
nor U7647 (N_7647,N_6661,N_6306);
nand U7648 (N_7648,N_5466,N_5428);
xnor U7649 (N_7649,N_6137,N_6222);
nor U7650 (N_7650,N_6814,N_6238);
and U7651 (N_7651,N_6117,N_6511);
or U7652 (N_7652,N_5268,N_5825);
or U7653 (N_7653,N_6175,N_6596);
or U7654 (N_7654,N_5430,N_6402);
nor U7655 (N_7655,N_6666,N_6284);
nand U7656 (N_7656,N_6400,N_5079);
and U7657 (N_7657,N_5698,N_7239);
nor U7658 (N_7658,N_7366,N_5161);
xnor U7659 (N_7659,N_5137,N_5654);
nor U7660 (N_7660,N_5417,N_6257);
nand U7661 (N_7661,N_7139,N_5538);
and U7662 (N_7662,N_5928,N_6927);
and U7663 (N_7663,N_5445,N_6330);
or U7664 (N_7664,N_7013,N_6456);
nor U7665 (N_7665,N_7319,N_6213);
nor U7666 (N_7666,N_5332,N_6538);
and U7667 (N_7667,N_5939,N_5979);
or U7668 (N_7668,N_7373,N_5421);
xor U7669 (N_7669,N_6722,N_7211);
and U7670 (N_7670,N_6061,N_6631);
or U7671 (N_7671,N_6833,N_6788);
nand U7672 (N_7672,N_6038,N_6894);
xor U7673 (N_7673,N_6723,N_5378);
xor U7674 (N_7674,N_7484,N_5660);
or U7675 (N_7675,N_7011,N_7158);
nor U7676 (N_7676,N_5784,N_5044);
or U7677 (N_7677,N_5499,N_6252);
nand U7678 (N_7678,N_7209,N_5793);
nand U7679 (N_7679,N_6208,N_6138);
xor U7680 (N_7680,N_5055,N_5111);
or U7681 (N_7681,N_6639,N_5922);
and U7682 (N_7682,N_5361,N_7475);
and U7683 (N_7683,N_6684,N_5359);
or U7684 (N_7684,N_6846,N_6946);
and U7685 (N_7685,N_7275,N_5611);
xnor U7686 (N_7686,N_7128,N_7415);
nor U7687 (N_7687,N_5962,N_5187);
nor U7688 (N_7688,N_5953,N_5762);
or U7689 (N_7689,N_6689,N_5789);
and U7690 (N_7690,N_5536,N_5115);
nand U7691 (N_7691,N_5866,N_6211);
and U7692 (N_7692,N_6085,N_6114);
nor U7693 (N_7693,N_7144,N_7053);
and U7694 (N_7694,N_5132,N_5081);
xor U7695 (N_7695,N_6630,N_6191);
and U7696 (N_7696,N_6906,N_5303);
and U7697 (N_7697,N_6704,N_5069);
nor U7698 (N_7698,N_6575,N_5769);
and U7699 (N_7699,N_7476,N_5678);
xor U7700 (N_7700,N_5402,N_6622);
or U7701 (N_7701,N_7257,N_5639);
and U7702 (N_7702,N_7297,N_6104);
nand U7703 (N_7703,N_7151,N_5965);
nor U7704 (N_7704,N_6424,N_6107);
nor U7705 (N_7705,N_7224,N_5327);
or U7706 (N_7706,N_7294,N_6427);
and U7707 (N_7707,N_6897,N_6750);
nand U7708 (N_7708,N_5584,N_7120);
nor U7709 (N_7709,N_6985,N_7442);
nor U7710 (N_7710,N_5557,N_7109);
or U7711 (N_7711,N_7110,N_7429);
nor U7712 (N_7712,N_7237,N_6316);
nor U7713 (N_7713,N_6153,N_6769);
nor U7714 (N_7714,N_5530,N_7400);
nand U7715 (N_7715,N_7443,N_5150);
and U7716 (N_7716,N_5821,N_6965);
and U7717 (N_7717,N_6701,N_7049);
nor U7718 (N_7718,N_6389,N_5929);
and U7719 (N_7719,N_6911,N_6215);
and U7720 (N_7720,N_5517,N_5451);
or U7721 (N_7721,N_7352,N_6597);
nand U7722 (N_7722,N_7452,N_7081);
xor U7723 (N_7723,N_5223,N_5443);
or U7724 (N_7724,N_5000,N_6790);
nor U7725 (N_7725,N_5463,N_5447);
nand U7726 (N_7726,N_7291,N_7339);
or U7727 (N_7727,N_5856,N_6580);
and U7728 (N_7728,N_5068,N_5544);
nor U7729 (N_7729,N_6197,N_6230);
or U7730 (N_7730,N_6669,N_5845);
nand U7731 (N_7731,N_6463,N_5984);
or U7732 (N_7732,N_5418,N_6349);
or U7733 (N_7733,N_6308,N_6692);
and U7734 (N_7734,N_6767,N_5326);
and U7735 (N_7735,N_5258,N_6173);
nand U7736 (N_7736,N_6922,N_5976);
nor U7737 (N_7737,N_7320,N_5133);
and U7738 (N_7738,N_7042,N_6942);
xnor U7739 (N_7739,N_5395,N_5414);
and U7740 (N_7740,N_5666,N_6533);
and U7741 (N_7741,N_5508,N_6078);
xor U7742 (N_7742,N_6813,N_6100);
or U7743 (N_7743,N_5952,N_5663);
nor U7744 (N_7744,N_7396,N_7377);
and U7745 (N_7745,N_6232,N_6544);
nor U7746 (N_7746,N_5846,N_5444);
or U7747 (N_7747,N_7267,N_6745);
nor U7748 (N_7748,N_7421,N_6550);
nand U7749 (N_7749,N_6874,N_5533);
or U7750 (N_7750,N_5691,N_6811);
xor U7751 (N_7751,N_6585,N_6785);
or U7752 (N_7752,N_6559,N_5982);
and U7753 (N_7753,N_6512,N_5785);
xnor U7754 (N_7754,N_6490,N_5048);
or U7755 (N_7755,N_5738,N_5930);
xnor U7756 (N_7756,N_6092,N_5259);
nand U7757 (N_7757,N_6210,N_5279);
and U7758 (N_7758,N_7186,N_7046);
xor U7759 (N_7759,N_6338,N_5651);
or U7760 (N_7760,N_7178,N_6934);
xnor U7761 (N_7761,N_7242,N_5278);
nor U7762 (N_7762,N_6262,N_6070);
and U7763 (N_7763,N_5748,N_6992);
and U7764 (N_7764,N_6524,N_6124);
xor U7765 (N_7765,N_6357,N_6850);
nand U7766 (N_7766,N_7337,N_6432);
and U7767 (N_7767,N_5272,N_5449);
and U7768 (N_7768,N_5320,N_6872);
and U7769 (N_7769,N_6164,N_6558);
nand U7770 (N_7770,N_5114,N_5318);
nor U7771 (N_7771,N_6624,N_6298);
or U7772 (N_7772,N_5649,N_6123);
nor U7773 (N_7773,N_5794,N_5289);
and U7774 (N_7774,N_6568,N_6327);
or U7775 (N_7775,N_5198,N_7157);
nand U7776 (N_7776,N_5234,N_7351);
or U7777 (N_7777,N_5024,N_6313);
and U7778 (N_7778,N_7431,N_6081);
and U7779 (N_7779,N_6824,N_7401);
nand U7780 (N_7780,N_6154,N_5168);
nand U7781 (N_7781,N_7301,N_5532);
and U7782 (N_7782,N_6177,N_6373);
nor U7783 (N_7783,N_7188,N_6727);
nor U7784 (N_7784,N_5423,N_7325);
or U7785 (N_7785,N_5915,N_6925);
xor U7786 (N_7786,N_5248,N_5147);
nand U7787 (N_7787,N_6638,N_7298);
and U7788 (N_7788,N_6099,N_6258);
or U7789 (N_7789,N_6026,N_5919);
or U7790 (N_7790,N_5594,N_5503);
xor U7791 (N_7791,N_5467,N_5260);
or U7792 (N_7792,N_6266,N_6118);
and U7793 (N_7793,N_5250,N_6546);
or U7794 (N_7794,N_7427,N_5620);
and U7795 (N_7795,N_6781,N_5732);
and U7796 (N_7796,N_5095,N_7077);
and U7797 (N_7797,N_5632,N_7093);
xor U7798 (N_7798,N_5392,N_7482);
and U7799 (N_7799,N_7226,N_6469);
or U7800 (N_7800,N_6119,N_5432);
and U7801 (N_7801,N_6671,N_5407);
nand U7802 (N_7802,N_5707,N_6008);
nor U7803 (N_7803,N_5512,N_6369);
nand U7804 (N_7804,N_5102,N_5236);
or U7805 (N_7805,N_6648,N_5067);
nand U7806 (N_7806,N_6120,N_6768);
nand U7807 (N_7807,N_6002,N_6698);
xnor U7808 (N_7808,N_6467,N_5076);
nand U7809 (N_7809,N_6329,N_7462);
and U7810 (N_7810,N_7439,N_7149);
and U7811 (N_7811,N_5720,N_7392);
or U7812 (N_7812,N_5398,N_7261);
and U7813 (N_7813,N_5894,N_5814);
or U7814 (N_7814,N_7222,N_6292);
nor U7815 (N_7815,N_6729,N_5961);
or U7816 (N_7816,N_6941,N_5959);
xor U7817 (N_7817,N_5039,N_7370);
nand U7818 (N_7818,N_7265,N_6202);
nor U7819 (N_7819,N_6724,N_6699);
nor U7820 (N_7820,N_5209,N_6378);
or U7821 (N_7821,N_6129,N_5799);
or U7822 (N_7822,N_5749,N_5206);
and U7823 (N_7823,N_5744,N_7384);
nor U7824 (N_7824,N_6494,N_6969);
nor U7825 (N_7825,N_5439,N_6807);
nand U7826 (N_7826,N_6655,N_7048);
nand U7827 (N_7827,N_7194,N_5586);
or U7828 (N_7828,N_7030,N_5583);
nand U7829 (N_7829,N_6050,N_6381);
nand U7830 (N_7830,N_6112,N_6012);
nor U7831 (N_7831,N_5857,N_5631);
and U7832 (N_7832,N_7094,N_7314);
xor U7833 (N_7833,N_5110,N_5803);
xor U7834 (N_7834,N_5970,N_6361);
and U7835 (N_7835,N_5409,N_5170);
and U7836 (N_7836,N_5400,N_7474);
and U7837 (N_7837,N_6335,N_6972);
and U7838 (N_7838,N_5766,N_5975);
or U7839 (N_7839,N_7258,N_5143);
xnor U7840 (N_7840,N_7397,N_5992);
nand U7841 (N_7841,N_6505,N_5829);
xor U7842 (N_7842,N_6543,N_7283);
nand U7843 (N_7843,N_5177,N_6964);
and U7844 (N_7844,N_5101,N_6482);
nor U7845 (N_7845,N_6281,N_6076);
and U7846 (N_7846,N_6685,N_6383);
or U7847 (N_7847,N_6291,N_5214);
nand U7848 (N_7848,N_5901,N_6006);
or U7849 (N_7849,N_6127,N_5456);
nand U7850 (N_7850,N_5693,N_6522);
or U7851 (N_7851,N_5756,N_5873);
or U7852 (N_7852,N_7425,N_5498);
or U7853 (N_7853,N_7413,N_6149);
nor U7854 (N_7854,N_5945,N_6654);
nand U7855 (N_7855,N_5118,N_5711);
or U7856 (N_7856,N_6665,N_5298);
nor U7857 (N_7857,N_6226,N_7195);
or U7858 (N_7858,N_6834,N_5942);
nand U7859 (N_7859,N_6509,N_5786);
or U7860 (N_7860,N_5365,N_5644);
and U7861 (N_7861,N_7493,N_6388);
xor U7862 (N_7862,N_6730,N_6928);
or U7863 (N_7863,N_5801,N_5795);
nand U7864 (N_7864,N_6068,N_7164);
nand U7865 (N_7865,N_5242,N_5954);
nor U7866 (N_7866,N_6320,N_7001);
nor U7867 (N_7867,N_7485,N_5811);
or U7868 (N_7868,N_6244,N_5190);
and U7869 (N_7869,N_6031,N_6064);
and U7870 (N_7870,N_6421,N_5525);
or U7871 (N_7871,N_5387,N_7318);
nor U7872 (N_7872,N_5295,N_6454);
and U7873 (N_7873,N_5040,N_6789);
nand U7874 (N_7874,N_5454,N_6779);
nand U7875 (N_7875,N_6106,N_5587);
and U7876 (N_7876,N_7303,N_6111);
nor U7877 (N_7877,N_6216,N_6042);
nor U7878 (N_7878,N_5202,N_5888);
xnor U7879 (N_7879,N_5094,N_5049);
nand U7880 (N_7880,N_7076,N_5741);
and U7881 (N_7881,N_6819,N_5001);
and U7882 (N_7882,N_7406,N_6938);
nor U7883 (N_7883,N_5153,N_7099);
or U7884 (N_7884,N_5135,N_5612);
nand U7885 (N_7885,N_6347,N_6425);
or U7886 (N_7886,N_7031,N_5624);
or U7887 (N_7887,N_6908,N_5841);
nand U7888 (N_7888,N_7448,N_5057);
nand U7889 (N_7889,N_6739,N_6829);
nor U7890 (N_7890,N_5054,N_6599);
nand U7891 (N_7891,N_6994,N_7098);
xor U7892 (N_7892,N_5290,N_6474);
or U7893 (N_7893,N_6358,N_7470);
and U7894 (N_7894,N_7281,N_5077);
xor U7895 (N_7895,N_7469,N_5796);
and U7896 (N_7896,N_7016,N_6324);
and U7897 (N_7897,N_6155,N_5770);
nand U7898 (N_7898,N_6401,N_6270);
or U7899 (N_7899,N_6231,N_5677);
nor U7900 (N_7900,N_6771,N_5108);
and U7901 (N_7901,N_5241,N_7299);
nand U7902 (N_7902,N_5779,N_6838);
nor U7903 (N_7903,N_6600,N_5900);
nor U7904 (N_7904,N_6832,N_5972);
and U7905 (N_7905,N_6958,N_5399);
nand U7906 (N_7906,N_5078,N_6968);
nor U7907 (N_7907,N_5697,N_5802);
or U7908 (N_7908,N_6370,N_6020);
and U7909 (N_7909,N_6594,N_5345);
nand U7910 (N_7910,N_5507,N_5495);
and U7911 (N_7911,N_5005,N_5379);
xnor U7912 (N_7912,N_5485,N_5285);
and U7913 (N_7913,N_5656,N_6652);
nor U7914 (N_7914,N_5694,N_6880);
and U7915 (N_7915,N_5045,N_6670);
or U7916 (N_7916,N_7175,N_6122);
or U7917 (N_7917,N_5021,N_6949);
or U7918 (N_7918,N_5450,N_5588);
or U7919 (N_7919,N_6140,N_6434);
or U7920 (N_7920,N_7035,N_5247);
nand U7921 (N_7921,N_5434,N_5307);
nor U7922 (N_7922,N_5288,N_6525);
nor U7923 (N_7923,N_7371,N_7169);
and U7924 (N_7924,N_5130,N_6879);
nand U7925 (N_7925,N_5740,N_5136);
nand U7926 (N_7926,N_5637,N_7436);
xnor U7927 (N_7927,N_7408,N_7286);
and U7928 (N_7928,N_6206,N_6209);
nand U7929 (N_7929,N_6839,N_6097);
or U7930 (N_7930,N_5410,N_6653);
nor U7931 (N_7931,N_7134,N_7170);
and U7932 (N_7932,N_5980,N_5840);
and U7933 (N_7933,N_5554,N_5684);
or U7934 (N_7934,N_5457,N_5681);
and U7935 (N_7935,N_5047,N_6139);
nand U7936 (N_7936,N_5924,N_6952);
or U7937 (N_7937,N_7122,N_6756);
nor U7938 (N_7938,N_6916,N_6805);
and U7939 (N_7939,N_6478,N_6682);
nor U7940 (N_7940,N_5366,N_5310);
nand U7941 (N_7941,N_6878,N_5323);
xnor U7942 (N_7942,N_6611,N_7084);
and U7943 (N_7943,N_7054,N_6249);
or U7944 (N_7944,N_5863,N_5837);
and U7945 (N_7945,N_6608,N_6679);
or U7946 (N_7946,N_5348,N_5537);
xnor U7947 (N_7947,N_6527,N_5944);
or U7948 (N_7948,N_7328,N_6962);
or U7949 (N_7949,N_6625,N_6025);
xnor U7950 (N_7950,N_5887,N_7363);
and U7951 (N_7951,N_6903,N_6255);
or U7952 (N_7952,N_6560,N_7203);
or U7953 (N_7953,N_6636,N_5702);
or U7954 (N_7954,N_6981,N_5382);
nor U7955 (N_7955,N_5589,N_6690);
xor U7956 (N_7956,N_6515,N_6351);
nand U7957 (N_7957,N_6950,N_6438);
nor U7958 (N_7958,N_7486,N_5983);
and U7959 (N_7959,N_5215,N_6019);
and U7960 (N_7960,N_5925,N_5117);
nand U7961 (N_7961,N_5743,N_6742);
and U7962 (N_7962,N_6561,N_5705);
nand U7963 (N_7963,N_5771,N_5878);
and U7964 (N_7964,N_6674,N_6913);
nor U7965 (N_7965,N_7385,N_6668);
and U7966 (N_7966,N_5380,N_7414);
xnor U7967 (N_7967,N_6673,N_7150);
nor U7968 (N_7968,N_6504,N_6418);
nand U7969 (N_7969,N_7179,N_6614);
xor U7970 (N_7970,N_6269,N_6863);
nand U7971 (N_7971,N_5733,N_5213);
or U7972 (N_7972,N_6825,N_5932);
and U7973 (N_7973,N_5516,N_5630);
xnor U7974 (N_7974,N_6815,N_5360);
or U7975 (N_7975,N_5687,N_7165);
nor U7976 (N_7976,N_5364,N_5633);
and U7977 (N_7977,N_7497,N_6821);
nand U7978 (N_7978,N_5221,N_6657);
nor U7979 (N_7979,N_7457,N_7066);
xnor U7980 (N_7980,N_7409,N_6214);
and U7981 (N_7981,N_5180,N_7107);
or U7982 (N_7982,N_5416,N_6059);
nor U7983 (N_7983,N_6713,N_7219);
xnor U7984 (N_7984,N_6786,N_6084);
nor U7985 (N_7985,N_5319,N_6296);
and U7986 (N_7986,N_6300,N_5908);
and U7987 (N_7987,N_5265,N_7231);
nand U7988 (N_7988,N_6453,N_5032);
xnor U7989 (N_7989,N_5438,N_5640);
nand U7990 (N_7990,N_5165,N_5264);
and U7991 (N_7991,N_6772,N_5073);
nand U7992 (N_7992,N_7273,N_5717);
or U7993 (N_7993,N_6495,N_5035);
or U7994 (N_7994,N_7285,N_7480);
nor U7995 (N_7995,N_5715,N_5314);
nand U7996 (N_7996,N_5146,N_6696);
and U7997 (N_7997,N_6873,N_6647);
or U7998 (N_7998,N_5494,N_6634);
and U7999 (N_7999,N_6337,N_6344);
nor U8000 (N_8000,N_6835,N_6498);
xnor U8001 (N_8001,N_5968,N_6433);
nand U8002 (N_8002,N_5907,N_6590);
or U8003 (N_8003,N_6562,N_5317);
nand U8004 (N_8004,N_6620,N_5598);
nand U8005 (N_8005,N_7471,N_6204);
or U8006 (N_8006,N_6299,N_6738);
and U8007 (N_8007,N_5185,N_6067);
and U8008 (N_8008,N_5905,N_7353);
nor U8009 (N_8009,N_5994,N_6393);
nand U8010 (N_8010,N_5818,N_5699);
nand U8011 (N_8011,N_6302,N_6086);
nor U8012 (N_8012,N_6340,N_5396);
or U8013 (N_8013,N_5514,N_5489);
or U8014 (N_8014,N_5497,N_6613);
and U8015 (N_8015,N_5832,N_5227);
nand U8016 (N_8016,N_5844,N_6793);
or U8017 (N_8017,N_5257,N_5385);
or U8018 (N_8018,N_5501,N_7079);
and U8019 (N_8019,N_7307,N_7097);
nor U8020 (N_8020,N_7491,N_7118);
or U8021 (N_8021,N_5562,N_5127);
xnor U8022 (N_8022,N_7326,N_6322);
nand U8023 (N_8023,N_6374,N_7140);
or U8024 (N_8024,N_7216,N_5425);
xnor U8025 (N_8025,N_6379,N_7317);
nand U8026 (N_8026,N_5981,N_7495);
and U8027 (N_8027,N_7472,N_5910);
xor U8028 (N_8028,N_5822,N_6131);
xnor U8029 (N_8029,N_5574,N_6113);
or U8030 (N_8030,N_6862,N_6458);
nor U8031 (N_8031,N_7354,N_7083);
or U8032 (N_8032,N_5240,N_7088);
xor U8033 (N_8033,N_5496,N_6691);
nor U8034 (N_8034,N_5487,N_6518);
or U8035 (N_8035,N_5550,N_5013);
and U8036 (N_8036,N_5712,N_7037);
or U8037 (N_8037,N_5662,N_5595);
or U8038 (N_8038,N_5949,N_6053);
or U8039 (N_8039,N_5898,N_6978);
xnor U8040 (N_8040,N_6553,N_6776);
or U8041 (N_8041,N_6700,N_6023);
or U8042 (N_8042,N_6283,N_5216);
or U8043 (N_8043,N_6184,N_7368);
and U8044 (N_8044,N_5556,N_6984);
nand U8045 (N_8045,N_6676,N_6382);
nand U8046 (N_8046,N_5231,N_5254);
xnor U8047 (N_8047,N_5883,N_6246);
nor U8048 (N_8048,N_6063,N_5125);
xor U8049 (N_8049,N_6923,N_5783);
nand U8050 (N_8050,N_5534,N_6555);
xor U8051 (N_8051,N_7256,N_5867);
nand U8052 (N_8052,N_5355,N_6521);
or U8053 (N_8053,N_6587,N_6664);
and U8054 (N_8054,N_6172,N_6534);
or U8055 (N_8055,N_6810,N_6753);
xnor U8056 (N_8056,N_7420,N_5442);
nor U8057 (N_8057,N_5019,N_6318);
and U8058 (N_8058,N_5273,N_5472);
nand U8059 (N_8059,N_7130,N_5033);
nand U8060 (N_8060,N_6621,N_5504);
nand U8061 (N_8061,N_5482,N_5810);
nand U8062 (N_8062,N_6801,N_6497);
and U8063 (N_8063,N_5597,N_5338);
nand U8064 (N_8064,N_7220,N_6413);
and U8065 (N_8065,N_6795,N_6589);
nand U8066 (N_8066,N_6286,N_5617);
or U8067 (N_8067,N_5977,N_5608);
nand U8068 (N_8068,N_5436,N_6010);
xor U8069 (N_8069,N_6404,N_6899);
nor U8070 (N_8070,N_6180,N_6765);
nor U8071 (N_8071,N_5555,N_6030);
nor U8072 (N_8072,N_5324,N_6708);
xor U8073 (N_8073,N_6168,N_7335);
or U8074 (N_8074,N_7477,N_6236);
and U8075 (N_8075,N_5090,N_6289);
xnor U8076 (N_8076,N_6319,N_7260);
nand U8077 (N_8077,N_6932,N_7191);
xor U8078 (N_8078,N_6397,N_5986);
nand U8079 (N_8079,N_7355,N_6261);
or U8080 (N_8080,N_5578,N_7020);
and U8081 (N_8081,N_6851,N_5243);
xnor U8082 (N_8082,N_5157,N_6093);
or U8083 (N_8083,N_7459,N_5592);
and U8084 (N_8084,N_7341,N_6535);
nor U8085 (N_8085,N_6277,N_5614);
or U8086 (N_8086,N_5686,N_6065);
nand U8087 (N_8087,N_5315,N_7494);
xor U8088 (N_8088,N_5758,N_6577);
nor U8089 (N_8089,N_7225,N_6339);
nor U8090 (N_8090,N_6054,N_6931);
or U8091 (N_8091,N_6224,N_5322);
nand U8092 (N_8092,N_6885,N_5853);
or U8093 (N_8093,N_5551,N_6356);
nand U8094 (N_8094,N_5377,N_7126);
and U8095 (N_8095,N_5331,N_6314);
xnor U8096 (N_8096,N_6719,N_5119);
or U8097 (N_8097,N_5351,N_7075);
and U8098 (N_8098,N_6717,N_5513);
xor U8099 (N_8099,N_6735,N_5230);
and U8100 (N_8100,N_5813,N_5156);
or U8101 (N_8101,N_5606,N_6882);
nor U8102 (N_8102,N_5724,N_6419);
or U8103 (N_8103,N_6966,N_5368);
and U8104 (N_8104,N_6290,N_5559);
nor U8105 (N_8105,N_6588,N_5478);
nor U8106 (N_8106,N_5646,N_6241);
nor U8107 (N_8107,N_5816,N_5228);
nand U8108 (N_8108,N_6196,N_5842);
and U8109 (N_8109,N_7402,N_5778);
or U8110 (N_8110,N_6733,N_7051);
nor U8111 (N_8111,N_6212,N_7419);
nor U8112 (N_8112,N_7454,N_5860);
xor U8113 (N_8113,N_7111,N_6757);
nor U8114 (N_8114,N_6390,N_7202);
nand U8115 (N_8115,N_7358,N_5765);
nand U8116 (N_8116,N_5164,N_7374);
and U8117 (N_8117,N_7135,N_6034);
or U8118 (N_8118,N_7270,N_5861);
nand U8119 (N_8119,N_6239,N_5726);
or U8120 (N_8120,N_5627,N_6881);
xnor U8121 (N_8121,N_6426,N_6430);
nor U8122 (N_8122,N_7050,N_7014);
and U8123 (N_8123,N_7340,N_6728);
nand U8124 (N_8124,N_5600,N_7289);
nor U8125 (N_8125,N_7302,N_5411);
nand U8126 (N_8126,N_6939,N_7057);
and U8127 (N_8127,N_6510,N_6248);
or U8128 (N_8128,N_5098,N_7333);
xor U8129 (N_8129,N_5148,N_5222);
nor U8130 (N_8130,N_7101,N_6711);
and U8131 (N_8131,N_7123,N_6157);
nand U8132 (N_8132,N_5043,N_6641);
xor U8133 (N_8133,N_6784,N_5747);
and U8134 (N_8134,N_5776,N_7213);
and U8135 (N_8135,N_6461,N_6501);
and U8136 (N_8136,N_6552,N_5388);
nor U8137 (N_8137,N_6250,N_6506);
and U8138 (N_8138,N_7026,N_6830);
nand U8139 (N_8139,N_5563,N_5328);
and U8140 (N_8140,N_5375,N_5526);
nor U8141 (N_8141,N_6132,N_6702);
and U8142 (N_8142,N_5807,N_5511);
nand U8143 (N_8143,N_7246,N_7106);
nand U8144 (N_8144,N_5891,N_7193);
and U8145 (N_8145,N_5211,N_6520);
nor U8146 (N_8146,N_5619,N_5312);
or U8147 (N_8147,N_6761,N_5025);
nand U8148 (N_8148,N_5082,N_7036);
nor U8149 (N_8149,N_5629,N_5764);
or U8150 (N_8150,N_7259,N_5325);
or U8151 (N_8151,N_5232,N_5100);
or U8152 (N_8152,N_6995,N_6265);
nor U8153 (N_8153,N_6264,N_7021);
xnor U8154 (N_8154,N_7156,N_5390);
nor U8155 (N_8155,N_7155,N_5141);
xnor U8156 (N_8156,N_7437,N_7438);
nor U8157 (N_8157,N_7124,N_7117);
nand U8158 (N_8158,N_6416,N_5718);
and U8159 (N_8159,N_5435,N_5296);
and U8160 (N_8160,N_6570,N_7422);
nand U8161 (N_8161,N_7376,N_5897);
nor U8162 (N_8162,N_5710,N_7263);
and U8163 (N_8163,N_5201,N_6667);
xor U8164 (N_8164,N_7334,N_5623);
nand U8165 (N_8165,N_6101,N_5086);
nor U8166 (N_8166,N_6847,N_7210);
nor U8167 (N_8167,N_5775,N_6901);
nor U8168 (N_8168,N_7271,N_6342);
and U8169 (N_8169,N_6380,N_5142);
nor U8170 (N_8170,N_7487,N_5973);
and U8171 (N_8171,N_6884,N_7455);
and U8172 (N_8172,N_5352,N_6459);
or U8173 (N_8173,N_5728,N_5301);
and U8174 (N_8174,N_7252,N_5854);
and U8175 (N_8175,N_6633,N_5091);
nand U8176 (N_8176,N_5713,N_7160);
nand U8177 (N_8177,N_7424,N_6091);
or U8178 (N_8178,N_5899,N_6317);
or U8179 (N_8179,N_7003,N_7172);
nand U8180 (N_8180,N_5415,N_7218);
nand U8181 (N_8181,N_7114,N_7490);
and U8182 (N_8182,N_5245,N_7346);
nor U8183 (N_8183,N_5616,N_5031);
nand U8184 (N_8184,N_5208,N_6460);
or U8185 (N_8185,N_7102,N_7248);
nand U8186 (N_8186,N_6429,N_6276);
nand U8187 (N_8187,N_5145,N_7423);
nor U8188 (N_8188,N_5759,N_6080);
nand U8189 (N_8189,N_7032,N_7190);
xor U8190 (N_8190,N_7171,N_5066);
nor U8191 (N_8191,N_7018,N_7241);
and U8192 (N_8192,N_5474,N_6866);
nand U8193 (N_8193,N_7069,N_5868);
or U8194 (N_8194,N_6736,N_5850);
nor U8195 (N_8195,N_6615,N_6718);
and U8196 (N_8196,N_5028,N_5812);
and U8197 (N_8197,N_6110,N_7047);
and U8198 (N_8198,N_6841,N_5052);
or U8199 (N_8199,N_7264,N_5183);
and U8200 (N_8200,N_5912,N_5007);
xnor U8201 (N_8201,N_6423,N_6583);
or U8202 (N_8202,N_5113,N_7300);
xnor U8203 (N_8203,N_7276,N_7187);
nor U8204 (N_8204,N_7007,N_6940);
and U8205 (N_8205,N_7238,N_7112);
nor U8206 (N_8206,N_7389,N_5419);
nor U8207 (N_8207,N_7372,N_6519);
xor U8208 (N_8208,N_5281,N_5349);
xor U8209 (N_8209,N_5484,N_5096);
or U8210 (N_8210,N_6332,N_6158);
or U8211 (N_8211,N_5657,N_7488);
and U8212 (N_8212,N_5336,N_5112);
nand U8213 (N_8213,N_6003,N_5505);
or U8214 (N_8214,N_6492,N_6646);
nand U8215 (N_8215,N_5292,N_5576);
or U8216 (N_8216,N_7176,N_6780);
and U8217 (N_8217,N_5564,N_5971);
xnor U8218 (N_8218,N_6409,N_5672);
and U8219 (N_8219,N_6549,N_5404);
and U8220 (N_8220,N_6472,N_7039);
and U8221 (N_8221,N_6087,N_5403);
nand U8222 (N_8222,N_7201,N_5987);
or U8223 (N_8223,N_6394,N_5476);
nand U8224 (N_8224,N_5539,N_6145);
or U8225 (N_8225,N_6499,N_6809);
nor U8226 (N_8226,N_6816,N_6488);
nor U8227 (N_8227,N_6632,N_5913);
nor U8228 (N_8228,N_6408,N_6909);
xnor U8229 (N_8229,N_5287,N_5316);
and U8230 (N_8230,N_6162,N_7215);
nor U8231 (N_8231,N_7173,N_5459);
nand U8232 (N_8232,N_6603,N_5493);
nand U8233 (N_8233,N_6074,N_6861);
and U8234 (N_8234,N_5335,N_6752);
and U8235 (N_8235,N_6446,N_5904);
or U8236 (N_8236,N_6079,N_7432);
or U8237 (N_8237,N_7284,N_5140);
or U8238 (N_8238,N_6975,N_6802);
xor U8239 (N_8239,N_6758,N_7253);
or U8240 (N_8240,N_5831,N_7321);
nor U8241 (N_8241,N_5302,N_5704);
and U8242 (N_8242,N_6004,N_6539);
nand U8243 (N_8243,N_6937,N_7105);
nor U8244 (N_8244,N_5304,N_6875);
nor U8245 (N_8245,N_5023,N_5792);
nand U8246 (N_8246,N_5219,N_5820);
and U8247 (N_8247,N_5552,N_5408);
and U8248 (N_8248,N_5060,N_6052);
nand U8249 (N_8249,N_6440,N_5452);
nor U8250 (N_8250,N_7010,N_7458);
and U8251 (N_8251,N_6189,N_6274);
and U8252 (N_8252,N_7479,N_6601);
or U8253 (N_8253,N_7381,N_6355);
nor U8254 (N_8254,N_5203,N_7103);
nor U8255 (N_8255,N_7217,N_5903);
nor U8256 (N_8256,N_6887,N_6439);
or U8257 (N_8257,N_5636,N_6001);
and U8258 (N_8258,N_6731,N_6889);
and U8259 (N_8259,N_7364,N_5950);
nand U8260 (N_8260,N_6643,N_6831);
nor U8261 (N_8261,N_7311,N_6582);
nor U8262 (N_8262,N_6973,N_7349);
and U8263 (N_8263,N_6465,N_6876);
nor U8264 (N_8264,N_5916,N_5881);
or U8265 (N_8265,N_6147,N_6697);
nor U8266 (N_8266,N_6014,N_5569);
nor U8267 (N_8267,N_6280,N_6970);
xnor U8268 (N_8268,N_5581,N_7082);
or U8269 (N_8269,N_5601,N_6480);
or U8270 (N_8270,N_6693,N_7254);
and U8271 (N_8271,N_6449,N_6743);
nor U8272 (N_8272,N_6716,N_6890);
nor U8273 (N_8273,N_6366,N_6960);
and U8274 (N_8274,N_7045,N_6377);
or U8275 (N_8275,N_6485,N_6628);
and U8276 (N_8276,N_5027,N_5167);
or U8277 (N_8277,N_6763,N_5277);
nand U8278 (N_8278,N_6746,N_5343);
or U8279 (N_8279,N_6487,N_7233);
and U8280 (N_8280,N_6642,N_5991);
or U8281 (N_8281,N_6376,N_5376);
xor U8282 (N_8282,N_6345,N_6726);
or U8283 (N_8283,N_7028,N_6627);
or U8284 (N_8284,N_6333,N_5798);
nand U8285 (N_8285,N_5543,N_7449);
nand U8286 (N_8286,N_6060,N_5835);
or U8287 (N_8287,N_6954,N_7279);
nor U8288 (N_8288,N_6569,N_6143);
or U8289 (N_8289,N_7359,N_6528);
or U8290 (N_8290,N_5546,N_6171);
and U8291 (N_8291,N_7433,N_6891);
nand U8292 (N_8292,N_6979,N_7087);
and U8293 (N_8293,N_7394,N_6576);
and U8294 (N_8294,N_7282,N_5849);
nor U8295 (N_8295,N_5607,N_6867);
or U8296 (N_8296,N_6102,N_7492);
nand U8297 (N_8297,N_5063,N_6326);
nand U8298 (N_8298,N_6759,N_6254);
nand U8299 (N_8299,N_6961,N_5291);
nand U8300 (N_8300,N_5297,N_6986);
nor U8301 (N_8301,N_6953,N_6747);
nor U8302 (N_8302,N_5362,N_7204);
nor U8303 (N_8303,N_6869,N_6853);
nand U8304 (N_8304,N_6077,N_5871);
and U8305 (N_8305,N_5648,N_6016);
or U8306 (N_8306,N_5354,N_6399);
xnor U8307 (N_8307,N_6017,N_5906);
or U8308 (N_8308,N_6564,N_5226);
nor U8309 (N_8309,N_7182,N_7460);
and U8310 (N_8310,N_7331,N_6912);
or U8311 (N_8311,N_5571,N_5313);
or U8312 (N_8312,N_6920,N_5688);
nor U8313 (N_8313,N_7430,N_6967);
or U8314 (N_8314,N_7356,N_5780);
and U8315 (N_8315,N_7161,N_7174);
or U8316 (N_8316,N_6865,N_5689);
and U8317 (N_8317,N_6818,N_6503);
and U8318 (N_8318,N_6572,N_6375);
nor U8319 (N_8319,N_5464,N_6812);
and U8320 (N_8320,N_7148,N_7229);
nand U8321 (N_8321,N_5545,N_6395);
and U8322 (N_8322,N_5692,N_5746);
and U8323 (N_8323,N_6075,N_7305);
xnor U8324 (N_8324,N_7290,N_5572);
nor U8325 (N_8325,N_6295,N_5050);
nand U8326 (N_8326,N_6792,N_7086);
and U8327 (N_8327,N_6331,N_6945);
and U8328 (N_8328,N_5253,N_7146);
nor U8329 (N_8329,N_6982,N_7395);
and U8330 (N_8330,N_7228,N_7312);
nor U8331 (N_8331,N_5486,N_5955);
or U8332 (N_8332,N_7159,N_5229);
nand U8333 (N_8333,N_6977,N_6680);
xnor U8334 (N_8334,N_6579,N_6870);
and U8335 (N_8335,N_7287,N_7214);
nand U8336 (N_8336,N_6411,N_5089);
xnor U8337 (N_8337,N_5989,N_5461);
or U8338 (N_8338,N_6445,N_5767);
and U8339 (N_8339,N_6256,N_6473);
nor U8340 (N_8340,N_6387,N_5956);
and U8341 (N_8341,N_5431,N_5679);
nor U8342 (N_8342,N_5591,N_5999);
nand U8343 (N_8343,N_6919,N_5128);
and U8344 (N_8344,N_6362,N_6303);
nor U8345 (N_8345,N_7061,N_5565);
nand U8346 (N_8346,N_5575,N_6926);
and U8347 (N_8347,N_5103,N_5220);
xnor U8348 (N_8348,N_7055,N_6412);
or U8349 (N_8349,N_5003,N_7043);
nor U8350 (N_8350,N_5477,N_7295);
and U8351 (N_8351,N_5016,N_5622);
nor U8352 (N_8352,N_6161,N_6924);
and U8353 (N_8353,N_6242,N_6007);
and U8354 (N_8354,N_6537,N_5817);
or U8355 (N_8355,N_7059,N_7306);
nor U8356 (N_8356,N_7483,N_6517);
xor U8357 (N_8357,N_6705,N_5967);
nor U8358 (N_8358,N_5824,N_7015);
nor U8359 (N_8359,N_6857,N_6237);
nand U8360 (N_8360,N_7234,N_5269);
nand U8361 (N_8361,N_6165,N_6868);
and U8362 (N_8362,N_5966,N_5064);
nand U8363 (N_8363,N_6477,N_6486);
nor U8364 (N_8364,N_5652,N_5834);
or U8365 (N_8365,N_7091,N_7288);
nor U8366 (N_8366,N_5683,N_7280);
xnor U8367 (N_8367,N_5255,N_5384);
nand U8368 (N_8368,N_6253,N_6703);
and U8369 (N_8369,N_7461,N_6046);
nor U8370 (N_8370,N_6341,N_6871);
nor U8371 (N_8371,N_7192,N_6476);
or U8372 (N_8372,N_5568,N_7313);
nand U8373 (N_8373,N_6548,N_6396);
and U8374 (N_8374,N_5696,N_6417);
nor U8375 (N_8375,N_6526,N_5618);
or U8376 (N_8376,N_5008,N_5267);
or U8377 (N_8377,N_6951,N_6414);
or U8378 (N_8378,N_5311,N_5200);
or U8379 (N_8379,N_5030,N_5879);
nand U8380 (N_8380,N_7108,N_5978);
and U8381 (N_8381,N_5641,N_6755);
nand U8382 (N_8382,N_6783,N_5006);
nand U8383 (N_8383,N_5406,N_5902);
and U8384 (N_8384,N_6027,N_6936);
or U8385 (N_8385,N_7350,N_7168);
nor U8386 (N_8386,N_6637,N_6749);
nor U8387 (N_8387,N_5714,N_5329);
or U8388 (N_8388,N_5655,N_7451);
and U8389 (N_8389,N_5635,N_5122);
xnor U8390 (N_8390,N_5531,N_6644);
or U8391 (N_8391,N_7407,N_5540);
and U8392 (N_8392,N_5731,N_6574);
or U8393 (N_8393,N_7137,N_5875);
and U8394 (N_8394,N_6860,N_7060);
and U8395 (N_8395,N_5957,N_6072);
or U8396 (N_8396,N_5191,N_5155);
or U8397 (N_8397,N_5440,N_6563);
and U8398 (N_8398,N_6066,N_7347);
and U8399 (N_8399,N_7095,N_5865);
nand U8400 (N_8400,N_5519,N_6005);
and U8401 (N_8401,N_6372,N_7177);
and U8402 (N_8402,N_5669,N_5851);
and U8403 (N_8403,N_5985,N_6859);
nand U8404 (N_8404,N_5848,N_5058);
nand U8405 (N_8405,N_6170,N_6148);
or U8406 (N_8406,N_6715,N_7445);
and U8407 (N_8407,N_7044,N_5524);
or U8408 (N_8408,N_5266,N_5522);
nor U8409 (N_8409,N_7464,N_6301);
nor U8410 (N_8410,N_6000,N_5680);
nand U8411 (N_8411,N_5665,N_5433);
nor U8412 (N_8412,N_5750,N_6754);
or U8413 (N_8413,N_7189,N_6297);
nor U8414 (N_8414,N_7236,N_5615);
or U8415 (N_8415,N_5561,N_6791);
and U8416 (N_8416,N_5869,N_7250);
nor U8417 (N_8417,N_7064,N_6144);
nand U8418 (N_8418,N_6135,N_6029);
xnor U8419 (N_8419,N_6321,N_6447);
nor U8420 (N_8420,N_7345,N_7323);
nor U8421 (N_8421,N_7240,N_5757);
nor U8422 (N_8422,N_7428,N_5777);
nor U8423 (N_8423,N_7369,N_5890);
nand U8424 (N_8424,N_6271,N_6840);
xor U8425 (N_8425,N_5917,N_7008);
and U8426 (N_8426,N_6479,N_5674);
or U8427 (N_8427,N_5996,N_5911);
nor U8428 (N_8428,N_5462,N_5401);
nand U8429 (N_8429,N_6198,N_6895);
xnor U8430 (N_8430,N_5070,N_6905);
nor U8431 (N_8431,N_5321,N_5276);
or U8432 (N_8432,N_7136,N_5299);
nand U8433 (N_8433,N_5582,N_7405);
or U8434 (N_8434,N_7207,N_5727);
and U8435 (N_8435,N_5059,N_7041);
nor U8436 (N_8436,N_5199,N_6496);
and U8437 (N_8437,N_5026,N_6804);
nand U8438 (N_8438,N_7235,N_6686);
nand U8439 (N_8439,N_7272,N_5806);
or U8440 (N_8440,N_6744,N_6929);
nand U8441 (N_8441,N_7360,N_5889);
nand U8442 (N_8442,N_6179,N_7023);
and U8443 (N_8443,N_5626,N_5998);
nor U8444 (N_8444,N_6822,N_6797);
or U8445 (N_8445,N_7027,N_7330);
nand U8446 (N_8446,N_6598,N_6407);
nor U8447 (N_8447,N_6062,N_5363);
and U8448 (N_8448,N_6187,N_6228);
nand U8449 (N_8449,N_7416,N_5393);
or U8450 (N_8450,N_7052,N_6893);
or U8451 (N_8451,N_7005,N_7153);
nor U8452 (N_8452,N_5358,N_5080);
and U8453 (N_8453,N_7440,N_5596);
and U8454 (N_8454,N_5340,N_5129);
nand U8455 (N_8455,N_5405,N_7029);
nand U8456 (N_8456,N_7183,N_5549);
and U8457 (N_8457,N_6036,N_6220);
and U8458 (N_8458,N_6223,N_6386);
and U8459 (N_8459,N_5990,N_5701);
nand U8460 (N_8460,N_7100,N_6626);
nor U8461 (N_8461,N_7447,N_6471);
and U8462 (N_8462,N_6451,N_5964);
nor U8463 (N_8463,N_7268,N_7167);
xnor U8464 (N_8464,N_7344,N_5197);
nand U8465 (N_8465,N_5424,N_6181);
nor U8466 (N_8466,N_6623,N_6854);
nand U8467 (N_8467,N_6363,N_6516);
nand U8468 (N_8468,N_5144,N_5739);
and U8469 (N_8469,N_5931,N_7342);
or U8470 (N_8470,N_7244,N_7310);
nor U8471 (N_8471,N_7197,N_6808);
and U8472 (N_8472,N_6436,N_6288);
or U8473 (N_8473,N_7365,N_6182);
nand U8474 (N_8474,N_7090,N_6595);
nand U8475 (N_8475,N_6293,N_5809);
and U8476 (N_8476,N_6888,N_7247);
or U8477 (N_8477,N_7398,N_5131);
nor U8478 (N_8478,N_7141,N_5092);
nor U8479 (N_8479,N_6166,N_6721);
nand U8480 (N_8480,N_5528,N_6190);
nor U8481 (N_8481,N_5797,N_7410);
or U8482 (N_8482,N_6635,N_5558);
or U8483 (N_8483,N_5579,N_7196);
nand U8484 (N_8484,N_5261,N_6096);
xor U8485 (N_8485,N_6201,N_6823);
and U8486 (N_8486,N_5182,N_5936);
or U8487 (N_8487,N_7089,N_5723);
and U8488 (N_8488,N_5337,N_7292);
nand U8489 (N_8489,N_5638,N_6441);
nor U8490 (N_8490,N_7367,N_5941);
nand U8491 (N_8491,N_5121,N_5342);
nand U8492 (N_8492,N_5736,N_5270);
nor U8493 (N_8493,N_7444,N_5263);
or U8494 (N_8494,N_5074,N_5448);
and U8495 (N_8495,N_7489,N_5065);
and U8496 (N_8496,N_5280,N_5237);
nand U8497 (N_8497,N_5995,N_5943);
or U8498 (N_8498,N_6826,N_6195);
nor U8499 (N_8499,N_6976,N_5500);
nand U8500 (N_8500,N_7078,N_5506);
or U8501 (N_8501,N_5754,N_5036);
xor U8502 (N_8502,N_5381,N_6403);
and U8503 (N_8503,N_5653,N_7357);
and U8504 (N_8504,N_5175,N_5947);
and U8505 (N_8505,N_6406,N_5602);
and U8506 (N_8506,N_5011,N_6240);
or U8507 (N_8507,N_5235,N_7434);
nor U8508 (N_8508,N_6128,N_5012);
nand U8509 (N_8509,N_6987,N_6217);
and U8510 (N_8510,N_5176,N_5722);
xor U8511 (N_8511,N_5371,N_5529);
xor U8512 (N_8512,N_6405,N_5341);
and U8513 (N_8513,N_6532,N_7309);
nand U8514 (N_8514,N_6514,N_6444);
nand U8515 (N_8515,N_7468,N_5178);
and U8516 (N_8516,N_5490,N_6493);
nand U8517 (N_8517,N_6304,N_6178);
nand U8518 (N_8518,N_5708,N_5819);
nor U8519 (N_8519,N_5535,N_5350);
nand U8520 (N_8520,N_5864,N_6663);
nor U8521 (N_8521,N_6845,N_6999);
and U8522 (N_8522,N_6013,N_6593);
nor U8523 (N_8523,N_5300,N_6545);
nand U8524 (N_8524,N_7329,N_5212);
nand U8525 (N_8525,N_7293,N_6616);
and U8526 (N_8526,N_6348,N_6043);
nand U8527 (N_8527,N_5394,N_5479);
nor U8528 (N_8528,N_7085,N_6787);
or U8529 (N_8529,N_5763,N_6466);
nor U8530 (N_8530,N_7426,N_7205);
and U8531 (N_8531,N_7163,N_5152);
or U8532 (N_8532,N_7404,N_5585);
xnor U8533 (N_8533,N_6904,N_5018);
nand U8534 (N_8534,N_7274,N_6606);
nand U8535 (N_8535,N_6336,N_5120);
xnor U8536 (N_8536,N_6777,N_6567);
and U8537 (N_8537,N_7304,N_5294);
nand U8538 (N_8538,N_6207,N_7322);
nor U8539 (N_8539,N_6192,N_7465);
and U8540 (N_8540,N_5735,N_7473);
or U8541 (N_8541,N_5083,N_7453);
or U8542 (N_8542,N_7162,N_6541);
nor U8543 (N_8543,N_5647,N_7000);
nor U8544 (N_8544,N_6855,N_5166);
or U8545 (N_8545,N_5009,N_6462);
nor U8546 (N_8546,N_7125,N_5502);
nor U8547 (N_8547,N_7022,N_5826);
or U8548 (N_8548,N_5333,N_5650);
or U8549 (N_8549,N_7382,N_5719);
nor U8550 (N_8550,N_5334,N_6656);
and U8551 (N_8551,N_5160,N_7024);
and U8552 (N_8552,N_7245,N_5951);
and U8553 (N_8553,N_5610,N_7104);
and U8554 (N_8554,N_7184,N_6858);
nor U8555 (N_8555,N_7391,N_5356);
nor U8556 (N_8556,N_6775,N_5173);
nand U8557 (N_8557,N_6422,N_6203);
nand U8558 (N_8558,N_6205,N_7435);
nand U8559 (N_8559,N_5725,N_7467);
nor U8560 (N_8560,N_6083,N_6200);
and U8561 (N_8561,N_6235,N_6837);
or U8562 (N_8562,N_7251,N_5171);
xor U8563 (N_8563,N_6989,N_5293);
nor U8564 (N_8564,N_6307,N_6263);
or U8565 (N_8565,N_5700,N_5344);
or U8566 (N_8566,N_5839,N_7388);
and U8567 (N_8567,N_7147,N_6710);
xor U8568 (N_8568,N_7004,N_6188);
xnor U8569 (N_8569,N_5751,N_6681);
nor U8570 (N_8570,N_7056,N_6955);
nor U8571 (N_8571,N_6194,N_6741);
and U8572 (N_8572,N_6199,N_5752);
nor U8573 (N_8573,N_6384,N_5195);
and U8574 (N_8574,N_5658,N_5833);
or U8575 (N_8575,N_6602,N_7199);
nand U8576 (N_8576,N_5567,N_5880);
and U8577 (N_8577,N_5804,N_7412);
nand U8578 (N_8578,N_6612,N_5520);
nand U8579 (N_8579,N_7152,N_6803);
and U8580 (N_8580,N_5593,N_5993);
nor U8581 (N_8581,N_6287,N_7463);
or U8582 (N_8582,N_6762,N_6146);
nor U8583 (N_8583,N_6571,N_5473);
nor U8584 (N_8584,N_6022,N_5397);
xor U8585 (N_8585,N_7411,N_6273);
or U8586 (N_8586,N_6902,N_5800);
nand U8587 (N_8587,N_7383,N_7361);
nand U8588 (N_8588,N_6917,N_6828);
nor U8589 (N_8589,N_5510,N_7009);
xor U8590 (N_8590,N_6443,N_5599);
nor U8591 (N_8591,N_5391,N_5172);
nor U8592 (N_8592,N_7348,N_5087);
nand U8593 (N_8593,N_5239,N_7277);
nor U8594 (N_8594,N_6245,N_7243);
and U8595 (N_8595,N_5022,N_6090);
or U8596 (N_8596,N_6933,N_5116);
and U8597 (N_8597,N_6442,N_6056);
nand U8598 (N_8598,N_6584,N_5570);
xor U8599 (N_8599,N_5877,N_5017);
nor U8600 (N_8600,N_7096,N_7316);
nor U8601 (N_8601,N_6963,N_5072);
nor U8602 (N_8602,N_5224,N_5162);
or U8603 (N_8603,N_6071,N_6687);
nand U8604 (N_8604,N_5138,N_5553);
or U8605 (N_8605,N_6896,N_7378);
nand U8606 (N_8606,N_7119,N_5874);
nor U8607 (N_8607,N_5207,N_5634);
nand U8608 (N_8608,N_6098,N_6617);
nor U8609 (N_8609,N_6604,N_5184);
or U8610 (N_8610,N_7185,N_6566);
xnor U8611 (N_8611,N_5468,N_5085);
and U8612 (N_8612,N_6185,N_5892);
xor U8613 (N_8613,N_5051,N_7418);
nand U8614 (N_8614,N_6174,N_5859);
xor U8615 (N_8615,N_7386,N_6094);
or U8616 (N_8616,N_6591,N_5149);
nor U8617 (N_8617,N_5305,N_5104);
and U8618 (N_8618,N_6353,N_5643);
nand U8619 (N_8619,N_6260,N_6186);
nor U8620 (N_8620,N_7206,N_6167);
and U8621 (N_8621,N_5523,N_6360);
or U8622 (N_8622,N_7070,N_6343);
nor U8623 (N_8623,N_5029,N_5642);
and U8624 (N_8624,N_6770,N_5346);
or U8625 (N_8625,N_6581,N_6760);
or U8626 (N_8626,N_5921,N_6935);
xor U8627 (N_8627,N_6134,N_5286);
nand U8628 (N_8628,N_6947,N_5923);
nor U8629 (N_8629,N_5339,N_6350);
nor U8630 (N_8630,N_5895,N_5667);
nor U8631 (N_8631,N_5205,N_5827);
nor U8632 (N_8632,N_6662,N_6037);
xnor U8633 (N_8633,N_5675,N_5838);
nand U8634 (N_8634,N_7038,N_5233);
xor U8635 (N_8635,N_6268,N_6279);
xor U8636 (N_8636,N_5855,N_6450);
nor U8637 (N_8637,N_5625,N_7227);
nand U8638 (N_8638,N_6956,N_6605);
xor U8639 (N_8639,N_7255,N_6368);
or U8640 (N_8640,N_5933,N_6930);
nor U8641 (N_8641,N_6229,N_6057);
nand U8642 (N_8642,N_7379,N_5682);
or U8643 (N_8643,N_5790,N_7142);
and U8644 (N_8644,N_5774,N_7121);
and U8645 (N_8645,N_6225,N_6219);
and U8646 (N_8646,N_6311,N_7478);
or U8647 (N_8647,N_5628,N_5960);
nand U8648 (N_8648,N_5084,N_6554);
or U8649 (N_8649,N_6849,N_6233);
and U8650 (N_8650,N_6983,N_5383);
or U8651 (N_8651,N_7230,N_5884);
and U8652 (N_8652,N_5188,N_5453);
and U8653 (N_8653,N_5690,N_6683);
nor U8654 (N_8654,N_7499,N_6049);
and U8655 (N_8655,N_6773,N_6130);
or U8656 (N_8656,N_6997,N_6365);
nand U8657 (N_8657,N_5357,N_6039);
nor U8658 (N_8658,N_5238,N_6677);
and U8659 (N_8659,N_6468,N_7380);
xnor U8660 (N_8660,N_6455,N_6732);
and U8661 (N_8661,N_5062,N_5609);
nor U8662 (N_8662,N_6048,N_5194);
or U8663 (N_8663,N_6041,N_7115);
nor U8664 (N_8664,N_7113,N_7127);
and U8665 (N_8665,N_6748,N_5920);
xor U8666 (N_8666,N_6918,N_6218);
xor U8667 (N_8667,N_5737,N_6592);
and U8668 (N_8668,N_5742,N_7249);
nor U8669 (N_8669,N_5604,N_5123);
nand U8670 (N_8670,N_6864,N_5262);
and U8671 (N_8671,N_6470,N_5862);
and U8672 (N_8672,N_6251,N_5772);
nor U8673 (N_8673,N_7131,N_6751);
or U8674 (N_8674,N_6234,N_6044);
or U8675 (N_8675,N_6089,N_5676);
nor U8676 (N_8676,N_5963,N_6073);
nor U8677 (N_8677,N_5109,N_6542);
and U8678 (N_8678,N_5480,N_5573);
nor U8679 (N_8679,N_7269,N_6900);
nor U8680 (N_8680,N_5099,N_6848);
nand U8681 (N_8681,N_5745,N_6259);
nand U8682 (N_8682,N_7296,N_6282);
nor U8683 (N_8683,N_5527,N_5613);
and U8684 (N_8684,N_5664,N_5580);
nor U8685 (N_8685,N_6278,N_6011);
nor U8686 (N_8686,N_6328,N_5948);
or U8687 (N_8687,N_6309,N_5020);
and U8688 (N_8688,N_6033,N_6764);
nand U8689 (N_8689,N_6028,N_6367);
nor U8690 (N_8690,N_6420,N_5703);
nor U8691 (N_8691,N_6325,N_7387);
xor U8692 (N_8692,N_6709,N_6660);
nand U8693 (N_8693,N_5958,N_6675);
and U8694 (N_8694,N_5010,N_5353);
nor U8695 (N_8695,N_6428,N_6712);
or U8696 (N_8696,N_6150,N_5306);
and U8697 (N_8697,N_5413,N_6650);
or U8698 (N_8698,N_7025,N_7012);
or U8699 (N_8699,N_6678,N_6892);
or U8700 (N_8700,N_7058,N_6557);
and U8701 (N_8701,N_5420,N_5969);
and U8702 (N_8702,N_6141,N_7375);
nand U8703 (N_8703,N_6115,N_5755);
nor U8704 (N_8704,N_7006,N_7073);
and U8705 (N_8705,N_5367,N_7208);
and U8706 (N_8706,N_6720,N_5154);
nand U8707 (N_8707,N_6645,N_6500);
or U8708 (N_8708,N_6990,N_5927);
nor U8709 (N_8709,N_7266,N_5760);
nor U8710 (N_8710,N_5858,N_6272);
nand U8711 (N_8711,N_5730,N_7017);
xor U8712 (N_8712,N_5828,N_7343);
nor U8713 (N_8713,N_5169,N_6536);
nor U8714 (N_8714,N_6018,N_6484);
and U8715 (N_8715,N_5483,N_6843);
and U8716 (N_8716,N_5515,N_5455);
and U8717 (N_8717,N_5661,N_6943);
or U8718 (N_8718,N_6069,N_6778);
and U8719 (N_8719,N_6392,N_5386);
or U8720 (N_8720,N_6483,N_6694);
nand U8721 (N_8721,N_7466,N_6944);
xnor U8722 (N_8722,N_7074,N_5446);
or U8723 (N_8723,N_6475,N_5909);
or U8724 (N_8724,N_5347,N_5460);
and U8725 (N_8725,N_6243,N_6221);
or U8726 (N_8726,N_6082,N_6323);
or U8727 (N_8727,N_7450,N_5134);
and U8728 (N_8728,N_6714,N_5412);
and U8729 (N_8729,N_6907,N_5603);
or U8730 (N_8730,N_6659,N_5159);
nor U8731 (N_8731,N_6431,N_5560);
or U8732 (N_8732,N_5282,N_7336);
nor U8733 (N_8733,N_5014,N_5876);
or U8734 (N_8734,N_5940,N_7143);
xor U8735 (N_8735,N_6193,N_5491);
or U8736 (N_8736,N_6794,N_6618);
nor U8737 (N_8737,N_6798,N_6774);
and U8738 (N_8738,N_6836,N_6706);
nand U8739 (N_8739,N_6410,N_6133);
and U8740 (N_8740,N_6021,N_5106);
nand U8741 (N_8741,N_5621,N_7441);
nor U8742 (N_8742,N_7129,N_6088);
nor U8743 (N_8743,N_6877,N_7496);
and U8744 (N_8744,N_6176,N_5788);
nand U8745 (N_8745,N_6883,N_6993);
nand U8746 (N_8746,N_7362,N_6334);
and U8747 (N_8747,N_6540,N_6163);
nor U8748 (N_8748,N_7327,N_7180);
nand U8749 (N_8749,N_6359,N_5852);
and U8750 (N_8750,N_7190,N_5247);
nor U8751 (N_8751,N_5203,N_7356);
nand U8752 (N_8752,N_6407,N_5492);
and U8753 (N_8753,N_7040,N_6854);
and U8754 (N_8754,N_6697,N_5412);
xor U8755 (N_8755,N_7434,N_5867);
xnor U8756 (N_8756,N_6579,N_6284);
and U8757 (N_8757,N_5897,N_7247);
and U8758 (N_8758,N_6912,N_7460);
and U8759 (N_8759,N_7129,N_7222);
or U8760 (N_8760,N_7293,N_5158);
xnor U8761 (N_8761,N_7300,N_6155);
nand U8762 (N_8762,N_5120,N_5738);
nand U8763 (N_8763,N_6807,N_6670);
nand U8764 (N_8764,N_5506,N_6566);
or U8765 (N_8765,N_5750,N_5337);
xnor U8766 (N_8766,N_5557,N_7063);
nor U8767 (N_8767,N_6665,N_6371);
nand U8768 (N_8768,N_7159,N_6143);
nand U8769 (N_8769,N_5823,N_6697);
nor U8770 (N_8770,N_6440,N_5878);
and U8771 (N_8771,N_5233,N_6511);
and U8772 (N_8772,N_5259,N_6659);
nor U8773 (N_8773,N_6943,N_7343);
nand U8774 (N_8774,N_5783,N_6790);
or U8775 (N_8775,N_6666,N_6787);
nand U8776 (N_8776,N_6852,N_6827);
and U8777 (N_8777,N_7437,N_6784);
and U8778 (N_8778,N_5668,N_6577);
nand U8779 (N_8779,N_6888,N_7023);
and U8780 (N_8780,N_6649,N_7392);
or U8781 (N_8781,N_6445,N_5730);
and U8782 (N_8782,N_5120,N_6265);
and U8783 (N_8783,N_5611,N_5153);
nor U8784 (N_8784,N_5458,N_6132);
and U8785 (N_8785,N_5636,N_6697);
nor U8786 (N_8786,N_7018,N_7221);
and U8787 (N_8787,N_5671,N_6038);
and U8788 (N_8788,N_6004,N_7263);
nor U8789 (N_8789,N_5570,N_5631);
and U8790 (N_8790,N_6150,N_7123);
nor U8791 (N_8791,N_7091,N_6282);
and U8792 (N_8792,N_7069,N_7009);
and U8793 (N_8793,N_6408,N_5450);
or U8794 (N_8794,N_5433,N_5839);
nor U8795 (N_8795,N_6292,N_7084);
and U8796 (N_8796,N_6875,N_6340);
or U8797 (N_8797,N_5921,N_7465);
xnor U8798 (N_8798,N_6938,N_6907);
and U8799 (N_8799,N_7431,N_5702);
and U8800 (N_8800,N_7331,N_6177);
xnor U8801 (N_8801,N_7359,N_5405);
and U8802 (N_8802,N_6502,N_5738);
nor U8803 (N_8803,N_5252,N_7083);
or U8804 (N_8804,N_6953,N_6858);
xor U8805 (N_8805,N_6023,N_5056);
or U8806 (N_8806,N_7110,N_5435);
and U8807 (N_8807,N_5198,N_5243);
xor U8808 (N_8808,N_7313,N_5669);
nand U8809 (N_8809,N_6550,N_7139);
nand U8810 (N_8810,N_5213,N_6184);
xor U8811 (N_8811,N_6094,N_5657);
and U8812 (N_8812,N_6488,N_7338);
and U8813 (N_8813,N_6250,N_7218);
nor U8814 (N_8814,N_5593,N_7041);
nor U8815 (N_8815,N_5146,N_5321);
nor U8816 (N_8816,N_5587,N_6042);
nor U8817 (N_8817,N_5708,N_6742);
and U8818 (N_8818,N_5732,N_5546);
nor U8819 (N_8819,N_5019,N_5955);
and U8820 (N_8820,N_5271,N_6495);
and U8821 (N_8821,N_7484,N_6867);
or U8822 (N_8822,N_6553,N_6701);
nor U8823 (N_8823,N_7123,N_7108);
nand U8824 (N_8824,N_7351,N_6731);
and U8825 (N_8825,N_6977,N_7107);
nor U8826 (N_8826,N_6487,N_6907);
nor U8827 (N_8827,N_6964,N_6175);
nor U8828 (N_8828,N_7434,N_5619);
nor U8829 (N_8829,N_5927,N_7288);
or U8830 (N_8830,N_7206,N_6012);
or U8831 (N_8831,N_7304,N_7456);
xor U8832 (N_8832,N_5981,N_7291);
or U8833 (N_8833,N_5668,N_5079);
nand U8834 (N_8834,N_7239,N_5736);
and U8835 (N_8835,N_7208,N_7417);
nand U8836 (N_8836,N_6408,N_7485);
and U8837 (N_8837,N_6838,N_5728);
nor U8838 (N_8838,N_6770,N_5096);
or U8839 (N_8839,N_5703,N_7038);
nand U8840 (N_8840,N_7055,N_6418);
and U8841 (N_8841,N_6556,N_5842);
nand U8842 (N_8842,N_6166,N_7246);
nand U8843 (N_8843,N_7102,N_5601);
nand U8844 (N_8844,N_5800,N_7446);
or U8845 (N_8845,N_7053,N_5764);
or U8846 (N_8846,N_5969,N_6443);
xnor U8847 (N_8847,N_7054,N_5650);
nand U8848 (N_8848,N_6658,N_6991);
nor U8849 (N_8849,N_5856,N_6667);
and U8850 (N_8850,N_5931,N_5642);
and U8851 (N_8851,N_5593,N_5421);
or U8852 (N_8852,N_5802,N_5805);
xnor U8853 (N_8853,N_7037,N_5121);
or U8854 (N_8854,N_5868,N_5062);
nand U8855 (N_8855,N_6445,N_5860);
nor U8856 (N_8856,N_6078,N_6456);
nand U8857 (N_8857,N_5244,N_5517);
and U8858 (N_8858,N_5415,N_6015);
and U8859 (N_8859,N_5076,N_5531);
nor U8860 (N_8860,N_6104,N_5949);
nand U8861 (N_8861,N_5381,N_7093);
and U8862 (N_8862,N_6357,N_5534);
xnor U8863 (N_8863,N_7381,N_6607);
and U8864 (N_8864,N_5804,N_5409);
nand U8865 (N_8865,N_6617,N_5387);
nor U8866 (N_8866,N_5828,N_5590);
or U8867 (N_8867,N_6922,N_5310);
nand U8868 (N_8868,N_5731,N_5192);
or U8869 (N_8869,N_5958,N_5814);
or U8870 (N_8870,N_6046,N_5440);
and U8871 (N_8871,N_7050,N_5639);
or U8872 (N_8872,N_7424,N_5015);
or U8873 (N_8873,N_6370,N_6296);
nor U8874 (N_8874,N_7347,N_5151);
and U8875 (N_8875,N_5893,N_5800);
and U8876 (N_8876,N_5273,N_5529);
nor U8877 (N_8877,N_6914,N_7229);
nor U8878 (N_8878,N_6326,N_5622);
nand U8879 (N_8879,N_7166,N_5598);
or U8880 (N_8880,N_6481,N_5354);
nand U8881 (N_8881,N_5597,N_5562);
nor U8882 (N_8882,N_7264,N_5718);
nand U8883 (N_8883,N_6535,N_6490);
and U8884 (N_8884,N_6241,N_5469);
or U8885 (N_8885,N_7420,N_5564);
and U8886 (N_8886,N_6210,N_5422);
and U8887 (N_8887,N_6901,N_6447);
and U8888 (N_8888,N_5154,N_5236);
nor U8889 (N_8889,N_7176,N_7112);
nor U8890 (N_8890,N_7310,N_5188);
or U8891 (N_8891,N_5765,N_5456);
nand U8892 (N_8892,N_5038,N_5284);
and U8893 (N_8893,N_5999,N_7417);
xnor U8894 (N_8894,N_6797,N_6949);
or U8895 (N_8895,N_6113,N_5965);
nand U8896 (N_8896,N_7089,N_5266);
or U8897 (N_8897,N_5087,N_6905);
nor U8898 (N_8898,N_7357,N_5334);
nand U8899 (N_8899,N_5839,N_6192);
nand U8900 (N_8900,N_6435,N_5447);
nand U8901 (N_8901,N_6214,N_7461);
nand U8902 (N_8902,N_7330,N_7245);
nor U8903 (N_8903,N_5448,N_6933);
and U8904 (N_8904,N_6465,N_6037);
and U8905 (N_8905,N_6998,N_6843);
nand U8906 (N_8906,N_5957,N_5381);
nand U8907 (N_8907,N_5731,N_6403);
nand U8908 (N_8908,N_7184,N_6216);
nor U8909 (N_8909,N_6953,N_6248);
nor U8910 (N_8910,N_6915,N_6593);
or U8911 (N_8911,N_6760,N_5485);
nor U8912 (N_8912,N_6715,N_7145);
or U8913 (N_8913,N_6087,N_5443);
nor U8914 (N_8914,N_6923,N_7218);
xor U8915 (N_8915,N_5231,N_6938);
and U8916 (N_8916,N_5725,N_6837);
nand U8917 (N_8917,N_5946,N_5258);
xnor U8918 (N_8918,N_5149,N_7226);
nand U8919 (N_8919,N_5641,N_5069);
nand U8920 (N_8920,N_5899,N_5244);
nor U8921 (N_8921,N_5638,N_6598);
nand U8922 (N_8922,N_6058,N_6701);
and U8923 (N_8923,N_6247,N_6402);
xor U8924 (N_8924,N_6297,N_5153);
and U8925 (N_8925,N_5022,N_5589);
nor U8926 (N_8926,N_7187,N_6398);
xor U8927 (N_8927,N_5064,N_7454);
nor U8928 (N_8928,N_5229,N_5114);
nor U8929 (N_8929,N_6203,N_5026);
xor U8930 (N_8930,N_5052,N_5218);
nor U8931 (N_8931,N_5406,N_5124);
nand U8932 (N_8932,N_6418,N_5502);
nor U8933 (N_8933,N_5165,N_7230);
or U8934 (N_8934,N_6326,N_5868);
nor U8935 (N_8935,N_6828,N_5478);
or U8936 (N_8936,N_5504,N_5204);
nor U8937 (N_8937,N_6066,N_6316);
nand U8938 (N_8938,N_5164,N_5660);
xor U8939 (N_8939,N_5212,N_6860);
and U8940 (N_8940,N_5246,N_5203);
or U8941 (N_8941,N_6350,N_5331);
nor U8942 (N_8942,N_7320,N_7378);
nand U8943 (N_8943,N_6430,N_7063);
or U8944 (N_8944,N_5380,N_5410);
nand U8945 (N_8945,N_6559,N_6157);
nor U8946 (N_8946,N_6905,N_5708);
and U8947 (N_8947,N_5404,N_6799);
and U8948 (N_8948,N_6242,N_7117);
nand U8949 (N_8949,N_5883,N_5436);
and U8950 (N_8950,N_6037,N_6979);
nand U8951 (N_8951,N_6665,N_6267);
nand U8952 (N_8952,N_7017,N_5624);
and U8953 (N_8953,N_6545,N_5872);
xor U8954 (N_8954,N_6002,N_5636);
nor U8955 (N_8955,N_5535,N_7144);
and U8956 (N_8956,N_7237,N_7221);
nor U8957 (N_8957,N_5769,N_6168);
nor U8958 (N_8958,N_5966,N_7225);
nand U8959 (N_8959,N_6614,N_6625);
xnor U8960 (N_8960,N_5772,N_5045);
nand U8961 (N_8961,N_6052,N_5638);
or U8962 (N_8962,N_5807,N_7106);
nor U8963 (N_8963,N_7475,N_5544);
or U8964 (N_8964,N_6505,N_5879);
or U8965 (N_8965,N_6047,N_5226);
nor U8966 (N_8966,N_7238,N_6314);
and U8967 (N_8967,N_5332,N_6163);
nor U8968 (N_8968,N_6397,N_6138);
and U8969 (N_8969,N_7499,N_5058);
nand U8970 (N_8970,N_7486,N_6373);
nor U8971 (N_8971,N_6888,N_5885);
nor U8972 (N_8972,N_5340,N_7037);
or U8973 (N_8973,N_7474,N_7370);
or U8974 (N_8974,N_6835,N_7018);
nor U8975 (N_8975,N_5738,N_5877);
and U8976 (N_8976,N_5356,N_6994);
xor U8977 (N_8977,N_6701,N_6298);
or U8978 (N_8978,N_6631,N_5229);
or U8979 (N_8979,N_7181,N_5599);
and U8980 (N_8980,N_7227,N_7411);
nor U8981 (N_8981,N_5393,N_5496);
and U8982 (N_8982,N_5515,N_5690);
or U8983 (N_8983,N_5474,N_6393);
or U8984 (N_8984,N_6616,N_6147);
or U8985 (N_8985,N_5975,N_6382);
nand U8986 (N_8986,N_6100,N_6182);
or U8987 (N_8987,N_6043,N_6809);
nand U8988 (N_8988,N_5823,N_6628);
and U8989 (N_8989,N_5203,N_6958);
nor U8990 (N_8990,N_6764,N_7218);
nand U8991 (N_8991,N_7111,N_6992);
or U8992 (N_8992,N_6184,N_6747);
and U8993 (N_8993,N_6933,N_5729);
or U8994 (N_8994,N_5706,N_7038);
or U8995 (N_8995,N_5221,N_6789);
nor U8996 (N_8996,N_5258,N_6969);
nand U8997 (N_8997,N_7434,N_6858);
or U8998 (N_8998,N_5911,N_5514);
nor U8999 (N_8999,N_7432,N_5887);
and U9000 (N_9000,N_5863,N_6041);
and U9001 (N_9001,N_7323,N_7409);
nor U9002 (N_9002,N_6903,N_7303);
or U9003 (N_9003,N_6749,N_7011);
nand U9004 (N_9004,N_5513,N_7047);
nand U9005 (N_9005,N_7490,N_5983);
or U9006 (N_9006,N_6741,N_7393);
nand U9007 (N_9007,N_6953,N_6600);
xnor U9008 (N_9008,N_5529,N_6659);
nor U9009 (N_9009,N_5637,N_5166);
xnor U9010 (N_9010,N_5239,N_5021);
nand U9011 (N_9011,N_7337,N_6663);
nand U9012 (N_9012,N_6817,N_5952);
nor U9013 (N_9013,N_5603,N_6665);
or U9014 (N_9014,N_6689,N_6389);
nand U9015 (N_9015,N_5859,N_5033);
xnor U9016 (N_9016,N_5947,N_5700);
and U9017 (N_9017,N_7394,N_5921);
or U9018 (N_9018,N_5912,N_7002);
nor U9019 (N_9019,N_6242,N_6726);
nor U9020 (N_9020,N_5256,N_6761);
nand U9021 (N_9021,N_5995,N_6412);
or U9022 (N_9022,N_5539,N_6898);
nor U9023 (N_9023,N_6766,N_6638);
and U9024 (N_9024,N_6951,N_7049);
nor U9025 (N_9025,N_7474,N_5051);
and U9026 (N_9026,N_6828,N_7326);
or U9027 (N_9027,N_7322,N_5961);
and U9028 (N_9028,N_6731,N_6354);
nor U9029 (N_9029,N_5789,N_5219);
nand U9030 (N_9030,N_5823,N_7282);
and U9031 (N_9031,N_6823,N_7031);
or U9032 (N_9032,N_6048,N_7359);
and U9033 (N_9033,N_7325,N_5775);
nor U9034 (N_9034,N_6850,N_6397);
and U9035 (N_9035,N_6443,N_7224);
nor U9036 (N_9036,N_5195,N_7192);
nand U9037 (N_9037,N_6240,N_6735);
nand U9038 (N_9038,N_5371,N_5913);
or U9039 (N_9039,N_5000,N_5589);
nor U9040 (N_9040,N_5720,N_5034);
and U9041 (N_9041,N_5387,N_5143);
nand U9042 (N_9042,N_5056,N_6708);
and U9043 (N_9043,N_5090,N_5335);
nand U9044 (N_9044,N_7259,N_6512);
or U9045 (N_9045,N_5896,N_6280);
and U9046 (N_9046,N_6063,N_5302);
or U9047 (N_9047,N_5007,N_6695);
and U9048 (N_9048,N_5399,N_5320);
nor U9049 (N_9049,N_6355,N_5214);
or U9050 (N_9050,N_6053,N_6192);
and U9051 (N_9051,N_5553,N_6212);
nand U9052 (N_9052,N_5539,N_6268);
and U9053 (N_9053,N_5363,N_7178);
or U9054 (N_9054,N_5064,N_6314);
or U9055 (N_9055,N_6083,N_6116);
or U9056 (N_9056,N_7087,N_7290);
xor U9057 (N_9057,N_7433,N_6039);
or U9058 (N_9058,N_6192,N_6244);
or U9059 (N_9059,N_5921,N_7114);
nor U9060 (N_9060,N_6972,N_7481);
nand U9061 (N_9061,N_6845,N_6045);
and U9062 (N_9062,N_6364,N_5428);
nor U9063 (N_9063,N_5256,N_5044);
nand U9064 (N_9064,N_6218,N_5601);
nand U9065 (N_9065,N_7227,N_6253);
xor U9066 (N_9066,N_5396,N_6856);
xnor U9067 (N_9067,N_6224,N_5555);
xnor U9068 (N_9068,N_6420,N_5890);
nand U9069 (N_9069,N_6978,N_5815);
and U9070 (N_9070,N_6051,N_7030);
nor U9071 (N_9071,N_7098,N_5098);
nor U9072 (N_9072,N_5982,N_6575);
and U9073 (N_9073,N_5069,N_6174);
and U9074 (N_9074,N_5685,N_6230);
nor U9075 (N_9075,N_7143,N_6590);
or U9076 (N_9076,N_6165,N_5445);
and U9077 (N_9077,N_6016,N_7279);
nor U9078 (N_9078,N_6724,N_5177);
and U9079 (N_9079,N_5102,N_6791);
nand U9080 (N_9080,N_5170,N_5926);
and U9081 (N_9081,N_6062,N_5725);
or U9082 (N_9082,N_6328,N_7385);
nor U9083 (N_9083,N_6008,N_5918);
and U9084 (N_9084,N_5483,N_6410);
and U9085 (N_9085,N_7401,N_5748);
nor U9086 (N_9086,N_5798,N_7105);
or U9087 (N_9087,N_5368,N_5390);
nand U9088 (N_9088,N_5537,N_5137);
nand U9089 (N_9089,N_7278,N_5109);
or U9090 (N_9090,N_7159,N_6798);
and U9091 (N_9091,N_7283,N_6251);
or U9092 (N_9092,N_6752,N_5590);
or U9093 (N_9093,N_6920,N_7100);
or U9094 (N_9094,N_5194,N_5491);
or U9095 (N_9095,N_5143,N_6200);
or U9096 (N_9096,N_6126,N_6594);
nor U9097 (N_9097,N_5790,N_6717);
or U9098 (N_9098,N_6723,N_7042);
and U9099 (N_9099,N_5696,N_5531);
nand U9100 (N_9100,N_5718,N_6475);
nor U9101 (N_9101,N_6770,N_6858);
or U9102 (N_9102,N_6542,N_6069);
nor U9103 (N_9103,N_5564,N_6392);
nor U9104 (N_9104,N_5653,N_5303);
nor U9105 (N_9105,N_7156,N_6094);
nand U9106 (N_9106,N_6952,N_7122);
and U9107 (N_9107,N_5143,N_6323);
nor U9108 (N_9108,N_5392,N_7060);
nand U9109 (N_9109,N_5056,N_7461);
and U9110 (N_9110,N_6102,N_7331);
and U9111 (N_9111,N_6728,N_6306);
or U9112 (N_9112,N_7033,N_6760);
nand U9113 (N_9113,N_6339,N_5795);
and U9114 (N_9114,N_5196,N_6627);
or U9115 (N_9115,N_6964,N_6319);
nand U9116 (N_9116,N_5803,N_6159);
nor U9117 (N_9117,N_5173,N_5400);
or U9118 (N_9118,N_6439,N_7302);
or U9119 (N_9119,N_5126,N_6875);
nor U9120 (N_9120,N_5538,N_7257);
and U9121 (N_9121,N_7103,N_6421);
xor U9122 (N_9122,N_6399,N_6430);
nor U9123 (N_9123,N_5510,N_6036);
nand U9124 (N_9124,N_6199,N_7165);
nor U9125 (N_9125,N_6643,N_5990);
or U9126 (N_9126,N_6498,N_6235);
nor U9127 (N_9127,N_5885,N_5660);
and U9128 (N_9128,N_6789,N_7018);
nand U9129 (N_9129,N_6042,N_6803);
and U9130 (N_9130,N_6414,N_6118);
and U9131 (N_9131,N_6872,N_6326);
or U9132 (N_9132,N_5442,N_5732);
and U9133 (N_9133,N_5869,N_6965);
nor U9134 (N_9134,N_6453,N_5401);
nor U9135 (N_9135,N_5355,N_7265);
nand U9136 (N_9136,N_5675,N_6505);
and U9137 (N_9137,N_5053,N_7473);
nand U9138 (N_9138,N_5949,N_7073);
nor U9139 (N_9139,N_6123,N_6887);
nand U9140 (N_9140,N_5823,N_6390);
or U9141 (N_9141,N_6392,N_5890);
or U9142 (N_9142,N_6663,N_7086);
nand U9143 (N_9143,N_6136,N_7077);
nor U9144 (N_9144,N_7062,N_5512);
nor U9145 (N_9145,N_5616,N_6333);
nand U9146 (N_9146,N_6965,N_6858);
nand U9147 (N_9147,N_5530,N_7375);
nor U9148 (N_9148,N_7230,N_6221);
xor U9149 (N_9149,N_5287,N_5480);
nor U9150 (N_9150,N_6203,N_5525);
nor U9151 (N_9151,N_6063,N_6202);
or U9152 (N_9152,N_5236,N_6406);
nand U9153 (N_9153,N_5285,N_5902);
nor U9154 (N_9154,N_6464,N_6482);
or U9155 (N_9155,N_6062,N_5201);
xor U9156 (N_9156,N_6565,N_5973);
nand U9157 (N_9157,N_5624,N_5186);
or U9158 (N_9158,N_6823,N_6568);
and U9159 (N_9159,N_5680,N_6219);
nand U9160 (N_9160,N_6990,N_5665);
nand U9161 (N_9161,N_7433,N_6998);
nor U9162 (N_9162,N_5874,N_5777);
and U9163 (N_9163,N_5978,N_6334);
or U9164 (N_9164,N_7363,N_6648);
nor U9165 (N_9165,N_5720,N_6716);
or U9166 (N_9166,N_7469,N_5634);
and U9167 (N_9167,N_5846,N_7400);
and U9168 (N_9168,N_5493,N_6403);
or U9169 (N_9169,N_6579,N_6721);
or U9170 (N_9170,N_5005,N_7490);
and U9171 (N_9171,N_5569,N_6990);
xnor U9172 (N_9172,N_7427,N_5885);
nand U9173 (N_9173,N_7206,N_7320);
or U9174 (N_9174,N_5266,N_7464);
nor U9175 (N_9175,N_6077,N_5228);
and U9176 (N_9176,N_7110,N_7079);
nor U9177 (N_9177,N_6426,N_5821);
nand U9178 (N_9178,N_6837,N_7257);
and U9179 (N_9179,N_7218,N_5918);
xor U9180 (N_9180,N_7299,N_5554);
or U9181 (N_9181,N_5835,N_6737);
and U9182 (N_9182,N_5516,N_5272);
nand U9183 (N_9183,N_5784,N_7067);
nor U9184 (N_9184,N_5614,N_6112);
xor U9185 (N_9185,N_6453,N_6390);
or U9186 (N_9186,N_7049,N_6745);
or U9187 (N_9187,N_7494,N_5672);
and U9188 (N_9188,N_6832,N_7464);
and U9189 (N_9189,N_7147,N_5435);
nand U9190 (N_9190,N_5753,N_7094);
nand U9191 (N_9191,N_6264,N_7369);
and U9192 (N_9192,N_6948,N_6800);
nor U9193 (N_9193,N_5141,N_6833);
or U9194 (N_9194,N_6455,N_7033);
nor U9195 (N_9195,N_7444,N_5424);
and U9196 (N_9196,N_7416,N_6711);
nand U9197 (N_9197,N_5745,N_6400);
nor U9198 (N_9198,N_5968,N_5618);
and U9199 (N_9199,N_5305,N_5592);
and U9200 (N_9200,N_5195,N_5240);
xor U9201 (N_9201,N_7365,N_5517);
xnor U9202 (N_9202,N_5904,N_7051);
and U9203 (N_9203,N_7338,N_5574);
or U9204 (N_9204,N_6972,N_5091);
and U9205 (N_9205,N_6880,N_6562);
and U9206 (N_9206,N_7320,N_6519);
nand U9207 (N_9207,N_6420,N_7412);
nand U9208 (N_9208,N_5025,N_5351);
or U9209 (N_9209,N_5471,N_6677);
or U9210 (N_9210,N_6977,N_6891);
and U9211 (N_9211,N_5807,N_5135);
nand U9212 (N_9212,N_7127,N_6492);
nand U9213 (N_9213,N_5890,N_5566);
and U9214 (N_9214,N_7089,N_5102);
nand U9215 (N_9215,N_6366,N_5630);
and U9216 (N_9216,N_6177,N_6980);
or U9217 (N_9217,N_7237,N_5787);
nand U9218 (N_9218,N_6700,N_6368);
nand U9219 (N_9219,N_5383,N_6396);
nand U9220 (N_9220,N_6516,N_5047);
and U9221 (N_9221,N_6834,N_5599);
xor U9222 (N_9222,N_5493,N_5763);
nor U9223 (N_9223,N_7084,N_6696);
nor U9224 (N_9224,N_5375,N_6065);
nand U9225 (N_9225,N_5245,N_7482);
nand U9226 (N_9226,N_5748,N_5422);
and U9227 (N_9227,N_5921,N_6640);
nor U9228 (N_9228,N_5875,N_7354);
and U9229 (N_9229,N_6872,N_7242);
or U9230 (N_9230,N_5118,N_5861);
and U9231 (N_9231,N_6476,N_5538);
xnor U9232 (N_9232,N_6955,N_5722);
nand U9233 (N_9233,N_7138,N_6977);
nor U9234 (N_9234,N_5435,N_6471);
nor U9235 (N_9235,N_6558,N_6559);
nor U9236 (N_9236,N_7199,N_6175);
nand U9237 (N_9237,N_6365,N_5981);
nor U9238 (N_9238,N_6435,N_6327);
nor U9239 (N_9239,N_6280,N_6920);
or U9240 (N_9240,N_6977,N_6256);
nand U9241 (N_9241,N_6801,N_5708);
nand U9242 (N_9242,N_5524,N_6910);
or U9243 (N_9243,N_6378,N_5810);
xor U9244 (N_9244,N_7412,N_6641);
nor U9245 (N_9245,N_7258,N_5175);
and U9246 (N_9246,N_6863,N_7007);
nand U9247 (N_9247,N_6819,N_7193);
and U9248 (N_9248,N_6448,N_5524);
or U9249 (N_9249,N_6364,N_6607);
or U9250 (N_9250,N_5951,N_5997);
nand U9251 (N_9251,N_5014,N_6064);
and U9252 (N_9252,N_6488,N_5078);
nor U9253 (N_9253,N_5179,N_6813);
nor U9254 (N_9254,N_5003,N_5183);
and U9255 (N_9255,N_6043,N_6495);
or U9256 (N_9256,N_7468,N_6841);
or U9257 (N_9257,N_5153,N_5496);
or U9258 (N_9258,N_5136,N_5472);
or U9259 (N_9259,N_6812,N_6517);
nand U9260 (N_9260,N_7285,N_6506);
nand U9261 (N_9261,N_5963,N_5506);
or U9262 (N_9262,N_7227,N_6361);
and U9263 (N_9263,N_5037,N_7282);
or U9264 (N_9264,N_5045,N_7416);
nor U9265 (N_9265,N_6245,N_6513);
nand U9266 (N_9266,N_6387,N_7306);
nor U9267 (N_9267,N_5404,N_7203);
nor U9268 (N_9268,N_5349,N_7417);
or U9269 (N_9269,N_5004,N_6707);
and U9270 (N_9270,N_5240,N_6265);
nor U9271 (N_9271,N_5720,N_7409);
and U9272 (N_9272,N_7354,N_6593);
or U9273 (N_9273,N_5769,N_5365);
nand U9274 (N_9274,N_5266,N_5264);
nor U9275 (N_9275,N_6698,N_5621);
and U9276 (N_9276,N_6008,N_5820);
nor U9277 (N_9277,N_7468,N_7240);
nand U9278 (N_9278,N_7462,N_5455);
xnor U9279 (N_9279,N_5473,N_7299);
nor U9280 (N_9280,N_5456,N_6622);
nand U9281 (N_9281,N_5249,N_5283);
or U9282 (N_9282,N_5793,N_7373);
nor U9283 (N_9283,N_6455,N_7462);
xor U9284 (N_9284,N_5829,N_5533);
nor U9285 (N_9285,N_5263,N_5606);
nand U9286 (N_9286,N_7186,N_6807);
and U9287 (N_9287,N_6862,N_6012);
or U9288 (N_9288,N_5539,N_6832);
nand U9289 (N_9289,N_7185,N_6463);
or U9290 (N_9290,N_5667,N_6519);
or U9291 (N_9291,N_5317,N_5250);
nand U9292 (N_9292,N_6933,N_6986);
or U9293 (N_9293,N_5814,N_5260);
or U9294 (N_9294,N_6059,N_6588);
nand U9295 (N_9295,N_6029,N_7052);
nand U9296 (N_9296,N_6197,N_5993);
or U9297 (N_9297,N_6629,N_6437);
nor U9298 (N_9298,N_5280,N_5330);
and U9299 (N_9299,N_6816,N_6198);
and U9300 (N_9300,N_6824,N_7118);
and U9301 (N_9301,N_6366,N_6957);
and U9302 (N_9302,N_5570,N_7095);
xnor U9303 (N_9303,N_6825,N_6141);
or U9304 (N_9304,N_5249,N_6716);
and U9305 (N_9305,N_6932,N_6914);
nand U9306 (N_9306,N_6199,N_5539);
nand U9307 (N_9307,N_5513,N_6819);
or U9308 (N_9308,N_6766,N_5287);
and U9309 (N_9309,N_6344,N_7397);
nand U9310 (N_9310,N_6651,N_7356);
or U9311 (N_9311,N_5026,N_7347);
xor U9312 (N_9312,N_5333,N_6925);
or U9313 (N_9313,N_6839,N_6456);
xor U9314 (N_9314,N_5882,N_5563);
and U9315 (N_9315,N_7020,N_7060);
nor U9316 (N_9316,N_6966,N_5429);
nand U9317 (N_9317,N_5302,N_7009);
or U9318 (N_9318,N_7245,N_6740);
nor U9319 (N_9319,N_5164,N_5559);
and U9320 (N_9320,N_6654,N_7118);
nand U9321 (N_9321,N_5692,N_7429);
or U9322 (N_9322,N_6657,N_5677);
nor U9323 (N_9323,N_7218,N_6584);
and U9324 (N_9324,N_5752,N_6277);
xor U9325 (N_9325,N_6053,N_5101);
or U9326 (N_9326,N_6373,N_5547);
nor U9327 (N_9327,N_6050,N_5751);
or U9328 (N_9328,N_6614,N_6896);
nand U9329 (N_9329,N_6323,N_5487);
or U9330 (N_9330,N_6774,N_7036);
or U9331 (N_9331,N_6424,N_5074);
or U9332 (N_9332,N_7432,N_6289);
nor U9333 (N_9333,N_5446,N_5411);
xnor U9334 (N_9334,N_7037,N_5491);
xor U9335 (N_9335,N_5282,N_5286);
or U9336 (N_9336,N_5582,N_6721);
xnor U9337 (N_9337,N_6023,N_6555);
nand U9338 (N_9338,N_7228,N_7034);
xor U9339 (N_9339,N_5926,N_7129);
nor U9340 (N_9340,N_5095,N_6762);
nand U9341 (N_9341,N_6405,N_7326);
nand U9342 (N_9342,N_7459,N_7189);
xor U9343 (N_9343,N_5479,N_6883);
nand U9344 (N_9344,N_6627,N_6941);
and U9345 (N_9345,N_7403,N_6038);
or U9346 (N_9346,N_5799,N_7400);
nand U9347 (N_9347,N_6717,N_6570);
nor U9348 (N_9348,N_6611,N_5107);
nor U9349 (N_9349,N_5674,N_6337);
or U9350 (N_9350,N_5514,N_7176);
nand U9351 (N_9351,N_5577,N_5326);
xnor U9352 (N_9352,N_7231,N_5984);
nor U9353 (N_9353,N_5422,N_6319);
nand U9354 (N_9354,N_6781,N_5903);
or U9355 (N_9355,N_5565,N_5148);
nor U9356 (N_9356,N_5304,N_7120);
and U9357 (N_9357,N_6755,N_5387);
nand U9358 (N_9358,N_5440,N_5053);
nand U9359 (N_9359,N_6888,N_6088);
or U9360 (N_9360,N_7262,N_5521);
or U9361 (N_9361,N_6838,N_6811);
nand U9362 (N_9362,N_6117,N_6286);
nand U9363 (N_9363,N_6666,N_6835);
nand U9364 (N_9364,N_5132,N_5292);
nor U9365 (N_9365,N_6675,N_7411);
nand U9366 (N_9366,N_6932,N_7355);
xor U9367 (N_9367,N_6007,N_6154);
nand U9368 (N_9368,N_7465,N_6775);
and U9369 (N_9369,N_6222,N_7018);
or U9370 (N_9370,N_5727,N_5399);
nand U9371 (N_9371,N_6767,N_6334);
nand U9372 (N_9372,N_6433,N_5859);
xnor U9373 (N_9373,N_6933,N_5537);
nor U9374 (N_9374,N_5803,N_6333);
and U9375 (N_9375,N_5874,N_5080);
or U9376 (N_9376,N_6691,N_5636);
and U9377 (N_9377,N_5571,N_6044);
nand U9378 (N_9378,N_6364,N_5122);
nor U9379 (N_9379,N_6087,N_6421);
xor U9380 (N_9380,N_5502,N_6247);
and U9381 (N_9381,N_6056,N_6801);
nand U9382 (N_9382,N_7458,N_7238);
and U9383 (N_9383,N_6437,N_7181);
and U9384 (N_9384,N_6583,N_6619);
and U9385 (N_9385,N_7111,N_7071);
nor U9386 (N_9386,N_5114,N_5773);
and U9387 (N_9387,N_7442,N_7484);
and U9388 (N_9388,N_6527,N_6493);
and U9389 (N_9389,N_5888,N_6084);
and U9390 (N_9390,N_7026,N_6062);
and U9391 (N_9391,N_6182,N_6330);
and U9392 (N_9392,N_7048,N_7002);
and U9393 (N_9393,N_6959,N_7365);
or U9394 (N_9394,N_5877,N_6138);
and U9395 (N_9395,N_6892,N_5891);
nor U9396 (N_9396,N_5682,N_5789);
and U9397 (N_9397,N_6177,N_5852);
nor U9398 (N_9398,N_6001,N_6761);
xnor U9399 (N_9399,N_7121,N_7497);
or U9400 (N_9400,N_6702,N_6763);
nand U9401 (N_9401,N_6623,N_6406);
xnor U9402 (N_9402,N_5812,N_6461);
nand U9403 (N_9403,N_6826,N_6236);
nor U9404 (N_9404,N_7496,N_7208);
nor U9405 (N_9405,N_5286,N_7081);
nor U9406 (N_9406,N_5172,N_7492);
nor U9407 (N_9407,N_7151,N_5800);
nand U9408 (N_9408,N_5488,N_6456);
or U9409 (N_9409,N_5691,N_5548);
or U9410 (N_9410,N_6389,N_7421);
and U9411 (N_9411,N_7153,N_6889);
or U9412 (N_9412,N_7444,N_6607);
nor U9413 (N_9413,N_7339,N_6541);
nand U9414 (N_9414,N_5143,N_6472);
xnor U9415 (N_9415,N_7332,N_5390);
and U9416 (N_9416,N_6679,N_5268);
or U9417 (N_9417,N_5517,N_7068);
or U9418 (N_9418,N_5068,N_5231);
nand U9419 (N_9419,N_5737,N_5376);
and U9420 (N_9420,N_6986,N_7355);
and U9421 (N_9421,N_6231,N_6846);
or U9422 (N_9422,N_7082,N_5559);
nor U9423 (N_9423,N_5995,N_5090);
and U9424 (N_9424,N_5231,N_6001);
nand U9425 (N_9425,N_5494,N_5263);
or U9426 (N_9426,N_6940,N_5663);
and U9427 (N_9427,N_7485,N_6444);
or U9428 (N_9428,N_5786,N_6255);
or U9429 (N_9429,N_5920,N_7062);
xor U9430 (N_9430,N_5837,N_7097);
nor U9431 (N_9431,N_5123,N_6991);
nand U9432 (N_9432,N_7040,N_7399);
or U9433 (N_9433,N_6697,N_6223);
and U9434 (N_9434,N_6578,N_7452);
and U9435 (N_9435,N_6515,N_5704);
or U9436 (N_9436,N_5770,N_6372);
nand U9437 (N_9437,N_5557,N_7207);
nor U9438 (N_9438,N_5373,N_6797);
and U9439 (N_9439,N_6572,N_5548);
and U9440 (N_9440,N_5636,N_6462);
nand U9441 (N_9441,N_5577,N_6691);
nor U9442 (N_9442,N_5899,N_6665);
or U9443 (N_9443,N_7107,N_7438);
nor U9444 (N_9444,N_5233,N_6608);
or U9445 (N_9445,N_6758,N_6873);
nand U9446 (N_9446,N_5871,N_6087);
and U9447 (N_9447,N_6677,N_5773);
or U9448 (N_9448,N_7304,N_5133);
nor U9449 (N_9449,N_7231,N_5040);
or U9450 (N_9450,N_5857,N_6893);
or U9451 (N_9451,N_6025,N_6140);
and U9452 (N_9452,N_5742,N_6881);
or U9453 (N_9453,N_6308,N_7013);
and U9454 (N_9454,N_5329,N_6961);
or U9455 (N_9455,N_5516,N_6194);
and U9456 (N_9456,N_6662,N_6613);
nor U9457 (N_9457,N_5413,N_5252);
nand U9458 (N_9458,N_7480,N_5642);
nor U9459 (N_9459,N_5729,N_6935);
and U9460 (N_9460,N_7209,N_7475);
nor U9461 (N_9461,N_5908,N_5970);
nand U9462 (N_9462,N_5895,N_6543);
nor U9463 (N_9463,N_6281,N_7028);
nor U9464 (N_9464,N_6370,N_5870);
nand U9465 (N_9465,N_6203,N_7131);
and U9466 (N_9466,N_5060,N_7181);
nand U9467 (N_9467,N_5713,N_5718);
and U9468 (N_9468,N_7246,N_5791);
nor U9469 (N_9469,N_7111,N_5865);
or U9470 (N_9470,N_7215,N_6860);
nor U9471 (N_9471,N_5465,N_6251);
or U9472 (N_9472,N_5920,N_6226);
nand U9473 (N_9473,N_5765,N_6084);
nor U9474 (N_9474,N_5167,N_5638);
and U9475 (N_9475,N_7129,N_6337);
and U9476 (N_9476,N_5328,N_5405);
nand U9477 (N_9477,N_7365,N_6772);
nand U9478 (N_9478,N_5578,N_5626);
and U9479 (N_9479,N_6430,N_5469);
nand U9480 (N_9480,N_5350,N_5983);
nor U9481 (N_9481,N_5962,N_7391);
nand U9482 (N_9482,N_7412,N_6699);
nand U9483 (N_9483,N_7328,N_5171);
nand U9484 (N_9484,N_6622,N_6050);
and U9485 (N_9485,N_5520,N_6547);
or U9486 (N_9486,N_7324,N_6814);
or U9487 (N_9487,N_5809,N_5618);
and U9488 (N_9488,N_6571,N_5300);
and U9489 (N_9489,N_6569,N_6025);
nand U9490 (N_9490,N_6861,N_6506);
nand U9491 (N_9491,N_5193,N_7470);
and U9492 (N_9492,N_5699,N_5618);
nand U9493 (N_9493,N_5224,N_7337);
and U9494 (N_9494,N_6858,N_6409);
or U9495 (N_9495,N_7352,N_5937);
nor U9496 (N_9496,N_6029,N_6605);
nand U9497 (N_9497,N_7034,N_5878);
xnor U9498 (N_9498,N_6845,N_5391);
nor U9499 (N_9499,N_6818,N_5802);
and U9500 (N_9500,N_5809,N_7105);
or U9501 (N_9501,N_6433,N_6289);
xnor U9502 (N_9502,N_5035,N_5388);
nor U9503 (N_9503,N_6963,N_5555);
and U9504 (N_9504,N_6312,N_6520);
and U9505 (N_9505,N_7198,N_5142);
nor U9506 (N_9506,N_5292,N_5273);
xor U9507 (N_9507,N_7441,N_7208);
and U9508 (N_9508,N_6926,N_6017);
xor U9509 (N_9509,N_5014,N_5221);
and U9510 (N_9510,N_5964,N_5435);
and U9511 (N_9511,N_5745,N_6822);
nand U9512 (N_9512,N_5345,N_5576);
and U9513 (N_9513,N_5635,N_7336);
and U9514 (N_9514,N_7331,N_6205);
or U9515 (N_9515,N_6760,N_6961);
and U9516 (N_9516,N_5867,N_5099);
and U9517 (N_9517,N_7318,N_5667);
nand U9518 (N_9518,N_6907,N_7262);
xor U9519 (N_9519,N_6930,N_5664);
or U9520 (N_9520,N_6798,N_6320);
nor U9521 (N_9521,N_6822,N_6518);
nand U9522 (N_9522,N_6643,N_6621);
nor U9523 (N_9523,N_6348,N_7198);
nor U9524 (N_9524,N_6317,N_5183);
and U9525 (N_9525,N_7010,N_6222);
xor U9526 (N_9526,N_6158,N_5699);
xnor U9527 (N_9527,N_6619,N_6176);
nand U9528 (N_9528,N_6475,N_5526);
and U9529 (N_9529,N_7113,N_7116);
or U9530 (N_9530,N_6016,N_6561);
nand U9531 (N_9531,N_6008,N_7370);
and U9532 (N_9532,N_7475,N_5340);
and U9533 (N_9533,N_6779,N_5769);
xnor U9534 (N_9534,N_5637,N_6386);
and U9535 (N_9535,N_5938,N_6203);
nor U9536 (N_9536,N_5961,N_6235);
or U9537 (N_9537,N_6132,N_5435);
nor U9538 (N_9538,N_6269,N_5375);
and U9539 (N_9539,N_6721,N_5149);
and U9540 (N_9540,N_6393,N_7082);
nor U9541 (N_9541,N_5764,N_5850);
or U9542 (N_9542,N_6086,N_6407);
or U9543 (N_9543,N_5582,N_5293);
nor U9544 (N_9544,N_7445,N_7265);
xor U9545 (N_9545,N_6479,N_5911);
and U9546 (N_9546,N_5289,N_6956);
nand U9547 (N_9547,N_7160,N_6929);
or U9548 (N_9548,N_6952,N_6212);
xor U9549 (N_9549,N_7229,N_5711);
xnor U9550 (N_9550,N_6862,N_6006);
xnor U9551 (N_9551,N_5574,N_6659);
and U9552 (N_9552,N_5311,N_5134);
and U9553 (N_9553,N_7094,N_5739);
and U9554 (N_9554,N_6100,N_5349);
and U9555 (N_9555,N_5310,N_6249);
or U9556 (N_9556,N_7419,N_5163);
or U9557 (N_9557,N_5130,N_5098);
nor U9558 (N_9558,N_5141,N_7480);
xor U9559 (N_9559,N_5725,N_5490);
and U9560 (N_9560,N_6061,N_6071);
nand U9561 (N_9561,N_6332,N_7246);
and U9562 (N_9562,N_6654,N_6628);
or U9563 (N_9563,N_6505,N_7497);
or U9564 (N_9564,N_5955,N_7134);
xnor U9565 (N_9565,N_6200,N_6315);
nor U9566 (N_9566,N_7001,N_5165);
xnor U9567 (N_9567,N_5161,N_6562);
nand U9568 (N_9568,N_6372,N_6231);
or U9569 (N_9569,N_5517,N_5073);
nand U9570 (N_9570,N_6851,N_6427);
xor U9571 (N_9571,N_5352,N_6269);
or U9572 (N_9572,N_6093,N_7022);
nor U9573 (N_9573,N_5953,N_6993);
xnor U9574 (N_9574,N_5214,N_6672);
nor U9575 (N_9575,N_6542,N_5659);
or U9576 (N_9576,N_7206,N_6823);
nor U9577 (N_9577,N_5782,N_7379);
or U9578 (N_9578,N_7449,N_7450);
nor U9579 (N_9579,N_5660,N_5560);
and U9580 (N_9580,N_5306,N_5075);
nor U9581 (N_9581,N_5621,N_7400);
or U9582 (N_9582,N_5284,N_5175);
and U9583 (N_9583,N_5049,N_7468);
nor U9584 (N_9584,N_5613,N_5210);
xnor U9585 (N_9585,N_5950,N_6297);
nor U9586 (N_9586,N_5025,N_5536);
and U9587 (N_9587,N_6283,N_5071);
nand U9588 (N_9588,N_6876,N_6076);
and U9589 (N_9589,N_5114,N_5798);
xor U9590 (N_9590,N_6283,N_5400);
and U9591 (N_9591,N_7112,N_7004);
nor U9592 (N_9592,N_6537,N_6766);
and U9593 (N_9593,N_5217,N_6985);
or U9594 (N_9594,N_6155,N_6307);
nand U9595 (N_9595,N_7278,N_6340);
nor U9596 (N_9596,N_5470,N_6770);
and U9597 (N_9597,N_5756,N_5012);
nor U9598 (N_9598,N_5463,N_5476);
or U9599 (N_9599,N_6061,N_6765);
and U9600 (N_9600,N_6622,N_5261);
and U9601 (N_9601,N_5299,N_7258);
nor U9602 (N_9602,N_7076,N_6507);
nand U9603 (N_9603,N_5286,N_5369);
nor U9604 (N_9604,N_6271,N_6729);
or U9605 (N_9605,N_5380,N_5871);
and U9606 (N_9606,N_7047,N_5286);
nand U9607 (N_9607,N_7100,N_6458);
nor U9608 (N_9608,N_5171,N_5956);
xor U9609 (N_9609,N_5643,N_5420);
and U9610 (N_9610,N_6021,N_5799);
xor U9611 (N_9611,N_7020,N_6576);
nand U9612 (N_9612,N_6832,N_7328);
nor U9613 (N_9613,N_5003,N_6783);
or U9614 (N_9614,N_7225,N_5546);
xor U9615 (N_9615,N_5836,N_6477);
nand U9616 (N_9616,N_6716,N_6115);
and U9617 (N_9617,N_6623,N_6257);
nand U9618 (N_9618,N_6637,N_6484);
or U9619 (N_9619,N_6346,N_6149);
nor U9620 (N_9620,N_5529,N_6268);
or U9621 (N_9621,N_5996,N_7353);
nand U9622 (N_9622,N_7360,N_5157);
and U9623 (N_9623,N_6691,N_6873);
nor U9624 (N_9624,N_5295,N_5970);
nor U9625 (N_9625,N_7478,N_7243);
and U9626 (N_9626,N_6812,N_6749);
and U9627 (N_9627,N_5651,N_5849);
and U9628 (N_9628,N_7247,N_5048);
xnor U9629 (N_9629,N_5322,N_5866);
and U9630 (N_9630,N_5995,N_6668);
nand U9631 (N_9631,N_5068,N_7020);
nor U9632 (N_9632,N_5242,N_7099);
nand U9633 (N_9633,N_7144,N_6659);
or U9634 (N_9634,N_6843,N_6261);
nor U9635 (N_9635,N_6264,N_5044);
nor U9636 (N_9636,N_7054,N_5158);
nand U9637 (N_9637,N_6203,N_6426);
xnor U9638 (N_9638,N_6952,N_5170);
xnor U9639 (N_9639,N_6216,N_6416);
nor U9640 (N_9640,N_5498,N_7430);
nand U9641 (N_9641,N_5604,N_5485);
nor U9642 (N_9642,N_5962,N_7189);
nor U9643 (N_9643,N_6887,N_5786);
nand U9644 (N_9644,N_6142,N_7052);
and U9645 (N_9645,N_7001,N_5323);
xnor U9646 (N_9646,N_6054,N_5851);
or U9647 (N_9647,N_7024,N_6098);
nand U9648 (N_9648,N_6953,N_5087);
and U9649 (N_9649,N_7199,N_7191);
or U9650 (N_9650,N_7260,N_5250);
and U9651 (N_9651,N_6903,N_5931);
and U9652 (N_9652,N_5295,N_5706);
xnor U9653 (N_9653,N_6965,N_7436);
nand U9654 (N_9654,N_6788,N_6144);
nand U9655 (N_9655,N_6377,N_6703);
and U9656 (N_9656,N_5542,N_6759);
or U9657 (N_9657,N_5122,N_6458);
nand U9658 (N_9658,N_5509,N_6898);
and U9659 (N_9659,N_5363,N_6509);
or U9660 (N_9660,N_5487,N_7486);
nor U9661 (N_9661,N_5647,N_7017);
nand U9662 (N_9662,N_5350,N_5130);
nor U9663 (N_9663,N_6748,N_5106);
nor U9664 (N_9664,N_5009,N_5896);
or U9665 (N_9665,N_5263,N_5128);
and U9666 (N_9666,N_5541,N_6500);
and U9667 (N_9667,N_5625,N_6811);
or U9668 (N_9668,N_5741,N_5456);
or U9669 (N_9669,N_5304,N_5292);
nand U9670 (N_9670,N_5084,N_5961);
nor U9671 (N_9671,N_5157,N_6868);
nor U9672 (N_9672,N_6760,N_6828);
and U9673 (N_9673,N_7453,N_5029);
nor U9674 (N_9674,N_6017,N_6252);
nand U9675 (N_9675,N_6583,N_5057);
nand U9676 (N_9676,N_7038,N_7027);
or U9677 (N_9677,N_5043,N_7220);
and U9678 (N_9678,N_6745,N_6742);
and U9679 (N_9679,N_7301,N_6311);
xor U9680 (N_9680,N_6036,N_5034);
nand U9681 (N_9681,N_5865,N_6475);
nand U9682 (N_9682,N_5705,N_6896);
and U9683 (N_9683,N_5894,N_5229);
or U9684 (N_9684,N_5774,N_5872);
or U9685 (N_9685,N_5844,N_6744);
xor U9686 (N_9686,N_6069,N_7284);
or U9687 (N_9687,N_7100,N_6891);
nor U9688 (N_9688,N_6508,N_5735);
nor U9689 (N_9689,N_6471,N_5605);
nand U9690 (N_9690,N_6921,N_5264);
nor U9691 (N_9691,N_5766,N_5082);
nand U9692 (N_9692,N_7005,N_6330);
and U9693 (N_9693,N_5256,N_7343);
and U9694 (N_9694,N_6371,N_7429);
or U9695 (N_9695,N_5157,N_7228);
xnor U9696 (N_9696,N_5554,N_5034);
nor U9697 (N_9697,N_6890,N_7352);
nor U9698 (N_9698,N_5279,N_5062);
nand U9699 (N_9699,N_6951,N_6867);
nand U9700 (N_9700,N_6665,N_5896);
and U9701 (N_9701,N_6936,N_7304);
or U9702 (N_9702,N_6150,N_5661);
and U9703 (N_9703,N_6754,N_7375);
and U9704 (N_9704,N_5148,N_5373);
or U9705 (N_9705,N_7103,N_6706);
nor U9706 (N_9706,N_6796,N_7364);
xnor U9707 (N_9707,N_7078,N_6233);
nand U9708 (N_9708,N_5157,N_6794);
and U9709 (N_9709,N_5986,N_6366);
xnor U9710 (N_9710,N_6143,N_5872);
or U9711 (N_9711,N_6682,N_6388);
nand U9712 (N_9712,N_5682,N_7496);
or U9713 (N_9713,N_6394,N_5522);
nor U9714 (N_9714,N_5156,N_7180);
and U9715 (N_9715,N_7021,N_6065);
xnor U9716 (N_9716,N_6316,N_5238);
nor U9717 (N_9717,N_6913,N_5767);
and U9718 (N_9718,N_5110,N_6211);
nand U9719 (N_9719,N_6031,N_5571);
and U9720 (N_9720,N_5903,N_6492);
or U9721 (N_9721,N_7428,N_5903);
and U9722 (N_9722,N_5357,N_5713);
nand U9723 (N_9723,N_6719,N_6460);
and U9724 (N_9724,N_7366,N_5041);
or U9725 (N_9725,N_6647,N_5808);
nand U9726 (N_9726,N_6260,N_5558);
nor U9727 (N_9727,N_6044,N_7470);
and U9728 (N_9728,N_5930,N_7306);
xor U9729 (N_9729,N_7193,N_7333);
or U9730 (N_9730,N_5727,N_6956);
nand U9731 (N_9731,N_5178,N_5537);
nor U9732 (N_9732,N_6402,N_5127);
nand U9733 (N_9733,N_7265,N_5920);
nor U9734 (N_9734,N_7463,N_6212);
and U9735 (N_9735,N_5295,N_5087);
or U9736 (N_9736,N_5152,N_7044);
and U9737 (N_9737,N_6277,N_6926);
nor U9738 (N_9738,N_5297,N_5885);
nor U9739 (N_9739,N_5803,N_6557);
nand U9740 (N_9740,N_6892,N_7328);
nand U9741 (N_9741,N_5567,N_5790);
nand U9742 (N_9742,N_6985,N_5112);
and U9743 (N_9743,N_6240,N_7224);
or U9744 (N_9744,N_6611,N_6734);
nand U9745 (N_9745,N_6295,N_5655);
or U9746 (N_9746,N_6550,N_6293);
nand U9747 (N_9747,N_5606,N_5553);
nor U9748 (N_9748,N_6889,N_6078);
and U9749 (N_9749,N_5234,N_7280);
nor U9750 (N_9750,N_6697,N_7106);
nor U9751 (N_9751,N_5905,N_7410);
or U9752 (N_9752,N_6790,N_5134);
or U9753 (N_9753,N_7340,N_6365);
xor U9754 (N_9754,N_6536,N_6791);
and U9755 (N_9755,N_7261,N_6395);
nor U9756 (N_9756,N_7062,N_6419);
or U9757 (N_9757,N_5127,N_6699);
nand U9758 (N_9758,N_6864,N_6378);
nor U9759 (N_9759,N_6214,N_5187);
nor U9760 (N_9760,N_6235,N_6365);
nand U9761 (N_9761,N_7335,N_7296);
nand U9762 (N_9762,N_6086,N_6068);
or U9763 (N_9763,N_6410,N_6674);
nor U9764 (N_9764,N_6774,N_7136);
nand U9765 (N_9765,N_6244,N_6485);
and U9766 (N_9766,N_6170,N_6419);
and U9767 (N_9767,N_7288,N_6939);
or U9768 (N_9768,N_7144,N_7474);
nand U9769 (N_9769,N_6048,N_5371);
nor U9770 (N_9770,N_5610,N_5779);
nor U9771 (N_9771,N_6392,N_6636);
nand U9772 (N_9772,N_5274,N_7429);
xnor U9773 (N_9773,N_5802,N_6589);
nand U9774 (N_9774,N_6984,N_6448);
and U9775 (N_9775,N_5225,N_6882);
or U9776 (N_9776,N_6006,N_6019);
nor U9777 (N_9777,N_5341,N_5466);
xnor U9778 (N_9778,N_6165,N_5291);
xnor U9779 (N_9779,N_7145,N_5852);
nor U9780 (N_9780,N_5296,N_6687);
nand U9781 (N_9781,N_6329,N_6589);
and U9782 (N_9782,N_6886,N_6404);
and U9783 (N_9783,N_6714,N_5828);
and U9784 (N_9784,N_5656,N_5653);
nor U9785 (N_9785,N_6809,N_6994);
nand U9786 (N_9786,N_6936,N_6906);
nand U9787 (N_9787,N_6297,N_6852);
nor U9788 (N_9788,N_5286,N_5868);
nor U9789 (N_9789,N_6923,N_7161);
or U9790 (N_9790,N_7413,N_5444);
or U9791 (N_9791,N_6115,N_7439);
xnor U9792 (N_9792,N_6897,N_6719);
nor U9793 (N_9793,N_6128,N_5723);
xor U9794 (N_9794,N_6301,N_6786);
nand U9795 (N_9795,N_5811,N_7161);
xnor U9796 (N_9796,N_6218,N_6837);
nand U9797 (N_9797,N_6161,N_7079);
and U9798 (N_9798,N_5680,N_7199);
nor U9799 (N_9799,N_7173,N_5976);
nor U9800 (N_9800,N_6383,N_5155);
xnor U9801 (N_9801,N_7426,N_6157);
or U9802 (N_9802,N_6168,N_5844);
and U9803 (N_9803,N_6184,N_6661);
and U9804 (N_9804,N_6478,N_7343);
and U9805 (N_9805,N_6333,N_6774);
or U9806 (N_9806,N_7031,N_5136);
and U9807 (N_9807,N_6960,N_6066);
and U9808 (N_9808,N_7300,N_5322);
and U9809 (N_9809,N_7044,N_7187);
nand U9810 (N_9810,N_6909,N_7439);
nor U9811 (N_9811,N_6365,N_6869);
nor U9812 (N_9812,N_7336,N_5594);
or U9813 (N_9813,N_7140,N_6847);
nor U9814 (N_9814,N_5842,N_5116);
or U9815 (N_9815,N_5591,N_5718);
nand U9816 (N_9816,N_6710,N_5685);
or U9817 (N_9817,N_5213,N_5137);
nand U9818 (N_9818,N_5625,N_6386);
nand U9819 (N_9819,N_6973,N_5583);
and U9820 (N_9820,N_5169,N_6846);
nor U9821 (N_9821,N_6321,N_5218);
xor U9822 (N_9822,N_6097,N_7472);
and U9823 (N_9823,N_5215,N_7376);
xor U9824 (N_9824,N_6069,N_7159);
nor U9825 (N_9825,N_6331,N_6464);
nor U9826 (N_9826,N_7279,N_5532);
nor U9827 (N_9827,N_6971,N_7070);
xnor U9828 (N_9828,N_5978,N_5558);
nor U9829 (N_9829,N_7307,N_7255);
or U9830 (N_9830,N_6331,N_5411);
or U9831 (N_9831,N_5300,N_6791);
and U9832 (N_9832,N_6448,N_7174);
nor U9833 (N_9833,N_6103,N_5545);
or U9834 (N_9834,N_6080,N_6913);
and U9835 (N_9835,N_6669,N_6041);
nand U9836 (N_9836,N_5165,N_5429);
or U9837 (N_9837,N_6592,N_7389);
nor U9838 (N_9838,N_7343,N_7179);
nor U9839 (N_9839,N_6659,N_6977);
and U9840 (N_9840,N_6615,N_5554);
and U9841 (N_9841,N_5300,N_5279);
or U9842 (N_9842,N_6155,N_6229);
nand U9843 (N_9843,N_5824,N_6434);
or U9844 (N_9844,N_5433,N_5600);
xnor U9845 (N_9845,N_5945,N_7471);
and U9846 (N_9846,N_6908,N_7291);
nor U9847 (N_9847,N_6072,N_6481);
nand U9848 (N_9848,N_6427,N_6266);
nand U9849 (N_9849,N_5690,N_6645);
or U9850 (N_9850,N_6967,N_6846);
nand U9851 (N_9851,N_6086,N_6603);
or U9852 (N_9852,N_5694,N_7108);
and U9853 (N_9853,N_6387,N_6306);
nand U9854 (N_9854,N_6208,N_5405);
nand U9855 (N_9855,N_5114,N_6998);
or U9856 (N_9856,N_7100,N_6579);
and U9857 (N_9857,N_7128,N_6257);
nand U9858 (N_9858,N_6270,N_6028);
and U9859 (N_9859,N_5125,N_7013);
nor U9860 (N_9860,N_6807,N_5228);
nand U9861 (N_9861,N_5354,N_6895);
nor U9862 (N_9862,N_5497,N_7050);
nor U9863 (N_9863,N_7072,N_5652);
xnor U9864 (N_9864,N_6629,N_7119);
and U9865 (N_9865,N_6406,N_7428);
nor U9866 (N_9866,N_6341,N_6603);
nand U9867 (N_9867,N_5195,N_5394);
or U9868 (N_9868,N_6432,N_6049);
and U9869 (N_9869,N_7011,N_6977);
nand U9870 (N_9870,N_5670,N_6558);
nand U9871 (N_9871,N_5142,N_5569);
nor U9872 (N_9872,N_5639,N_5822);
or U9873 (N_9873,N_6889,N_6433);
or U9874 (N_9874,N_7498,N_5595);
xnor U9875 (N_9875,N_6081,N_5492);
nand U9876 (N_9876,N_5236,N_6893);
nor U9877 (N_9877,N_7338,N_7270);
nand U9878 (N_9878,N_7480,N_7012);
or U9879 (N_9879,N_6598,N_6520);
nor U9880 (N_9880,N_6576,N_5415);
or U9881 (N_9881,N_6453,N_5289);
nor U9882 (N_9882,N_5362,N_5229);
nand U9883 (N_9883,N_5955,N_6155);
nand U9884 (N_9884,N_6953,N_5376);
or U9885 (N_9885,N_5268,N_6189);
xor U9886 (N_9886,N_7174,N_7218);
or U9887 (N_9887,N_5010,N_6142);
and U9888 (N_9888,N_7094,N_7277);
or U9889 (N_9889,N_5291,N_6837);
or U9890 (N_9890,N_7036,N_6463);
nor U9891 (N_9891,N_7383,N_6477);
nand U9892 (N_9892,N_5334,N_5998);
nand U9893 (N_9893,N_7377,N_7444);
nand U9894 (N_9894,N_6114,N_5678);
xnor U9895 (N_9895,N_5178,N_5325);
or U9896 (N_9896,N_7221,N_6771);
and U9897 (N_9897,N_6301,N_7232);
or U9898 (N_9898,N_7063,N_7247);
or U9899 (N_9899,N_7393,N_5937);
and U9900 (N_9900,N_6904,N_7473);
or U9901 (N_9901,N_5160,N_5804);
nor U9902 (N_9902,N_7203,N_5297);
or U9903 (N_9903,N_5898,N_5164);
or U9904 (N_9904,N_6048,N_5902);
xnor U9905 (N_9905,N_5432,N_5131);
nand U9906 (N_9906,N_7394,N_5924);
xnor U9907 (N_9907,N_6162,N_6441);
and U9908 (N_9908,N_6455,N_5522);
and U9909 (N_9909,N_7052,N_5635);
and U9910 (N_9910,N_5219,N_7282);
xnor U9911 (N_9911,N_6995,N_6631);
nand U9912 (N_9912,N_6236,N_5248);
xor U9913 (N_9913,N_6478,N_5517);
and U9914 (N_9914,N_7115,N_6001);
or U9915 (N_9915,N_6904,N_7115);
and U9916 (N_9916,N_6567,N_7076);
or U9917 (N_9917,N_6476,N_5286);
nand U9918 (N_9918,N_6083,N_5065);
nor U9919 (N_9919,N_6395,N_7404);
xor U9920 (N_9920,N_5020,N_5600);
or U9921 (N_9921,N_6719,N_7166);
or U9922 (N_9922,N_5445,N_5722);
and U9923 (N_9923,N_5266,N_5763);
nor U9924 (N_9924,N_5767,N_5540);
nor U9925 (N_9925,N_6649,N_6647);
xor U9926 (N_9926,N_6080,N_6022);
nor U9927 (N_9927,N_7447,N_5020);
xnor U9928 (N_9928,N_6202,N_6269);
and U9929 (N_9929,N_5835,N_7488);
or U9930 (N_9930,N_5012,N_7132);
nand U9931 (N_9931,N_6012,N_6245);
or U9932 (N_9932,N_6392,N_6672);
nand U9933 (N_9933,N_5884,N_6936);
and U9934 (N_9934,N_7363,N_7399);
nor U9935 (N_9935,N_5331,N_7069);
or U9936 (N_9936,N_6857,N_5760);
nand U9937 (N_9937,N_5142,N_6256);
nor U9938 (N_9938,N_7088,N_5673);
nand U9939 (N_9939,N_6427,N_7208);
or U9940 (N_9940,N_6077,N_5153);
nand U9941 (N_9941,N_5792,N_5999);
and U9942 (N_9942,N_5177,N_5202);
or U9943 (N_9943,N_6925,N_6607);
nor U9944 (N_9944,N_5285,N_7157);
nor U9945 (N_9945,N_6517,N_6616);
or U9946 (N_9946,N_5597,N_6595);
nand U9947 (N_9947,N_7002,N_6394);
xnor U9948 (N_9948,N_5167,N_7187);
and U9949 (N_9949,N_5581,N_7205);
xnor U9950 (N_9950,N_6518,N_7129);
and U9951 (N_9951,N_7394,N_5950);
and U9952 (N_9952,N_5989,N_7216);
nand U9953 (N_9953,N_6652,N_6486);
nand U9954 (N_9954,N_7459,N_5822);
nand U9955 (N_9955,N_5908,N_6418);
or U9956 (N_9956,N_6055,N_6100);
xnor U9957 (N_9957,N_7400,N_6809);
or U9958 (N_9958,N_7486,N_6319);
or U9959 (N_9959,N_7136,N_6288);
or U9960 (N_9960,N_6930,N_6532);
nor U9961 (N_9961,N_6895,N_7380);
and U9962 (N_9962,N_5960,N_5922);
nand U9963 (N_9963,N_7366,N_6914);
nor U9964 (N_9964,N_5787,N_7300);
nor U9965 (N_9965,N_6092,N_7229);
or U9966 (N_9966,N_7312,N_5846);
nor U9967 (N_9967,N_6849,N_5286);
nor U9968 (N_9968,N_5657,N_6613);
nor U9969 (N_9969,N_5547,N_5191);
nand U9970 (N_9970,N_6903,N_6971);
nor U9971 (N_9971,N_7430,N_5379);
nor U9972 (N_9972,N_7130,N_6011);
nor U9973 (N_9973,N_7354,N_5475);
xor U9974 (N_9974,N_6443,N_5921);
and U9975 (N_9975,N_5599,N_6075);
nand U9976 (N_9976,N_6188,N_6360);
and U9977 (N_9977,N_7042,N_6088);
or U9978 (N_9978,N_5523,N_5712);
nor U9979 (N_9979,N_6460,N_5202);
and U9980 (N_9980,N_5137,N_5374);
nand U9981 (N_9981,N_6719,N_6082);
xor U9982 (N_9982,N_6718,N_6304);
nand U9983 (N_9983,N_7304,N_6094);
nand U9984 (N_9984,N_5841,N_5023);
nor U9985 (N_9985,N_5172,N_6763);
or U9986 (N_9986,N_7097,N_7321);
and U9987 (N_9987,N_6522,N_6122);
nand U9988 (N_9988,N_7116,N_6962);
nor U9989 (N_9989,N_6901,N_6972);
nand U9990 (N_9990,N_7254,N_7005);
nor U9991 (N_9991,N_5617,N_7440);
nor U9992 (N_9992,N_6271,N_7413);
nor U9993 (N_9993,N_7454,N_6843);
or U9994 (N_9994,N_6091,N_6192);
or U9995 (N_9995,N_5904,N_6561);
xnor U9996 (N_9996,N_6428,N_6549);
and U9997 (N_9997,N_6834,N_5252);
and U9998 (N_9998,N_6647,N_6493);
or U9999 (N_9999,N_6073,N_6193);
and UO_0 (O_0,N_8788,N_9633);
nor UO_1 (O_1,N_8109,N_9221);
nor UO_2 (O_2,N_8884,N_9629);
or UO_3 (O_3,N_8458,N_9570);
nand UO_4 (O_4,N_7856,N_9678);
or UO_5 (O_5,N_7896,N_8329);
or UO_6 (O_6,N_8463,N_9946);
nor UO_7 (O_7,N_8644,N_9029);
or UO_8 (O_8,N_8722,N_9701);
xor UO_9 (O_9,N_8478,N_8831);
or UO_10 (O_10,N_8557,N_7905);
nor UO_11 (O_11,N_8743,N_8712);
nor UO_12 (O_12,N_9515,N_7547);
and UO_13 (O_13,N_9735,N_9256);
nand UO_14 (O_14,N_8508,N_8550);
nand UO_15 (O_15,N_9422,N_8257);
nand UO_16 (O_16,N_7992,N_8032);
or UO_17 (O_17,N_9310,N_7651);
nand UO_18 (O_18,N_9144,N_8039);
nor UO_19 (O_19,N_9942,N_7505);
nand UO_20 (O_20,N_9922,N_8830);
and UO_21 (O_21,N_9242,N_9383);
or UO_22 (O_22,N_8866,N_8872);
and UO_23 (O_23,N_9008,N_8229);
and UO_24 (O_24,N_8612,N_9333);
and UO_25 (O_25,N_7944,N_7987);
or UO_26 (O_26,N_9547,N_7846);
and UO_27 (O_27,N_9913,N_9795);
nor UO_28 (O_28,N_8649,N_8771);
nor UO_29 (O_29,N_7707,N_7590);
xnor UO_30 (O_30,N_9666,N_9831);
and UO_31 (O_31,N_8756,N_9694);
nor UO_32 (O_32,N_8286,N_9757);
and UO_33 (O_33,N_8947,N_8427);
nor UO_34 (O_34,N_9075,N_8887);
nor UO_35 (O_35,N_9183,N_9905);
nand UO_36 (O_36,N_7709,N_9484);
nand UO_37 (O_37,N_9382,N_8922);
and UO_38 (O_38,N_8952,N_8152);
or UO_39 (O_39,N_9035,N_8966);
and UO_40 (O_40,N_7870,N_9263);
nand UO_41 (O_41,N_8358,N_8620);
nand UO_42 (O_42,N_9005,N_7776);
nand UO_43 (O_43,N_8927,N_7514);
and UO_44 (O_44,N_8816,N_9281);
and UO_45 (O_45,N_8851,N_8894);
or UO_46 (O_46,N_9385,N_8399);
or UO_47 (O_47,N_9684,N_8706);
and UO_48 (O_48,N_7558,N_8531);
or UO_49 (O_49,N_9402,N_8052);
nor UO_50 (O_50,N_7711,N_8323);
xor UO_51 (O_51,N_9821,N_8536);
or UO_52 (O_52,N_9488,N_9377);
nand UO_53 (O_53,N_9345,N_9343);
or UO_54 (O_54,N_9954,N_8078);
and UO_55 (O_55,N_8034,N_9725);
and UO_56 (O_56,N_9365,N_8086);
and UO_57 (O_57,N_9911,N_8356);
or UO_58 (O_58,N_9313,N_8361);
and UO_59 (O_59,N_7762,N_7704);
or UO_60 (O_60,N_8325,N_8689);
nand UO_61 (O_61,N_9110,N_9948);
xnor UO_62 (O_62,N_7812,N_7605);
and UO_63 (O_63,N_9537,N_9391);
and UO_64 (O_64,N_8912,N_8605);
nand UO_65 (O_65,N_7942,N_8727);
xor UO_66 (O_66,N_9732,N_7678);
xor UO_67 (O_67,N_9424,N_8247);
and UO_68 (O_68,N_9850,N_7562);
nor UO_69 (O_69,N_8559,N_7694);
nand UO_70 (O_70,N_8203,N_8138);
nand UO_71 (O_71,N_7512,N_9827);
xnor UO_72 (O_72,N_9909,N_7719);
xnor UO_73 (O_73,N_8583,N_8123);
and UO_74 (O_74,N_8470,N_9775);
xor UO_75 (O_75,N_8455,N_9455);
xnor UO_76 (O_76,N_8719,N_8501);
nand UO_77 (O_77,N_9705,N_9425);
nor UO_78 (O_78,N_9977,N_8310);
or UO_79 (O_79,N_9497,N_7802);
xnor UO_80 (O_80,N_9606,N_9135);
nand UO_81 (O_81,N_9438,N_7873);
xor UO_82 (O_82,N_9072,N_9454);
xor UO_83 (O_83,N_9236,N_7831);
or UO_84 (O_84,N_8210,N_7765);
xnor UO_85 (O_85,N_9293,N_7527);
or UO_86 (O_86,N_9607,N_9415);
and UO_87 (O_87,N_8466,N_8429);
and UO_88 (O_88,N_9786,N_9591);
xnor UO_89 (O_89,N_9906,N_7923);
and UO_90 (O_90,N_8379,N_8079);
nor UO_91 (O_91,N_9625,N_8219);
and UO_92 (O_92,N_7926,N_8277);
nand UO_93 (O_93,N_9037,N_7933);
and UO_94 (O_94,N_8849,N_9134);
nand UO_95 (O_95,N_7890,N_9397);
nand UO_96 (O_96,N_9091,N_7985);
or UO_97 (O_97,N_9957,N_9372);
nor UO_98 (O_98,N_9217,N_9380);
nand UO_99 (O_99,N_7978,N_9118);
and UO_100 (O_100,N_8163,N_8858);
and UO_101 (O_101,N_8755,N_8986);
nor UO_102 (O_102,N_8741,N_9900);
and UO_103 (O_103,N_8116,N_8994);
nor UO_104 (O_104,N_7895,N_8024);
nor UO_105 (O_105,N_9604,N_7677);
nor UO_106 (O_106,N_8418,N_7876);
nor UO_107 (O_107,N_8198,N_9342);
xnor UO_108 (O_108,N_7687,N_7949);
nor UO_109 (O_109,N_8593,N_8139);
nand UO_110 (O_110,N_9514,N_7929);
nand UO_111 (O_111,N_8616,N_9318);
and UO_112 (O_112,N_7872,N_9620);
or UO_113 (O_113,N_8029,N_8119);
nand UO_114 (O_114,N_9930,N_8217);
nor UO_115 (O_115,N_9754,N_9704);
nor UO_116 (O_116,N_7570,N_7750);
or UO_117 (O_117,N_7782,N_8594);
xnor UO_118 (O_118,N_7549,N_9811);
and UO_119 (O_119,N_8129,N_9619);
or UO_120 (O_120,N_9239,N_8068);
nor UO_121 (O_121,N_7954,N_8386);
nor UO_122 (O_122,N_8443,N_9332);
nand UO_123 (O_123,N_9583,N_8506);
nand UO_124 (O_124,N_9806,N_9561);
nand UO_125 (O_125,N_8193,N_9100);
nor UO_126 (O_126,N_7675,N_7518);
xor UO_127 (O_127,N_9522,N_8005);
nand UO_128 (O_128,N_8081,N_9452);
and UO_129 (O_129,N_7986,N_7946);
nand UO_130 (O_130,N_8855,N_8744);
or UO_131 (O_131,N_9554,N_9159);
nand UO_132 (O_132,N_7758,N_8118);
nor UO_133 (O_133,N_9011,N_8638);
xnor UO_134 (O_134,N_8456,N_8579);
or UO_135 (O_135,N_9578,N_9737);
nand UO_136 (O_136,N_8045,N_9612);
nor UO_137 (O_137,N_9112,N_9637);
xnor UO_138 (O_138,N_9172,N_7533);
nor UO_139 (O_139,N_9020,N_8882);
nand UO_140 (O_140,N_9138,N_8273);
xor UO_141 (O_141,N_9745,N_9241);
or UO_142 (O_142,N_8664,N_8950);
and UO_143 (O_143,N_8209,N_7959);
nor UO_144 (O_144,N_9535,N_8975);
or UO_145 (O_145,N_9171,N_8225);
xor UO_146 (O_146,N_8342,N_8993);
xnor UO_147 (O_147,N_9892,N_8497);
or UO_148 (O_148,N_8328,N_9416);
nand UO_149 (O_149,N_9658,N_8474);
nor UO_150 (O_150,N_9350,N_9190);
and UO_151 (O_151,N_9067,N_9609);
and UO_152 (O_152,N_8535,N_9104);
nor UO_153 (O_153,N_9918,N_9300);
xnor UO_154 (O_154,N_8683,N_8651);
nor UO_155 (O_155,N_9045,N_8933);
or UO_156 (O_156,N_7703,N_8959);
nand UO_157 (O_157,N_8835,N_7768);
and UO_158 (O_158,N_8697,N_8023);
nor UO_159 (O_159,N_8235,N_8935);
nand UO_160 (O_160,N_9436,N_9574);
or UO_161 (O_161,N_8956,N_8428);
and UO_162 (O_162,N_9750,N_8588);
and UO_163 (O_163,N_9177,N_9682);
or UO_164 (O_164,N_8069,N_8174);
nand UO_165 (O_165,N_9558,N_8955);
nand UO_166 (O_166,N_8367,N_7577);
nand UO_167 (O_167,N_8269,N_8949);
xor UO_168 (O_168,N_7948,N_9053);
and UO_169 (O_169,N_9854,N_7685);
nor UO_170 (O_170,N_9407,N_9487);
or UO_171 (O_171,N_9687,N_7725);
and UO_172 (O_172,N_8663,N_9568);
and UO_173 (O_173,N_9841,N_9081);
nor UO_174 (O_174,N_7508,N_9133);
nor UO_175 (O_175,N_8666,N_9700);
nand UO_176 (O_176,N_8703,N_9411);
nand UO_177 (O_177,N_9501,N_7778);
xnor UO_178 (O_178,N_9245,N_8025);
and UO_179 (O_179,N_9778,N_8505);
and UO_180 (O_180,N_9917,N_9148);
nand UO_181 (O_181,N_8084,N_9240);
nand UO_182 (O_182,N_8658,N_8014);
or UO_183 (O_183,N_9214,N_8360);
nand UO_184 (O_184,N_9655,N_9399);
and UO_185 (O_185,N_8004,N_9567);
or UO_186 (O_186,N_8717,N_9675);
xor UO_187 (O_187,N_9193,N_9941);
nand UO_188 (O_188,N_8691,N_7983);
and UO_189 (O_189,N_9587,N_7920);
nand UO_190 (O_190,N_7860,N_7803);
nand UO_191 (O_191,N_8914,N_8962);
nand UO_192 (O_192,N_8404,N_9871);
and UO_193 (O_193,N_9767,N_9379);
nand UO_194 (O_194,N_9640,N_8553);
or UO_195 (O_195,N_8001,N_9042);
nand UO_196 (O_196,N_7600,N_8905);
nor UO_197 (O_197,N_7511,N_8224);
xnor UO_198 (O_198,N_9553,N_9228);
nand UO_199 (O_199,N_8077,N_9987);
and UO_200 (O_200,N_7767,N_9769);
nand UO_201 (O_201,N_9610,N_7847);
and UO_202 (O_202,N_7915,N_7658);
xnor UO_203 (O_203,N_7951,N_9462);
nand UO_204 (O_204,N_8041,N_8312);
or UO_205 (O_205,N_8292,N_9481);
nand UO_206 (O_206,N_8287,N_8022);
nor UO_207 (O_207,N_7808,N_8801);
nand UO_208 (O_208,N_9471,N_7692);
nand UO_209 (O_209,N_9276,N_9914);
nor UO_210 (O_210,N_9070,N_9614);
nor UO_211 (O_211,N_8473,N_8746);
nor UO_212 (O_212,N_9791,N_9124);
nand UO_213 (O_213,N_9373,N_8963);
or UO_214 (O_214,N_9920,N_8218);
nor UO_215 (O_215,N_8708,N_8874);
or UO_216 (O_216,N_8660,N_8177);
and UO_217 (O_217,N_8643,N_8941);
and UO_218 (O_218,N_7774,N_8645);
or UO_219 (O_219,N_7764,N_9782);
nand UO_220 (O_220,N_9187,N_7780);
or UO_221 (O_221,N_9468,N_8441);
or UO_222 (O_222,N_9621,N_9294);
or UO_223 (O_223,N_8685,N_7727);
nand UO_224 (O_224,N_8406,N_9055);
nand UO_225 (O_225,N_8781,N_8684);
and UO_226 (O_226,N_7720,N_8421);
nor UO_227 (O_227,N_8817,N_8538);
or UO_228 (O_228,N_7543,N_9290);
and UO_229 (O_229,N_8566,N_8058);
nor UO_230 (O_230,N_8483,N_9404);
xnor UO_231 (O_231,N_8270,N_9309);
or UO_232 (O_232,N_8031,N_9996);
nand UO_233 (O_233,N_7937,N_8982);
nand UO_234 (O_234,N_7927,N_9036);
xor UO_235 (O_235,N_8969,N_8699);
and UO_236 (O_236,N_8648,N_9079);
xor UO_237 (O_237,N_9085,N_8143);
and UO_238 (O_238,N_9809,N_9460);
or UO_239 (O_239,N_7688,N_7749);
nand UO_240 (O_240,N_8751,N_8716);
and UO_241 (O_241,N_8281,N_7855);
or UO_242 (O_242,N_7947,N_7880);
xnor UO_243 (O_243,N_8033,N_7906);
or UO_244 (O_244,N_7519,N_8339);
or UO_245 (O_245,N_7918,N_9302);
nand UO_246 (O_246,N_7664,N_9155);
nor UO_247 (O_247,N_7894,N_7628);
xnor UO_248 (O_248,N_8056,N_8814);
or UO_249 (O_249,N_8980,N_8591);
and UO_250 (O_250,N_9600,N_9647);
or UO_251 (O_251,N_9789,N_8798);
xnor UO_252 (O_252,N_7838,N_9393);
or UO_253 (O_253,N_9213,N_9504);
and UO_254 (O_254,N_7775,N_9836);
or UO_255 (O_255,N_9232,N_8586);
or UO_256 (O_256,N_8534,N_8839);
nor UO_257 (O_257,N_7783,N_8070);
or UO_258 (O_258,N_9226,N_7886);
and UO_259 (O_259,N_8237,N_7702);
or UO_260 (O_260,N_7631,N_8322);
nor UO_261 (O_261,N_9021,N_8194);
xnor UO_262 (O_262,N_9971,N_9864);
nand UO_263 (O_263,N_8826,N_7500);
and UO_264 (O_264,N_7633,N_8330);
and UO_265 (O_265,N_7943,N_8173);
nand UO_266 (O_266,N_9165,N_8636);
or UO_267 (O_267,N_8797,N_9780);
xor UO_268 (O_268,N_9325,N_7958);
xnor UO_269 (O_269,N_8942,N_8695);
and UO_270 (O_270,N_9087,N_9819);
and UO_271 (O_271,N_9288,N_9137);
and UO_272 (O_272,N_9009,N_8002);
and UO_273 (O_273,N_9319,N_9368);
or UO_274 (O_274,N_9622,N_7585);
and UO_275 (O_275,N_7612,N_9002);
nor UO_276 (O_276,N_8772,N_9758);
nand UO_277 (O_277,N_7607,N_8364);
nand UO_278 (O_278,N_8373,N_9483);
and UO_279 (O_279,N_9802,N_8195);
nand UO_280 (O_280,N_9576,N_8484);
or UO_281 (O_281,N_8157,N_9868);
nand UO_282 (O_282,N_8422,N_9538);
nor UO_283 (O_283,N_8010,N_9949);
or UO_284 (O_284,N_9152,N_9933);
and UO_285 (O_285,N_8048,N_8168);
nand UO_286 (O_286,N_9145,N_9163);
xor UO_287 (O_287,N_8037,N_8562);
nand UO_288 (O_288,N_8375,N_8315);
nand UO_289 (O_289,N_9039,N_9825);
nor UO_290 (O_290,N_7548,N_8140);
or UO_291 (O_291,N_9878,N_9505);
and UO_292 (O_292,N_9673,N_7935);
xnor UO_293 (O_293,N_7857,N_9995);
nor UO_294 (O_294,N_9928,N_9715);
or UO_295 (O_295,N_8674,N_7551);
nor UO_296 (O_296,N_9550,N_9244);
and UO_297 (O_297,N_7801,N_9916);
or UO_298 (O_298,N_8657,N_7790);
and UO_299 (O_299,N_9446,N_8232);
nand UO_300 (O_300,N_9650,N_7795);
or UO_301 (O_301,N_9798,N_8197);
and UO_302 (O_302,N_9511,N_8979);
and UO_303 (O_303,N_7579,N_9109);
and UO_304 (O_304,N_7741,N_9477);
nor UO_305 (O_305,N_8598,N_7829);
nor UO_306 (O_306,N_8750,N_8042);
or UO_307 (O_307,N_9233,N_8633);
xor UO_308 (O_308,N_8667,N_9936);
nor UO_309 (O_309,N_7523,N_9392);
and UO_310 (O_310,N_7861,N_9270);
or UO_311 (O_311,N_7635,N_9595);
nor UO_312 (O_312,N_9787,N_8714);
and UO_313 (O_313,N_9141,N_8321);
or UO_314 (O_314,N_9102,N_7834);
and UO_315 (O_315,N_9727,N_8394);
or UO_316 (O_316,N_9461,N_9980);
and UO_317 (O_317,N_9351,N_9699);
or UO_318 (O_318,N_8696,N_8600);
nor UO_319 (O_319,N_9613,N_9156);
xor UO_320 (O_320,N_9433,N_7836);
xnor UO_321 (O_321,N_8264,N_9589);
or UO_322 (O_322,N_8692,N_9566);
or UO_323 (O_323,N_8450,N_9453);
and UO_324 (O_324,N_9781,N_8347);
nand UO_325 (O_325,N_8383,N_9139);
nor UO_326 (O_326,N_9096,N_8641);
nor UO_327 (O_327,N_7591,N_9349);
xor UO_328 (O_328,N_7571,N_7921);
nand UO_329 (O_329,N_8477,N_8752);
or UO_330 (O_330,N_8834,N_7645);
xnor UO_331 (O_331,N_8494,N_8868);
or UO_332 (O_332,N_9608,N_8211);
nor UO_333 (O_333,N_9533,N_9001);
xor UO_334 (O_334,N_8540,N_7567);
xor UO_335 (O_335,N_8888,N_8778);
or UO_336 (O_336,N_7849,N_8552);
and UO_337 (O_337,N_8460,N_9508);
or UO_338 (O_338,N_8745,N_9975);
xor UO_339 (O_339,N_9863,N_8655);
or UO_340 (O_340,N_8688,N_9099);
or UO_341 (O_341,N_8036,N_7841);
nand UO_342 (O_342,N_8791,N_8804);
nor UO_343 (O_343,N_8300,N_7648);
nand UO_344 (O_344,N_9466,N_7736);
and UO_345 (O_345,N_8578,N_8350);
nor UO_346 (O_346,N_9966,N_7657);
nor UO_347 (O_347,N_7968,N_9330);
nor UO_348 (O_348,N_8498,N_8385);
and UO_349 (O_349,N_9237,N_7824);
or UO_350 (O_350,N_8027,N_9847);
or UO_351 (O_351,N_9255,N_8230);
xnor UO_352 (O_352,N_8160,N_7934);
and UO_353 (O_353,N_9797,N_9115);
and UO_354 (O_354,N_8523,N_7854);
or UO_355 (O_355,N_8028,N_7820);
or UO_356 (O_356,N_8976,N_8548);
nand UO_357 (O_357,N_7842,N_9931);
or UO_358 (O_358,N_8654,N_9119);
or UO_359 (O_359,N_9321,N_9421);
xor UO_360 (O_360,N_8913,N_8928);
or UO_361 (O_361,N_9014,N_9268);
or UO_362 (O_362,N_8125,N_8192);
and UO_363 (O_363,N_7524,N_8970);
nand UO_364 (O_364,N_8946,N_8522);
xnor UO_365 (O_365,N_9518,N_9185);
nand UO_366 (O_366,N_7544,N_8739);
or UO_367 (O_367,N_9026,N_8191);
nor UO_368 (O_368,N_7536,N_7907);
nor UO_369 (O_369,N_7738,N_8981);
nand UO_370 (O_370,N_9495,N_7592);
nand UO_371 (O_371,N_8596,N_8800);
and UO_372 (O_372,N_9273,N_8398);
nand UO_373 (O_373,N_8391,N_8865);
and UO_374 (O_374,N_7785,N_7932);
nand UO_375 (O_375,N_9485,N_9128);
and UO_376 (O_376,N_9248,N_9285);
or UO_377 (O_377,N_9788,N_9486);
and UO_378 (O_378,N_9677,N_9662);
nor UO_379 (O_379,N_7910,N_7990);
or UO_380 (O_380,N_9006,N_9891);
nand UO_381 (O_381,N_8121,N_7811);
and UO_382 (O_382,N_9969,N_9759);
nor UO_383 (O_383,N_8646,N_9867);
or UO_384 (O_384,N_8833,N_8721);
and UO_385 (O_385,N_8464,N_9523);
or UO_386 (O_386,N_8561,N_9817);
or UO_387 (O_387,N_8189,N_9603);
xnor UO_388 (O_388,N_8449,N_7654);
nor UO_389 (O_389,N_7596,N_8690);
or UO_390 (O_390,N_8249,N_8491);
or UO_391 (O_391,N_8120,N_9683);
or UO_392 (O_392,N_8783,N_9052);
or UO_393 (O_393,N_8362,N_8926);
nor UO_394 (O_394,N_7914,N_7723);
and UO_395 (O_395,N_8803,N_9275);
xor UO_396 (O_396,N_9186,N_9189);
or UO_397 (O_397,N_8246,N_7724);
nor UO_398 (O_398,N_9489,N_9929);
or UO_399 (O_399,N_7588,N_7881);
and UO_400 (O_400,N_8742,N_9066);
and UO_401 (O_401,N_9509,N_7871);
or UO_402 (O_402,N_7630,N_8931);
and UO_403 (O_403,N_9443,N_8278);
and UO_404 (O_404,N_9154,N_7650);
or UO_405 (O_405,N_9266,N_9470);
nand UO_406 (O_406,N_9912,N_8920);
nand UO_407 (O_407,N_9113,N_9828);
nor UO_408 (O_408,N_9061,N_9569);
xor UO_409 (O_409,N_8440,N_8779);
nor UO_410 (O_410,N_8091,N_7893);
and UO_411 (O_411,N_8298,N_7832);
and UO_412 (O_412,N_9264,N_7627);
or UO_413 (O_413,N_9116,N_7690);
or UO_414 (O_414,N_9989,N_9136);
nand UO_415 (O_415,N_8202,N_8971);
or UO_416 (O_416,N_9652,N_8439);
and UO_417 (O_417,N_7815,N_8013);
nand UO_418 (O_418,N_9586,N_9303);
or UO_419 (O_419,N_9327,N_8038);
or UO_420 (O_420,N_7599,N_9857);
and UO_421 (O_421,N_7902,N_9341);
and UO_422 (O_422,N_9370,N_7644);
and UO_423 (O_423,N_7898,N_9361);
or UO_424 (O_424,N_9741,N_8568);
and UO_425 (O_425,N_7634,N_9639);
nor UO_426 (O_426,N_9950,N_9979);
nor UO_427 (O_427,N_9360,N_9175);
or UO_428 (O_428,N_9108,N_9755);
or UO_429 (O_429,N_8702,N_7560);
or UO_430 (O_430,N_8546,N_7626);
nand UO_431 (O_431,N_8585,N_9651);
nor UO_432 (O_432,N_7826,N_9356);
nand UO_433 (O_433,N_7740,N_8402);
or UO_434 (O_434,N_9888,N_9896);
or UO_435 (O_435,N_7900,N_7960);
or UO_436 (O_436,N_9178,N_8977);
or UO_437 (O_437,N_8802,N_9284);
nor UO_438 (O_438,N_8539,N_9763);
and UO_439 (O_439,N_9976,N_7797);
and UO_440 (O_440,N_9921,N_8901);
nand UO_441 (O_441,N_9494,N_9668);
nor UO_442 (O_442,N_7862,N_9335);
and UO_443 (O_443,N_8629,N_7742);
and UO_444 (O_444,N_9708,N_8919);
and UO_445 (O_445,N_7839,N_8650);
or UO_446 (O_446,N_8984,N_8765);
and UO_447 (O_447,N_9959,N_8500);
nand UO_448 (O_448,N_8479,N_9858);
nand UO_449 (O_449,N_9320,N_8661);
or UO_450 (O_450,N_8789,N_8419);
nor UO_451 (O_451,N_9364,N_8652);
nor UO_452 (O_452,N_9179,N_9230);
and UO_453 (O_453,N_7521,N_8496);
nand UO_454 (O_454,N_9747,N_8293);
nor UO_455 (O_455,N_9180,N_8737);
nor UO_456 (O_456,N_9150,N_9901);
nor UO_457 (O_457,N_9674,N_7745);
nor UO_458 (O_458,N_9845,N_8572);
and UO_459 (O_459,N_9555,N_8843);
or UO_460 (O_460,N_7903,N_9785);
nand UO_461 (O_461,N_9602,N_8212);
or UO_462 (O_462,N_8414,N_9030);
and UO_463 (O_463,N_7979,N_8821);
nor UO_464 (O_464,N_9157,N_8824);
nor UO_465 (O_465,N_7615,N_9225);
nand UO_466 (O_466,N_8340,N_9103);
nand UO_467 (O_467,N_8723,N_7813);
nor UO_468 (O_468,N_9751,N_7755);
nand UO_469 (O_469,N_8255,N_9915);
nand UO_470 (O_470,N_7563,N_9659);
nand UO_471 (O_471,N_9935,N_9296);
nand UO_472 (O_472,N_9592,N_9322);
and UO_473 (O_473,N_8451,N_7682);
nor UO_474 (O_474,N_8873,N_9564);
and UO_475 (O_475,N_9084,N_9050);
nand UO_476 (O_476,N_8521,N_8881);
nor UO_477 (O_477,N_7636,N_7601);
or UO_478 (O_478,N_9679,N_9852);
nand UO_479 (O_479,N_9525,N_7976);
nand UO_480 (O_480,N_8499,N_9790);
nor UO_481 (O_481,N_8726,N_8408);
or UO_482 (O_482,N_7806,N_9644);
and UO_483 (O_483,N_7580,N_9712);
nor UO_484 (O_484,N_9161,N_9846);
or UO_485 (O_485,N_8381,N_8770);
and UO_486 (O_486,N_7728,N_8348);
nor UO_487 (O_487,N_7502,N_7516);
nand UO_488 (O_488,N_9267,N_9482);
xor UO_489 (O_489,N_8879,N_8575);
or UO_490 (O_490,N_8186,N_8592);
nor UO_491 (O_491,N_7538,N_7743);
nand UO_492 (O_492,N_9210,N_9196);
nor UO_493 (O_493,N_9069,N_8049);
nor UO_494 (O_494,N_8607,N_8335);
nor UO_495 (O_495,N_9835,N_8054);
nand UO_496 (O_496,N_8961,N_7509);
nand UO_497 (O_497,N_9998,N_9347);
and UO_498 (O_498,N_9882,N_8390);
or UO_499 (O_499,N_9601,N_8774);
nand UO_500 (O_500,N_8363,N_8459);
or UO_501 (O_501,N_7950,N_8886);
nand UO_502 (O_502,N_9317,N_9714);
and UO_503 (O_503,N_9252,N_9292);
nand UO_504 (O_504,N_8892,N_7679);
nand UO_505 (O_505,N_8185,N_9464);
nand UO_506 (O_506,N_7680,N_8438);
and UO_507 (O_507,N_8149,N_8231);
and UO_508 (O_508,N_7924,N_8828);
nor UO_509 (O_509,N_9534,N_7568);
nor UO_510 (O_510,N_7535,N_9090);
nor UO_511 (O_511,N_8861,N_8990);
or UO_512 (O_512,N_8542,N_9463);
nand UO_513 (O_513,N_8476,N_8732);
and UO_514 (O_514,N_7611,N_8009);
and UO_515 (O_515,N_8766,N_7706);
or UO_516 (O_516,N_8631,N_9247);
nor UO_517 (O_517,N_8196,N_8220);
and UO_518 (O_518,N_9311,N_8628);
nand UO_519 (O_519,N_9902,N_8528);
xor UO_520 (O_520,N_9095,N_8448);
or UO_521 (O_521,N_7550,N_9068);
nor UO_522 (O_522,N_7779,N_7928);
and UO_523 (O_523,N_8812,N_8724);
nand UO_524 (O_524,N_8244,N_7646);
and UO_525 (O_525,N_7788,N_7866);
and UO_526 (O_526,N_7957,N_7529);
or UO_527 (O_527,N_8260,N_9885);
or UO_528 (O_528,N_8319,N_7730);
nor UO_529 (O_529,N_7659,N_8094);
or UO_530 (O_530,N_7970,N_9898);
and UO_531 (O_531,N_7525,N_7830);
and UO_532 (O_532,N_8854,N_8167);
or UO_533 (O_533,N_9886,N_7887);
nand UO_534 (O_534,N_8640,N_9952);
and UO_535 (O_535,N_8113,N_8388);
and UO_536 (O_536,N_7589,N_7504);
or UO_537 (O_537,N_8280,N_8625);
nand UO_538 (O_538,N_8958,N_7721);
or UO_539 (O_539,N_9316,N_8805);
or UO_540 (O_540,N_9078,N_7618);
nand UO_541 (O_541,N_8818,N_9040);
nand UO_542 (O_542,N_7796,N_7530);
and UO_543 (O_543,N_9810,N_7748);
nor UO_544 (O_544,N_9286,N_7822);
or UO_545 (O_545,N_8275,N_8876);
or UO_546 (O_546,N_8852,N_9703);
nand UO_547 (O_547,N_9043,N_9323);
xnor UO_548 (O_548,N_8622,N_9632);
nand UO_549 (O_549,N_7552,N_8846);
or UO_550 (O_550,N_8595,N_8475);
and UO_551 (O_551,N_9743,N_9423);
and UO_552 (O_552,N_9870,N_8718);
or UO_553 (O_553,N_8297,N_7770);
or UO_554 (O_554,N_9681,N_9271);
nor UO_555 (O_555,N_7583,N_9376);
and UO_556 (O_556,N_8468,N_8581);
nand UO_557 (O_557,N_8214,N_9895);
nand UO_558 (O_558,N_8911,N_9837);
and UO_559 (O_559,N_9277,N_7697);
and UO_560 (O_560,N_8518,N_8488);
or UO_561 (O_561,N_9897,N_8681);
nand UO_562 (O_562,N_9657,N_8953);
nor UO_563 (O_563,N_8758,N_8840);
xnor UO_564 (O_564,N_9132,N_8345);
nand UO_565 (O_565,N_9702,N_7513);
or UO_566 (O_566,N_9046,N_9693);
nand UO_567 (O_567,N_8563,N_8847);
nor UO_568 (O_568,N_9605,N_8604);
and UO_569 (O_569,N_7556,N_7956);
nand UO_570 (O_570,N_7773,N_7908);
or UO_571 (O_571,N_8964,N_7674);
nand UO_572 (O_572,N_9216,N_8517);
and UO_573 (O_573,N_8917,N_8613);
and UO_574 (O_574,N_7734,N_8271);
nand UO_575 (O_575,N_8701,N_9164);
or UO_576 (O_576,N_8908,N_8096);
xor UO_577 (O_577,N_8359,N_9054);
or UO_578 (O_578,N_8509,N_9691);
and UO_579 (O_579,N_7586,N_9733);
nor UO_580 (O_580,N_8100,N_8815);
or UO_581 (O_581,N_9654,N_9474);
nor UO_582 (O_582,N_9738,N_8480);
or UO_583 (O_583,N_9340,N_9401);
or UO_584 (O_584,N_8216,N_9355);
nor UO_585 (O_585,N_9660,N_8067);
nand UO_586 (O_586,N_9176,N_7647);
xor UO_587 (O_587,N_9532,N_8136);
nand UO_588 (O_588,N_7877,N_8316);
and UO_589 (O_589,N_8796,N_9667);
nand UO_590 (O_590,N_8387,N_7699);
xor UO_591 (O_591,N_8662,N_9204);
or UO_592 (O_592,N_9686,N_8453);
xor UO_593 (O_593,N_9167,N_9304);
or UO_594 (O_594,N_8085,N_7974);
nand UO_595 (O_595,N_8472,N_7982);
or UO_596 (O_596,N_8150,N_7975);
nand UO_597 (O_597,N_8263,N_8603);
and UO_598 (O_598,N_9815,N_9429);
nand UO_599 (O_599,N_9512,N_8939);
or UO_600 (O_600,N_8845,N_7660);
nor UO_601 (O_601,N_9563,N_9756);
nand UO_602 (O_602,N_9480,N_9999);
and UO_603 (O_603,N_7610,N_8763);
nor UO_604 (O_604,N_7593,N_9105);
xnor UO_605 (O_605,N_9988,N_8965);
nand UO_606 (O_606,N_8733,N_8573);
nor UO_607 (O_607,N_9027,N_9130);
nand UO_608 (O_608,N_7686,N_9269);
or UO_609 (O_609,N_9158,N_8093);
nand UO_610 (O_610,N_7526,N_7619);
or UO_611 (O_611,N_8288,N_8893);
or UO_612 (O_612,N_7989,N_7805);
nor UO_613 (O_613,N_9513,N_9923);
nand UO_614 (O_614,N_8425,N_8923);
nand UO_615 (O_615,N_9004,N_9209);
and UO_616 (O_616,N_9584,N_9123);
nand UO_617 (O_617,N_8272,N_8682);
nor UO_618 (O_618,N_8072,N_9120);
and UO_619 (O_619,N_9968,N_9541);
nor UO_620 (O_620,N_9181,N_8074);
or UO_621 (O_621,N_8951,N_8610);
or UO_622 (O_622,N_8680,N_9510);
nor UO_623 (O_623,N_8524,N_7581);
nor UO_624 (O_624,N_9963,N_7807);
and UO_625 (O_625,N_9643,N_8161);
nor UO_626 (O_626,N_8065,N_7823);
or UO_627 (O_627,N_8171,N_7884);
or UO_628 (O_628,N_9635,N_9649);
xor UO_629 (O_629,N_9848,N_9146);
nand UO_630 (O_630,N_8279,N_9459);
and UO_631 (O_631,N_8555,N_7501);
nand UO_632 (O_632,N_7574,N_8925);
and UO_633 (O_633,N_8735,N_9218);
or UO_634 (O_634,N_9458,N_8792);
or UO_635 (O_635,N_8374,N_9997);
xor UO_636 (O_636,N_9842,N_9974);
or UO_637 (O_637,N_8354,N_8529);
nand UO_638 (O_638,N_8223,N_8469);
and UO_639 (O_639,N_7792,N_8985);
xor UO_640 (O_640,N_9358,N_8446);
nor UO_641 (O_641,N_7614,N_9381);
and UO_642 (O_642,N_8158,N_9215);
or UO_643 (O_643,N_9017,N_8864);
nand UO_644 (O_644,N_9951,N_8533);
or UO_645 (O_645,N_9794,N_9696);
nand UO_646 (O_646,N_8142,N_8482);
or UO_647 (O_647,N_7840,N_7613);
and UO_648 (O_648,N_8169,N_9628);
xor UO_649 (O_649,N_8290,N_8462);
or UO_650 (O_650,N_8261,N_8199);
nand UO_651 (O_651,N_8276,N_7997);
xor UO_652 (O_652,N_7864,N_9246);
and UO_653 (O_653,N_9529,N_9016);
or UO_654 (O_654,N_9348,N_7708);
or UO_655 (O_655,N_8011,N_8910);
nor UO_656 (O_656,N_8978,N_9106);
nor UO_657 (O_657,N_9697,N_7911);
or UO_658 (O_658,N_7714,N_9736);
and UO_659 (O_659,N_8842,N_7769);
or UO_660 (O_660,N_7718,N_8165);
nand UO_661 (O_661,N_8885,N_8602);
nor UO_662 (O_662,N_9645,N_7681);
nor UO_663 (O_663,N_7901,N_7763);
or UO_664 (O_664,N_9710,N_8380);
or UO_665 (O_665,N_9274,N_7710);
and UO_666 (O_666,N_8172,N_8233);
or UO_667 (O_667,N_8015,N_8097);
nor UO_668 (O_668,N_9492,N_8236);
nor UO_669 (O_669,N_9062,N_8794);
and UO_670 (O_670,N_9993,N_8515);
and UO_671 (O_671,N_8114,N_7967);
nor UO_672 (O_672,N_8008,N_8164);
xor UO_673 (O_673,N_9387,N_7874);
and UO_674 (O_674,N_8334,N_8526);
or UO_675 (O_675,N_8987,N_9502);
xor UO_676 (O_676,N_7827,N_7625);
nand UO_677 (O_677,N_9531,N_8382);
and UO_678 (O_678,N_8669,N_8960);
or UO_679 (O_679,N_7553,N_8092);
nand UO_680 (O_680,N_9491,N_9972);
nand UO_681 (O_681,N_7977,N_7503);
nor UO_682 (O_682,N_7899,N_8311);
xor UO_683 (O_683,N_8504,N_9430);
or UO_684 (O_684,N_8432,N_9890);
nor UO_685 (O_685,N_7994,N_9669);
xor UO_686 (O_686,N_9773,N_7666);
nand UO_687 (O_687,N_7809,N_8871);
nand UO_688 (O_688,N_7696,N_9879);
nor UO_689 (O_689,N_9260,N_9184);
xor UO_690 (O_690,N_8050,N_8213);
nand UO_691 (O_691,N_8200,N_8576);
nor UO_692 (O_692,N_8637,N_8431);
or UO_693 (O_693,N_7981,N_8106);
nor UO_694 (O_694,N_8710,N_7850);
or UO_695 (O_695,N_8713,N_9223);
and UO_696 (O_696,N_8624,N_8424);
and UO_697 (O_697,N_9572,N_8731);
and UO_698 (O_698,N_9394,N_9219);
and UO_699 (O_699,N_8577,N_9089);
nand UO_700 (O_700,N_8883,N_8410);
and UO_701 (O_701,N_8393,N_8415);
xnor UO_702 (O_702,N_9143,N_9565);
and UO_703 (O_703,N_9983,N_7665);
nor UO_704 (O_704,N_9729,N_8103);
and UO_705 (O_705,N_9243,N_9688);
nand UO_706 (O_706,N_8609,N_9212);
or UO_707 (O_707,N_9749,N_9445);
xor UO_708 (O_708,N_7566,N_8998);
nor UO_709 (O_709,N_8860,N_9074);
nor UO_710 (O_710,N_8569,N_9707);
and UO_711 (O_711,N_8207,N_7848);
and UO_712 (O_712,N_8902,N_9556);
nor UO_713 (O_713,N_8228,N_7772);
and UO_714 (O_714,N_8915,N_9851);
nand UO_715 (O_715,N_8493,N_7973);
nor UO_716 (O_716,N_7961,N_9388);
nand UO_717 (O_717,N_8389,N_9713);
or UO_718 (O_718,N_7663,N_9770);
nand UO_719 (O_719,N_9229,N_8527);
xor UO_720 (O_720,N_8679,N_9297);
or UO_721 (O_721,N_7587,N_9559);
nor UO_722 (O_722,N_8808,N_8392);
nand UO_723 (O_723,N_8188,N_7540);
or UO_724 (O_724,N_8930,N_9822);
nand UO_725 (O_725,N_9201,N_8793);
or UO_726 (O_726,N_7953,N_8753);
or UO_727 (O_727,N_8862,N_7885);
or UO_728 (O_728,N_9279,N_9540);
nand UO_729 (O_729,N_9003,N_8043);
and UO_730 (O_730,N_8799,N_8112);
and UO_731 (O_731,N_9690,N_9598);
nand UO_732 (O_732,N_9656,N_9420);
nor UO_733 (O_733,N_9664,N_8176);
nand UO_734 (O_734,N_8968,N_8995);
or UO_735 (O_735,N_9295,N_9173);
and UO_736 (O_736,N_7988,N_7941);
nand UO_737 (O_737,N_9362,N_8426);
xor UO_738 (O_738,N_9441,N_9964);
or UO_739 (O_739,N_8525,N_9834);
or UO_740 (O_740,N_9195,N_8162);
xor UO_741 (O_741,N_9618,N_8903);
xnor UO_742 (O_742,N_8513,N_9434);
xor UO_743 (O_743,N_7641,N_7597);
and UO_744 (O_744,N_7603,N_8837);
nor UO_745 (O_745,N_8795,N_7629);
xor UO_746 (O_746,N_8021,N_8486);
or UO_747 (O_747,N_8988,N_8349);
nor UO_748 (O_748,N_9205,N_7594);
and UO_749 (O_749,N_9287,N_8215);
xnor UO_750 (O_750,N_8698,N_9577);
nand UO_751 (O_751,N_8938,N_9444);
nor UO_752 (O_752,N_8151,N_8331);
and UO_753 (O_753,N_9627,N_9328);
nor UO_754 (O_754,N_9543,N_9861);
nand UO_755 (O_755,N_8327,N_7653);
nor UO_756 (O_756,N_9331,N_7828);
or UO_757 (O_757,N_8659,N_7810);
nand UO_758 (O_758,N_9503,N_8944);
nor UO_759 (O_759,N_9590,N_8259);
nor UO_760 (O_760,N_8762,N_9197);
nor UO_761 (O_761,N_8423,N_9919);
and UO_762 (O_762,N_9615,N_7716);
and UO_763 (O_763,N_9022,N_8416);
nand UO_764 (O_764,N_7859,N_8099);
nand UO_765 (O_765,N_8853,N_8863);
xor UO_766 (O_766,N_8686,N_9730);
and UO_767 (O_767,N_7667,N_9594);
xor UO_768 (O_768,N_7569,N_9956);
and UO_769 (O_769,N_8647,N_9410);
and UO_770 (O_770,N_9772,N_7640);
nor UO_771 (O_771,N_8740,N_7622);
nand UO_772 (O_772,N_9893,N_7917);
or UO_773 (O_773,N_8782,N_8063);
nor UO_774 (O_774,N_9829,N_7751);
nor UO_775 (O_775,N_8972,N_9940);
or UO_776 (O_776,N_7564,N_8251);
or UO_777 (O_777,N_8677,N_8376);
nand UO_778 (O_778,N_7760,N_7620);
or UO_779 (O_779,N_9395,N_7800);
and UO_780 (O_780,N_7798,N_8999);
nand UO_781 (O_781,N_9887,N_9671);
nand UO_782 (O_782,N_8945,N_8064);
nand UO_783 (O_783,N_7888,N_9437);
and UO_784 (O_784,N_9728,N_9585);
nand UO_785 (O_785,N_9843,N_7617);
nand UO_786 (O_786,N_7825,N_7791);
and UO_787 (O_787,N_8709,N_8204);
and UO_788 (O_788,N_9934,N_9299);
nand UO_789 (O_789,N_8075,N_9369);
and UO_790 (O_790,N_9400,N_8126);
or UO_791 (O_791,N_7938,N_8378);
nor UO_792 (O_792,N_9685,N_9149);
nand UO_793 (O_793,N_8006,N_9641);
nand UO_794 (O_794,N_8549,N_9262);
nor UO_795 (O_795,N_9812,N_9127);
and UO_796 (O_796,N_8082,N_7698);
nand UO_797 (O_797,N_7656,N_8206);
nor UO_798 (O_798,N_9720,N_8487);
nand UO_799 (O_799,N_9884,N_9063);
or UO_800 (O_800,N_8355,N_9065);
nor UO_801 (O_801,N_9783,N_8435);
xnor UO_802 (O_802,N_8729,N_7693);
or UO_803 (O_803,N_9191,N_9025);
nand UO_804 (O_804,N_8102,N_9926);
and UO_805 (O_805,N_9876,N_7852);
xor UO_806 (O_806,N_8973,N_9991);
nand UO_807 (O_807,N_9412,N_8282);
nand UO_808 (O_808,N_7882,N_7541);
and UO_809 (O_809,N_9866,N_9824);
or UO_810 (O_810,N_9938,N_8904);
nand UO_811 (O_811,N_8556,N_9719);
nand UO_812 (O_812,N_9908,N_9314);
and UO_813 (O_813,N_9498,N_8020);
nor UO_814 (O_814,N_8974,N_7962);
nand UO_815 (O_815,N_8623,N_9599);
or UO_816 (O_816,N_9058,N_7715);
nand UO_817 (O_817,N_9634,N_9717);
or UO_818 (O_818,N_9500,N_9200);
nand UO_819 (O_819,N_8614,N_9985);
or UO_820 (O_820,N_9334,N_8098);
nand UO_821 (O_821,N_8201,N_8234);
or UO_822 (O_822,N_9192,N_8940);
nand UO_823 (O_823,N_9642,N_9910);
and UO_824 (O_824,N_8768,N_8317);
or UO_825 (O_825,N_8343,N_8630);
and UO_826 (O_826,N_9636,N_7555);
and UO_827 (O_827,N_9283,N_9814);
or UO_828 (O_828,N_9023,N_9235);
nor UO_829 (O_829,N_8372,N_8035);
and UO_830 (O_830,N_8254,N_8352);
or UO_831 (O_831,N_7754,N_9475);
nor UO_832 (O_832,N_8377,N_8047);
nand UO_833 (O_833,N_8080,N_9992);
or UO_834 (O_834,N_7673,N_9259);
nor UO_835 (O_835,N_9862,N_8621);
nor UO_836 (O_836,N_8989,N_7717);
nand UO_837 (O_837,N_8878,N_7705);
nand UO_838 (O_838,N_8829,N_7752);
nand UO_839 (O_839,N_7996,N_9194);
or UO_840 (O_840,N_9257,N_7528);
nor UO_841 (O_841,N_8720,N_9961);
and UO_842 (O_842,N_9631,N_8353);
nand UO_843 (O_843,N_9408,N_7931);
nand UO_844 (O_844,N_7668,N_7781);
or UO_845 (O_845,N_8252,N_8848);
nand UO_846 (O_846,N_8182,N_9041);
and UO_847 (O_847,N_7534,N_8409);
nand UO_848 (O_848,N_7964,N_9611);
nand UO_849 (O_849,N_9440,N_9251);
and UO_850 (O_850,N_8159,N_9560);
nor UO_851 (O_851,N_8243,N_9552);
or UO_852 (O_852,N_8627,N_9428);
xor UO_853 (O_853,N_7662,N_8083);
and UO_854 (O_854,N_9044,N_8619);
and UO_855 (O_855,N_7510,N_9844);
xnor UO_856 (O_856,N_8606,N_9581);
nand UO_857 (O_857,N_8653,N_9077);
nand UO_858 (O_858,N_9984,N_8337);
nor UO_859 (O_859,N_8258,N_9336);
nand UO_860 (O_860,N_7759,N_9308);
and UO_861 (O_861,N_9676,N_8026);
nand UO_862 (O_862,N_9807,N_8777);
and UO_863 (O_863,N_8827,N_7897);
nor UO_864 (O_864,N_7546,N_8166);
nor UO_865 (O_865,N_7793,N_8239);
nor UO_866 (O_866,N_9766,N_8148);
or UO_867 (O_867,N_8208,N_9366);
or UO_868 (O_868,N_9315,N_9932);
nand UO_869 (O_869,N_8457,N_9469);
or UO_870 (O_870,N_8867,N_9855);
or UO_871 (O_871,N_9718,N_9943);
nand UO_872 (O_872,N_8761,N_8541);
nor UO_873 (O_873,N_9012,N_7814);
nand UO_874 (O_874,N_7573,N_9689);
nor UO_875 (O_875,N_8543,N_9796);
nor UO_876 (O_876,N_9580,N_8738);
nor UO_877 (O_877,N_8532,N_7984);
and UO_878 (O_878,N_9973,N_8537);
xor UO_879 (O_879,N_7726,N_7922);
and UO_880 (O_880,N_7655,N_7584);
nand UO_881 (O_881,N_8656,N_8304);
nand UO_882 (O_882,N_8672,N_9131);
nor UO_883 (O_883,N_8632,N_9306);
nor UO_884 (O_884,N_9955,N_8111);
nand UO_885 (O_885,N_9506,N_9528);
nor UO_886 (O_886,N_9097,N_9253);
nand UO_887 (O_887,N_9374,N_8018);
nand UO_888 (O_888,N_8012,N_8511);
and UO_889 (O_889,N_7784,N_8512);
or UO_890 (O_890,N_8599,N_9234);
and UO_891 (O_891,N_9439,N_8564);
nor UO_892 (O_892,N_8016,N_8407);
nor UO_893 (O_893,N_8295,N_8442);
and UO_894 (O_894,N_8302,N_8700);
nor UO_895 (O_895,N_9094,N_9031);
or UO_896 (O_896,N_9386,N_8324);
nor UO_897 (O_897,N_7816,N_7604);
and UO_898 (O_898,N_9744,N_9573);
nand UO_899 (O_899,N_9748,N_7835);
nor UO_900 (O_900,N_9764,N_8813);
nand UO_901 (O_901,N_9588,N_9384);
or UO_902 (O_902,N_7642,N_9761);
or UO_903 (O_903,N_9258,N_8530);
nand UO_904 (O_904,N_9427,N_8296);
xor UO_905 (O_905,N_9160,N_9517);
nand UO_906 (O_906,N_9338,N_9451);
and UO_907 (O_907,N_9760,N_8400);
nand UO_908 (O_908,N_9626,N_9432);
xnor UO_909 (O_909,N_9353,N_9034);
nor UO_910 (O_910,N_8291,N_9856);
or UO_911 (O_911,N_9962,N_8895);
nand UO_912 (O_912,N_7532,N_7701);
nand UO_913 (O_913,N_9816,N_9776);
nand UO_914 (O_914,N_7557,N_7771);
nor UO_915 (O_915,N_9803,N_8051);
nor UO_916 (O_916,N_9945,N_8107);
nor UO_917 (O_917,N_7909,N_7575);
or UO_918 (O_918,N_9711,N_8869);
nor UO_919 (O_919,N_8130,N_8076);
and UO_920 (O_920,N_9519,N_8283);
and UO_921 (O_921,N_9823,N_9153);
nor UO_922 (O_922,N_7863,N_8673);
nor UO_923 (O_923,N_8516,N_8184);
nand UO_924 (O_924,N_8019,N_8875);
nand UO_925 (O_925,N_9449,N_7845);
or UO_926 (O_926,N_9114,N_8877);
nand UO_927 (O_927,N_8642,N_9860);
nand UO_928 (O_928,N_8823,N_8122);
nor UO_929 (O_929,N_8128,N_8369);
nand UO_930 (O_930,N_8492,N_9777);
or UO_931 (O_931,N_8891,N_7554);
nand UO_932 (O_932,N_9753,N_9059);
nand UO_933 (O_933,N_8371,N_9524);
or UO_934 (O_934,N_7561,N_7980);
nor UO_935 (O_935,N_8294,N_9298);
nor UO_936 (O_936,N_7661,N_7595);
or UO_937 (O_937,N_9142,N_9291);
nand UO_938 (O_938,N_9254,N_9853);
or UO_939 (O_939,N_9231,N_8135);
and UO_940 (O_940,N_8844,N_8147);
and UO_941 (O_941,N_9431,N_8850);
nand UO_942 (O_942,N_7916,N_9249);
nor UO_943 (O_943,N_7609,N_9739);
or UO_944 (O_944,N_9648,N_9990);
and UO_945 (O_945,N_7966,N_9597);
or UO_946 (O_946,N_8954,N_8748);
or UO_947 (O_947,N_9818,N_7787);
nor UO_948 (O_948,N_8725,N_7676);
or UO_949 (O_949,N_8983,N_9472);
or UO_950 (O_950,N_9060,N_8153);
and UO_951 (O_951,N_9354,N_9049);
nand UO_952 (O_952,N_8467,N_8436);
nand UO_953 (O_953,N_8222,N_9448);
and UO_954 (O_954,N_9203,N_8618);
nand UO_955 (O_955,N_9307,N_9709);
nand UO_956 (O_956,N_9670,N_8403);
or UO_957 (O_957,N_8825,N_9579);
nand UO_958 (O_958,N_9663,N_9418);
nand UO_959 (O_959,N_9056,N_8396);
xor UO_960 (O_960,N_9994,N_8705);
or UO_961 (O_961,N_7729,N_7522);
xnor UO_962 (O_962,N_7695,N_9048);
nand UO_963 (O_963,N_9672,N_8790);
and UO_964 (O_964,N_8059,N_9740);
or UO_965 (O_965,N_7766,N_8132);
nor UO_966 (O_966,N_9801,N_9378);
xnor UO_967 (O_967,N_9526,N_8170);
nor UO_968 (O_968,N_8759,N_9038);
or UO_969 (O_969,N_8227,N_8519);
or UO_970 (O_970,N_8639,N_8238);
nand UO_971 (O_971,N_8997,N_7995);
or UO_972 (O_972,N_9779,N_9830);
nand UO_973 (O_973,N_7883,N_8250);
or UO_974 (O_974,N_8857,N_9881);
nand UO_975 (O_975,N_7889,N_8711);
and UO_976 (O_976,N_9883,N_9282);
nand UO_977 (O_977,N_7582,N_9057);
or UO_978 (O_978,N_9122,N_8413);
and UO_979 (O_979,N_8900,N_8634);
and UO_980 (O_980,N_8590,N_7735);
or UO_981 (O_981,N_7670,N_9478);
nor UO_982 (O_982,N_8906,N_7621);
nand UO_983 (O_983,N_7722,N_7598);
xnor UO_984 (O_984,N_9419,N_7891);
and UO_985 (O_985,N_8053,N_7689);
and UO_986 (O_986,N_9546,N_9496);
or UO_987 (O_987,N_9646,N_7537);
nand UO_988 (O_988,N_8145,N_9182);
nor UO_989 (O_989,N_9880,N_9413);
xor UO_990 (O_990,N_7818,N_8967);
nor UO_991 (O_991,N_8916,N_8786);
nand UO_992 (O_992,N_8190,N_9086);
xnor UO_993 (O_993,N_8306,N_9033);
and UO_994 (O_994,N_8155,N_7747);
xor UO_995 (O_995,N_7919,N_9925);
or UO_996 (O_996,N_8370,N_7520);
nor UO_997 (O_997,N_7731,N_8178);
or UO_998 (O_998,N_9414,N_9222);
and UO_999 (O_999,N_9101,N_9493);
nor UO_1000 (O_1000,N_8809,N_8267);
nand UO_1001 (O_1001,N_7637,N_9706);
and UO_1002 (O_1002,N_8554,N_9211);
or UO_1003 (O_1003,N_9272,N_9406);
nand UO_1004 (O_1004,N_8062,N_9359);
nand UO_1005 (O_1005,N_8309,N_9937);
and UO_1006 (O_1006,N_7939,N_7837);
xnor UO_1007 (O_1007,N_8764,N_8934);
and UO_1008 (O_1008,N_8503,N_9174);
nand UO_1009 (O_1009,N_8670,N_9220);
nand UO_1010 (O_1010,N_9329,N_7858);
nor UO_1011 (O_1011,N_7539,N_8314);
nand UO_1012 (O_1012,N_9722,N_7936);
nor UO_1013 (O_1013,N_8992,N_9849);
nor UO_1014 (O_1014,N_9227,N_9093);
or UO_1015 (O_1015,N_7817,N_9170);
nor UO_1016 (O_1016,N_7972,N_9771);
or UO_1017 (O_1017,N_9575,N_7971);
nand UO_1018 (O_1018,N_7669,N_8156);
nand UO_1019 (O_1019,N_7684,N_9762);
and UO_1020 (O_1020,N_9140,N_8909);
xnor UO_1021 (O_1021,N_8366,N_9092);
and UO_1022 (O_1022,N_7507,N_7875);
and UO_1023 (O_1023,N_9417,N_8003);
nand UO_1024 (O_1024,N_7913,N_9389);
or UO_1025 (O_1025,N_9616,N_8205);
nand UO_1026 (O_1026,N_7865,N_8617);
and UO_1027 (O_1027,N_8754,N_8570);
or UO_1028 (O_1028,N_7739,N_8088);
xnor UO_1029 (O_1029,N_9367,N_9630);
nand UO_1030 (O_1030,N_8320,N_8597);
nor UO_1031 (O_1031,N_7999,N_9774);
nand UO_1032 (O_1032,N_9907,N_8560);
nor UO_1033 (O_1033,N_9924,N_9865);
nand UO_1034 (O_1034,N_8452,N_8336);
nand UO_1035 (O_1035,N_9516,N_8890);
and UO_1036 (O_1036,N_8898,N_7606);
or UO_1037 (O_1037,N_9859,N_8936);
and UO_1038 (O_1038,N_8454,N_8924);
nand UO_1039 (O_1039,N_7789,N_8544);
nand UO_1040 (O_1040,N_8127,N_8405);
and UO_1041 (O_1041,N_9542,N_9371);
or UO_1042 (O_1042,N_8678,N_9826);
xnor UO_1043 (O_1043,N_7649,N_8836);
nand UO_1044 (O_1044,N_7867,N_9623);
and UO_1045 (O_1045,N_7712,N_9947);
xor UO_1046 (O_1046,N_9301,N_9544);
or UO_1047 (O_1047,N_8807,N_7868);
nand UO_1048 (O_1048,N_8780,N_8175);
or UO_1049 (O_1049,N_9064,N_9562);
xnor UO_1050 (O_1050,N_9289,N_9799);
nand UO_1051 (O_1051,N_8420,N_9792);
or UO_1052 (O_1052,N_7744,N_9013);
nor UO_1053 (O_1053,N_8344,N_9530);
nand UO_1054 (O_1054,N_8507,N_9337);
nand UO_1055 (O_1055,N_8757,N_7853);
or UO_1056 (O_1056,N_8061,N_9833);
and UO_1057 (O_1057,N_8838,N_9151);
xor UO_1058 (O_1058,N_8071,N_9978);
nor UO_1059 (O_1059,N_9125,N_9724);
nor UO_1060 (O_1060,N_9746,N_9121);
and UO_1061 (O_1061,N_9840,N_9499);
nand UO_1062 (O_1062,N_8545,N_8769);
xor UO_1063 (O_1063,N_8090,N_8180);
and UO_1064 (O_1064,N_8357,N_7624);
and UO_1065 (O_1065,N_8957,N_8105);
nand UO_1066 (O_1066,N_7878,N_9944);
nor UO_1067 (O_1067,N_9958,N_8582);
and UO_1068 (O_1068,N_8510,N_8401);
nor UO_1069 (O_1069,N_9545,N_9793);
nor UO_1070 (O_1070,N_9051,N_9765);
and UO_1071 (O_1071,N_9467,N_9967);
nand UO_1072 (O_1072,N_8747,N_8417);
or UO_1073 (O_1073,N_7746,N_8520);
nor UO_1074 (O_1074,N_8248,N_8000);
nor UO_1075 (O_1075,N_8465,N_8044);
xnor UO_1076 (O_1076,N_8671,N_9939);
or UO_1077 (O_1077,N_9661,N_9894);
nand UO_1078 (O_1078,N_8918,N_7506);
xor UO_1079 (O_1079,N_7559,N_8608);
nor UO_1080 (O_1080,N_8785,N_7652);
nor UO_1081 (O_1081,N_8365,N_9169);
xor UO_1082 (O_1082,N_8461,N_9375);
nor UO_1083 (O_1083,N_9073,N_8574);
nor UO_1084 (O_1084,N_7843,N_9265);
or UO_1085 (O_1085,N_7844,N_7879);
nor UO_1086 (O_1086,N_7794,N_8007);
or UO_1087 (O_1087,N_8707,N_7945);
xor UO_1088 (O_1088,N_9638,N_7517);
xor UO_1089 (O_1089,N_8565,N_8437);
nor UO_1090 (O_1090,N_8253,N_8820);
nor UO_1091 (O_1091,N_9010,N_8117);
and UO_1092 (O_1092,N_8146,N_9088);
and UO_1093 (O_1093,N_9832,N_8471);
and UO_1094 (O_1094,N_7904,N_8040);
and UO_1095 (O_1095,N_8571,N_9390);
or UO_1096 (O_1096,N_9398,N_9716);
or UO_1097 (O_1097,N_8299,N_9551);
and UO_1098 (O_1098,N_8773,N_9224);
and UO_1099 (O_1099,N_9206,N_8558);
nor UO_1100 (O_1100,N_8089,N_8784);
nor UO_1101 (O_1101,N_9076,N_8601);
nor UO_1102 (O_1102,N_7952,N_8242);
or UO_1103 (O_1103,N_9199,N_8736);
and UO_1104 (O_1104,N_9083,N_8587);
nor UO_1105 (O_1105,N_8368,N_9363);
or UO_1106 (O_1106,N_8626,N_9457);
and UO_1107 (O_1107,N_8502,N_9960);
xor UO_1108 (O_1108,N_8937,N_7777);
nand UO_1109 (O_1109,N_9726,N_8776);
nor UO_1110 (O_1110,N_7963,N_9653);
nand UO_1111 (O_1111,N_7572,N_8635);
nor UO_1112 (O_1112,N_8806,N_8395);
and UO_1113 (O_1113,N_7683,N_8181);
nand UO_1114 (O_1114,N_7737,N_9442);
and UO_1115 (O_1115,N_8284,N_9280);
or UO_1116 (O_1116,N_8495,N_7671);
or UO_1117 (O_1117,N_8154,N_8341);
and UO_1118 (O_1118,N_7700,N_8338);
and UO_1119 (O_1119,N_9476,N_8551);
or UO_1120 (O_1120,N_8749,N_7930);
and UO_1121 (O_1121,N_9981,N_8547);
or UO_1122 (O_1122,N_7576,N_8567);
and UO_1123 (O_1123,N_9396,N_8101);
nand UO_1124 (O_1124,N_7616,N_8104);
and UO_1125 (O_1125,N_9028,N_9450);
and UO_1126 (O_1126,N_8332,N_7732);
nor UO_1127 (O_1127,N_8313,N_8318);
and UO_1128 (O_1128,N_8245,N_8880);
nor UO_1129 (O_1129,N_9507,N_9479);
or UO_1130 (O_1130,N_9107,N_8921);
nor UO_1131 (O_1131,N_9742,N_9549);
and UO_1132 (O_1132,N_7691,N_8665);
nand UO_1133 (O_1133,N_9250,N_7638);
or UO_1134 (O_1134,N_8268,N_9813);
or UO_1135 (O_1135,N_8611,N_8087);
nand UO_1136 (O_1136,N_9082,N_9838);
or UO_1137 (O_1137,N_8141,N_8760);
and UO_1138 (O_1138,N_8589,N_8991);
or UO_1139 (O_1139,N_7821,N_8485);
nand UO_1140 (O_1140,N_9904,N_9024);
and UO_1141 (O_1141,N_7940,N_8489);
or UO_1142 (O_1142,N_8676,N_8017);
and UO_1143 (O_1143,N_9548,N_8108);
xor UO_1144 (O_1144,N_8704,N_8095);
and UO_1145 (O_1145,N_8262,N_7639);
or UO_1146 (O_1146,N_7608,N_9305);
nand UO_1147 (O_1147,N_9986,N_8303);
nand UO_1148 (O_1148,N_8384,N_8351);
nand UO_1149 (O_1149,N_9582,N_7565);
nand UO_1150 (O_1150,N_9344,N_8221);
nor UO_1151 (O_1151,N_9456,N_9261);
nor UO_1152 (O_1152,N_9166,N_7869);
and UO_1153 (O_1153,N_7965,N_7925);
nor UO_1154 (O_1154,N_8514,N_8179);
or UO_1155 (O_1155,N_7799,N_8274);
or UO_1156 (O_1156,N_9473,N_8397);
nor UO_1157 (O_1157,N_7757,N_8787);
or UO_1158 (O_1158,N_8694,N_8066);
and UO_1159 (O_1159,N_8819,N_9278);
nor UO_1160 (O_1160,N_9188,N_8730);
nand UO_1161 (O_1161,N_8183,N_8434);
or UO_1162 (O_1162,N_8346,N_8433);
and UO_1163 (O_1163,N_8444,N_8841);
nand UO_1164 (O_1164,N_8333,N_9015);
nor UO_1165 (O_1165,N_9129,N_8133);
xnor UO_1166 (O_1166,N_7753,N_8811);
and UO_1167 (O_1167,N_8240,N_9000);
and UO_1168 (O_1168,N_7993,N_9877);
nand UO_1169 (O_1169,N_9873,N_9520);
or UO_1170 (O_1170,N_9208,N_9680);
or UO_1171 (O_1171,N_7892,N_8256);
or UO_1172 (O_1172,N_8030,N_7713);
nand UO_1173 (O_1173,N_9324,N_9571);
xnor UO_1174 (O_1174,N_8907,N_8055);
nand UO_1175 (O_1175,N_7632,N_7643);
nand UO_1176 (O_1176,N_9874,N_8693);
and UO_1177 (O_1177,N_8266,N_9447);
or UO_1178 (O_1178,N_9521,N_9768);
nor UO_1179 (O_1179,N_8057,N_8615);
and UO_1180 (O_1180,N_9527,N_7733);
or UO_1181 (O_1181,N_9800,N_9808);
nor UO_1182 (O_1182,N_7991,N_9617);
nor UO_1183 (O_1183,N_9889,N_9426);
nor UO_1184 (O_1184,N_9805,N_8899);
nor UO_1185 (O_1185,N_7515,N_8734);
nand UO_1186 (O_1186,N_9207,N_9018);
nand UO_1187 (O_1187,N_9071,N_9465);
and UO_1188 (O_1188,N_9405,N_8285);
and UO_1189 (O_1189,N_8144,N_8856);
nand UO_1190 (O_1190,N_7672,N_8308);
and UO_1191 (O_1191,N_9147,N_8948);
or UO_1192 (O_1192,N_8481,N_9731);
or UO_1193 (O_1193,N_7602,N_8073);
nand UO_1194 (O_1194,N_8929,N_9080);
xor UO_1195 (O_1195,N_9982,N_9723);
nor UO_1196 (O_1196,N_8046,N_7578);
or UO_1197 (O_1197,N_8187,N_9168);
nand UO_1198 (O_1198,N_9162,N_9126);
or UO_1199 (O_1199,N_8430,N_9536);
nor UO_1200 (O_1200,N_8445,N_9839);
nor UO_1201 (O_1201,N_8115,N_9111);
nand UO_1202 (O_1202,N_8584,N_7851);
nand UO_1203 (O_1203,N_8326,N_9804);
and UO_1204 (O_1204,N_7761,N_9117);
nand UO_1205 (O_1205,N_9339,N_9098);
nor UO_1206 (O_1206,N_9899,N_8289);
or UO_1207 (O_1207,N_8226,N_8767);
or UO_1208 (O_1208,N_8668,N_8896);
and UO_1209 (O_1209,N_8687,N_8775);
and UO_1210 (O_1210,N_9403,N_9875);
and UO_1211 (O_1211,N_9752,N_9007);
and UO_1212 (O_1212,N_9953,N_8447);
and UO_1213 (O_1213,N_9557,N_9596);
nor UO_1214 (O_1214,N_8943,N_7545);
xnor UO_1215 (O_1215,N_9435,N_8859);
nand UO_1216 (O_1216,N_9927,N_8996);
nand UO_1217 (O_1217,N_9784,N_8411);
nand UO_1218 (O_1218,N_8307,N_9352);
and UO_1219 (O_1219,N_9965,N_7969);
or UO_1220 (O_1220,N_8265,N_8822);
nand UO_1221 (O_1221,N_8241,N_9238);
nand UO_1222 (O_1222,N_8137,N_8897);
nand UO_1223 (O_1223,N_9872,N_8301);
nand UO_1224 (O_1224,N_8675,N_7955);
nor UO_1225 (O_1225,N_8110,N_8715);
and UO_1226 (O_1226,N_9357,N_8305);
and UO_1227 (O_1227,N_8870,N_8889);
and UO_1228 (O_1228,N_7819,N_9692);
nand UO_1229 (O_1229,N_7623,N_7804);
nor UO_1230 (O_1230,N_8932,N_9665);
or UO_1231 (O_1231,N_9019,N_9970);
nor UO_1232 (O_1232,N_9698,N_8131);
and UO_1233 (O_1233,N_7531,N_8060);
nor UO_1234 (O_1234,N_9695,N_9198);
nand UO_1235 (O_1235,N_7998,N_9869);
nand UO_1236 (O_1236,N_8832,N_7833);
nand UO_1237 (O_1237,N_9490,N_9624);
and UO_1238 (O_1238,N_9047,N_7756);
nor UO_1239 (O_1239,N_8728,N_8490);
nor UO_1240 (O_1240,N_9734,N_7786);
nor UO_1241 (O_1241,N_9202,N_8412);
xnor UO_1242 (O_1242,N_9820,N_9409);
nand UO_1243 (O_1243,N_9903,N_8810);
xnor UO_1244 (O_1244,N_9593,N_7542);
xor UO_1245 (O_1245,N_9346,N_8134);
nor UO_1246 (O_1246,N_8124,N_9032);
nor UO_1247 (O_1247,N_9326,N_9539);
nor UO_1248 (O_1248,N_9312,N_8580);
or UO_1249 (O_1249,N_7912,N_9721);
nand UO_1250 (O_1250,N_8471,N_9535);
nand UO_1251 (O_1251,N_7985,N_9277);
and UO_1252 (O_1252,N_7542,N_8100);
nor UO_1253 (O_1253,N_9377,N_9570);
nor UO_1254 (O_1254,N_8846,N_7589);
nor UO_1255 (O_1255,N_9295,N_8845);
xor UO_1256 (O_1256,N_7851,N_8509);
xor UO_1257 (O_1257,N_9572,N_8692);
xor UO_1258 (O_1258,N_9414,N_7586);
nand UO_1259 (O_1259,N_7931,N_9383);
and UO_1260 (O_1260,N_7650,N_8473);
and UO_1261 (O_1261,N_9700,N_8621);
xor UO_1262 (O_1262,N_8893,N_8810);
or UO_1263 (O_1263,N_8269,N_9624);
or UO_1264 (O_1264,N_8841,N_9299);
and UO_1265 (O_1265,N_9379,N_8314);
and UO_1266 (O_1266,N_8129,N_8075);
xor UO_1267 (O_1267,N_7742,N_7572);
nor UO_1268 (O_1268,N_9450,N_8565);
nor UO_1269 (O_1269,N_9222,N_8771);
and UO_1270 (O_1270,N_8868,N_9682);
or UO_1271 (O_1271,N_8795,N_9464);
nand UO_1272 (O_1272,N_8055,N_8786);
nor UO_1273 (O_1273,N_8545,N_9119);
nor UO_1274 (O_1274,N_8121,N_8146);
nand UO_1275 (O_1275,N_8011,N_8662);
and UO_1276 (O_1276,N_8950,N_8185);
nand UO_1277 (O_1277,N_9287,N_8282);
nor UO_1278 (O_1278,N_9067,N_9669);
and UO_1279 (O_1279,N_9657,N_8471);
and UO_1280 (O_1280,N_7736,N_9236);
and UO_1281 (O_1281,N_8361,N_8493);
and UO_1282 (O_1282,N_9179,N_9980);
or UO_1283 (O_1283,N_8920,N_9394);
nand UO_1284 (O_1284,N_8314,N_9473);
or UO_1285 (O_1285,N_9232,N_8227);
nand UO_1286 (O_1286,N_8389,N_9878);
nand UO_1287 (O_1287,N_7996,N_7896);
or UO_1288 (O_1288,N_9606,N_9182);
or UO_1289 (O_1289,N_8467,N_7747);
nand UO_1290 (O_1290,N_8513,N_8955);
nor UO_1291 (O_1291,N_8232,N_9086);
xor UO_1292 (O_1292,N_9830,N_7655);
nand UO_1293 (O_1293,N_9965,N_8446);
nand UO_1294 (O_1294,N_9681,N_9356);
nor UO_1295 (O_1295,N_9533,N_9399);
xnor UO_1296 (O_1296,N_8460,N_9206);
or UO_1297 (O_1297,N_9571,N_8455);
and UO_1298 (O_1298,N_9272,N_8103);
nor UO_1299 (O_1299,N_7998,N_8252);
or UO_1300 (O_1300,N_8495,N_9214);
and UO_1301 (O_1301,N_8908,N_8149);
or UO_1302 (O_1302,N_9382,N_8237);
and UO_1303 (O_1303,N_9369,N_9391);
and UO_1304 (O_1304,N_9688,N_9284);
or UO_1305 (O_1305,N_8613,N_9290);
or UO_1306 (O_1306,N_9791,N_9265);
xor UO_1307 (O_1307,N_8357,N_7541);
and UO_1308 (O_1308,N_9473,N_8477);
and UO_1309 (O_1309,N_8896,N_8267);
and UO_1310 (O_1310,N_9893,N_9257);
nor UO_1311 (O_1311,N_8728,N_8755);
nor UO_1312 (O_1312,N_8024,N_9480);
xnor UO_1313 (O_1313,N_8726,N_8263);
and UO_1314 (O_1314,N_7921,N_9067);
nor UO_1315 (O_1315,N_9518,N_9478);
and UO_1316 (O_1316,N_9499,N_9256);
xnor UO_1317 (O_1317,N_9184,N_8462);
xor UO_1318 (O_1318,N_9684,N_7874);
xnor UO_1319 (O_1319,N_9298,N_9527);
nand UO_1320 (O_1320,N_8122,N_8199);
nor UO_1321 (O_1321,N_8678,N_9077);
or UO_1322 (O_1322,N_9803,N_7882);
and UO_1323 (O_1323,N_9946,N_8369);
nor UO_1324 (O_1324,N_7616,N_9972);
and UO_1325 (O_1325,N_9679,N_8958);
nor UO_1326 (O_1326,N_9635,N_9378);
or UO_1327 (O_1327,N_9325,N_9691);
or UO_1328 (O_1328,N_9962,N_9956);
or UO_1329 (O_1329,N_7812,N_8627);
nor UO_1330 (O_1330,N_8023,N_9566);
and UO_1331 (O_1331,N_8105,N_7940);
nand UO_1332 (O_1332,N_8188,N_7782);
nand UO_1333 (O_1333,N_7844,N_9051);
nor UO_1334 (O_1334,N_7792,N_8854);
nor UO_1335 (O_1335,N_8156,N_8723);
xnor UO_1336 (O_1336,N_9702,N_8079);
and UO_1337 (O_1337,N_9903,N_8313);
and UO_1338 (O_1338,N_9552,N_9635);
nand UO_1339 (O_1339,N_9123,N_8452);
and UO_1340 (O_1340,N_8837,N_8955);
or UO_1341 (O_1341,N_9962,N_8500);
nor UO_1342 (O_1342,N_8417,N_7657);
and UO_1343 (O_1343,N_9308,N_9900);
or UO_1344 (O_1344,N_9120,N_8640);
nand UO_1345 (O_1345,N_7673,N_9699);
nor UO_1346 (O_1346,N_8010,N_9957);
nand UO_1347 (O_1347,N_8762,N_8495);
nor UO_1348 (O_1348,N_8143,N_9820);
nor UO_1349 (O_1349,N_9668,N_8764);
nand UO_1350 (O_1350,N_7542,N_9837);
or UO_1351 (O_1351,N_8351,N_8856);
nand UO_1352 (O_1352,N_8601,N_8712);
or UO_1353 (O_1353,N_9405,N_9904);
or UO_1354 (O_1354,N_9230,N_9605);
nand UO_1355 (O_1355,N_8405,N_9380);
xor UO_1356 (O_1356,N_9797,N_8446);
or UO_1357 (O_1357,N_7875,N_8991);
or UO_1358 (O_1358,N_8057,N_7570);
and UO_1359 (O_1359,N_9870,N_9212);
and UO_1360 (O_1360,N_8843,N_7662);
nor UO_1361 (O_1361,N_9495,N_7634);
or UO_1362 (O_1362,N_8356,N_9353);
xor UO_1363 (O_1363,N_9954,N_8881);
nand UO_1364 (O_1364,N_9121,N_9114);
nor UO_1365 (O_1365,N_8565,N_9434);
and UO_1366 (O_1366,N_8636,N_7613);
and UO_1367 (O_1367,N_8535,N_9654);
or UO_1368 (O_1368,N_8022,N_7702);
or UO_1369 (O_1369,N_8472,N_9880);
or UO_1370 (O_1370,N_9525,N_9273);
nand UO_1371 (O_1371,N_9771,N_9976);
and UO_1372 (O_1372,N_8830,N_9023);
and UO_1373 (O_1373,N_8521,N_7754);
nand UO_1374 (O_1374,N_9751,N_8697);
nor UO_1375 (O_1375,N_8694,N_9984);
nand UO_1376 (O_1376,N_9469,N_7945);
and UO_1377 (O_1377,N_8992,N_9923);
or UO_1378 (O_1378,N_8035,N_9316);
nand UO_1379 (O_1379,N_9146,N_8683);
nor UO_1380 (O_1380,N_9601,N_8029);
xor UO_1381 (O_1381,N_9209,N_9570);
xor UO_1382 (O_1382,N_8181,N_9379);
and UO_1383 (O_1383,N_9010,N_8830);
and UO_1384 (O_1384,N_8020,N_7897);
nand UO_1385 (O_1385,N_8357,N_8136);
nand UO_1386 (O_1386,N_9553,N_8429);
and UO_1387 (O_1387,N_7668,N_9949);
or UO_1388 (O_1388,N_7714,N_7835);
or UO_1389 (O_1389,N_8984,N_9644);
nand UO_1390 (O_1390,N_8920,N_9501);
or UO_1391 (O_1391,N_8119,N_8888);
or UO_1392 (O_1392,N_9501,N_7812);
nor UO_1393 (O_1393,N_9118,N_9960);
nand UO_1394 (O_1394,N_9883,N_8691);
and UO_1395 (O_1395,N_9889,N_9739);
or UO_1396 (O_1396,N_9007,N_9264);
nand UO_1397 (O_1397,N_8450,N_8151);
nor UO_1398 (O_1398,N_9514,N_8786);
nand UO_1399 (O_1399,N_9842,N_8635);
nand UO_1400 (O_1400,N_8443,N_9512);
and UO_1401 (O_1401,N_9796,N_8411);
xnor UO_1402 (O_1402,N_9814,N_7556);
nand UO_1403 (O_1403,N_9055,N_8287);
or UO_1404 (O_1404,N_9245,N_8276);
or UO_1405 (O_1405,N_9963,N_9063);
nand UO_1406 (O_1406,N_9936,N_9871);
nand UO_1407 (O_1407,N_9054,N_7549);
and UO_1408 (O_1408,N_9908,N_8262);
xor UO_1409 (O_1409,N_8150,N_9876);
nor UO_1410 (O_1410,N_8021,N_9424);
and UO_1411 (O_1411,N_9355,N_7575);
or UO_1412 (O_1412,N_8180,N_8843);
or UO_1413 (O_1413,N_8517,N_8966);
or UO_1414 (O_1414,N_9917,N_8700);
or UO_1415 (O_1415,N_9149,N_8452);
nor UO_1416 (O_1416,N_9608,N_9969);
nor UO_1417 (O_1417,N_9776,N_8256);
or UO_1418 (O_1418,N_8904,N_7653);
nor UO_1419 (O_1419,N_9345,N_8909);
xor UO_1420 (O_1420,N_9836,N_8632);
and UO_1421 (O_1421,N_9315,N_8862);
nor UO_1422 (O_1422,N_8771,N_8870);
and UO_1423 (O_1423,N_8636,N_9463);
and UO_1424 (O_1424,N_8755,N_9310);
nor UO_1425 (O_1425,N_9140,N_9713);
nor UO_1426 (O_1426,N_8803,N_8829);
and UO_1427 (O_1427,N_7954,N_7635);
nor UO_1428 (O_1428,N_7552,N_7677);
or UO_1429 (O_1429,N_8104,N_8106);
and UO_1430 (O_1430,N_7578,N_9195);
nand UO_1431 (O_1431,N_9317,N_9419);
or UO_1432 (O_1432,N_8743,N_9054);
or UO_1433 (O_1433,N_8320,N_8489);
and UO_1434 (O_1434,N_9602,N_8652);
or UO_1435 (O_1435,N_9537,N_8676);
nand UO_1436 (O_1436,N_8000,N_9869);
nand UO_1437 (O_1437,N_8116,N_9603);
and UO_1438 (O_1438,N_8997,N_8051);
nand UO_1439 (O_1439,N_9671,N_7822);
nand UO_1440 (O_1440,N_9364,N_8671);
and UO_1441 (O_1441,N_8112,N_9807);
or UO_1442 (O_1442,N_7634,N_9869);
nor UO_1443 (O_1443,N_7716,N_9872);
nor UO_1444 (O_1444,N_8502,N_7667);
xor UO_1445 (O_1445,N_9433,N_8717);
xor UO_1446 (O_1446,N_9557,N_8140);
nor UO_1447 (O_1447,N_9015,N_9922);
nor UO_1448 (O_1448,N_8761,N_9995);
nand UO_1449 (O_1449,N_8627,N_8480);
nand UO_1450 (O_1450,N_8831,N_8357);
nor UO_1451 (O_1451,N_8064,N_9149);
and UO_1452 (O_1452,N_8833,N_7974);
nand UO_1453 (O_1453,N_9394,N_9734);
nand UO_1454 (O_1454,N_7646,N_7858);
nor UO_1455 (O_1455,N_9031,N_7732);
nor UO_1456 (O_1456,N_7943,N_9067);
or UO_1457 (O_1457,N_8819,N_9672);
nand UO_1458 (O_1458,N_9412,N_7895);
xnor UO_1459 (O_1459,N_8610,N_9022);
nand UO_1460 (O_1460,N_9968,N_9092);
or UO_1461 (O_1461,N_9755,N_8780);
xor UO_1462 (O_1462,N_9468,N_9810);
and UO_1463 (O_1463,N_7691,N_9481);
and UO_1464 (O_1464,N_8572,N_9338);
or UO_1465 (O_1465,N_9954,N_8765);
nor UO_1466 (O_1466,N_8637,N_9811);
xnor UO_1467 (O_1467,N_9172,N_8750);
and UO_1468 (O_1468,N_7810,N_7709);
nand UO_1469 (O_1469,N_9409,N_9633);
or UO_1470 (O_1470,N_8173,N_7669);
or UO_1471 (O_1471,N_8138,N_9005);
nor UO_1472 (O_1472,N_7610,N_8573);
nand UO_1473 (O_1473,N_8744,N_7706);
or UO_1474 (O_1474,N_8576,N_7561);
or UO_1475 (O_1475,N_8200,N_9716);
and UO_1476 (O_1476,N_8142,N_9902);
and UO_1477 (O_1477,N_9757,N_9138);
nor UO_1478 (O_1478,N_9778,N_9197);
and UO_1479 (O_1479,N_7558,N_9142);
nand UO_1480 (O_1480,N_9893,N_7944);
nand UO_1481 (O_1481,N_9901,N_9266);
or UO_1482 (O_1482,N_9640,N_8992);
or UO_1483 (O_1483,N_8727,N_9729);
and UO_1484 (O_1484,N_8508,N_8678);
nand UO_1485 (O_1485,N_8518,N_9478);
nand UO_1486 (O_1486,N_7547,N_8712);
and UO_1487 (O_1487,N_9091,N_9252);
nand UO_1488 (O_1488,N_9858,N_8365);
nand UO_1489 (O_1489,N_9076,N_9155);
nand UO_1490 (O_1490,N_7960,N_8243);
nand UO_1491 (O_1491,N_8532,N_8386);
and UO_1492 (O_1492,N_9342,N_7822);
or UO_1493 (O_1493,N_9439,N_8819);
xor UO_1494 (O_1494,N_9818,N_9263);
nor UO_1495 (O_1495,N_7720,N_8020);
or UO_1496 (O_1496,N_9241,N_8603);
nor UO_1497 (O_1497,N_8904,N_7766);
nor UO_1498 (O_1498,N_8922,N_7889);
nor UO_1499 (O_1499,N_9477,N_9289);
endmodule