module basic_500_3000_500_3_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_482,In_322);
xnor U1 (N_1,In_391,In_433);
nor U2 (N_2,In_270,In_308);
nor U3 (N_3,In_455,In_244);
and U4 (N_4,In_379,In_128);
nand U5 (N_5,In_3,In_36);
nand U6 (N_6,In_269,In_30);
nor U7 (N_7,In_319,In_441);
nor U8 (N_8,In_69,In_54);
nor U9 (N_9,In_486,In_43);
nand U10 (N_10,In_144,In_227);
and U11 (N_11,In_68,In_323);
or U12 (N_12,In_428,In_293);
and U13 (N_13,In_337,In_204);
or U14 (N_14,In_496,In_449);
or U15 (N_15,In_38,In_429);
xor U16 (N_16,In_76,In_414);
and U17 (N_17,In_468,In_422);
nand U18 (N_18,In_45,In_330);
nor U19 (N_19,In_488,In_56);
nor U20 (N_20,In_116,In_312);
nand U21 (N_21,In_368,In_487);
nand U22 (N_22,In_230,In_196);
or U23 (N_23,In_29,In_396);
or U24 (N_24,In_154,In_62);
nor U25 (N_25,In_387,In_370);
or U26 (N_26,In_303,In_124);
or U27 (N_27,In_137,In_106);
nand U28 (N_28,In_127,In_341);
nor U29 (N_29,In_434,In_181);
or U30 (N_30,In_232,In_363);
and U31 (N_31,In_9,In_286);
and U32 (N_32,In_499,In_267);
nand U33 (N_33,In_7,In_409);
nand U34 (N_34,In_194,In_346);
nor U35 (N_35,In_132,In_453);
or U36 (N_36,In_444,In_343);
nor U37 (N_37,In_167,In_281);
or U38 (N_38,In_225,In_413);
and U39 (N_39,In_313,In_222);
and U40 (N_40,In_81,In_331);
xor U41 (N_41,In_259,In_411);
and U42 (N_42,In_140,In_390);
nand U43 (N_43,In_431,In_284);
and U44 (N_44,In_419,In_205);
xor U45 (N_45,In_220,In_34);
nor U46 (N_46,In_41,In_288);
or U47 (N_47,In_383,In_478);
and U48 (N_48,In_130,In_394);
and U49 (N_49,In_171,In_160);
xor U50 (N_50,In_299,In_82);
or U51 (N_51,In_406,In_125);
xnor U52 (N_52,In_493,In_275);
and U53 (N_53,In_242,In_374);
xnor U54 (N_54,In_161,In_283);
xnor U55 (N_55,In_276,In_64);
nor U56 (N_56,In_102,In_121);
nor U57 (N_57,In_479,In_287);
nand U58 (N_58,In_297,In_342);
or U59 (N_59,In_321,In_329);
nand U60 (N_60,In_377,In_19);
or U61 (N_61,In_345,In_354);
xnor U62 (N_62,In_21,In_178);
or U63 (N_63,In_129,In_233);
and U64 (N_64,In_101,In_265);
nand U65 (N_65,In_192,In_358);
nand U66 (N_66,In_97,In_136);
nand U67 (N_67,In_2,In_268);
nor U68 (N_68,In_122,In_236);
and U69 (N_69,In_96,In_350);
nor U70 (N_70,In_6,In_445);
or U71 (N_71,In_469,In_235);
and U72 (N_72,In_89,In_498);
nand U73 (N_73,In_495,In_214);
nor U74 (N_74,In_381,In_364);
and U75 (N_75,In_91,In_494);
nand U76 (N_76,In_70,In_53);
and U77 (N_77,In_65,In_114);
or U78 (N_78,In_367,In_172);
nor U79 (N_79,In_474,In_271);
nor U80 (N_80,In_351,In_485);
nor U81 (N_81,In_17,In_376);
and U82 (N_82,In_423,In_247);
nor U83 (N_83,In_158,In_75);
nor U84 (N_84,In_209,In_246);
nand U85 (N_85,In_272,In_111);
nor U86 (N_86,In_292,In_382);
xor U87 (N_87,In_46,In_371);
and U88 (N_88,In_256,In_52);
and U89 (N_89,In_226,In_15);
or U90 (N_90,In_476,In_177);
and U91 (N_91,In_88,In_249);
and U92 (N_92,In_285,In_145);
xor U93 (N_93,In_25,In_85);
or U94 (N_94,In_440,In_59);
or U95 (N_95,In_380,In_176);
xor U96 (N_96,In_173,In_179);
or U97 (N_97,In_55,In_94);
or U98 (N_98,In_13,In_8);
or U99 (N_99,In_170,In_373);
nor U100 (N_100,In_12,In_245);
nor U101 (N_101,In_67,In_400);
xnor U102 (N_102,In_415,In_378);
or U103 (N_103,In_120,In_134);
and U104 (N_104,In_456,In_118);
and U105 (N_105,In_186,In_426);
and U106 (N_106,In_32,In_325);
and U107 (N_107,In_10,In_483);
and U108 (N_108,In_99,In_250);
or U109 (N_109,In_159,In_105);
nor U110 (N_110,In_165,In_490);
xnor U111 (N_111,In_335,In_141);
nor U112 (N_112,In_215,In_31);
nor U113 (N_113,In_78,In_131);
and U114 (N_114,In_182,In_115);
nand U115 (N_115,In_255,In_221);
nor U116 (N_116,In_307,In_188);
nor U117 (N_117,In_277,In_344);
nor U118 (N_118,In_135,In_403);
or U119 (N_119,In_309,In_274);
nand U120 (N_120,In_138,In_44);
nor U121 (N_121,In_163,In_149);
and U122 (N_122,In_318,In_466);
nor U123 (N_123,In_86,In_16);
or U124 (N_124,In_266,In_39);
or U125 (N_125,In_446,In_336);
nor U126 (N_126,In_458,In_326);
and U127 (N_127,In_107,In_48);
nor U128 (N_128,In_295,In_80);
nor U129 (N_129,In_454,In_35);
and U130 (N_130,In_180,In_332);
and U131 (N_131,In_185,In_470);
or U132 (N_132,In_305,In_50);
nand U133 (N_133,In_310,In_27);
and U134 (N_134,In_234,In_407);
or U135 (N_135,In_430,In_304);
or U136 (N_136,In_388,In_448);
and U137 (N_137,In_229,In_366);
and U138 (N_138,In_110,In_328);
and U139 (N_139,In_484,In_42);
and U140 (N_140,In_334,In_216);
nor U141 (N_141,In_477,In_14);
or U142 (N_142,In_0,In_262);
and U143 (N_143,In_77,In_280);
nor U144 (N_144,In_23,In_211);
or U145 (N_145,In_210,In_393);
nand U146 (N_146,In_100,In_156);
nor U147 (N_147,In_147,In_218);
nand U148 (N_148,In_207,In_253);
nor U149 (N_149,In_324,In_20);
and U150 (N_150,In_489,In_152);
xor U151 (N_151,In_195,In_40);
nand U152 (N_152,In_260,In_93);
nor U153 (N_153,In_392,In_347);
nand U154 (N_154,In_162,In_384);
and U155 (N_155,In_133,In_389);
nor U156 (N_156,In_98,In_47);
nor U157 (N_157,In_150,In_404);
or U158 (N_158,In_333,In_432);
or U159 (N_159,In_74,In_164);
nand U160 (N_160,In_1,In_103);
or U161 (N_161,In_237,In_224);
nor U162 (N_162,In_278,In_157);
nor U163 (N_163,In_240,In_475);
xnor U164 (N_164,In_294,In_258);
nor U165 (N_165,In_357,In_208);
or U166 (N_166,In_349,In_356);
and U167 (N_167,In_264,In_375);
and U168 (N_168,In_187,In_372);
nand U169 (N_169,In_348,In_200);
and U170 (N_170,In_11,In_459);
nand U171 (N_171,In_241,In_203);
nand U172 (N_172,In_340,In_213);
xnor U173 (N_173,In_184,In_320);
nor U174 (N_174,In_28,In_83);
or U175 (N_175,In_123,In_315);
xnor U176 (N_176,In_51,In_175);
nand U177 (N_177,In_442,In_497);
and U178 (N_178,In_155,In_327);
xnor U179 (N_179,In_362,In_438);
and U180 (N_180,In_174,In_104);
or U181 (N_181,In_61,In_261);
and U182 (N_182,In_359,In_311);
or U183 (N_183,In_316,In_228);
or U184 (N_184,In_151,In_231);
xnor U185 (N_185,In_212,In_143);
xnor U186 (N_186,In_18,In_464);
or U187 (N_187,In_84,In_153);
and U188 (N_188,In_416,In_338);
nand U189 (N_189,In_168,In_339);
or U190 (N_190,In_113,In_399);
nor U191 (N_191,In_169,In_425);
and U192 (N_192,In_71,In_427);
or U193 (N_193,In_451,In_37);
or U194 (N_194,In_139,In_24);
nand U195 (N_195,In_95,In_360);
and U196 (N_196,In_206,In_443);
xnor U197 (N_197,In_398,In_298);
xnor U198 (N_198,In_296,In_257);
and U199 (N_199,In_421,In_462);
or U200 (N_200,In_290,In_420);
nor U201 (N_201,In_273,In_217);
or U202 (N_202,In_439,In_219);
or U203 (N_203,In_435,In_243);
nor U204 (N_204,In_4,In_263);
and U205 (N_205,In_418,In_405);
nor U206 (N_206,In_199,In_457);
nand U207 (N_207,In_119,In_291);
and U208 (N_208,In_467,In_190);
nor U209 (N_209,In_481,In_386);
nor U210 (N_210,In_412,In_279);
and U211 (N_211,In_26,In_142);
nand U212 (N_212,In_146,In_395);
or U213 (N_213,In_417,In_452);
and U214 (N_214,In_5,In_166);
nand U215 (N_215,In_126,In_66);
or U216 (N_216,In_189,In_22);
or U217 (N_217,In_251,In_197);
nand U218 (N_218,In_397,In_385);
and U219 (N_219,In_437,In_480);
nor U220 (N_220,In_108,In_90);
or U221 (N_221,In_58,In_73);
nor U222 (N_222,In_289,In_408);
and U223 (N_223,In_463,In_369);
and U224 (N_224,In_239,In_447);
xnor U225 (N_225,In_148,In_60);
nand U226 (N_226,In_79,In_223);
and U227 (N_227,In_353,In_202);
and U228 (N_228,In_401,In_492);
nor U229 (N_229,In_450,In_87);
nor U230 (N_230,In_352,In_117);
nand U231 (N_231,In_473,In_201);
or U232 (N_232,In_57,In_254);
nor U233 (N_233,In_461,In_300);
or U234 (N_234,In_306,In_365);
nor U235 (N_235,In_191,In_282);
or U236 (N_236,In_355,In_402);
or U237 (N_237,In_460,In_112);
nor U238 (N_238,In_193,In_472);
nand U239 (N_239,In_33,In_301);
or U240 (N_240,In_471,In_198);
nand U241 (N_241,In_317,In_252);
nand U242 (N_242,In_424,In_465);
or U243 (N_243,In_314,In_248);
nand U244 (N_244,In_361,In_49);
and U245 (N_245,In_410,In_491);
or U246 (N_246,In_92,In_238);
nor U247 (N_247,In_302,In_183);
nor U248 (N_248,In_109,In_72);
nor U249 (N_249,In_436,In_63);
or U250 (N_250,In_305,In_234);
xor U251 (N_251,In_496,In_413);
xor U252 (N_252,In_25,In_417);
nor U253 (N_253,In_246,In_9);
and U254 (N_254,In_322,In_479);
nor U255 (N_255,In_67,In_488);
and U256 (N_256,In_298,In_337);
nand U257 (N_257,In_282,In_459);
nor U258 (N_258,In_112,In_75);
xor U259 (N_259,In_3,In_294);
nor U260 (N_260,In_55,In_105);
nor U261 (N_261,In_360,In_10);
or U262 (N_262,In_467,In_441);
nor U263 (N_263,In_206,In_6);
xor U264 (N_264,In_190,In_9);
nor U265 (N_265,In_249,In_480);
or U266 (N_266,In_483,In_80);
nand U267 (N_267,In_299,In_197);
nand U268 (N_268,In_128,In_37);
nand U269 (N_269,In_306,In_477);
nor U270 (N_270,In_285,In_387);
and U271 (N_271,In_353,In_118);
or U272 (N_272,In_116,In_250);
or U273 (N_273,In_454,In_7);
or U274 (N_274,In_303,In_268);
or U275 (N_275,In_296,In_181);
nand U276 (N_276,In_258,In_301);
nor U277 (N_277,In_464,In_306);
nand U278 (N_278,In_56,In_175);
and U279 (N_279,In_382,In_495);
nand U280 (N_280,In_463,In_118);
and U281 (N_281,In_368,In_451);
nand U282 (N_282,In_112,In_252);
or U283 (N_283,In_26,In_240);
or U284 (N_284,In_472,In_458);
nand U285 (N_285,In_391,In_299);
nand U286 (N_286,In_69,In_182);
or U287 (N_287,In_241,In_11);
or U288 (N_288,In_175,In_359);
or U289 (N_289,In_79,In_291);
nand U290 (N_290,In_49,In_225);
or U291 (N_291,In_125,In_35);
nand U292 (N_292,In_125,In_374);
nand U293 (N_293,In_380,In_1);
or U294 (N_294,In_359,In_229);
nand U295 (N_295,In_283,In_357);
nand U296 (N_296,In_302,In_106);
and U297 (N_297,In_481,In_252);
and U298 (N_298,In_98,In_330);
nand U299 (N_299,In_387,In_348);
or U300 (N_300,In_66,In_499);
or U301 (N_301,In_72,In_341);
and U302 (N_302,In_390,In_289);
nor U303 (N_303,In_496,In_300);
nor U304 (N_304,In_312,In_381);
and U305 (N_305,In_103,In_33);
and U306 (N_306,In_208,In_11);
xor U307 (N_307,In_74,In_115);
and U308 (N_308,In_301,In_216);
and U309 (N_309,In_330,In_166);
or U310 (N_310,In_195,In_429);
and U311 (N_311,In_158,In_396);
nand U312 (N_312,In_463,In_149);
and U313 (N_313,In_381,In_165);
and U314 (N_314,In_396,In_225);
nor U315 (N_315,In_425,In_345);
or U316 (N_316,In_364,In_369);
and U317 (N_317,In_432,In_67);
nor U318 (N_318,In_438,In_397);
or U319 (N_319,In_3,In_134);
nand U320 (N_320,In_186,In_158);
and U321 (N_321,In_238,In_461);
xnor U322 (N_322,In_223,In_46);
and U323 (N_323,In_192,In_10);
or U324 (N_324,In_237,In_453);
nor U325 (N_325,In_349,In_116);
or U326 (N_326,In_22,In_324);
and U327 (N_327,In_423,In_360);
xnor U328 (N_328,In_208,In_79);
and U329 (N_329,In_71,In_247);
xor U330 (N_330,In_291,In_257);
or U331 (N_331,In_133,In_469);
nand U332 (N_332,In_406,In_34);
nor U333 (N_333,In_115,In_54);
or U334 (N_334,In_101,In_102);
nand U335 (N_335,In_343,In_451);
nor U336 (N_336,In_318,In_379);
and U337 (N_337,In_167,In_65);
xor U338 (N_338,In_490,In_422);
xnor U339 (N_339,In_225,In_183);
or U340 (N_340,In_418,In_381);
and U341 (N_341,In_429,In_422);
nor U342 (N_342,In_432,In_248);
nand U343 (N_343,In_109,In_342);
nor U344 (N_344,In_153,In_498);
or U345 (N_345,In_128,In_287);
nand U346 (N_346,In_396,In_116);
or U347 (N_347,In_78,In_199);
nor U348 (N_348,In_487,In_335);
or U349 (N_349,In_319,In_265);
nor U350 (N_350,In_496,In_141);
nand U351 (N_351,In_71,In_273);
or U352 (N_352,In_242,In_260);
nor U353 (N_353,In_248,In_72);
nor U354 (N_354,In_189,In_7);
or U355 (N_355,In_430,In_241);
and U356 (N_356,In_231,In_311);
xnor U357 (N_357,In_411,In_401);
nand U358 (N_358,In_110,In_364);
and U359 (N_359,In_153,In_130);
nor U360 (N_360,In_31,In_297);
and U361 (N_361,In_413,In_113);
and U362 (N_362,In_216,In_328);
xnor U363 (N_363,In_124,In_54);
nand U364 (N_364,In_343,In_280);
nand U365 (N_365,In_383,In_261);
nand U366 (N_366,In_87,In_100);
and U367 (N_367,In_151,In_49);
nor U368 (N_368,In_327,In_260);
nor U369 (N_369,In_402,In_124);
nor U370 (N_370,In_187,In_184);
xor U371 (N_371,In_295,In_56);
nor U372 (N_372,In_275,In_44);
nor U373 (N_373,In_210,In_300);
xnor U374 (N_374,In_104,In_444);
xor U375 (N_375,In_203,In_458);
nand U376 (N_376,In_137,In_71);
nor U377 (N_377,In_150,In_173);
nor U378 (N_378,In_14,In_90);
nand U379 (N_379,In_329,In_278);
and U380 (N_380,In_299,In_320);
nand U381 (N_381,In_57,In_458);
and U382 (N_382,In_121,In_460);
xnor U383 (N_383,In_467,In_397);
nor U384 (N_384,In_155,In_415);
nand U385 (N_385,In_338,In_110);
and U386 (N_386,In_458,In_395);
nand U387 (N_387,In_303,In_279);
and U388 (N_388,In_344,In_215);
nand U389 (N_389,In_190,In_455);
nand U390 (N_390,In_416,In_126);
and U391 (N_391,In_249,In_276);
nand U392 (N_392,In_202,In_22);
and U393 (N_393,In_100,In_348);
nand U394 (N_394,In_487,In_333);
nand U395 (N_395,In_305,In_382);
nor U396 (N_396,In_231,In_30);
nor U397 (N_397,In_117,In_386);
nor U398 (N_398,In_237,In_219);
or U399 (N_399,In_47,In_458);
nand U400 (N_400,In_79,In_230);
or U401 (N_401,In_211,In_310);
nor U402 (N_402,In_377,In_463);
nand U403 (N_403,In_297,In_204);
or U404 (N_404,In_7,In_268);
nand U405 (N_405,In_453,In_126);
xor U406 (N_406,In_148,In_175);
nand U407 (N_407,In_284,In_238);
or U408 (N_408,In_384,In_436);
or U409 (N_409,In_250,In_405);
nor U410 (N_410,In_320,In_420);
or U411 (N_411,In_261,In_301);
nand U412 (N_412,In_112,In_435);
xnor U413 (N_413,In_225,In_419);
xor U414 (N_414,In_319,In_12);
or U415 (N_415,In_470,In_74);
or U416 (N_416,In_293,In_452);
nor U417 (N_417,In_0,In_104);
or U418 (N_418,In_346,In_273);
nand U419 (N_419,In_368,In_342);
nor U420 (N_420,In_400,In_91);
nor U421 (N_421,In_389,In_61);
nor U422 (N_422,In_281,In_464);
nand U423 (N_423,In_113,In_129);
and U424 (N_424,In_445,In_66);
nand U425 (N_425,In_424,In_447);
and U426 (N_426,In_127,In_24);
nor U427 (N_427,In_240,In_495);
and U428 (N_428,In_185,In_210);
nor U429 (N_429,In_491,In_129);
or U430 (N_430,In_424,In_287);
nor U431 (N_431,In_113,In_317);
and U432 (N_432,In_145,In_142);
nor U433 (N_433,In_325,In_75);
or U434 (N_434,In_205,In_61);
or U435 (N_435,In_17,In_433);
or U436 (N_436,In_479,In_68);
and U437 (N_437,In_71,In_167);
or U438 (N_438,In_28,In_123);
nand U439 (N_439,In_273,In_35);
nand U440 (N_440,In_267,In_182);
or U441 (N_441,In_477,In_116);
and U442 (N_442,In_458,In_11);
nor U443 (N_443,In_33,In_53);
or U444 (N_444,In_125,In_386);
xnor U445 (N_445,In_116,In_102);
or U446 (N_446,In_399,In_218);
nand U447 (N_447,In_406,In_463);
or U448 (N_448,In_30,In_246);
nor U449 (N_449,In_439,In_316);
nor U450 (N_450,In_194,In_217);
nand U451 (N_451,In_212,In_146);
xor U452 (N_452,In_264,In_311);
or U453 (N_453,In_234,In_327);
or U454 (N_454,In_283,In_355);
and U455 (N_455,In_146,In_206);
and U456 (N_456,In_463,In_471);
nand U457 (N_457,In_160,In_465);
nand U458 (N_458,In_326,In_399);
nor U459 (N_459,In_267,In_458);
xor U460 (N_460,In_452,In_153);
nor U461 (N_461,In_319,In_399);
and U462 (N_462,In_134,In_79);
nor U463 (N_463,In_453,In_479);
or U464 (N_464,In_160,In_486);
or U465 (N_465,In_328,In_26);
nor U466 (N_466,In_382,In_214);
and U467 (N_467,In_331,In_268);
nand U468 (N_468,In_298,In_49);
xnor U469 (N_469,In_314,In_189);
and U470 (N_470,In_418,In_219);
nor U471 (N_471,In_76,In_243);
nand U472 (N_472,In_385,In_84);
xor U473 (N_473,In_338,In_42);
nand U474 (N_474,In_428,In_47);
nand U475 (N_475,In_454,In_345);
or U476 (N_476,In_40,In_34);
nand U477 (N_477,In_412,In_106);
nor U478 (N_478,In_310,In_147);
or U479 (N_479,In_410,In_479);
or U480 (N_480,In_475,In_235);
or U481 (N_481,In_409,In_146);
and U482 (N_482,In_287,In_1);
nor U483 (N_483,In_293,In_150);
xor U484 (N_484,In_393,In_465);
and U485 (N_485,In_197,In_379);
nor U486 (N_486,In_331,In_380);
or U487 (N_487,In_188,In_409);
nor U488 (N_488,In_212,In_157);
or U489 (N_489,In_110,In_70);
and U490 (N_490,In_53,In_310);
nand U491 (N_491,In_449,In_195);
xor U492 (N_492,In_6,In_355);
or U493 (N_493,In_83,In_498);
nand U494 (N_494,In_17,In_115);
xnor U495 (N_495,In_164,In_413);
nand U496 (N_496,In_156,In_427);
nand U497 (N_497,In_471,In_174);
xor U498 (N_498,In_117,In_324);
nor U499 (N_499,In_346,In_467);
xor U500 (N_500,In_368,In_416);
and U501 (N_501,In_116,In_373);
nor U502 (N_502,In_325,In_226);
nor U503 (N_503,In_108,In_109);
nor U504 (N_504,In_438,In_196);
or U505 (N_505,In_184,In_86);
nor U506 (N_506,In_311,In_219);
and U507 (N_507,In_128,In_423);
nand U508 (N_508,In_55,In_421);
nand U509 (N_509,In_203,In_476);
nand U510 (N_510,In_6,In_40);
nand U511 (N_511,In_390,In_93);
nor U512 (N_512,In_289,In_345);
nor U513 (N_513,In_94,In_454);
nor U514 (N_514,In_98,In_261);
nor U515 (N_515,In_275,In_137);
nor U516 (N_516,In_168,In_226);
or U517 (N_517,In_347,In_274);
and U518 (N_518,In_89,In_339);
nand U519 (N_519,In_213,In_221);
or U520 (N_520,In_476,In_88);
and U521 (N_521,In_268,In_81);
and U522 (N_522,In_160,In_323);
and U523 (N_523,In_447,In_33);
nand U524 (N_524,In_451,In_41);
nor U525 (N_525,In_123,In_417);
or U526 (N_526,In_479,In_84);
and U527 (N_527,In_162,In_222);
nand U528 (N_528,In_246,In_459);
or U529 (N_529,In_127,In_197);
nand U530 (N_530,In_148,In_56);
or U531 (N_531,In_211,In_285);
nor U532 (N_532,In_261,In_156);
nand U533 (N_533,In_153,In_289);
nor U534 (N_534,In_200,In_103);
nor U535 (N_535,In_443,In_490);
or U536 (N_536,In_114,In_103);
and U537 (N_537,In_226,In_83);
or U538 (N_538,In_367,In_345);
nand U539 (N_539,In_72,In_169);
nor U540 (N_540,In_350,In_272);
and U541 (N_541,In_413,In_224);
nand U542 (N_542,In_70,In_327);
nor U543 (N_543,In_431,In_127);
or U544 (N_544,In_81,In_447);
and U545 (N_545,In_159,In_289);
and U546 (N_546,In_348,In_332);
and U547 (N_547,In_398,In_345);
nand U548 (N_548,In_266,In_381);
xnor U549 (N_549,In_6,In_491);
nand U550 (N_550,In_92,In_445);
nor U551 (N_551,In_390,In_251);
nand U552 (N_552,In_118,In_268);
nand U553 (N_553,In_297,In_7);
and U554 (N_554,In_97,In_138);
nand U555 (N_555,In_56,In_293);
nand U556 (N_556,In_206,In_357);
and U557 (N_557,In_257,In_134);
nor U558 (N_558,In_171,In_486);
xnor U559 (N_559,In_244,In_95);
and U560 (N_560,In_437,In_335);
nand U561 (N_561,In_416,In_59);
and U562 (N_562,In_416,In_10);
nand U563 (N_563,In_88,In_108);
nor U564 (N_564,In_251,In_367);
nand U565 (N_565,In_340,In_453);
or U566 (N_566,In_374,In_348);
and U567 (N_567,In_380,In_463);
or U568 (N_568,In_203,In_99);
xnor U569 (N_569,In_489,In_415);
nor U570 (N_570,In_303,In_460);
and U571 (N_571,In_327,In_298);
nor U572 (N_572,In_142,In_224);
nor U573 (N_573,In_38,In_341);
nor U574 (N_574,In_25,In_92);
nor U575 (N_575,In_369,In_423);
nand U576 (N_576,In_468,In_486);
nand U577 (N_577,In_40,In_332);
nand U578 (N_578,In_37,In_199);
nor U579 (N_579,In_166,In_223);
nand U580 (N_580,In_79,In_59);
nand U581 (N_581,In_199,In_287);
nand U582 (N_582,In_361,In_65);
and U583 (N_583,In_240,In_258);
nor U584 (N_584,In_153,In_134);
or U585 (N_585,In_478,In_494);
nand U586 (N_586,In_209,In_249);
nand U587 (N_587,In_466,In_311);
nand U588 (N_588,In_350,In_415);
nor U589 (N_589,In_466,In_373);
or U590 (N_590,In_222,In_229);
nor U591 (N_591,In_440,In_88);
nor U592 (N_592,In_116,In_333);
nor U593 (N_593,In_148,In_38);
and U594 (N_594,In_468,In_392);
xor U595 (N_595,In_324,In_212);
nand U596 (N_596,In_230,In_227);
nand U597 (N_597,In_340,In_228);
or U598 (N_598,In_160,In_467);
or U599 (N_599,In_317,In_271);
nand U600 (N_600,In_184,In_348);
nand U601 (N_601,In_394,In_335);
or U602 (N_602,In_32,In_451);
xor U603 (N_603,In_190,In_369);
xnor U604 (N_604,In_447,In_71);
nand U605 (N_605,In_480,In_347);
or U606 (N_606,In_135,In_487);
nand U607 (N_607,In_295,In_189);
nand U608 (N_608,In_297,In_349);
and U609 (N_609,In_344,In_191);
xor U610 (N_610,In_332,In_387);
xnor U611 (N_611,In_407,In_428);
nand U612 (N_612,In_408,In_175);
and U613 (N_613,In_406,In_83);
and U614 (N_614,In_85,In_437);
nor U615 (N_615,In_464,In_3);
and U616 (N_616,In_234,In_337);
nand U617 (N_617,In_115,In_53);
and U618 (N_618,In_269,In_339);
or U619 (N_619,In_74,In_403);
and U620 (N_620,In_291,In_208);
nand U621 (N_621,In_306,In_41);
and U622 (N_622,In_391,In_105);
or U623 (N_623,In_270,In_173);
nand U624 (N_624,In_211,In_239);
nand U625 (N_625,In_444,In_143);
and U626 (N_626,In_178,In_405);
nor U627 (N_627,In_166,In_266);
nand U628 (N_628,In_112,In_111);
or U629 (N_629,In_302,In_346);
nor U630 (N_630,In_88,In_152);
or U631 (N_631,In_200,In_183);
or U632 (N_632,In_436,In_139);
and U633 (N_633,In_261,In_3);
xor U634 (N_634,In_303,In_221);
and U635 (N_635,In_298,In_308);
or U636 (N_636,In_101,In_32);
nand U637 (N_637,In_367,In_3);
nand U638 (N_638,In_279,In_409);
or U639 (N_639,In_274,In_398);
nor U640 (N_640,In_292,In_162);
nor U641 (N_641,In_203,In_186);
xor U642 (N_642,In_462,In_186);
nand U643 (N_643,In_267,In_200);
and U644 (N_644,In_411,In_367);
and U645 (N_645,In_428,In_247);
and U646 (N_646,In_425,In_295);
nor U647 (N_647,In_379,In_395);
or U648 (N_648,In_72,In_269);
nand U649 (N_649,In_262,In_421);
xnor U650 (N_650,In_413,In_182);
nor U651 (N_651,In_236,In_244);
or U652 (N_652,In_287,In_385);
and U653 (N_653,In_351,In_425);
and U654 (N_654,In_389,In_39);
xnor U655 (N_655,In_297,In_254);
xnor U656 (N_656,In_280,In_335);
nor U657 (N_657,In_166,In_226);
nand U658 (N_658,In_289,In_88);
or U659 (N_659,In_459,In_325);
or U660 (N_660,In_252,In_417);
nand U661 (N_661,In_96,In_326);
and U662 (N_662,In_7,In_462);
nor U663 (N_663,In_415,In_209);
nand U664 (N_664,In_349,In_319);
and U665 (N_665,In_14,In_492);
and U666 (N_666,In_49,In_253);
xnor U667 (N_667,In_189,In_161);
nand U668 (N_668,In_311,In_33);
nor U669 (N_669,In_135,In_161);
and U670 (N_670,In_70,In_324);
or U671 (N_671,In_389,In_120);
and U672 (N_672,In_258,In_71);
nand U673 (N_673,In_152,In_405);
xor U674 (N_674,In_1,In_46);
nor U675 (N_675,In_466,In_209);
or U676 (N_676,In_114,In_158);
nor U677 (N_677,In_20,In_11);
nand U678 (N_678,In_53,In_119);
and U679 (N_679,In_82,In_192);
nand U680 (N_680,In_393,In_226);
or U681 (N_681,In_273,In_423);
or U682 (N_682,In_132,In_121);
nor U683 (N_683,In_318,In_463);
nor U684 (N_684,In_422,In_228);
or U685 (N_685,In_64,In_82);
nor U686 (N_686,In_61,In_315);
xor U687 (N_687,In_63,In_454);
or U688 (N_688,In_338,In_263);
nor U689 (N_689,In_382,In_294);
nor U690 (N_690,In_419,In_401);
or U691 (N_691,In_449,In_198);
nand U692 (N_692,In_463,In_465);
and U693 (N_693,In_84,In_43);
and U694 (N_694,In_466,In_230);
and U695 (N_695,In_110,In_138);
and U696 (N_696,In_307,In_413);
nor U697 (N_697,In_31,In_16);
xor U698 (N_698,In_124,In_0);
and U699 (N_699,In_31,In_201);
nor U700 (N_700,In_340,In_169);
nor U701 (N_701,In_351,In_267);
or U702 (N_702,In_479,In_296);
and U703 (N_703,In_143,In_281);
and U704 (N_704,In_16,In_108);
nand U705 (N_705,In_430,In_367);
or U706 (N_706,In_153,In_82);
xor U707 (N_707,In_244,In_302);
or U708 (N_708,In_306,In_379);
nor U709 (N_709,In_173,In_70);
and U710 (N_710,In_377,In_130);
nor U711 (N_711,In_355,In_196);
and U712 (N_712,In_211,In_215);
or U713 (N_713,In_301,In_184);
or U714 (N_714,In_204,In_332);
nor U715 (N_715,In_286,In_431);
or U716 (N_716,In_33,In_96);
and U717 (N_717,In_31,In_46);
nor U718 (N_718,In_442,In_47);
or U719 (N_719,In_422,In_280);
or U720 (N_720,In_184,In_99);
or U721 (N_721,In_430,In_324);
or U722 (N_722,In_103,In_259);
nand U723 (N_723,In_312,In_31);
nor U724 (N_724,In_350,In_370);
and U725 (N_725,In_120,In_2);
and U726 (N_726,In_357,In_244);
nor U727 (N_727,In_338,In_197);
nor U728 (N_728,In_109,In_13);
and U729 (N_729,In_335,In_30);
nor U730 (N_730,In_207,In_480);
and U731 (N_731,In_120,In_135);
nand U732 (N_732,In_45,In_53);
and U733 (N_733,In_226,In_165);
nor U734 (N_734,In_324,In_105);
and U735 (N_735,In_439,In_430);
nand U736 (N_736,In_178,In_123);
or U737 (N_737,In_458,In_16);
or U738 (N_738,In_132,In_375);
or U739 (N_739,In_299,In_301);
and U740 (N_740,In_10,In_386);
nand U741 (N_741,In_214,In_294);
and U742 (N_742,In_198,In_165);
and U743 (N_743,In_172,In_29);
and U744 (N_744,In_154,In_466);
nor U745 (N_745,In_224,In_46);
nand U746 (N_746,In_305,In_228);
nor U747 (N_747,In_77,In_95);
and U748 (N_748,In_345,In_201);
and U749 (N_749,In_111,In_172);
or U750 (N_750,In_464,In_235);
nor U751 (N_751,In_445,In_406);
nor U752 (N_752,In_404,In_488);
and U753 (N_753,In_137,In_142);
and U754 (N_754,In_386,In_68);
nand U755 (N_755,In_484,In_354);
and U756 (N_756,In_111,In_14);
and U757 (N_757,In_103,In_212);
nand U758 (N_758,In_233,In_454);
nand U759 (N_759,In_308,In_396);
nand U760 (N_760,In_386,In_240);
nor U761 (N_761,In_171,In_443);
or U762 (N_762,In_337,In_15);
nor U763 (N_763,In_242,In_24);
nor U764 (N_764,In_348,In_485);
nor U765 (N_765,In_79,In_491);
or U766 (N_766,In_433,In_92);
and U767 (N_767,In_155,In_358);
nor U768 (N_768,In_101,In_247);
and U769 (N_769,In_429,In_248);
or U770 (N_770,In_405,In_2);
and U771 (N_771,In_363,In_284);
and U772 (N_772,In_372,In_7);
nor U773 (N_773,In_192,In_434);
nand U774 (N_774,In_332,In_15);
nor U775 (N_775,In_323,In_45);
or U776 (N_776,In_494,In_345);
nor U777 (N_777,In_138,In_213);
xnor U778 (N_778,In_165,In_115);
nor U779 (N_779,In_393,In_445);
or U780 (N_780,In_131,In_237);
nand U781 (N_781,In_111,In_211);
and U782 (N_782,In_179,In_138);
nand U783 (N_783,In_213,In_484);
and U784 (N_784,In_309,In_129);
or U785 (N_785,In_179,In_123);
or U786 (N_786,In_80,In_214);
nor U787 (N_787,In_230,In_183);
nor U788 (N_788,In_53,In_256);
nor U789 (N_789,In_300,In_247);
nor U790 (N_790,In_340,In_255);
or U791 (N_791,In_146,In_327);
nor U792 (N_792,In_365,In_206);
and U793 (N_793,In_236,In_195);
nand U794 (N_794,In_65,In_438);
nand U795 (N_795,In_198,In_461);
nand U796 (N_796,In_163,In_385);
nand U797 (N_797,In_492,In_399);
or U798 (N_798,In_412,In_237);
nor U799 (N_799,In_478,In_21);
and U800 (N_800,In_176,In_28);
nand U801 (N_801,In_434,In_30);
xor U802 (N_802,In_278,In_383);
nor U803 (N_803,In_426,In_494);
xor U804 (N_804,In_292,In_138);
nand U805 (N_805,In_461,In_84);
and U806 (N_806,In_320,In_239);
nand U807 (N_807,In_198,In_235);
nand U808 (N_808,In_365,In_236);
nand U809 (N_809,In_223,In_416);
nor U810 (N_810,In_176,In_216);
nor U811 (N_811,In_233,In_419);
nor U812 (N_812,In_485,In_56);
xnor U813 (N_813,In_213,In_78);
and U814 (N_814,In_260,In_126);
or U815 (N_815,In_434,In_41);
nand U816 (N_816,In_398,In_15);
xor U817 (N_817,In_281,In_232);
nor U818 (N_818,In_267,In_437);
nor U819 (N_819,In_379,In_328);
nor U820 (N_820,In_384,In_131);
nand U821 (N_821,In_29,In_153);
or U822 (N_822,In_32,In_41);
nand U823 (N_823,In_188,In_43);
and U824 (N_824,In_455,In_365);
nand U825 (N_825,In_102,In_456);
nand U826 (N_826,In_108,In_277);
xor U827 (N_827,In_416,In_449);
nand U828 (N_828,In_494,In_24);
and U829 (N_829,In_126,In_495);
nor U830 (N_830,In_98,In_185);
nand U831 (N_831,In_326,In_218);
or U832 (N_832,In_201,In_251);
nand U833 (N_833,In_255,In_487);
nor U834 (N_834,In_123,In_406);
and U835 (N_835,In_162,In_457);
nand U836 (N_836,In_187,In_338);
nand U837 (N_837,In_74,In_343);
and U838 (N_838,In_468,In_226);
xnor U839 (N_839,In_262,In_274);
nand U840 (N_840,In_431,In_401);
and U841 (N_841,In_134,In_278);
nand U842 (N_842,In_317,In_217);
and U843 (N_843,In_273,In_73);
nor U844 (N_844,In_98,In_366);
nor U845 (N_845,In_317,In_295);
nand U846 (N_846,In_256,In_302);
nor U847 (N_847,In_114,In_473);
xnor U848 (N_848,In_25,In_257);
nand U849 (N_849,In_11,In_400);
nand U850 (N_850,In_109,In_314);
xnor U851 (N_851,In_85,In_32);
and U852 (N_852,In_15,In_71);
nand U853 (N_853,In_480,In_165);
nor U854 (N_854,In_394,In_209);
nand U855 (N_855,In_27,In_489);
or U856 (N_856,In_254,In_337);
nand U857 (N_857,In_133,In_356);
nand U858 (N_858,In_231,In_398);
nor U859 (N_859,In_273,In_288);
nor U860 (N_860,In_420,In_409);
or U861 (N_861,In_309,In_273);
nor U862 (N_862,In_130,In_298);
or U863 (N_863,In_462,In_56);
nand U864 (N_864,In_333,In_380);
xor U865 (N_865,In_108,In_380);
nand U866 (N_866,In_249,In_101);
nand U867 (N_867,In_102,In_152);
and U868 (N_868,In_449,In_297);
nor U869 (N_869,In_32,In_14);
and U870 (N_870,In_6,In_428);
nor U871 (N_871,In_28,In_347);
and U872 (N_872,In_457,In_23);
and U873 (N_873,In_180,In_186);
and U874 (N_874,In_412,In_398);
nand U875 (N_875,In_224,In_462);
nor U876 (N_876,In_51,In_239);
nor U877 (N_877,In_276,In_372);
xor U878 (N_878,In_464,In_399);
nand U879 (N_879,In_425,In_89);
and U880 (N_880,In_104,In_183);
and U881 (N_881,In_496,In_292);
xor U882 (N_882,In_377,In_198);
or U883 (N_883,In_244,In_167);
nand U884 (N_884,In_476,In_375);
or U885 (N_885,In_53,In_271);
nand U886 (N_886,In_237,In_147);
or U887 (N_887,In_20,In_3);
nor U888 (N_888,In_95,In_435);
xor U889 (N_889,In_244,In_15);
and U890 (N_890,In_491,In_416);
nand U891 (N_891,In_242,In_218);
and U892 (N_892,In_426,In_131);
and U893 (N_893,In_372,In_245);
and U894 (N_894,In_474,In_390);
nor U895 (N_895,In_241,In_54);
and U896 (N_896,In_420,In_473);
and U897 (N_897,In_448,In_422);
and U898 (N_898,In_135,In_382);
or U899 (N_899,In_202,In_122);
nor U900 (N_900,In_340,In_417);
and U901 (N_901,In_436,In_242);
or U902 (N_902,In_130,In_289);
nand U903 (N_903,In_61,In_203);
nand U904 (N_904,In_420,In_340);
nor U905 (N_905,In_139,In_78);
xor U906 (N_906,In_292,In_103);
or U907 (N_907,In_450,In_474);
nor U908 (N_908,In_459,In_97);
and U909 (N_909,In_168,In_445);
nor U910 (N_910,In_461,In_259);
nor U911 (N_911,In_301,In_14);
nand U912 (N_912,In_86,In_12);
and U913 (N_913,In_367,In_256);
nand U914 (N_914,In_404,In_147);
and U915 (N_915,In_61,In_330);
and U916 (N_916,In_472,In_191);
and U917 (N_917,In_287,In_480);
and U918 (N_918,In_433,In_235);
nor U919 (N_919,In_131,In_359);
nand U920 (N_920,In_473,In_440);
or U921 (N_921,In_466,In_382);
and U922 (N_922,In_41,In_300);
and U923 (N_923,In_50,In_121);
xnor U924 (N_924,In_251,In_300);
xnor U925 (N_925,In_420,In_389);
or U926 (N_926,In_323,In_267);
or U927 (N_927,In_463,In_57);
nand U928 (N_928,In_455,In_430);
or U929 (N_929,In_124,In_192);
and U930 (N_930,In_186,In_76);
nor U931 (N_931,In_110,In_90);
and U932 (N_932,In_462,In_377);
and U933 (N_933,In_60,In_493);
or U934 (N_934,In_261,In_136);
and U935 (N_935,In_178,In_275);
nand U936 (N_936,In_105,In_153);
nor U937 (N_937,In_471,In_305);
nor U938 (N_938,In_143,In_471);
or U939 (N_939,In_473,In_168);
or U940 (N_940,In_326,In_69);
xor U941 (N_941,In_170,In_188);
or U942 (N_942,In_330,In_464);
and U943 (N_943,In_7,In_392);
or U944 (N_944,In_427,In_67);
or U945 (N_945,In_307,In_249);
nand U946 (N_946,In_412,In_413);
nor U947 (N_947,In_248,In_454);
and U948 (N_948,In_157,In_217);
or U949 (N_949,In_390,In_197);
and U950 (N_950,In_373,In_304);
nand U951 (N_951,In_18,In_401);
or U952 (N_952,In_312,In_274);
or U953 (N_953,In_307,In_410);
nand U954 (N_954,In_149,In_116);
nor U955 (N_955,In_162,In_131);
nor U956 (N_956,In_344,In_179);
nor U957 (N_957,In_339,In_201);
nor U958 (N_958,In_3,In_497);
nand U959 (N_959,In_387,In_95);
nand U960 (N_960,In_244,In_21);
nand U961 (N_961,In_497,In_458);
xor U962 (N_962,In_195,In_159);
nand U963 (N_963,In_199,In_305);
and U964 (N_964,In_157,In_353);
or U965 (N_965,In_264,In_3);
and U966 (N_966,In_71,In_91);
nor U967 (N_967,In_381,In_7);
or U968 (N_968,In_297,In_238);
or U969 (N_969,In_73,In_15);
nor U970 (N_970,In_299,In_494);
nor U971 (N_971,In_457,In_125);
xor U972 (N_972,In_280,In_277);
nand U973 (N_973,In_199,In_206);
nor U974 (N_974,In_242,In_150);
or U975 (N_975,In_483,In_424);
nor U976 (N_976,In_42,In_381);
or U977 (N_977,In_87,In_494);
and U978 (N_978,In_417,In_328);
nand U979 (N_979,In_240,In_278);
or U980 (N_980,In_12,In_173);
or U981 (N_981,In_128,In_275);
and U982 (N_982,In_442,In_228);
nor U983 (N_983,In_291,In_356);
nand U984 (N_984,In_289,In_192);
nand U985 (N_985,In_351,In_279);
nand U986 (N_986,In_319,In_453);
nand U987 (N_987,In_197,In_388);
nand U988 (N_988,In_178,In_286);
nand U989 (N_989,In_53,In_446);
and U990 (N_990,In_318,In_372);
and U991 (N_991,In_494,In_465);
or U992 (N_992,In_230,In_242);
nand U993 (N_993,In_357,In_103);
nor U994 (N_994,In_2,In_178);
or U995 (N_995,In_347,In_236);
or U996 (N_996,In_291,In_64);
and U997 (N_997,In_425,In_220);
nor U998 (N_998,In_418,In_299);
or U999 (N_999,In_165,In_43);
and U1000 (N_1000,N_12,N_250);
or U1001 (N_1001,N_621,N_249);
and U1002 (N_1002,N_633,N_143);
nand U1003 (N_1003,N_54,N_996);
nor U1004 (N_1004,N_320,N_152);
nor U1005 (N_1005,N_408,N_614);
nand U1006 (N_1006,N_316,N_115);
and U1007 (N_1007,N_948,N_11);
or U1008 (N_1008,N_596,N_718);
or U1009 (N_1009,N_288,N_314);
or U1010 (N_1010,N_65,N_333);
and U1011 (N_1011,N_912,N_615);
or U1012 (N_1012,N_88,N_925);
nand U1013 (N_1013,N_165,N_432);
or U1014 (N_1014,N_370,N_50);
and U1015 (N_1015,N_375,N_185);
and U1016 (N_1016,N_772,N_368);
and U1017 (N_1017,N_737,N_608);
nor U1018 (N_1018,N_167,N_95);
and U1019 (N_1019,N_955,N_892);
and U1020 (N_1020,N_496,N_889);
nor U1021 (N_1021,N_819,N_295);
and U1022 (N_1022,N_126,N_939);
nor U1023 (N_1023,N_349,N_319);
nor U1024 (N_1024,N_949,N_10);
nand U1025 (N_1025,N_733,N_758);
nand U1026 (N_1026,N_776,N_492);
and U1027 (N_1027,N_373,N_573);
nand U1028 (N_1028,N_240,N_273);
and U1029 (N_1029,N_936,N_961);
and U1030 (N_1030,N_312,N_37);
and U1031 (N_1031,N_460,N_548);
and U1032 (N_1032,N_636,N_729);
or U1033 (N_1033,N_383,N_588);
nor U1034 (N_1034,N_982,N_626);
nor U1035 (N_1035,N_875,N_235);
and U1036 (N_1036,N_26,N_637);
or U1037 (N_1037,N_331,N_799);
and U1038 (N_1038,N_566,N_645);
or U1039 (N_1039,N_157,N_278);
and U1040 (N_1040,N_967,N_751);
nand U1041 (N_1041,N_199,N_835);
xnor U1042 (N_1042,N_502,N_505);
nor U1043 (N_1043,N_14,N_63);
or U1044 (N_1044,N_180,N_710);
nand U1045 (N_1045,N_29,N_155);
nor U1046 (N_1046,N_785,N_988);
and U1047 (N_1047,N_68,N_494);
or U1048 (N_1048,N_840,N_914);
nand U1049 (N_1049,N_653,N_591);
or U1050 (N_1050,N_145,N_438);
nand U1051 (N_1051,N_31,N_742);
and U1052 (N_1052,N_711,N_267);
or U1053 (N_1053,N_787,N_469);
nor U1054 (N_1054,N_233,N_191);
and U1055 (N_1055,N_509,N_232);
and U1056 (N_1056,N_123,N_0);
or U1057 (N_1057,N_499,N_523);
or U1058 (N_1058,N_649,N_693);
or U1059 (N_1059,N_485,N_226);
or U1060 (N_1060,N_407,N_89);
nor U1061 (N_1061,N_462,N_382);
and U1062 (N_1062,N_995,N_39);
nand U1063 (N_1063,N_38,N_582);
or U1064 (N_1064,N_218,N_625);
nor U1065 (N_1065,N_482,N_87);
nor U1066 (N_1066,N_285,N_946);
nor U1067 (N_1067,N_47,N_928);
nor U1068 (N_1068,N_823,N_712);
and U1069 (N_1069,N_13,N_365);
xor U1070 (N_1070,N_170,N_577);
nand U1071 (N_1071,N_24,N_203);
and U1072 (N_1072,N_471,N_28);
or U1073 (N_1073,N_215,N_581);
or U1074 (N_1074,N_397,N_513);
nand U1075 (N_1075,N_102,N_683);
or U1076 (N_1076,N_611,N_9);
xor U1077 (N_1077,N_586,N_998);
or U1078 (N_1078,N_966,N_77);
and U1079 (N_1079,N_868,N_725);
xor U1080 (N_1080,N_217,N_389);
nand U1081 (N_1081,N_832,N_275);
or U1082 (N_1082,N_325,N_94);
or U1083 (N_1083,N_594,N_488);
and U1084 (N_1084,N_197,N_16);
xnor U1085 (N_1085,N_585,N_357);
and U1086 (N_1086,N_470,N_72);
or U1087 (N_1087,N_701,N_562);
nand U1088 (N_1088,N_980,N_794);
and U1089 (N_1089,N_107,N_335);
nand U1090 (N_1090,N_527,N_259);
and U1091 (N_1091,N_71,N_74);
nand U1092 (N_1092,N_284,N_108);
xor U1093 (N_1093,N_866,N_779);
or U1094 (N_1094,N_67,N_981);
nor U1095 (N_1095,N_940,N_757);
nand U1096 (N_1096,N_668,N_714);
nand U1097 (N_1097,N_196,N_878);
nor U1098 (N_1098,N_907,N_650);
nand U1099 (N_1099,N_474,N_112);
nand U1100 (N_1100,N_193,N_436);
and U1101 (N_1101,N_337,N_330);
and U1102 (N_1102,N_334,N_392);
and U1103 (N_1103,N_201,N_628);
and U1104 (N_1104,N_703,N_506);
nor U1105 (N_1105,N_261,N_831);
or U1106 (N_1106,N_51,N_211);
and U1107 (N_1107,N_192,N_959);
nand U1108 (N_1108,N_526,N_796);
nor U1109 (N_1109,N_209,N_321);
or U1110 (N_1110,N_516,N_773);
and U1111 (N_1111,N_713,N_913);
nand U1112 (N_1112,N_789,N_704);
and U1113 (N_1113,N_223,N_539);
and U1114 (N_1114,N_290,N_243);
nand U1115 (N_1115,N_378,N_778);
nand U1116 (N_1116,N_663,N_834);
or U1117 (N_1117,N_416,N_457);
and U1118 (N_1118,N_876,N_410);
xnor U1119 (N_1119,N_696,N_919);
and U1120 (N_1120,N_991,N_260);
nor U1121 (N_1121,N_752,N_700);
or U1122 (N_1122,N_227,N_916);
or U1123 (N_1123,N_859,N_161);
or U1124 (N_1124,N_962,N_141);
nand U1125 (N_1125,N_935,N_113);
xnor U1126 (N_1126,N_297,N_134);
nand U1127 (N_1127,N_437,N_555);
xnor U1128 (N_1128,N_672,N_427);
or U1129 (N_1129,N_993,N_390);
xnor U1130 (N_1130,N_786,N_4);
nor U1131 (N_1131,N_43,N_403);
and U1132 (N_1132,N_453,N_556);
or U1133 (N_1133,N_184,N_651);
nand U1134 (N_1134,N_323,N_497);
or U1135 (N_1135,N_564,N_27);
nand U1136 (N_1136,N_56,N_309);
nand U1137 (N_1137,N_873,N_906);
nand U1138 (N_1138,N_341,N_424);
nor U1139 (N_1139,N_932,N_271);
or U1140 (N_1140,N_887,N_620);
or U1141 (N_1141,N_520,N_244);
nor U1142 (N_1142,N_746,N_613);
nand U1143 (N_1143,N_533,N_118);
or U1144 (N_1144,N_781,N_854);
nand U1145 (N_1145,N_396,N_768);
nor U1146 (N_1146,N_446,N_345);
and U1147 (N_1147,N_754,N_419);
and U1148 (N_1148,N_874,N_549);
and U1149 (N_1149,N_968,N_904);
nand U1150 (N_1150,N_190,N_810);
nor U1151 (N_1151,N_673,N_182);
or U1152 (N_1152,N_300,N_521);
nor U1153 (N_1153,N_36,N_519);
nor U1154 (N_1154,N_992,N_229);
xnor U1155 (N_1155,N_158,N_133);
xnor U1156 (N_1156,N_797,N_830);
nor U1157 (N_1157,N_138,N_40);
nand U1158 (N_1158,N_739,N_336);
or U1159 (N_1159,N_144,N_160);
nor U1160 (N_1160,N_524,N_52);
or U1161 (N_1161,N_719,N_281);
and U1162 (N_1162,N_164,N_808);
and U1163 (N_1163,N_2,N_366);
or U1164 (N_1164,N_553,N_332);
or U1165 (N_1165,N_542,N_986);
xor U1166 (N_1166,N_400,N_671);
nor U1167 (N_1167,N_247,N_872);
or U1168 (N_1168,N_895,N_25);
nor U1169 (N_1169,N_771,N_537);
nor U1170 (N_1170,N_142,N_237);
xnor U1171 (N_1171,N_764,N_412);
nor U1172 (N_1172,N_150,N_617);
and U1173 (N_1173,N_792,N_589);
or U1174 (N_1174,N_305,N_879);
or U1175 (N_1175,N_486,N_514);
nand U1176 (N_1176,N_805,N_265);
nand U1177 (N_1177,N_641,N_547);
and U1178 (N_1178,N_702,N_579);
xor U1179 (N_1179,N_230,N_745);
xor U1180 (N_1180,N_952,N_618);
or U1181 (N_1181,N_707,N_536);
and U1182 (N_1182,N_634,N_81);
nor U1183 (N_1183,N_747,N_691);
nand U1184 (N_1184,N_163,N_865);
and U1185 (N_1185,N_350,N_353);
nor U1186 (N_1186,N_664,N_210);
nand U1187 (N_1187,N_688,N_19);
nand U1188 (N_1188,N_224,N_97);
nor U1189 (N_1189,N_256,N_116);
nor U1190 (N_1190,N_607,N_443);
nor U1191 (N_1191,N_911,N_489);
and U1192 (N_1192,N_421,N_58);
or U1193 (N_1193,N_558,N_45);
xor U1194 (N_1194,N_395,N_544);
nor U1195 (N_1195,N_769,N_23);
nor U1196 (N_1196,N_682,N_66);
or U1197 (N_1197,N_156,N_624);
nor U1198 (N_1198,N_643,N_705);
nor U1199 (N_1199,N_803,N_99);
or U1200 (N_1200,N_84,N_299);
nor U1201 (N_1201,N_827,N_855);
nand U1202 (N_1202,N_619,N_128);
nand U1203 (N_1203,N_136,N_61);
nor U1204 (N_1204,N_724,N_857);
and U1205 (N_1205,N_379,N_780);
or U1206 (N_1206,N_678,N_263);
xor U1207 (N_1207,N_79,N_110);
nor U1208 (N_1208,N_820,N_606);
nand U1209 (N_1209,N_600,N_900);
and U1210 (N_1210,N_388,N_644);
or U1211 (N_1211,N_372,N_902);
and U1212 (N_1212,N_604,N_293);
or U1213 (N_1213,N_983,N_756);
nor U1214 (N_1214,N_569,N_475);
nor U1215 (N_1215,N_816,N_638);
nand U1216 (N_1216,N_730,N_91);
nor U1217 (N_1217,N_572,N_120);
or U1218 (N_1218,N_565,N_871);
or U1219 (N_1219,N_49,N_694);
or U1220 (N_1220,N_270,N_225);
or U1221 (N_1221,N_698,N_795);
nor U1222 (N_1222,N_124,N_103);
xnor U1223 (N_1223,N_491,N_930);
nor U1224 (N_1224,N_863,N_317);
or U1225 (N_1225,N_838,N_257);
or U1226 (N_1226,N_447,N_266);
nor U1227 (N_1227,N_53,N_80);
xor U1228 (N_1228,N_287,N_194);
or U1229 (N_1229,N_896,N_846);
and U1230 (N_1230,N_122,N_836);
nand U1231 (N_1231,N_105,N_692);
or U1232 (N_1232,N_169,N_958);
nor U1233 (N_1233,N_528,N_276);
or U1234 (N_1234,N_356,N_950);
and U1235 (N_1235,N_119,N_440);
nand U1236 (N_1236,N_655,N_583);
nand U1237 (N_1237,N_931,N_175);
nor U1238 (N_1238,N_951,N_479);
or U1239 (N_1239,N_851,N_759);
nor U1240 (N_1240,N_717,N_347);
and U1241 (N_1241,N_748,N_439);
nand U1242 (N_1242,N_723,N_953);
nor U1243 (N_1243,N_22,N_393);
nor U1244 (N_1244,N_377,N_352);
nor U1245 (N_1245,N_699,N_8);
nand U1246 (N_1246,N_363,N_550);
and U1247 (N_1247,N_679,N_587);
nor U1248 (N_1248,N_522,N_60);
and U1249 (N_1249,N_493,N_315);
nand U1250 (N_1250,N_367,N_695);
or U1251 (N_1251,N_977,N_64);
nor U1252 (N_1252,N_844,N_777);
nor U1253 (N_1253,N_860,N_665);
nor U1254 (N_1254,N_517,N_741);
or U1255 (N_1255,N_411,N_599);
or U1256 (N_1256,N_384,N_590);
or U1257 (N_1257,N_279,N_921);
and U1258 (N_1258,N_984,N_195);
or U1259 (N_1259,N_463,N_770);
nand U1260 (N_1260,N_34,N_697);
and U1261 (N_1261,N_861,N_114);
nor U1262 (N_1262,N_616,N_231);
xor U1263 (N_1263,N_455,N_924);
nand U1264 (N_1264,N_530,N_503);
nor U1265 (N_1265,N_578,N_46);
or U1266 (N_1266,N_391,N_570);
or U1267 (N_1267,N_121,N_677);
or U1268 (N_1268,N_510,N_749);
or U1269 (N_1269,N_632,N_883);
and U1270 (N_1270,N_728,N_277);
nand U1271 (N_1271,N_405,N_371);
or U1272 (N_1272,N_800,N_21);
or U1273 (N_1273,N_534,N_867);
nor U1274 (N_1274,N_918,N_426);
or U1275 (N_1275,N_675,N_82);
or U1276 (N_1276,N_812,N_721);
or U1277 (N_1277,N_85,N_690);
nor U1278 (N_1278,N_441,N_69);
or U1279 (N_1279,N_344,N_689);
or U1280 (N_1280,N_814,N_659);
and U1281 (N_1281,N_593,N_853);
and U1282 (N_1282,N_922,N_359);
nor U1283 (N_1283,N_401,N_971);
nand U1284 (N_1284,N_508,N_30);
or U1285 (N_1285,N_755,N_765);
xnor U1286 (N_1286,N_512,N_763);
nand U1287 (N_1287,N_686,N_822);
or U1288 (N_1288,N_923,N_848);
nor U1289 (N_1289,N_767,N_461);
and U1290 (N_1290,N_131,N_272);
or U1291 (N_1291,N_417,N_35);
nor U1292 (N_1292,N_465,N_760);
nand U1293 (N_1293,N_847,N_880);
nor U1294 (N_1294,N_662,N_456);
and U1295 (N_1295,N_652,N_434);
or U1296 (N_1296,N_228,N_858);
nand U1297 (N_1297,N_212,N_674);
nand U1298 (N_1298,N_829,N_938);
and U1299 (N_1299,N_444,N_654);
nand U1300 (N_1300,N_842,N_111);
nand U1301 (N_1301,N_669,N_850);
nor U1302 (N_1302,N_18,N_535);
nor U1303 (N_1303,N_478,N_660);
nand U1304 (N_1304,N_881,N_920);
nor U1305 (N_1305,N_648,N_62);
nor U1306 (N_1306,N_917,N_130);
nand U1307 (N_1307,N_109,N_430);
xor U1308 (N_1308,N_788,N_48);
nand U1309 (N_1309,N_135,N_162);
nor U1310 (N_1310,N_268,N_413);
xor U1311 (N_1311,N_623,N_198);
and U1312 (N_1312,N_525,N_908);
nand U1313 (N_1313,N_498,N_743);
nor U1314 (N_1314,N_732,N_355);
or U1315 (N_1315,N_687,N_464);
nor U1316 (N_1316,N_989,N_399);
and U1317 (N_1317,N_398,N_507);
or U1318 (N_1318,N_106,N_327);
nor U1319 (N_1319,N_20,N_804);
and U1320 (N_1320,N_269,N_59);
nor U1321 (N_1321,N_943,N_999);
or U1322 (N_1322,N_477,N_428);
and U1323 (N_1323,N_483,N_204);
or U1324 (N_1324,N_934,N_200);
nand U1325 (N_1325,N_964,N_845);
or U1326 (N_1326,N_234,N_258);
nor U1327 (N_1327,N_329,N_406);
nand U1328 (N_1328,N_985,N_100);
nor U1329 (N_1329,N_178,N_364);
nor U1330 (N_1330,N_560,N_839);
or U1331 (N_1331,N_956,N_969);
or U1332 (N_1332,N_775,N_639);
or U1333 (N_1333,N_744,N_450);
or U1334 (N_1334,N_214,N_610);
nor U1335 (N_1335,N_975,N_93);
nor U1336 (N_1336,N_96,N_394);
and U1337 (N_1337,N_283,N_709);
and U1338 (N_1338,N_843,N_90);
or U1339 (N_1339,N_6,N_905);
nor U1340 (N_1340,N_70,N_166);
or U1341 (N_1341,N_974,N_670);
and U1342 (N_1342,N_298,N_358);
nand U1343 (N_1343,N_891,N_997);
and U1344 (N_1344,N_117,N_442);
nand U1345 (N_1345,N_903,N_33);
and U1346 (N_1346,N_806,N_972);
xor U1347 (N_1347,N_540,N_168);
nor U1348 (N_1348,N_264,N_963);
and U1349 (N_1349,N_445,N_852);
nor U1350 (N_1350,N_484,N_973);
and U1351 (N_1351,N_627,N_206);
nand U1352 (N_1352,N_597,N_960);
nor U1353 (N_1353,N_481,N_708);
xnor U1354 (N_1354,N_149,N_612);
and U1355 (N_1355,N_304,N_76);
nor U1356 (N_1356,N_761,N_361);
nand U1357 (N_1357,N_125,N_947);
nor U1358 (N_1358,N_216,N_342);
or U1359 (N_1359,N_381,N_893);
nor U1360 (N_1360,N_140,N_684);
and U1361 (N_1361,N_584,N_807);
and U1362 (N_1362,N_657,N_177);
nand U1363 (N_1363,N_559,N_990);
nand U1364 (N_1364,N_734,N_55);
or U1365 (N_1365,N_374,N_369);
and U1366 (N_1366,N_176,N_531);
and U1367 (N_1367,N_576,N_159);
or U1368 (N_1368,N_1,N_504);
or U1369 (N_1369,N_574,N_255);
and U1370 (N_1370,N_976,N_837);
or U1371 (N_1371,N_793,N_236);
nand U1372 (N_1372,N_98,N_220);
and U1373 (N_1373,N_221,N_248);
nand U1374 (N_1374,N_825,N_245);
nor U1375 (N_1375,N_622,N_360);
nor U1376 (N_1376,N_635,N_385);
or U1377 (N_1377,N_821,N_862);
or U1378 (N_1378,N_127,N_41);
nor U1379 (N_1379,N_802,N_75);
nor U1380 (N_1380,N_941,N_899);
and U1381 (N_1381,N_720,N_459);
nor U1382 (N_1382,N_306,N_296);
nor U1383 (N_1383,N_318,N_376);
nor U1384 (N_1384,N_313,N_351);
or U1385 (N_1385,N_877,N_580);
nand U1386 (N_1386,N_605,N_292);
xnor U1387 (N_1387,N_529,N_307);
nand U1388 (N_1388,N_291,N_685);
nand U1389 (N_1389,N_640,N_246);
or U1390 (N_1390,N_104,N_824);
or U1391 (N_1391,N_811,N_557);
or U1392 (N_1392,N_929,N_894);
nor U1393 (N_1393,N_32,N_603);
or U1394 (N_1394,N_338,N_181);
or U1395 (N_1395,N_354,N_783);
and U1396 (N_1396,N_186,N_173);
nor U1397 (N_1397,N_801,N_809);
and U1398 (N_1398,N_595,N_568);
nand U1399 (N_1399,N_219,N_425);
nor U1400 (N_1400,N_954,N_841);
or U1401 (N_1401,N_42,N_602);
and U1402 (N_1402,N_994,N_910);
nor U1403 (N_1403,N_86,N_476);
or U1404 (N_1404,N_495,N_715);
and U1405 (N_1405,N_552,N_656);
nor U1406 (N_1406,N_926,N_44);
or U1407 (N_1407,N_241,N_500);
nor U1408 (N_1408,N_987,N_818);
nor U1409 (N_1409,N_592,N_137);
nor U1410 (N_1410,N_658,N_791);
nand U1411 (N_1411,N_680,N_187);
nor U1412 (N_1412,N_418,N_414);
nand U1413 (N_1413,N_251,N_945);
and U1414 (N_1414,N_601,N_890);
nand U1415 (N_1415,N_7,N_282);
and U1416 (N_1416,N_647,N_518);
or U1417 (N_1417,N_3,N_207);
or U1418 (N_1418,N_646,N_92);
nand U1419 (N_1419,N_833,N_466);
nand U1420 (N_1420,N_735,N_431);
or U1421 (N_1421,N_753,N_380);
nand U1422 (N_1422,N_172,N_609);
and U1423 (N_1423,N_815,N_253);
nor U1424 (N_1424,N_563,N_933);
nand U1425 (N_1425,N_490,N_362);
or U1426 (N_1426,N_189,N_454);
and U1427 (N_1427,N_629,N_151);
xnor U1428 (N_1428,N_409,N_501);
nand U1429 (N_1429,N_101,N_642);
nand U1430 (N_1430,N_979,N_681);
and U1431 (N_1431,N_179,N_885);
xor U1432 (N_1432,N_856,N_915);
xnor U1433 (N_1433,N_942,N_706);
nand U1434 (N_1434,N_554,N_965);
and U1435 (N_1435,N_551,N_139);
nand U1436 (N_1436,N_543,N_561);
and U1437 (N_1437,N_901,N_154);
nand U1438 (N_1438,N_449,N_864);
nand U1439 (N_1439,N_420,N_676);
nand U1440 (N_1440,N_541,N_262);
or U1441 (N_1441,N_458,N_452);
or U1442 (N_1442,N_302,N_386);
and U1443 (N_1443,N_826,N_937);
nor U1444 (N_1444,N_205,N_898);
nand U1445 (N_1445,N_340,N_736);
and U1446 (N_1446,N_15,N_762);
or U1447 (N_1447,N_666,N_433);
xor U1448 (N_1448,N_828,N_472);
and U1449 (N_1449,N_174,N_310);
and U1450 (N_1450,N_303,N_208);
nand U1451 (N_1451,N_897,N_239);
or U1452 (N_1452,N_132,N_222);
nor U1453 (N_1453,N_750,N_188);
or U1454 (N_1454,N_798,N_301);
and U1455 (N_1455,N_927,N_740);
or U1456 (N_1456,N_782,N_545);
or U1457 (N_1457,N_404,N_57);
xnor U1458 (N_1458,N_511,N_567);
or U1459 (N_1459,N_286,N_886);
or U1460 (N_1460,N_448,N_83);
and U1461 (N_1461,N_661,N_869);
nor U1462 (N_1462,N_348,N_451);
nand U1463 (N_1463,N_909,N_242);
nand U1464 (N_1464,N_978,N_343);
or U1465 (N_1465,N_402,N_5);
or U1466 (N_1466,N_716,N_727);
nand U1467 (N_1467,N_774,N_480);
and U1468 (N_1468,N_813,N_153);
or U1469 (N_1469,N_849,N_435);
nor U1470 (N_1470,N_429,N_346);
xor U1471 (N_1471,N_328,N_870);
xnor U1472 (N_1472,N_571,N_515);
and U1473 (N_1473,N_422,N_970);
or U1474 (N_1474,N_213,N_78);
nand U1475 (N_1475,N_294,N_238);
and U1476 (N_1476,N_731,N_129);
nand U1477 (N_1477,N_784,N_957);
and U1478 (N_1478,N_726,N_146);
nor U1479 (N_1479,N_148,N_630);
nand U1480 (N_1480,N_73,N_473);
nand U1481 (N_1481,N_888,N_468);
and U1482 (N_1482,N_147,N_326);
nand U1483 (N_1483,N_817,N_944);
nor U1484 (N_1484,N_254,N_17);
and U1485 (N_1485,N_538,N_308);
and U1486 (N_1486,N_667,N_423);
or U1487 (N_1487,N_280,N_202);
and U1488 (N_1488,N_339,N_738);
or U1489 (N_1489,N_790,N_289);
or U1490 (N_1490,N_274,N_882);
or U1491 (N_1491,N_467,N_252);
xnor U1492 (N_1492,N_884,N_598);
and U1493 (N_1493,N_322,N_766);
nand U1494 (N_1494,N_324,N_631);
or U1495 (N_1495,N_575,N_722);
and U1496 (N_1496,N_387,N_532);
and U1497 (N_1497,N_183,N_546);
nor U1498 (N_1498,N_171,N_415);
nand U1499 (N_1499,N_311,N_487);
nor U1500 (N_1500,N_891,N_506);
nor U1501 (N_1501,N_772,N_781);
nor U1502 (N_1502,N_200,N_881);
xnor U1503 (N_1503,N_910,N_730);
and U1504 (N_1504,N_341,N_76);
and U1505 (N_1505,N_809,N_125);
nor U1506 (N_1506,N_380,N_563);
or U1507 (N_1507,N_137,N_885);
nand U1508 (N_1508,N_560,N_999);
nand U1509 (N_1509,N_805,N_611);
nor U1510 (N_1510,N_567,N_672);
or U1511 (N_1511,N_915,N_23);
nand U1512 (N_1512,N_536,N_767);
nor U1513 (N_1513,N_800,N_176);
xnor U1514 (N_1514,N_690,N_248);
xor U1515 (N_1515,N_135,N_859);
nand U1516 (N_1516,N_672,N_867);
or U1517 (N_1517,N_653,N_914);
nand U1518 (N_1518,N_23,N_639);
and U1519 (N_1519,N_492,N_147);
nand U1520 (N_1520,N_411,N_132);
nor U1521 (N_1521,N_135,N_66);
and U1522 (N_1522,N_255,N_524);
nand U1523 (N_1523,N_955,N_640);
nor U1524 (N_1524,N_220,N_712);
and U1525 (N_1525,N_918,N_927);
and U1526 (N_1526,N_500,N_517);
or U1527 (N_1527,N_226,N_216);
nor U1528 (N_1528,N_349,N_61);
or U1529 (N_1529,N_951,N_425);
xor U1530 (N_1530,N_461,N_61);
and U1531 (N_1531,N_374,N_50);
nor U1532 (N_1532,N_206,N_34);
and U1533 (N_1533,N_206,N_192);
xnor U1534 (N_1534,N_264,N_954);
nor U1535 (N_1535,N_285,N_579);
and U1536 (N_1536,N_23,N_134);
or U1537 (N_1537,N_881,N_560);
nor U1538 (N_1538,N_467,N_876);
or U1539 (N_1539,N_845,N_809);
and U1540 (N_1540,N_424,N_952);
nand U1541 (N_1541,N_756,N_724);
and U1542 (N_1542,N_29,N_983);
and U1543 (N_1543,N_960,N_63);
nor U1544 (N_1544,N_6,N_241);
nand U1545 (N_1545,N_633,N_990);
nand U1546 (N_1546,N_353,N_945);
nand U1547 (N_1547,N_901,N_309);
nor U1548 (N_1548,N_974,N_504);
nand U1549 (N_1549,N_656,N_584);
xnor U1550 (N_1550,N_559,N_67);
nand U1551 (N_1551,N_576,N_285);
nand U1552 (N_1552,N_149,N_980);
and U1553 (N_1553,N_952,N_61);
nand U1554 (N_1554,N_374,N_927);
nor U1555 (N_1555,N_677,N_978);
or U1556 (N_1556,N_289,N_250);
xnor U1557 (N_1557,N_697,N_721);
or U1558 (N_1558,N_699,N_754);
or U1559 (N_1559,N_731,N_159);
nor U1560 (N_1560,N_896,N_574);
nor U1561 (N_1561,N_441,N_838);
nor U1562 (N_1562,N_77,N_339);
or U1563 (N_1563,N_3,N_629);
nand U1564 (N_1564,N_80,N_461);
xnor U1565 (N_1565,N_649,N_224);
and U1566 (N_1566,N_675,N_397);
or U1567 (N_1567,N_675,N_274);
or U1568 (N_1568,N_65,N_246);
or U1569 (N_1569,N_564,N_976);
or U1570 (N_1570,N_433,N_210);
or U1571 (N_1571,N_347,N_679);
nor U1572 (N_1572,N_655,N_185);
or U1573 (N_1573,N_423,N_504);
nor U1574 (N_1574,N_788,N_808);
or U1575 (N_1575,N_27,N_10);
nor U1576 (N_1576,N_141,N_473);
xnor U1577 (N_1577,N_662,N_158);
nor U1578 (N_1578,N_221,N_309);
xnor U1579 (N_1579,N_594,N_8);
and U1580 (N_1580,N_597,N_144);
nor U1581 (N_1581,N_825,N_575);
and U1582 (N_1582,N_376,N_259);
or U1583 (N_1583,N_249,N_784);
nor U1584 (N_1584,N_680,N_986);
nand U1585 (N_1585,N_394,N_325);
and U1586 (N_1586,N_408,N_501);
nand U1587 (N_1587,N_999,N_271);
nor U1588 (N_1588,N_508,N_907);
nand U1589 (N_1589,N_991,N_561);
xnor U1590 (N_1590,N_86,N_867);
xnor U1591 (N_1591,N_227,N_731);
and U1592 (N_1592,N_229,N_372);
or U1593 (N_1593,N_511,N_960);
and U1594 (N_1594,N_33,N_806);
nand U1595 (N_1595,N_142,N_111);
nor U1596 (N_1596,N_391,N_633);
nor U1597 (N_1597,N_43,N_601);
and U1598 (N_1598,N_427,N_905);
and U1599 (N_1599,N_750,N_419);
and U1600 (N_1600,N_73,N_213);
or U1601 (N_1601,N_278,N_103);
nand U1602 (N_1602,N_148,N_783);
nor U1603 (N_1603,N_331,N_18);
and U1604 (N_1604,N_745,N_855);
nor U1605 (N_1605,N_846,N_510);
and U1606 (N_1606,N_894,N_95);
nand U1607 (N_1607,N_241,N_71);
nor U1608 (N_1608,N_610,N_455);
nor U1609 (N_1609,N_945,N_589);
or U1610 (N_1610,N_775,N_563);
nand U1611 (N_1611,N_762,N_9);
or U1612 (N_1612,N_299,N_954);
xnor U1613 (N_1613,N_656,N_254);
nand U1614 (N_1614,N_60,N_67);
and U1615 (N_1615,N_38,N_167);
and U1616 (N_1616,N_863,N_961);
and U1617 (N_1617,N_522,N_400);
nor U1618 (N_1618,N_277,N_779);
nand U1619 (N_1619,N_931,N_721);
or U1620 (N_1620,N_696,N_477);
and U1621 (N_1621,N_443,N_462);
or U1622 (N_1622,N_269,N_781);
xor U1623 (N_1623,N_286,N_816);
and U1624 (N_1624,N_361,N_632);
and U1625 (N_1625,N_773,N_774);
nand U1626 (N_1626,N_118,N_782);
and U1627 (N_1627,N_444,N_667);
and U1628 (N_1628,N_148,N_678);
or U1629 (N_1629,N_968,N_419);
nor U1630 (N_1630,N_642,N_38);
or U1631 (N_1631,N_730,N_975);
and U1632 (N_1632,N_305,N_613);
and U1633 (N_1633,N_851,N_906);
and U1634 (N_1634,N_331,N_740);
xor U1635 (N_1635,N_744,N_642);
and U1636 (N_1636,N_533,N_679);
or U1637 (N_1637,N_144,N_850);
or U1638 (N_1638,N_372,N_295);
nor U1639 (N_1639,N_602,N_124);
or U1640 (N_1640,N_351,N_679);
nand U1641 (N_1641,N_297,N_296);
xor U1642 (N_1642,N_415,N_493);
or U1643 (N_1643,N_140,N_211);
xor U1644 (N_1644,N_710,N_163);
nor U1645 (N_1645,N_480,N_199);
and U1646 (N_1646,N_657,N_569);
or U1647 (N_1647,N_290,N_191);
nand U1648 (N_1648,N_119,N_42);
or U1649 (N_1649,N_79,N_274);
nand U1650 (N_1650,N_179,N_835);
nor U1651 (N_1651,N_413,N_345);
or U1652 (N_1652,N_824,N_446);
or U1653 (N_1653,N_679,N_28);
nor U1654 (N_1654,N_843,N_327);
and U1655 (N_1655,N_586,N_927);
nand U1656 (N_1656,N_190,N_558);
or U1657 (N_1657,N_663,N_896);
or U1658 (N_1658,N_697,N_392);
nand U1659 (N_1659,N_733,N_873);
nand U1660 (N_1660,N_391,N_187);
xnor U1661 (N_1661,N_937,N_841);
nor U1662 (N_1662,N_945,N_953);
xor U1663 (N_1663,N_175,N_694);
nor U1664 (N_1664,N_822,N_486);
nor U1665 (N_1665,N_177,N_737);
nand U1666 (N_1666,N_55,N_433);
or U1667 (N_1667,N_471,N_767);
or U1668 (N_1668,N_906,N_957);
nand U1669 (N_1669,N_40,N_650);
nor U1670 (N_1670,N_450,N_464);
or U1671 (N_1671,N_885,N_244);
or U1672 (N_1672,N_758,N_898);
or U1673 (N_1673,N_576,N_963);
xor U1674 (N_1674,N_389,N_648);
nor U1675 (N_1675,N_621,N_355);
nand U1676 (N_1676,N_44,N_946);
or U1677 (N_1677,N_944,N_764);
nand U1678 (N_1678,N_123,N_116);
nor U1679 (N_1679,N_902,N_693);
and U1680 (N_1680,N_756,N_260);
nor U1681 (N_1681,N_698,N_785);
nand U1682 (N_1682,N_430,N_817);
nor U1683 (N_1683,N_470,N_588);
and U1684 (N_1684,N_278,N_899);
nand U1685 (N_1685,N_347,N_406);
and U1686 (N_1686,N_0,N_981);
nor U1687 (N_1687,N_195,N_272);
or U1688 (N_1688,N_294,N_723);
and U1689 (N_1689,N_280,N_492);
and U1690 (N_1690,N_846,N_391);
or U1691 (N_1691,N_528,N_689);
and U1692 (N_1692,N_261,N_453);
and U1693 (N_1693,N_160,N_264);
or U1694 (N_1694,N_393,N_96);
xor U1695 (N_1695,N_832,N_417);
nand U1696 (N_1696,N_659,N_278);
or U1697 (N_1697,N_596,N_671);
or U1698 (N_1698,N_630,N_329);
nand U1699 (N_1699,N_603,N_709);
or U1700 (N_1700,N_287,N_525);
nor U1701 (N_1701,N_172,N_550);
xnor U1702 (N_1702,N_274,N_951);
or U1703 (N_1703,N_390,N_96);
or U1704 (N_1704,N_661,N_840);
or U1705 (N_1705,N_116,N_427);
and U1706 (N_1706,N_397,N_511);
nor U1707 (N_1707,N_733,N_502);
and U1708 (N_1708,N_179,N_782);
nand U1709 (N_1709,N_141,N_564);
nor U1710 (N_1710,N_8,N_836);
xor U1711 (N_1711,N_428,N_405);
and U1712 (N_1712,N_155,N_651);
nor U1713 (N_1713,N_651,N_941);
nor U1714 (N_1714,N_623,N_71);
nand U1715 (N_1715,N_54,N_350);
nand U1716 (N_1716,N_457,N_704);
nand U1717 (N_1717,N_649,N_980);
nand U1718 (N_1718,N_774,N_606);
nand U1719 (N_1719,N_68,N_985);
nor U1720 (N_1720,N_879,N_472);
xnor U1721 (N_1721,N_617,N_566);
and U1722 (N_1722,N_264,N_807);
or U1723 (N_1723,N_15,N_230);
and U1724 (N_1724,N_881,N_220);
and U1725 (N_1725,N_248,N_792);
nor U1726 (N_1726,N_641,N_199);
and U1727 (N_1727,N_255,N_717);
nand U1728 (N_1728,N_299,N_526);
and U1729 (N_1729,N_931,N_378);
and U1730 (N_1730,N_708,N_150);
xor U1731 (N_1731,N_276,N_567);
and U1732 (N_1732,N_746,N_659);
and U1733 (N_1733,N_162,N_141);
and U1734 (N_1734,N_217,N_288);
nand U1735 (N_1735,N_237,N_378);
nor U1736 (N_1736,N_483,N_698);
and U1737 (N_1737,N_481,N_777);
and U1738 (N_1738,N_84,N_408);
and U1739 (N_1739,N_1,N_694);
and U1740 (N_1740,N_661,N_908);
and U1741 (N_1741,N_998,N_316);
nor U1742 (N_1742,N_868,N_593);
nand U1743 (N_1743,N_248,N_131);
xnor U1744 (N_1744,N_186,N_336);
or U1745 (N_1745,N_19,N_778);
nor U1746 (N_1746,N_973,N_170);
xor U1747 (N_1747,N_587,N_318);
and U1748 (N_1748,N_522,N_378);
nor U1749 (N_1749,N_747,N_250);
nor U1750 (N_1750,N_951,N_406);
or U1751 (N_1751,N_368,N_150);
xnor U1752 (N_1752,N_904,N_146);
nand U1753 (N_1753,N_551,N_201);
and U1754 (N_1754,N_379,N_743);
nor U1755 (N_1755,N_215,N_384);
nand U1756 (N_1756,N_359,N_696);
nor U1757 (N_1757,N_883,N_983);
nor U1758 (N_1758,N_201,N_974);
nand U1759 (N_1759,N_891,N_364);
and U1760 (N_1760,N_408,N_541);
xnor U1761 (N_1761,N_582,N_99);
nand U1762 (N_1762,N_403,N_809);
or U1763 (N_1763,N_233,N_803);
and U1764 (N_1764,N_131,N_129);
nand U1765 (N_1765,N_355,N_773);
and U1766 (N_1766,N_302,N_246);
nand U1767 (N_1767,N_77,N_838);
xor U1768 (N_1768,N_572,N_430);
or U1769 (N_1769,N_816,N_663);
and U1770 (N_1770,N_607,N_251);
nand U1771 (N_1771,N_398,N_995);
nand U1772 (N_1772,N_461,N_379);
and U1773 (N_1773,N_451,N_201);
nand U1774 (N_1774,N_817,N_603);
nor U1775 (N_1775,N_696,N_491);
nand U1776 (N_1776,N_136,N_841);
nand U1777 (N_1777,N_262,N_886);
nor U1778 (N_1778,N_839,N_325);
nand U1779 (N_1779,N_762,N_304);
nor U1780 (N_1780,N_9,N_83);
nand U1781 (N_1781,N_345,N_411);
xor U1782 (N_1782,N_750,N_244);
or U1783 (N_1783,N_211,N_972);
nand U1784 (N_1784,N_132,N_448);
or U1785 (N_1785,N_474,N_469);
or U1786 (N_1786,N_5,N_313);
and U1787 (N_1787,N_169,N_992);
and U1788 (N_1788,N_479,N_366);
xnor U1789 (N_1789,N_153,N_1);
or U1790 (N_1790,N_541,N_824);
or U1791 (N_1791,N_211,N_943);
or U1792 (N_1792,N_199,N_33);
nand U1793 (N_1793,N_49,N_562);
nor U1794 (N_1794,N_915,N_796);
nor U1795 (N_1795,N_130,N_496);
nand U1796 (N_1796,N_960,N_381);
nor U1797 (N_1797,N_295,N_103);
and U1798 (N_1798,N_519,N_53);
nor U1799 (N_1799,N_300,N_804);
nor U1800 (N_1800,N_703,N_21);
xor U1801 (N_1801,N_259,N_391);
nand U1802 (N_1802,N_652,N_629);
or U1803 (N_1803,N_751,N_122);
nand U1804 (N_1804,N_225,N_209);
or U1805 (N_1805,N_236,N_512);
nor U1806 (N_1806,N_269,N_517);
and U1807 (N_1807,N_449,N_966);
or U1808 (N_1808,N_271,N_800);
nand U1809 (N_1809,N_115,N_455);
nor U1810 (N_1810,N_930,N_875);
xnor U1811 (N_1811,N_470,N_252);
and U1812 (N_1812,N_28,N_542);
and U1813 (N_1813,N_105,N_204);
and U1814 (N_1814,N_814,N_221);
nor U1815 (N_1815,N_87,N_863);
and U1816 (N_1816,N_147,N_819);
and U1817 (N_1817,N_820,N_798);
xor U1818 (N_1818,N_428,N_115);
nand U1819 (N_1819,N_393,N_882);
nor U1820 (N_1820,N_931,N_944);
and U1821 (N_1821,N_595,N_413);
and U1822 (N_1822,N_900,N_332);
or U1823 (N_1823,N_287,N_661);
nand U1824 (N_1824,N_837,N_417);
and U1825 (N_1825,N_791,N_612);
nor U1826 (N_1826,N_480,N_202);
or U1827 (N_1827,N_688,N_605);
nor U1828 (N_1828,N_529,N_479);
or U1829 (N_1829,N_63,N_954);
nand U1830 (N_1830,N_84,N_233);
nand U1831 (N_1831,N_685,N_627);
and U1832 (N_1832,N_569,N_490);
and U1833 (N_1833,N_973,N_699);
or U1834 (N_1834,N_215,N_948);
or U1835 (N_1835,N_827,N_136);
or U1836 (N_1836,N_311,N_344);
and U1837 (N_1837,N_816,N_385);
nor U1838 (N_1838,N_100,N_832);
nand U1839 (N_1839,N_868,N_388);
or U1840 (N_1840,N_302,N_631);
nand U1841 (N_1841,N_836,N_825);
nand U1842 (N_1842,N_70,N_301);
or U1843 (N_1843,N_307,N_76);
nor U1844 (N_1844,N_931,N_735);
or U1845 (N_1845,N_683,N_139);
nand U1846 (N_1846,N_442,N_301);
xnor U1847 (N_1847,N_448,N_732);
and U1848 (N_1848,N_439,N_644);
and U1849 (N_1849,N_38,N_321);
or U1850 (N_1850,N_979,N_367);
nor U1851 (N_1851,N_190,N_863);
nand U1852 (N_1852,N_549,N_115);
and U1853 (N_1853,N_826,N_455);
nand U1854 (N_1854,N_655,N_781);
or U1855 (N_1855,N_436,N_924);
or U1856 (N_1856,N_707,N_145);
nor U1857 (N_1857,N_84,N_29);
nor U1858 (N_1858,N_309,N_564);
nor U1859 (N_1859,N_297,N_337);
nor U1860 (N_1860,N_863,N_965);
and U1861 (N_1861,N_377,N_328);
nor U1862 (N_1862,N_399,N_819);
nor U1863 (N_1863,N_289,N_60);
and U1864 (N_1864,N_886,N_333);
xnor U1865 (N_1865,N_19,N_760);
xor U1866 (N_1866,N_498,N_848);
nand U1867 (N_1867,N_488,N_127);
or U1868 (N_1868,N_689,N_321);
and U1869 (N_1869,N_447,N_251);
or U1870 (N_1870,N_663,N_455);
and U1871 (N_1871,N_59,N_473);
or U1872 (N_1872,N_418,N_758);
nor U1873 (N_1873,N_815,N_449);
or U1874 (N_1874,N_330,N_946);
nor U1875 (N_1875,N_24,N_128);
and U1876 (N_1876,N_509,N_547);
and U1877 (N_1877,N_30,N_525);
or U1878 (N_1878,N_161,N_522);
xnor U1879 (N_1879,N_501,N_229);
nand U1880 (N_1880,N_567,N_72);
nand U1881 (N_1881,N_420,N_141);
nand U1882 (N_1882,N_700,N_890);
nor U1883 (N_1883,N_416,N_647);
nor U1884 (N_1884,N_131,N_921);
and U1885 (N_1885,N_929,N_982);
nand U1886 (N_1886,N_370,N_593);
nand U1887 (N_1887,N_31,N_331);
nand U1888 (N_1888,N_717,N_61);
xnor U1889 (N_1889,N_577,N_202);
nor U1890 (N_1890,N_995,N_178);
nand U1891 (N_1891,N_549,N_143);
or U1892 (N_1892,N_946,N_826);
nor U1893 (N_1893,N_628,N_538);
and U1894 (N_1894,N_235,N_69);
nand U1895 (N_1895,N_646,N_635);
nor U1896 (N_1896,N_81,N_577);
nor U1897 (N_1897,N_333,N_530);
or U1898 (N_1898,N_131,N_138);
or U1899 (N_1899,N_81,N_693);
or U1900 (N_1900,N_723,N_455);
or U1901 (N_1901,N_171,N_633);
or U1902 (N_1902,N_38,N_259);
nand U1903 (N_1903,N_952,N_192);
or U1904 (N_1904,N_917,N_283);
nor U1905 (N_1905,N_616,N_877);
nand U1906 (N_1906,N_67,N_21);
nand U1907 (N_1907,N_569,N_700);
or U1908 (N_1908,N_416,N_649);
xor U1909 (N_1909,N_483,N_540);
xnor U1910 (N_1910,N_474,N_356);
or U1911 (N_1911,N_949,N_953);
nand U1912 (N_1912,N_193,N_333);
nand U1913 (N_1913,N_518,N_639);
nor U1914 (N_1914,N_585,N_119);
or U1915 (N_1915,N_40,N_133);
and U1916 (N_1916,N_30,N_834);
or U1917 (N_1917,N_754,N_723);
and U1918 (N_1918,N_890,N_971);
nor U1919 (N_1919,N_335,N_125);
or U1920 (N_1920,N_908,N_246);
nand U1921 (N_1921,N_89,N_124);
nand U1922 (N_1922,N_370,N_77);
nor U1923 (N_1923,N_689,N_267);
or U1924 (N_1924,N_561,N_365);
nor U1925 (N_1925,N_587,N_469);
or U1926 (N_1926,N_10,N_596);
nor U1927 (N_1927,N_664,N_382);
or U1928 (N_1928,N_503,N_636);
or U1929 (N_1929,N_377,N_522);
and U1930 (N_1930,N_998,N_739);
nand U1931 (N_1931,N_575,N_470);
nor U1932 (N_1932,N_735,N_403);
or U1933 (N_1933,N_791,N_994);
and U1934 (N_1934,N_727,N_909);
xnor U1935 (N_1935,N_195,N_286);
nand U1936 (N_1936,N_135,N_759);
or U1937 (N_1937,N_428,N_620);
or U1938 (N_1938,N_644,N_265);
nor U1939 (N_1939,N_119,N_825);
or U1940 (N_1940,N_166,N_523);
nand U1941 (N_1941,N_889,N_630);
and U1942 (N_1942,N_370,N_982);
and U1943 (N_1943,N_796,N_392);
or U1944 (N_1944,N_419,N_159);
nor U1945 (N_1945,N_734,N_1);
nor U1946 (N_1946,N_865,N_522);
nand U1947 (N_1947,N_998,N_2);
and U1948 (N_1948,N_911,N_285);
and U1949 (N_1949,N_908,N_921);
nand U1950 (N_1950,N_519,N_510);
and U1951 (N_1951,N_360,N_881);
or U1952 (N_1952,N_108,N_291);
or U1953 (N_1953,N_851,N_45);
nor U1954 (N_1954,N_797,N_745);
nor U1955 (N_1955,N_359,N_279);
nand U1956 (N_1956,N_431,N_320);
nor U1957 (N_1957,N_584,N_738);
and U1958 (N_1958,N_946,N_299);
nor U1959 (N_1959,N_820,N_742);
nor U1960 (N_1960,N_461,N_27);
or U1961 (N_1961,N_355,N_216);
or U1962 (N_1962,N_448,N_467);
and U1963 (N_1963,N_122,N_936);
and U1964 (N_1964,N_152,N_167);
xor U1965 (N_1965,N_277,N_480);
and U1966 (N_1966,N_336,N_586);
and U1967 (N_1967,N_417,N_349);
and U1968 (N_1968,N_504,N_877);
nor U1969 (N_1969,N_774,N_685);
nor U1970 (N_1970,N_949,N_632);
nand U1971 (N_1971,N_249,N_806);
or U1972 (N_1972,N_429,N_111);
and U1973 (N_1973,N_271,N_785);
nor U1974 (N_1974,N_902,N_642);
nor U1975 (N_1975,N_138,N_600);
nand U1976 (N_1976,N_258,N_640);
or U1977 (N_1977,N_41,N_416);
and U1978 (N_1978,N_763,N_915);
and U1979 (N_1979,N_132,N_97);
nor U1980 (N_1980,N_753,N_212);
or U1981 (N_1981,N_542,N_450);
nor U1982 (N_1982,N_412,N_872);
and U1983 (N_1983,N_759,N_496);
or U1984 (N_1984,N_881,N_517);
and U1985 (N_1985,N_944,N_588);
and U1986 (N_1986,N_373,N_699);
nor U1987 (N_1987,N_46,N_910);
or U1988 (N_1988,N_917,N_616);
nand U1989 (N_1989,N_265,N_76);
nand U1990 (N_1990,N_66,N_481);
or U1991 (N_1991,N_450,N_469);
nand U1992 (N_1992,N_30,N_873);
xor U1993 (N_1993,N_982,N_784);
or U1994 (N_1994,N_38,N_515);
and U1995 (N_1995,N_735,N_371);
nand U1996 (N_1996,N_853,N_935);
nand U1997 (N_1997,N_692,N_537);
nand U1998 (N_1998,N_242,N_963);
nor U1999 (N_1999,N_885,N_544);
nor U2000 (N_2000,N_1761,N_1521);
and U2001 (N_2001,N_1211,N_1257);
nand U2002 (N_2002,N_1194,N_1205);
and U2003 (N_2003,N_1250,N_1534);
nor U2004 (N_2004,N_1291,N_1807);
nor U2005 (N_2005,N_1216,N_1861);
and U2006 (N_2006,N_1511,N_1971);
nand U2007 (N_2007,N_1667,N_1057);
and U2008 (N_2008,N_1497,N_1054);
or U2009 (N_2009,N_1372,N_1819);
nor U2010 (N_2010,N_1731,N_1662);
nor U2011 (N_2011,N_1188,N_1682);
nor U2012 (N_2012,N_1859,N_1849);
or U2013 (N_2013,N_1325,N_1994);
or U2014 (N_2014,N_1101,N_1953);
nor U2015 (N_2015,N_1890,N_1378);
or U2016 (N_2016,N_1705,N_1093);
or U2017 (N_2017,N_1597,N_1998);
or U2018 (N_2018,N_1190,N_1307);
or U2019 (N_2019,N_1400,N_1494);
nor U2020 (N_2020,N_1946,N_1388);
nor U2021 (N_2021,N_1742,N_1184);
or U2022 (N_2022,N_1229,N_1270);
nand U2023 (N_2023,N_1727,N_1745);
or U2024 (N_2024,N_1002,N_1919);
nand U2025 (N_2025,N_1676,N_1517);
nand U2026 (N_2026,N_1564,N_1814);
nand U2027 (N_2027,N_1384,N_1300);
and U2028 (N_2028,N_1851,N_1646);
nor U2029 (N_2029,N_1856,N_1656);
or U2030 (N_2030,N_1373,N_1556);
and U2031 (N_2031,N_1421,N_1450);
xnor U2032 (N_2032,N_1935,N_1603);
or U2033 (N_2033,N_1828,N_1830);
nor U2034 (N_2034,N_1850,N_1287);
nor U2035 (N_2035,N_1920,N_1255);
or U2036 (N_2036,N_1329,N_1258);
nor U2037 (N_2037,N_1275,N_1272);
or U2038 (N_2038,N_1724,N_1875);
and U2039 (N_2039,N_1631,N_1460);
nand U2040 (N_2040,N_1702,N_1126);
nor U2041 (N_2041,N_1066,N_1422);
xnor U2042 (N_2042,N_1672,N_1958);
nor U2043 (N_2043,N_1256,N_1296);
nor U2044 (N_2044,N_1537,N_1813);
xor U2045 (N_2045,N_1170,N_1472);
or U2046 (N_2046,N_1763,N_1728);
xor U2047 (N_2047,N_1929,N_1623);
nor U2048 (N_2048,N_1246,N_1453);
nand U2049 (N_2049,N_1000,N_1114);
nor U2050 (N_2050,N_1654,N_1166);
nor U2051 (N_2051,N_1367,N_1065);
nand U2052 (N_2052,N_1579,N_1226);
and U2053 (N_2053,N_1122,N_1345);
and U2054 (N_2054,N_1698,N_1019);
and U2055 (N_2055,N_1435,N_1303);
nand U2056 (N_2056,N_1679,N_1050);
nand U2057 (N_2057,N_1827,N_1797);
nand U2058 (N_2058,N_1868,N_1401);
or U2059 (N_2059,N_1286,N_1945);
or U2060 (N_2060,N_1034,N_1778);
xor U2061 (N_2061,N_1925,N_1684);
or U2062 (N_2062,N_1196,N_1173);
xor U2063 (N_2063,N_1559,N_1581);
nand U2064 (N_2064,N_1590,N_1112);
nor U2065 (N_2065,N_1722,N_1536);
and U2066 (N_2066,N_1647,N_1014);
nor U2067 (N_2067,N_1876,N_1833);
or U2068 (N_2068,N_1532,N_1940);
or U2069 (N_2069,N_1447,N_1897);
and U2070 (N_2070,N_1762,N_1455);
and U2071 (N_2071,N_1267,N_1094);
nand U2072 (N_2072,N_1750,N_1108);
xnor U2073 (N_2073,N_1706,N_1338);
or U2074 (N_2074,N_1515,N_1825);
nand U2075 (N_2075,N_1891,N_1733);
nand U2076 (N_2076,N_1200,N_1747);
and U2077 (N_2077,N_1448,N_1634);
or U2078 (N_2078,N_1549,N_1848);
or U2079 (N_2079,N_1077,N_1509);
xor U2080 (N_2080,N_1424,N_1941);
xor U2081 (N_2081,N_1955,N_1412);
nand U2082 (N_2082,N_1148,N_1817);
or U2083 (N_2083,N_1957,N_1324);
xnor U2084 (N_2084,N_1089,N_1587);
or U2085 (N_2085,N_1279,N_1409);
or U2086 (N_2086,N_1784,N_1067);
nand U2087 (N_2087,N_1803,N_1991);
or U2088 (N_2088,N_1349,N_1209);
nor U2089 (N_2089,N_1666,N_1873);
nand U2090 (N_2090,N_1723,N_1304);
nor U2091 (N_2091,N_1550,N_1467);
nor U2092 (N_2092,N_1443,N_1415);
nand U2093 (N_2093,N_1159,N_1691);
or U2094 (N_2094,N_1197,N_1042);
xor U2095 (N_2095,N_1525,N_1137);
nor U2096 (N_2096,N_1740,N_1210);
nand U2097 (N_2097,N_1181,N_1264);
or U2098 (N_2098,N_1241,N_1960);
nand U2099 (N_2099,N_1283,N_1468);
or U2100 (N_2100,N_1265,N_1852);
nor U2101 (N_2101,N_1117,N_1076);
nor U2102 (N_2102,N_1222,N_1075);
or U2103 (N_2103,N_1800,N_1083);
or U2104 (N_2104,N_1228,N_1410);
nand U2105 (N_2105,N_1193,N_1961);
or U2106 (N_2106,N_1127,N_1360);
and U2107 (N_2107,N_1463,N_1328);
nand U2108 (N_2108,N_1548,N_1572);
and U2109 (N_2109,N_1346,N_1554);
or U2110 (N_2110,N_1037,N_1038);
xnor U2111 (N_2111,N_1701,N_1476);
nand U2112 (N_2112,N_1175,N_1495);
and U2113 (N_2113,N_1821,N_1547);
nor U2114 (N_2114,N_1382,N_1700);
or U2115 (N_2115,N_1996,N_1978);
xnor U2116 (N_2116,N_1914,N_1072);
nor U2117 (N_2117,N_1674,N_1938);
and U2118 (N_2118,N_1474,N_1029);
or U2119 (N_2119,N_1759,N_1893);
nand U2120 (N_2120,N_1681,N_1119);
or U2121 (N_2121,N_1915,N_1863);
nand U2122 (N_2122,N_1316,N_1074);
or U2123 (N_2123,N_1504,N_1992);
nand U2124 (N_2124,N_1574,N_1614);
nor U2125 (N_2125,N_1744,N_1951);
nor U2126 (N_2126,N_1179,N_1232);
nor U2127 (N_2127,N_1737,N_1144);
nand U2128 (N_2128,N_1632,N_1273);
nand U2129 (N_2129,N_1295,N_1933);
nor U2130 (N_2130,N_1526,N_1792);
or U2131 (N_2131,N_1573,N_1353);
nand U2132 (N_2132,N_1952,N_1168);
nand U2133 (N_2133,N_1244,N_1398);
nor U2134 (N_2134,N_1558,N_1452);
nand U2135 (N_2135,N_1140,N_1428);
and U2136 (N_2136,N_1707,N_1294);
or U2137 (N_2137,N_1182,N_1206);
xnor U2138 (N_2138,N_1437,N_1386);
or U2139 (N_2139,N_1982,N_1418);
and U2140 (N_2140,N_1508,N_1326);
and U2141 (N_2141,N_1981,N_1688);
or U2142 (N_2142,N_1910,N_1266);
nor U2143 (N_2143,N_1485,N_1628);
nor U2144 (N_2144,N_1299,N_1165);
nand U2145 (N_2145,N_1489,N_1238);
or U2146 (N_2146,N_1816,N_1055);
and U2147 (N_2147,N_1610,N_1236);
nor U2148 (N_2148,N_1039,N_1823);
or U2149 (N_2149,N_1520,N_1125);
nor U2150 (N_2150,N_1393,N_1802);
or U2151 (N_2151,N_1649,N_1527);
nor U2152 (N_2152,N_1411,N_1732);
nor U2153 (N_2153,N_1913,N_1247);
xor U2154 (N_2154,N_1675,N_1027);
nand U2155 (N_2155,N_1845,N_1313);
xnor U2156 (N_2156,N_1260,N_1683);
and U2157 (N_2157,N_1909,N_1673);
or U2158 (N_2158,N_1539,N_1482);
nand U2159 (N_2159,N_1496,N_1098);
and U2160 (N_2160,N_1645,N_1446);
nand U2161 (N_2161,N_1668,N_1374);
nor U2162 (N_2162,N_1486,N_1726);
nor U2163 (N_2163,N_1630,N_1658);
and U2164 (N_2164,N_1595,N_1561);
nor U2165 (N_2165,N_1060,N_1358);
nand U2166 (N_2166,N_1626,N_1350);
or U2167 (N_2167,N_1967,N_1589);
xnor U2168 (N_2168,N_1853,N_1369);
or U2169 (N_2169,N_1231,N_1102);
nand U2170 (N_2170,N_1806,N_1020);
nor U2171 (N_2171,N_1187,N_1220);
xnor U2172 (N_2172,N_1147,N_1641);
xnor U2173 (N_2173,N_1237,N_1461);
and U2174 (N_2174,N_1135,N_1867);
and U2175 (N_2175,N_1576,N_1070);
xnor U2176 (N_2176,N_1633,N_1396);
nor U2177 (N_2177,N_1528,N_1756);
nand U2178 (N_2178,N_1134,N_1540);
or U2179 (N_2179,N_1301,N_1543);
nand U2180 (N_2180,N_1986,N_1051);
nand U2181 (N_2181,N_1145,N_1669);
nand U2182 (N_2182,N_1276,N_1846);
nand U2183 (N_2183,N_1354,N_1973);
and U2184 (N_2184,N_1282,N_1622);
nand U2185 (N_2185,N_1696,N_1908);
xor U2186 (N_2186,N_1703,N_1870);
xor U2187 (N_2187,N_1319,N_1627);
nand U2188 (N_2188,N_1047,N_1289);
and U2189 (N_2189,N_1298,N_1904);
or U2190 (N_2190,N_1591,N_1151);
nand U2191 (N_2191,N_1586,N_1417);
nor U2192 (N_2192,N_1028,N_1164);
nor U2193 (N_2193,N_1379,N_1001);
xor U2194 (N_2194,N_1605,N_1062);
xnor U2195 (N_2195,N_1330,N_1993);
or U2196 (N_2196,N_1715,N_1710);
nor U2197 (N_2197,N_1502,N_1071);
and U2198 (N_2198,N_1887,N_1189);
xor U2199 (N_2199,N_1533,N_1243);
nor U2200 (N_2200,N_1449,N_1397);
nand U2201 (N_2201,N_1871,N_1746);
nand U2202 (N_2202,N_1522,N_1213);
nand U2203 (N_2203,N_1760,N_1240);
or U2204 (N_2204,N_1619,N_1003);
or U2205 (N_2205,N_1033,N_1729);
nand U2206 (N_2206,N_1513,N_1245);
nor U2207 (N_2207,N_1161,N_1567);
nand U2208 (N_2208,N_1493,N_1847);
nor U2209 (N_2209,N_1713,N_1120);
nor U2210 (N_2210,N_1708,N_1481);
or U2211 (N_2211,N_1575,N_1963);
or U2212 (N_2212,N_1405,N_1092);
nor U2213 (N_2213,N_1433,N_1831);
nand U2214 (N_2214,N_1392,N_1201);
nand U2215 (N_2215,N_1928,N_1233);
and U2216 (N_2216,N_1560,N_1334);
nand U2217 (N_2217,N_1544,N_1441);
nand U2218 (N_2218,N_1898,N_1340);
nand U2219 (N_2219,N_1999,N_1894);
and U2220 (N_2220,N_1880,N_1796);
and U2221 (N_2221,N_1812,N_1478);
and U2222 (N_2222,N_1408,N_1390);
nor U2223 (N_2223,N_1529,N_1907);
and U2224 (N_2224,N_1389,N_1611);
nor U2225 (N_2225,N_1970,N_1090);
nand U2226 (N_2226,N_1288,N_1477);
nor U2227 (N_2227,N_1322,N_1139);
xor U2228 (N_2228,N_1862,N_1921);
nor U2229 (N_2229,N_1600,N_1416);
nand U2230 (N_2230,N_1557,N_1583);
xor U2231 (N_2231,N_1017,N_1592);
or U2232 (N_2232,N_1059,N_1180);
nand U2233 (N_2233,N_1458,N_1758);
or U2234 (N_2234,N_1342,N_1535);
nor U2235 (N_2235,N_1835,N_1638);
or U2236 (N_2236,N_1361,N_1088);
nor U2237 (N_2237,N_1568,N_1655);
nor U2238 (N_2238,N_1129,N_1053);
and U2239 (N_2239,N_1944,N_1121);
xnor U2240 (N_2240,N_1826,N_1290);
or U2241 (N_2241,N_1026,N_1766);
nor U2242 (N_2242,N_1271,N_1484);
nand U2243 (N_2243,N_1082,N_1230);
xnor U2244 (N_2244,N_1618,N_1588);
nor U2245 (N_2245,N_1906,N_1555);
nor U2246 (N_2246,N_1878,N_1212);
nand U2247 (N_2247,N_1006,N_1671);
xor U2248 (N_2248,N_1031,N_1106);
nor U2249 (N_2249,N_1172,N_1776);
and U2250 (N_2250,N_1874,N_1900);
or U2251 (N_2251,N_1444,N_1507);
and U2252 (N_2252,N_1843,N_1695);
or U2253 (N_2253,N_1749,N_1007);
xor U2254 (N_2254,N_1096,N_1785);
and U2255 (N_2255,N_1219,N_1036);
nand U2256 (N_2256,N_1406,N_1602);
xor U2257 (N_2257,N_1709,N_1984);
nand U2258 (N_2258,N_1451,N_1578);
nor U2259 (N_2259,N_1637,N_1505);
or U2260 (N_2260,N_1629,N_1297);
or U2261 (N_2261,N_1839,N_1068);
xnor U2262 (N_2262,N_1105,N_1764);
nor U2263 (N_2263,N_1162,N_1500);
nor U2264 (N_2264,N_1310,N_1085);
nand U2265 (N_2265,N_1217,N_1202);
nand U2266 (N_2266,N_1498,N_1199);
and U2267 (N_2267,N_1949,N_1399);
and U2268 (N_2268,N_1593,N_1010);
and U2269 (N_2269,N_1541,N_1652);
nor U2270 (N_2270,N_1154,N_1438);
nor U2271 (N_2271,N_1021,N_1782);
nand U2272 (N_2272,N_1768,N_1829);
and U2273 (N_2273,N_1538,N_1571);
and U2274 (N_2274,N_1371,N_1751);
and U2275 (N_2275,N_1043,N_1487);
nor U2276 (N_2276,N_1609,N_1832);
nor U2277 (N_2277,N_1881,N_1087);
nand U2278 (N_2278,N_1809,N_1918);
nand U2279 (N_2279,N_1158,N_1292);
nor U2280 (N_2280,N_1834,N_1128);
and U2281 (N_2281,N_1284,N_1176);
nand U2282 (N_2282,N_1153,N_1110);
nand U2283 (N_2283,N_1381,N_1368);
nor U2284 (N_2284,N_1058,N_1714);
nor U2285 (N_2285,N_1439,N_1254);
nand U2286 (N_2286,N_1136,N_1518);
nand U2287 (N_2287,N_1394,N_1252);
nor U2288 (N_2288,N_1670,N_1563);
nor U2289 (N_2289,N_1488,N_1142);
nor U2290 (N_2290,N_1312,N_1677);
or U2291 (N_2291,N_1351,N_1721);
or U2292 (N_2292,N_1889,N_1430);
and U2293 (N_2293,N_1968,N_1069);
nand U2294 (N_2294,N_1514,N_1403);
and U2295 (N_2295,N_1642,N_1734);
and U2296 (N_2296,N_1765,N_1171);
nor U2297 (N_2297,N_1787,N_1916);
or U2298 (N_2298,N_1789,N_1962);
and U2299 (N_2299,N_1318,N_1979);
or U2300 (N_2300,N_1895,N_1743);
xnor U2301 (N_2301,N_1280,N_1431);
nand U2302 (N_2302,N_1336,N_1757);
nor U2303 (N_2303,N_1391,N_1794);
or U2304 (N_2304,N_1262,N_1009);
xor U2305 (N_2305,N_1208,N_1344);
or U2306 (N_2306,N_1407,N_1738);
and U2307 (N_2307,N_1860,N_1869);
nor U2308 (N_2308,N_1224,N_1805);
and U2309 (N_2309,N_1490,N_1167);
and U2310 (N_2310,N_1902,N_1857);
or U2311 (N_2311,N_1073,N_1133);
nor U2312 (N_2312,N_1899,N_1598);
and U2313 (N_2313,N_1327,N_1820);
and U2314 (N_2314,N_1506,N_1005);
xnor U2315 (N_2315,N_1269,N_1183);
xnor U2316 (N_2316,N_1584,N_1221);
or U2317 (N_2317,N_1699,N_1364);
and U2318 (N_2318,N_1285,N_1132);
xor U2319 (N_2319,N_1169,N_1333);
nand U2320 (N_2320,N_1281,N_1775);
nand U2321 (N_2321,N_1442,N_1599);
and U2322 (N_2322,N_1056,N_1720);
or U2323 (N_2323,N_1531,N_1932);
nand U2324 (N_2324,N_1604,N_1818);
nand U2325 (N_2325,N_1109,N_1864);
xor U2326 (N_2326,N_1788,N_1657);
nand U2327 (N_2327,N_1694,N_1606);
nor U2328 (N_2328,N_1178,N_1046);
or U2329 (N_2329,N_1811,N_1516);
nand U2330 (N_2330,N_1032,N_1492);
or U2331 (N_2331,N_1022,N_1362);
and U2332 (N_2332,N_1964,N_1911);
nor U2333 (N_2333,N_1987,N_1580);
and U2334 (N_2334,N_1317,N_1064);
nand U2335 (N_2335,N_1711,N_1624);
nor U2336 (N_2336,N_1214,N_1608);
xor U2337 (N_2337,N_1357,N_1052);
nand U2338 (N_2338,N_1123,N_1239);
xnor U2339 (N_2339,N_1989,N_1473);
or U2340 (N_2340,N_1783,N_1427);
or U2341 (N_2341,N_1542,N_1988);
nor U2342 (N_2342,N_1983,N_1607);
nor U2343 (N_2343,N_1261,N_1293);
or U2344 (N_2344,N_1791,N_1277);
nand U2345 (N_2345,N_1152,N_1773);
xnor U2346 (N_2346,N_1717,N_1736);
nor U2347 (N_2347,N_1616,N_1966);
or U2348 (N_2348,N_1462,N_1767);
or U2349 (N_2349,N_1937,N_1546);
xnor U2350 (N_2350,N_1844,N_1772);
and U2351 (N_2351,N_1314,N_1824);
or U2352 (N_2352,N_1225,N_1355);
or U2353 (N_2353,N_1660,N_1565);
nor U2354 (N_2354,N_1552,N_1095);
xor U2355 (N_2355,N_1483,N_1769);
xor U2356 (N_2356,N_1923,N_1321);
or U2357 (N_2357,N_1086,N_1530);
nand U2358 (N_2358,N_1480,N_1615);
or U2359 (N_2359,N_1420,N_1582);
nor U2360 (N_2360,N_1259,N_1939);
or U2361 (N_2361,N_1815,N_1786);
or U2362 (N_2362,N_1922,N_1115);
xor U2363 (N_2363,N_1030,N_1471);
nor U2364 (N_2364,N_1934,N_1730);
nand U2365 (N_2365,N_1613,N_1084);
and U2366 (N_2366,N_1780,N_1013);
nand U2367 (N_2367,N_1302,N_1663);
nor U2368 (N_2368,N_1930,N_1570);
nor U2369 (N_2369,N_1440,N_1838);
or U2370 (N_2370,N_1836,N_1063);
nand U2371 (N_2371,N_1686,N_1207);
and U2372 (N_2372,N_1491,N_1997);
nand U2373 (N_2373,N_1693,N_1793);
nand U2374 (N_2374,N_1004,N_1917);
or U2375 (N_2375,N_1882,N_1596);
nor U2376 (N_2376,N_1061,N_1195);
nand U2377 (N_2377,N_1927,N_1204);
nor U2378 (N_2378,N_1690,N_1104);
nand U2379 (N_2379,N_1174,N_1687);
nand U2380 (N_2380,N_1545,N_1425);
nand U2381 (N_2381,N_1305,N_1116);
nand U2382 (N_2382,N_1323,N_1661);
or U2383 (N_2383,N_1113,N_1884);
or U2384 (N_2384,N_1841,N_1801);
nand U2385 (N_2385,N_1248,N_1359);
and U2386 (N_2386,N_1464,N_1886);
nand U2387 (N_2387,N_1370,N_1877);
nor U2388 (N_2388,N_1685,N_1948);
nand U2389 (N_2389,N_1770,N_1445);
nand U2390 (N_2390,N_1124,N_1936);
xnor U2391 (N_2391,N_1977,N_1377);
and U2392 (N_2392,N_1475,N_1192);
nand U2393 (N_2393,N_1643,N_1341);
nor U2394 (N_2394,N_1648,N_1423);
or U2395 (N_2395,N_1822,N_1779);
xnor U2396 (N_2396,N_1621,N_1650);
nor U2397 (N_2397,N_1015,N_1842);
nor U2398 (N_2398,N_1620,N_1956);
and U2399 (N_2399,N_1024,N_1249);
xor U2400 (N_2400,N_1888,N_1332);
or U2401 (N_2401,N_1959,N_1091);
and U2402 (N_2402,N_1146,N_1157);
nand U2403 (N_2403,N_1905,N_1739);
nand U2404 (N_2404,N_1885,N_1689);
xor U2405 (N_2405,N_1625,N_1653);
nand U2406 (N_2406,N_1429,N_1704);
nand U2407 (N_2407,N_1268,N_1459);
nand U2408 (N_2408,N_1659,N_1781);
nor U2409 (N_2409,N_1079,N_1748);
nand U2410 (N_2410,N_1138,N_1523);
nand U2411 (N_2411,N_1678,N_1426);
and U2412 (N_2412,N_1840,N_1111);
nor U2413 (N_2413,N_1078,N_1274);
nand U2414 (N_2414,N_1163,N_1156);
nor U2415 (N_2415,N_1311,N_1680);
or U2416 (N_2416,N_1718,N_1954);
or U2417 (N_2417,N_1617,N_1308);
and U2418 (N_2418,N_1735,N_1804);
nor U2419 (N_2419,N_1466,N_1218);
nor U2420 (N_2420,N_1866,N_1912);
nand U2421 (N_2421,N_1215,N_1456);
and U2422 (N_2422,N_1016,N_1810);
nor U2423 (N_2423,N_1501,N_1251);
nor U2424 (N_2424,N_1512,N_1253);
nand U2425 (N_2425,N_1242,N_1798);
nor U2426 (N_2426,N_1025,N_1436);
nand U2427 (N_2427,N_1223,N_1896);
or U2428 (N_2428,N_1434,N_1227);
nor U2429 (N_2429,N_1432,N_1012);
and U2430 (N_2430,N_1974,N_1049);
nand U2431 (N_2431,N_1040,N_1045);
nor U2432 (N_2432,N_1035,N_1865);
xnor U2433 (N_2433,N_1635,N_1018);
and U2434 (N_2434,N_1771,N_1931);
or U2435 (N_2435,N_1413,N_1081);
nand U2436 (N_2436,N_1376,N_1011);
and U2437 (N_2437,N_1777,N_1799);
and U2438 (N_2438,N_1404,N_1470);
nand U2439 (N_2439,N_1306,N_1665);
nor U2440 (N_2440,N_1048,N_1103);
or U2441 (N_2441,N_1808,N_1337);
nor U2442 (N_2442,N_1375,N_1185);
or U2443 (N_2443,N_1719,N_1524);
and U2444 (N_2444,N_1419,N_1395);
or U2445 (N_2445,N_1566,N_1562);
and U2446 (N_2446,N_1725,N_1837);
and U2447 (N_2447,N_1339,N_1234);
and U2448 (N_2448,N_1755,N_1995);
or U2449 (N_2449,N_1639,N_1479);
and U2450 (N_2450,N_1879,N_1741);
and U2451 (N_2451,N_1612,N_1872);
and U2452 (N_2452,N_1177,N_1186);
nor U2453 (N_2453,N_1363,N_1640);
and U2454 (N_2454,N_1569,N_1097);
nand U2455 (N_2455,N_1990,N_1414);
nor U2456 (N_2456,N_1601,N_1972);
nand U2457 (N_2457,N_1352,N_1644);
or U2458 (N_2458,N_1965,N_1585);
and U2459 (N_2459,N_1365,N_1969);
xor U2460 (N_2460,N_1383,N_1402);
or U2461 (N_2461,N_1883,N_1858);
and U2462 (N_2462,N_1141,N_1697);
nor U2463 (N_2463,N_1023,N_1278);
nor U2464 (N_2464,N_1712,N_1320);
nand U2465 (N_2465,N_1309,N_1754);
or U2466 (N_2466,N_1499,N_1790);
or U2467 (N_2467,N_1950,N_1465);
nor U2468 (N_2468,N_1980,N_1099);
and U2469 (N_2469,N_1903,N_1924);
xnor U2470 (N_2470,N_1753,N_1331);
and U2471 (N_2471,N_1107,N_1041);
and U2472 (N_2472,N_1553,N_1519);
and U2473 (N_2473,N_1457,N_1347);
xor U2474 (N_2474,N_1454,N_1348);
or U2475 (N_2475,N_1191,N_1795);
or U2476 (N_2476,N_1503,N_1080);
nand U2477 (N_2477,N_1130,N_1198);
nand U2478 (N_2478,N_1716,N_1356);
nor U2479 (N_2479,N_1118,N_1947);
nor U2480 (N_2480,N_1469,N_1366);
or U2481 (N_2481,N_1664,N_1976);
or U2482 (N_2482,N_1985,N_1577);
nor U2483 (N_2483,N_1387,N_1160);
xnor U2484 (N_2484,N_1551,N_1315);
xor U2485 (N_2485,N_1943,N_1235);
nand U2486 (N_2486,N_1942,N_1975);
and U2487 (N_2487,N_1510,N_1892);
and U2488 (N_2488,N_1143,N_1343);
or U2489 (N_2489,N_1155,N_1651);
and U2490 (N_2490,N_1044,N_1752);
and U2491 (N_2491,N_1203,N_1385);
nand U2492 (N_2492,N_1854,N_1100);
xor U2493 (N_2493,N_1926,N_1149);
nor U2494 (N_2494,N_1150,N_1131);
and U2495 (N_2495,N_1692,N_1774);
or U2496 (N_2496,N_1636,N_1263);
nor U2497 (N_2497,N_1335,N_1008);
xor U2498 (N_2498,N_1901,N_1855);
and U2499 (N_2499,N_1594,N_1380);
and U2500 (N_2500,N_1865,N_1605);
nand U2501 (N_2501,N_1793,N_1141);
nor U2502 (N_2502,N_1786,N_1468);
nand U2503 (N_2503,N_1196,N_1603);
and U2504 (N_2504,N_1580,N_1328);
nand U2505 (N_2505,N_1850,N_1532);
nand U2506 (N_2506,N_1683,N_1436);
nand U2507 (N_2507,N_1820,N_1705);
nor U2508 (N_2508,N_1181,N_1819);
or U2509 (N_2509,N_1507,N_1255);
and U2510 (N_2510,N_1824,N_1868);
and U2511 (N_2511,N_1403,N_1493);
nand U2512 (N_2512,N_1132,N_1438);
and U2513 (N_2513,N_1548,N_1827);
nand U2514 (N_2514,N_1773,N_1497);
and U2515 (N_2515,N_1663,N_1198);
and U2516 (N_2516,N_1616,N_1437);
and U2517 (N_2517,N_1081,N_1230);
xor U2518 (N_2518,N_1165,N_1977);
and U2519 (N_2519,N_1587,N_1235);
nand U2520 (N_2520,N_1654,N_1205);
nor U2521 (N_2521,N_1622,N_1026);
and U2522 (N_2522,N_1788,N_1894);
or U2523 (N_2523,N_1194,N_1193);
and U2524 (N_2524,N_1029,N_1957);
nand U2525 (N_2525,N_1858,N_1395);
nand U2526 (N_2526,N_1781,N_1050);
or U2527 (N_2527,N_1920,N_1108);
xor U2528 (N_2528,N_1106,N_1818);
or U2529 (N_2529,N_1076,N_1019);
nor U2530 (N_2530,N_1210,N_1513);
or U2531 (N_2531,N_1744,N_1047);
or U2532 (N_2532,N_1319,N_1614);
xor U2533 (N_2533,N_1046,N_1518);
and U2534 (N_2534,N_1090,N_1256);
nand U2535 (N_2535,N_1804,N_1590);
nor U2536 (N_2536,N_1023,N_1084);
or U2537 (N_2537,N_1509,N_1152);
or U2538 (N_2538,N_1097,N_1838);
and U2539 (N_2539,N_1641,N_1638);
xor U2540 (N_2540,N_1290,N_1884);
nor U2541 (N_2541,N_1548,N_1953);
or U2542 (N_2542,N_1798,N_1314);
xnor U2543 (N_2543,N_1736,N_1648);
or U2544 (N_2544,N_1949,N_1114);
xor U2545 (N_2545,N_1740,N_1123);
nor U2546 (N_2546,N_1796,N_1442);
and U2547 (N_2547,N_1048,N_1512);
and U2548 (N_2548,N_1411,N_1217);
xnor U2549 (N_2549,N_1230,N_1291);
and U2550 (N_2550,N_1343,N_1589);
nor U2551 (N_2551,N_1674,N_1773);
nand U2552 (N_2552,N_1893,N_1534);
or U2553 (N_2553,N_1008,N_1435);
nor U2554 (N_2554,N_1253,N_1810);
and U2555 (N_2555,N_1133,N_1545);
or U2556 (N_2556,N_1273,N_1865);
nor U2557 (N_2557,N_1861,N_1439);
or U2558 (N_2558,N_1211,N_1244);
or U2559 (N_2559,N_1457,N_1228);
nor U2560 (N_2560,N_1015,N_1159);
nor U2561 (N_2561,N_1068,N_1538);
and U2562 (N_2562,N_1361,N_1256);
nor U2563 (N_2563,N_1244,N_1245);
nand U2564 (N_2564,N_1073,N_1338);
xor U2565 (N_2565,N_1642,N_1580);
or U2566 (N_2566,N_1359,N_1529);
nand U2567 (N_2567,N_1103,N_1805);
nor U2568 (N_2568,N_1561,N_1329);
nand U2569 (N_2569,N_1781,N_1706);
xnor U2570 (N_2570,N_1148,N_1061);
nand U2571 (N_2571,N_1174,N_1293);
nor U2572 (N_2572,N_1317,N_1405);
and U2573 (N_2573,N_1010,N_1039);
and U2574 (N_2574,N_1281,N_1655);
and U2575 (N_2575,N_1078,N_1261);
or U2576 (N_2576,N_1794,N_1059);
and U2577 (N_2577,N_1639,N_1776);
nor U2578 (N_2578,N_1684,N_1076);
or U2579 (N_2579,N_1739,N_1263);
nand U2580 (N_2580,N_1048,N_1660);
nor U2581 (N_2581,N_1057,N_1221);
nand U2582 (N_2582,N_1983,N_1119);
nor U2583 (N_2583,N_1860,N_1421);
or U2584 (N_2584,N_1026,N_1568);
or U2585 (N_2585,N_1641,N_1876);
or U2586 (N_2586,N_1032,N_1075);
nor U2587 (N_2587,N_1217,N_1582);
or U2588 (N_2588,N_1079,N_1258);
nand U2589 (N_2589,N_1686,N_1593);
nor U2590 (N_2590,N_1425,N_1314);
or U2591 (N_2591,N_1034,N_1827);
and U2592 (N_2592,N_1284,N_1717);
nand U2593 (N_2593,N_1201,N_1474);
nor U2594 (N_2594,N_1457,N_1088);
nor U2595 (N_2595,N_1900,N_1635);
nor U2596 (N_2596,N_1218,N_1637);
or U2597 (N_2597,N_1581,N_1259);
and U2598 (N_2598,N_1390,N_1399);
nand U2599 (N_2599,N_1019,N_1378);
nand U2600 (N_2600,N_1961,N_1424);
nand U2601 (N_2601,N_1919,N_1875);
or U2602 (N_2602,N_1727,N_1329);
xnor U2603 (N_2603,N_1753,N_1440);
or U2604 (N_2604,N_1822,N_1834);
xnor U2605 (N_2605,N_1103,N_1517);
or U2606 (N_2606,N_1124,N_1707);
xnor U2607 (N_2607,N_1501,N_1247);
or U2608 (N_2608,N_1926,N_1035);
and U2609 (N_2609,N_1807,N_1580);
nor U2610 (N_2610,N_1508,N_1042);
nand U2611 (N_2611,N_1687,N_1389);
and U2612 (N_2612,N_1527,N_1742);
and U2613 (N_2613,N_1943,N_1178);
nor U2614 (N_2614,N_1339,N_1920);
nor U2615 (N_2615,N_1659,N_1628);
xnor U2616 (N_2616,N_1896,N_1911);
xnor U2617 (N_2617,N_1997,N_1887);
nand U2618 (N_2618,N_1914,N_1577);
nand U2619 (N_2619,N_1774,N_1366);
nand U2620 (N_2620,N_1698,N_1338);
and U2621 (N_2621,N_1617,N_1931);
xor U2622 (N_2622,N_1880,N_1837);
nor U2623 (N_2623,N_1549,N_1501);
or U2624 (N_2624,N_1308,N_1301);
xnor U2625 (N_2625,N_1852,N_1849);
xor U2626 (N_2626,N_1004,N_1400);
nor U2627 (N_2627,N_1625,N_1175);
xor U2628 (N_2628,N_1381,N_1017);
nand U2629 (N_2629,N_1510,N_1581);
or U2630 (N_2630,N_1944,N_1545);
and U2631 (N_2631,N_1714,N_1167);
xnor U2632 (N_2632,N_1530,N_1422);
nand U2633 (N_2633,N_1077,N_1689);
and U2634 (N_2634,N_1772,N_1571);
nand U2635 (N_2635,N_1540,N_1305);
and U2636 (N_2636,N_1373,N_1404);
xor U2637 (N_2637,N_1015,N_1388);
or U2638 (N_2638,N_1384,N_1205);
and U2639 (N_2639,N_1580,N_1667);
or U2640 (N_2640,N_1211,N_1709);
nand U2641 (N_2641,N_1319,N_1909);
and U2642 (N_2642,N_1944,N_1370);
or U2643 (N_2643,N_1286,N_1625);
nand U2644 (N_2644,N_1988,N_1442);
and U2645 (N_2645,N_1282,N_1947);
nor U2646 (N_2646,N_1464,N_1134);
nor U2647 (N_2647,N_1450,N_1373);
or U2648 (N_2648,N_1255,N_1900);
or U2649 (N_2649,N_1352,N_1754);
nand U2650 (N_2650,N_1824,N_1514);
nand U2651 (N_2651,N_1128,N_1872);
or U2652 (N_2652,N_1850,N_1200);
and U2653 (N_2653,N_1967,N_1200);
nor U2654 (N_2654,N_1052,N_1954);
nand U2655 (N_2655,N_1468,N_1186);
nand U2656 (N_2656,N_1954,N_1409);
and U2657 (N_2657,N_1331,N_1488);
or U2658 (N_2658,N_1172,N_1533);
nor U2659 (N_2659,N_1462,N_1060);
nand U2660 (N_2660,N_1770,N_1559);
nor U2661 (N_2661,N_1515,N_1881);
or U2662 (N_2662,N_1651,N_1096);
and U2663 (N_2663,N_1494,N_1523);
nor U2664 (N_2664,N_1994,N_1334);
nor U2665 (N_2665,N_1777,N_1341);
nor U2666 (N_2666,N_1367,N_1010);
nand U2667 (N_2667,N_1012,N_1653);
or U2668 (N_2668,N_1712,N_1775);
or U2669 (N_2669,N_1722,N_1171);
nand U2670 (N_2670,N_1506,N_1168);
or U2671 (N_2671,N_1120,N_1115);
or U2672 (N_2672,N_1784,N_1235);
and U2673 (N_2673,N_1295,N_1489);
nor U2674 (N_2674,N_1190,N_1906);
or U2675 (N_2675,N_1891,N_1453);
and U2676 (N_2676,N_1559,N_1207);
and U2677 (N_2677,N_1883,N_1124);
nand U2678 (N_2678,N_1257,N_1146);
nor U2679 (N_2679,N_1560,N_1322);
nor U2680 (N_2680,N_1072,N_1261);
and U2681 (N_2681,N_1339,N_1662);
or U2682 (N_2682,N_1444,N_1437);
and U2683 (N_2683,N_1443,N_1884);
and U2684 (N_2684,N_1012,N_1774);
and U2685 (N_2685,N_1902,N_1379);
nor U2686 (N_2686,N_1469,N_1835);
xnor U2687 (N_2687,N_1175,N_1517);
and U2688 (N_2688,N_1387,N_1865);
or U2689 (N_2689,N_1769,N_1775);
xnor U2690 (N_2690,N_1743,N_1156);
or U2691 (N_2691,N_1867,N_1188);
xnor U2692 (N_2692,N_1724,N_1561);
nor U2693 (N_2693,N_1862,N_1423);
nor U2694 (N_2694,N_1020,N_1660);
and U2695 (N_2695,N_1938,N_1300);
nor U2696 (N_2696,N_1938,N_1214);
nand U2697 (N_2697,N_1447,N_1482);
xnor U2698 (N_2698,N_1295,N_1622);
nand U2699 (N_2699,N_1021,N_1337);
or U2700 (N_2700,N_1824,N_1155);
or U2701 (N_2701,N_1514,N_1005);
and U2702 (N_2702,N_1635,N_1984);
or U2703 (N_2703,N_1048,N_1145);
and U2704 (N_2704,N_1990,N_1590);
or U2705 (N_2705,N_1231,N_1364);
and U2706 (N_2706,N_1234,N_1423);
nand U2707 (N_2707,N_1585,N_1525);
xor U2708 (N_2708,N_1869,N_1608);
or U2709 (N_2709,N_1033,N_1514);
xor U2710 (N_2710,N_1268,N_1316);
nor U2711 (N_2711,N_1921,N_1314);
nor U2712 (N_2712,N_1693,N_1047);
or U2713 (N_2713,N_1244,N_1482);
or U2714 (N_2714,N_1755,N_1381);
nand U2715 (N_2715,N_1996,N_1671);
and U2716 (N_2716,N_1449,N_1241);
or U2717 (N_2717,N_1902,N_1500);
nand U2718 (N_2718,N_1223,N_1593);
nor U2719 (N_2719,N_1815,N_1768);
nand U2720 (N_2720,N_1809,N_1787);
nor U2721 (N_2721,N_1536,N_1020);
and U2722 (N_2722,N_1492,N_1503);
and U2723 (N_2723,N_1275,N_1548);
nand U2724 (N_2724,N_1381,N_1418);
xor U2725 (N_2725,N_1117,N_1973);
or U2726 (N_2726,N_1915,N_1855);
and U2727 (N_2727,N_1807,N_1699);
and U2728 (N_2728,N_1364,N_1456);
nor U2729 (N_2729,N_1955,N_1499);
or U2730 (N_2730,N_1242,N_1331);
nand U2731 (N_2731,N_1357,N_1819);
and U2732 (N_2732,N_1047,N_1119);
nor U2733 (N_2733,N_1570,N_1328);
or U2734 (N_2734,N_1053,N_1446);
xnor U2735 (N_2735,N_1460,N_1792);
nor U2736 (N_2736,N_1581,N_1652);
xnor U2737 (N_2737,N_1544,N_1562);
nor U2738 (N_2738,N_1490,N_1332);
or U2739 (N_2739,N_1763,N_1218);
nand U2740 (N_2740,N_1410,N_1360);
nand U2741 (N_2741,N_1835,N_1699);
nor U2742 (N_2742,N_1647,N_1877);
nor U2743 (N_2743,N_1384,N_1991);
nor U2744 (N_2744,N_1657,N_1707);
nor U2745 (N_2745,N_1479,N_1750);
and U2746 (N_2746,N_1747,N_1426);
nand U2747 (N_2747,N_1716,N_1628);
or U2748 (N_2748,N_1124,N_1443);
xor U2749 (N_2749,N_1750,N_1001);
nor U2750 (N_2750,N_1681,N_1751);
or U2751 (N_2751,N_1105,N_1621);
and U2752 (N_2752,N_1314,N_1743);
nor U2753 (N_2753,N_1412,N_1387);
nor U2754 (N_2754,N_1394,N_1611);
or U2755 (N_2755,N_1609,N_1554);
xor U2756 (N_2756,N_1397,N_1332);
and U2757 (N_2757,N_1098,N_1222);
nor U2758 (N_2758,N_1530,N_1309);
or U2759 (N_2759,N_1908,N_1933);
nor U2760 (N_2760,N_1914,N_1204);
nor U2761 (N_2761,N_1938,N_1565);
and U2762 (N_2762,N_1352,N_1202);
or U2763 (N_2763,N_1846,N_1375);
or U2764 (N_2764,N_1377,N_1861);
and U2765 (N_2765,N_1054,N_1651);
nor U2766 (N_2766,N_1379,N_1614);
and U2767 (N_2767,N_1493,N_1228);
nand U2768 (N_2768,N_1857,N_1285);
nor U2769 (N_2769,N_1421,N_1521);
nor U2770 (N_2770,N_1861,N_1037);
nand U2771 (N_2771,N_1241,N_1976);
nand U2772 (N_2772,N_1200,N_1354);
nor U2773 (N_2773,N_1610,N_1883);
nor U2774 (N_2774,N_1174,N_1697);
xnor U2775 (N_2775,N_1185,N_1898);
and U2776 (N_2776,N_1467,N_1414);
nor U2777 (N_2777,N_1210,N_1348);
or U2778 (N_2778,N_1182,N_1632);
nand U2779 (N_2779,N_1225,N_1251);
nor U2780 (N_2780,N_1236,N_1269);
nor U2781 (N_2781,N_1164,N_1086);
nand U2782 (N_2782,N_1609,N_1272);
nand U2783 (N_2783,N_1597,N_1095);
xnor U2784 (N_2784,N_1342,N_1250);
nand U2785 (N_2785,N_1419,N_1087);
nand U2786 (N_2786,N_1505,N_1364);
and U2787 (N_2787,N_1950,N_1602);
nor U2788 (N_2788,N_1638,N_1495);
and U2789 (N_2789,N_1921,N_1190);
or U2790 (N_2790,N_1611,N_1665);
and U2791 (N_2791,N_1947,N_1310);
and U2792 (N_2792,N_1597,N_1002);
nor U2793 (N_2793,N_1763,N_1914);
and U2794 (N_2794,N_1123,N_1444);
nand U2795 (N_2795,N_1714,N_1405);
or U2796 (N_2796,N_1970,N_1385);
nand U2797 (N_2797,N_1639,N_1131);
nand U2798 (N_2798,N_1083,N_1395);
nor U2799 (N_2799,N_1000,N_1310);
or U2800 (N_2800,N_1170,N_1813);
or U2801 (N_2801,N_1578,N_1704);
or U2802 (N_2802,N_1406,N_1799);
nand U2803 (N_2803,N_1065,N_1940);
and U2804 (N_2804,N_1759,N_1772);
or U2805 (N_2805,N_1822,N_1197);
xnor U2806 (N_2806,N_1602,N_1943);
nor U2807 (N_2807,N_1364,N_1835);
nand U2808 (N_2808,N_1242,N_1900);
nor U2809 (N_2809,N_1408,N_1840);
nand U2810 (N_2810,N_1990,N_1578);
nand U2811 (N_2811,N_1199,N_1149);
nand U2812 (N_2812,N_1088,N_1718);
nor U2813 (N_2813,N_1876,N_1312);
nand U2814 (N_2814,N_1063,N_1234);
nor U2815 (N_2815,N_1897,N_1113);
nand U2816 (N_2816,N_1921,N_1760);
or U2817 (N_2817,N_1160,N_1546);
nand U2818 (N_2818,N_1670,N_1586);
nor U2819 (N_2819,N_1474,N_1572);
or U2820 (N_2820,N_1678,N_1775);
or U2821 (N_2821,N_1824,N_1798);
and U2822 (N_2822,N_1136,N_1251);
and U2823 (N_2823,N_1603,N_1929);
nand U2824 (N_2824,N_1134,N_1991);
nand U2825 (N_2825,N_1785,N_1451);
and U2826 (N_2826,N_1353,N_1400);
nor U2827 (N_2827,N_1347,N_1283);
and U2828 (N_2828,N_1550,N_1025);
or U2829 (N_2829,N_1201,N_1685);
nor U2830 (N_2830,N_1389,N_1195);
and U2831 (N_2831,N_1154,N_1379);
and U2832 (N_2832,N_1291,N_1528);
and U2833 (N_2833,N_1352,N_1560);
nor U2834 (N_2834,N_1166,N_1815);
or U2835 (N_2835,N_1018,N_1179);
nor U2836 (N_2836,N_1538,N_1329);
and U2837 (N_2837,N_1933,N_1810);
xor U2838 (N_2838,N_1618,N_1982);
nor U2839 (N_2839,N_1952,N_1626);
nor U2840 (N_2840,N_1132,N_1995);
or U2841 (N_2841,N_1174,N_1242);
or U2842 (N_2842,N_1288,N_1009);
or U2843 (N_2843,N_1229,N_1115);
or U2844 (N_2844,N_1121,N_1447);
and U2845 (N_2845,N_1204,N_1549);
nor U2846 (N_2846,N_1643,N_1023);
or U2847 (N_2847,N_1120,N_1368);
nand U2848 (N_2848,N_1578,N_1787);
xnor U2849 (N_2849,N_1299,N_1096);
nand U2850 (N_2850,N_1519,N_1312);
nand U2851 (N_2851,N_1281,N_1080);
nor U2852 (N_2852,N_1895,N_1002);
nand U2853 (N_2853,N_1030,N_1115);
xor U2854 (N_2854,N_1927,N_1961);
nand U2855 (N_2855,N_1895,N_1622);
and U2856 (N_2856,N_1473,N_1321);
nand U2857 (N_2857,N_1809,N_1474);
and U2858 (N_2858,N_1457,N_1318);
and U2859 (N_2859,N_1069,N_1983);
and U2860 (N_2860,N_1611,N_1303);
xor U2861 (N_2861,N_1031,N_1953);
nor U2862 (N_2862,N_1232,N_1307);
or U2863 (N_2863,N_1398,N_1001);
xnor U2864 (N_2864,N_1340,N_1256);
and U2865 (N_2865,N_1702,N_1517);
xor U2866 (N_2866,N_1199,N_1595);
and U2867 (N_2867,N_1465,N_1159);
and U2868 (N_2868,N_1110,N_1843);
xnor U2869 (N_2869,N_1367,N_1784);
nor U2870 (N_2870,N_1800,N_1943);
nand U2871 (N_2871,N_1785,N_1534);
nand U2872 (N_2872,N_1996,N_1454);
nand U2873 (N_2873,N_1666,N_1738);
or U2874 (N_2874,N_1922,N_1105);
and U2875 (N_2875,N_1020,N_1468);
and U2876 (N_2876,N_1853,N_1772);
nand U2877 (N_2877,N_1125,N_1072);
and U2878 (N_2878,N_1248,N_1092);
and U2879 (N_2879,N_1666,N_1572);
nor U2880 (N_2880,N_1660,N_1972);
and U2881 (N_2881,N_1168,N_1229);
nor U2882 (N_2882,N_1751,N_1913);
nand U2883 (N_2883,N_1402,N_1399);
or U2884 (N_2884,N_1699,N_1329);
or U2885 (N_2885,N_1634,N_1150);
and U2886 (N_2886,N_1424,N_1973);
xnor U2887 (N_2887,N_1760,N_1245);
xor U2888 (N_2888,N_1258,N_1180);
nor U2889 (N_2889,N_1612,N_1829);
or U2890 (N_2890,N_1519,N_1071);
xnor U2891 (N_2891,N_1891,N_1734);
nand U2892 (N_2892,N_1913,N_1603);
nor U2893 (N_2893,N_1498,N_1578);
or U2894 (N_2894,N_1099,N_1674);
or U2895 (N_2895,N_1120,N_1255);
nand U2896 (N_2896,N_1340,N_1325);
nor U2897 (N_2897,N_1893,N_1165);
nor U2898 (N_2898,N_1516,N_1373);
and U2899 (N_2899,N_1325,N_1936);
and U2900 (N_2900,N_1899,N_1474);
nand U2901 (N_2901,N_1605,N_1290);
nand U2902 (N_2902,N_1073,N_1632);
nand U2903 (N_2903,N_1183,N_1985);
and U2904 (N_2904,N_1835,N_1894);
and U2905 (N_2905,N_1342,N_1751);
nand U2906 (N_2906,N_1350,N_1005);
and U2907 (N_2907,N_1966,N_1238);
nand U2908 (N_2908,N_1641,N_1497);
or U2909 (N_2909,N_1700,N_1238);
or U2910 (N_2910,N_1066,N_1141);
nor U2911 (N_2911,N_1880,N_1400);
xor U2912 (N_2912,N_1650,N_1857);
nor U2913 (N_2913,N_1986,N_1868);
nand U2914 (N_2914,N_1810,N_1268);
nor U2915 (N_2915,N_1301,N_1871);
nor U2916 (N_2916,N_1444,N_1149);
or U2917 (N_2917,N_1409,N_1998);
nand U2918 (N_2918,N_1123,N_1545);
nor U2919 (N_2919,N_1766,N_1755);
and U2920 (N_2920,N_1905,N_1080);
or U2921 (N_2921,N_1740,N_1782);
and U2922 (N_2922,N_1790,N_1519);
and U2923 (N_2923,N_1263,N_1932);
and U2924 (N_2924,N_1833,N_1912);
nor U2925 (N_2925,N_1223,N_1097);
and U2926 (N_2926,N_1411,N_1395);
and U2927 (N_2927,N_1301,N_1833);
nor U2928 (N_2928,N_1147,N_1285);
nand U2929 (N_2929,N_1502,N_1647);
or U2930 (N_2930,N_1866,N_1737);
and U2931 (N_2931,N_1422,N_1006);
nand U2932 (N_2932,N_1191,N_1818);
nand U2933 (N_2933,N_1693,N_1415);
or U2934 (N_2934,N_1722,N_1944);
xor U2935 (N_2935,N_1096,N_1788);
nor U2936 (N_2936,N_1640,N_1062);
nand U2937 (N_2937,N_1830,N_1053);
nor U2938 (N_2938,N_1032,N_1911);
nand U2939 (N_2939,N_1359,N_1879);
nor U2940 (N_2940,N_1809,N_1674);
or U2941 (N_2941,N_1714,N_1213);
and U2942 (N_2942,N_1776,N_1680);
nor U2943 (N_2943,N_1638,N_1425);
or U2944 (N_2944,N_1260,N_1164);
nand U2945 (N_2945,N_1603,N_1234);
nor U2946 (N_2946,N_1459,N_1230);
nand U2947 (N_2947,N_1700,N_1866);
and U2948 (N_2948,N_1485,N_1276);
and U2949 (N_2949,N_1737,N_1455);
nor U2950 (N_2950,N_1229,N_1262);
and U2951 (N_2951,N_1393,N_1640);
nor U2952 (N_2952,N_1604,N_1263);
or U2953 (N_2953,N_1261,N_1041);
or U2954 (N_2954,N_1549,N_1526);
nand U2955 (N_2955,N_1703,N_1728);
nor U2956 (N_2956,N_1845,N_1764);
nor U2957 (N_2957,N_1070,N_1478);
xnor U2958 (N_2958,N_1154,N_1215);
xnor U2959 (N_2959,N_1358,N_1725);
or U2960 (N_2960,N_1667,N_1184);
and U2961 (N_2961,N_1824,N_1342);
or U2962 (N_2962,N_1534,N_1444);
xnor U2963 (N_2963,N_1834,N_1923);
nor U2964 (N_2964,N_1386,N_1681);
and U2965 (N_2965,N_1713,N_1377);
xor U2966 (N_2966,N_1631,N_1026);
and U2967 (N_2967,N_1898,N_1069);
and U2968 (N_2968,N_1326,N_1631);
nand U2969 (N_2969,N_1482,N_1643);
and U2970 (N_2970,N_1948,N_1233);
nor U2971 (N_2971,N_1783,N_1370);
nand U2972 (N_2972,N_1563,N_1241);
or U2973 (N_2973,N_1367,N_1722);
xor U2974 (N_2974,N_1198,N_1723);
or U2975 (N_2975,N_1921,N_1295);
nor U2976 (N_2976,N_1317,N_1810);
nand U2977 (N_2977,N_1803,N_1983);
or U2978 (N_2978,N_1869,N_1261);
nand U2979 (N_2979,N_1628,N_1562);
and U2980 (N_2980,N_1539,N_1004);
nand U2981 (N_2981,N_1523,N_1298);
nand U2982 (N_2982,N_1831,N_1083);
nand U2983 (N_2983,N_1539,N_1083);
nand U2984 (N_2984,N_1742,N_1404);
xnor U2985 (N_2985,N_1827,N_1441);
nand U2986 (N_2986,N_1230,N_1151);
and U2987 (N_2987,N_1568,N_1145);
nand U2988 (N_2988,N_1326,N_1932);
or U2989 (N_2989,N_1692,N_1649);
nand U2990 (N_2990,N_1628,N_1583);
nor U2991 (N_2991,N_1563,N_1631);
and U2992 (N_2992,N_1205,N_1077);
or U2993 (N_2993,N_1566,N_1810);
xnor U2994 (N_2994,N_1598,N_1777);
nor U2995 (N_2995,N_1007,N_1964);
nor U2996 (N_2996,N_1192,N_1611);
nand U2997 (N_2997,N_1767,N_1220);
nand U2998 (N_2998,N_1168,N_1542);
or U2999 (N_2999,N_1885,N_1654);
nand UO_0 (O_0,N_2515,N_2417);
or UO_1 (O_1,N_2864,N_2918);
and UO_2 (O_2,N_2104,N_2057);
nand UO_3 (O_3,N_2976,N_2763);
nand UO_4 (O_4,N_2937,N_2135);
and UO_5 (O_5,N_2053,N_2382);
nand UO_6 (O_6,N_2919,N_2565);
and UO_7 (O_7,N_2481,N_2905);
or UO_8 (O_8,N_2795,N_2004);
and UO_9 (O_9,N_2492,N_2815);
nand UO_10 (O_10,N_2758,N_2281);
and UO_11 (O_11,N_2608,N_2389);
nor UO_12 (O_12,N_2223,N_2519);
nor UO_13 (O_13,N_2764,N_2847);
or UO_14 (O_14,N_2371,N_2813);
xor UO_15 (O_15,N_2726,N_2476);
or UO_16 (O_16,N_2249,N_2468);
xnor UO_17 (O_17,N_2253,N_2091);
nand UO_18 (O_18,N_2036,N_2409);
xor UO_19 (O_19,N_2950,N_2451);
xor UO_20 (O_20,N_2830,N_2563);
and UO_21 (O_21,N_2202,N_2505);
nand UO_22 (O_22,N_2047,N_2376);
nand UO_23 (O_23,N_2616,N_2138);
nand UO_24 (O_24,N_2330,N_2752);
nor UO_25 (O_25,N_2353,N_2094);
xor UO_26 (O_26,N_2687,N_2248);
or UO_27 (O_27,N_2421,N_2835);
and UO_28 (O_28,N_2997,N_2020);
nand UO_29 (O_29,N_2979,N_2296);
and UO_30 (O_30,N_2879,N_2507);
or UO_31 (O_31,N_2911,N_2331);
and UO_32 (O_32,N_2454,N_2908);
or UO_33 (O_33,N_2518,N_2295);
nand UO_34 (O_34,N_2972,N_2705);
nor UO_35 (O_35,N_2803,N_2828);
or UO_36 (O_36,N_2786,N_2374);
and UO_37 (O_37,N_2147,N_2920);
nand UO_38 (O_38,N_2928,N_2289);
nand UO_39 (O_39,N_2048,N_2228);
nand UO_40 (O_40,N_2526,N_2931);
nor UO_41 (O_41,N_2595,N_2059);
and UO_42 (O_42,N_2050,N_2366);
or UO_43 (O_43,N_2743,N_2874);
nand UO_44 (O_44,N_2470,N_2955);
and UO_45 (O_45,N_2751,N_2079);
or UO_46 (O_46,N_2065,N_2863);
nand UO_47 (O_47,N_2493,N_2042);
nand UO_48 (O_48,N_2839,N_2986);
nand UO_49 (O_49,N_2842,N_2814);
or UO_50 (O_50,N_2346,N_2989);
nor UO_51 (O_51,N_2926,N_2506);
nand UO_52 (O_52,N_2142,N_2122);
nand UO_53 (O_53,N_2089,N_2106);
xnor UO_54 (O_54,N_2156,N_2818);
nor UO_55 (O_55,N_2647,N_2154);
nand UO_56 (O_56,N_2490,N_2210);
and UO_57 (O_57,N_2825,N_2218);
nor UO_58 (O_58,N_2153,N_2888);
nand UO_59 (O_59,N_2410,N_2232);
nand UO_60 (O_60,N_2582,N_2586);
nor UO_61 (O_61,N_2286,N_2824);
nor UO_62 (O_62,N_2163,N_2499);
or UO_63 (O_63,N_2599,N_2954);
nand UO_64 (O_64,N_2508,N_2539);
and UO_65 (O_65,N_2528,N_2822);
or UO_66 (O_66,N_2807,N_2870);
nand UO_67 (O_67,N_2385,N_2978);
nand UO_68 (O_68,N_2712,N_2112);
xor UO_69 (O_69,N_2173,N_2683);
nand UO_70 (O_70,N_2278,N_2244);
or UO_71 (O_71,N_2999,N_2922);
or UO_72 (O_72,N_2572,N_2808);
nand UO_73 (O_73,N_2140,N_2340);
and UO_74 (O_74,N_2061,N_2419);
and UO_75 (O_75,N_2766,N_2732);
or UO_76 (O_76,N_2692,N_2939);
or UO_77 (O_77,N_2548,N_2023);
nand UO_78 (O_78,N_2536,N_2541);
nor UO_79 (O_79,N_2898,N_2379);
or UO_80 (O_80,N_2985,N_2483);
or UO_81 (O_81,N_2715,N_2936);
nor UO_82 (O_82,N_2277,N_2642);
or UO_83 (O_83,N_2570,N_2949);
nand UO_84 (O_84,N_2229,N_2934);
xor UO_85 (O_85,N_2199,N_2471);
nand UO_86 (O_86,N_2355,N_2740);
xor UO_87 (O_87,N_2924,N_2022);
and UO_88 (O_88,N_2200,N_2373);
nand UO_89 (O_89,N_2625,N_2609);
nor UO_90 (O_90,N_2799,N_2110);
nand UO_91 (O_91,N_2427,N_2812);
nand UO_92 (O_92,N_2744,N_2323);
xor UO_93 (O_93,N_2660,N_2532);
nand UO_94 (O_94,N_2615,N_2524);
or UO_95 (O_95,N_2222,N_2995);
nor UO_96 (O_96,N_2266,N_2058);
xor UO_97 (O_97,N_2095,N_2845);
nand UO_98 (O_98,N_2258,N_2953);
and UO_99 (O_99,N_2361,N_2408);
nor UO_100 (O_100,N_2206,N_2378);
and UO_101 (O_101,N_2407,N_2975);
nor UO_102 (O_102,N_2363,N_2513);
nor UO_103 (O_103,N_2443,N_2733);
or UO_104 (O_104,N_2871,N_2968);
and UO_105 (O_105,N_2216,N_2884);
nor UO_106 (O_106,N_2334,N_2804);
or UO_107 (O_107,N_2170,N_2083);
xor UO_108 (O_108,N_2085,N_2875);
or UO_109 (O_109,N_2190,N_2587);
xnor UO_110 (O_110,N_2984,N_2321);
nand UO_111 (O_111,N_2956,N_2209);
nand UO_112 (O_112,N_2857,N_2194);
nor UO_113 (O_113,N_2891,N_2211);
nand UO_114 (O_114,N_2093,N_2257);
nand UO_115 (O_115,N_2246,N_2195);
and UO_116 (O_116,N_2298,N_2840);
and UO_117 (O_117,N_2991,N_2597);
and UO_118 (O_118,N_2500,N_2903);
nand UO_119 (O_119,N_2671,N_2957);
xnor UO_120 (O_120,N_2880,N_2052);
nand UO_121 (O_121,N_2482,N_2019);
or UO_122 (O_122,N_2598,N_2324);
and UO_123 (O_123,N_2622,N_2567);
nand UO_124 (O_124,N_2645,N_2876);
and UO_125 (O_125,N_2774,N_2486);
nand UO_126 (O_126,N_2546,N_2777);
nor UO_127 (O_127,N_2342,N_2648);
and UO_128 (O_128,N_2730,N_2855);
or UO_129 (O_129,N_2162,N_2082);
and UO_130 (O_130,N_2109,N_2203);
or UO_131 (O_131,N_2850,N_2425);
and UO_132 (O_132,N_2940,N_2463);
nor UO_133 (O_133,N_2489,N_2178);
or UO_134 (O_134,N_2259,N_2691);
nand UO_135 (O_135,N_2484,N_2894);
xor UO_136 (O_136,N_2575,N_2424);
nor UO_137 (O_137,N_2480,N_2204);
or UO_138 (O_138,N_2996,N_2478);
and UO_139 (O_139,N_2688,N_2741);
and UO_140 (O_140,N_2699,N_2593);
nand UO_141 (O_141,N_2086,N_2010);
nor UO_142 (O_142,N_2101,N_2717);
nor UO_143 (O_143,N_2551,N_2386);
and UO_144 (O_144,N_2959,N_2708);
nor UO_145 (O_145,N_2310,N_2064);
nand UO_146 (O_146,N_2237,N_2097);
and UO_147 (O_147,N_2588,N_2977);
or UO_148 (O_148,N_2196,N_2423);
and UO_149 (O_149,N_2654,N_2935);
or UO_150 (O_150,N_2242,N_2440);
xnor UO_151 (O_151,N_2714,N_2626);
or UO_152 (O_152,N_2562,N_2633);
and UO_153 (O_153,N_2365,N_2716);
nor UO_154 (O_154,N_2707,N_2983);
or UO_155 (O_155,N_2401,N_2779);
or UO_156 (O_156,N_2030,N_2697);
nand UO_157 (O_157,N_2092,N_2738);
nor UO_158 (O_158,N_2836,N_2723);
and UO_159 (O_159,N_2102,N_2148);
and UO_160 (O_160,N_2028,N_2711);
or UO_161 (O_161,N_2971,N_2273);
nand UO_162 (O_162,N_2474,N_2669);
or UO_163 (O_163,N_2873,N_2641);
or UO_164 (O_164,N_2487,N_2613);
nand UO_165 (O_165,N_2938,N_2472);
and UO_166 (O_166,N_2400,N_2369);
or UO_167 (O_167,N_2798,N_2554);
or UO_168 (O_168,N_2737,N_2987);
and UO_169 (O_169,N_2193,N_2848);
nand UO_170 (O_170,N_2317,N_2157);
nor UO_171 (O_171,N_2160,N_2638);
nor UO_172 (O_172,N_2927,N_2527);
and UO_173 (O_173,N_2322,N_2233);
and UO_174 (O_174,N_2351,N_2031);
nor UO_175 (O_175,N_2695,N_2702);
and UO_176 (O_176,N_2341,N_2542);
nor UO_177 (O_177,N_2428,N_2557);
nor UO_178 (O_178,N_2794,N_2458);
and UO_179 (O_179,N_2681,N_2267);
nor UO_180 (O_180,N_2914,N_2896);
and UO_181 (O_181,N_2414,N_2603);
nand UO_182 (O_182,N_2621,N_2854);
nand UO_183 (O_183,N_2358,N_2040);
or UO_184 (O_184,N_2168,N_2537);
and UO_185 (O_185,N_2159,N_2992);
nor UO_186 (O_186,N_2791,N_2618);
and UO_187 (O_187,N_2306,N_2449);
nand UO_188 (O_188,N_2769,N_2224);
xor UO_189 (O_189,N_2236,N_2074);
or UO_190 (O_190,N_2117,N_2139);
nor UO_191 (O_191,N_2653,N_2682);
nor UO_192 (O_192,N_2754,N_2912);
nor UO_193 (O_193,N_2447,N_2776);
and UO_194 (O_194,N_2217,N_2429);
nor UO_195 (O_195,N_2309,N_2114);
or UO_196 (O_196,N_2098,N_2559);
nand UO_197 (O_197,N_2982,N_2280);
xnor UO_198 (O_198,N_2496,N_2543);
nand UO_199 (O_199,N_2607,N_2166);
nand UO_200 (O_200,N_2651,N_2742);
nand UO_201 (O_201,N_2843,N_2069);
nand UO_202 (O_202,N_2547,N_2271);
nor UO_203 (O_203,N_2005,N_2747);
xor UO_204 (O_204,N_2326,N_2990);
nor UO_205 (O_205,N_2370,N_2788);
nand UO_206 (O_206,N_2132,N_2301);
or UO_207 (O_207,N_2580,N_2531);
nor UO_208 (O_208,N_2188,N_2319);
or UO_209 (O_209,N_2590,N_2491);
and UO_210 (O_210,N_2789,N_2197);
nand UO_211 (O_211,N_2823,N_2831);
and UO_212 (O_212,N_2853,N_2320);
or UO_213 (O_213,N_2214,N_2186);
or UO_214 (O_214,N_2055,N_2963);
nand UO_215 (O_215,N_2512,N_2314);
nor UO_216 (O_216,N_2039,N_2433);
or UO_217 (O_217,N_2335,N_2535);
nand UO_218 (O_218,N_2072,N_2383);
or UO_219 (O_219,N_2238,N_2285);
nor UO_220 (O_220,N_2413,N_2460);
or UO_221 (O_221,N_2591,N_2865);
and UO_222 (O_222,N_2727,N_2292);
or UO_223 (O_223,N_2388,N_2672);
nand UO_224 (O_224,N_2442,N_2096);
xnor UO_225 (O_225,N_2619,N_2269);
nand UO_226 (O_226,N_2029,N_2088);
nor UO_227 (O_227,N_2810,N_2377);
or UO_228 (O_228,N_2686,N_2834);
nand UO_229 (O_229,N_2315,N_2437);
or UO_230 (O_230,N_2600,N_2129);
nand UO_231 (O_231,N_2942,N_2930);
or UO_232 (O_232,N_2046,N_2631);
nor UO_233 (O_233,N_2966,N_2734);
nand UO_234 (O_234,N_2191,N_2165);
nand UO_235 (O_235,N_2304,N_2501);
or UO_236 (O_236,N_2384,N_2629);
nor UO_237 (O_237,N_2137,N_2063);
nand UO_238 (O_238,N_2602,N_2680);
nand UO_239 (O_239,N_2974,N_2455);
and UO_240 (O_240,N_2347,N_2494);
or UO_241 (O_241,N_2171,N_2418);
or UO_242 (O_242,N_2439,N_2951);
nand UO_243 (O_243,N_2650,N_2124);
and UO_244 (O_244,N_2525,N_2801);
nand UO_245 (O_245,N_2770,N_2674);
nand UO_246 (O_246,N_2014,N_2560);
and UO_247 (O_247,N_2430,N_2817);
or UO_248 (O_248,N_2806,N_2151);
nand UO_249 (O_249,N_2392,N_2504);
or UO_250 (O_250,N_2219,N_2820);
or UO_251 (O_251,N_2576,N_2704);
nand UO_252 (O_252,N_2375,N_2796);
or UO_253 (O_253,N_2829,N_2453);
nand UO_254 (O_254,N_2025,N_2231);
or UO_255 (O_255,N_2348,N_2540);
nor UO_256 (O_256,N_2062,N_2709);
nor UO_257 (O_257,N_2778,N_2144);
and UO_258 (O_258,N_2270,N_2364);
or UO_259 (O_259,N_2477,N_2108);
or UO_260 (O_260,N_2299,N_2033);
and UO_261 (O_261,N_2282,N_2946);
and UO_262 (O_262,N_2675,N_2878);
and UO_263 (O_263,N_2345,N_2890);
and UO_264 (O_264,N_2721,N_2900);
or UO_265 (O_265,N_2964,N_2422);
nand UO_266 (O_266,N_2561,N_2391);
nor UO_267 (O_267,N_2316,N_2397);
nand UO_268 (O_268,N_2338,N_2049);
xnor UO_269 (O_269,N_2658,N_2755);
nand UO_270 (O_270,N_2387,N_2533);
and UO_271 (O_271,N_2274,N_2509);
xnor UO_272 (O_272,N_2497,N_2811);
nor UO_273 (O_273,N_2416,N_2021);
xnor UO_274 (O_274,N_2256,N_2056);
nor UO_275 (O_275,N_2390,N_2993);
nand UO_276 (O_276,N_2511,N_2893);
nor UO_277 (O_277,N_2076,N_2923);
or UO_278 (O_278,N_2994,N_2434);
nor UO_279 (O_279,N_2556,N_2965);
and UO_280 (O_280,N_2724,N_2736);
and UO_281 (O_281,N_2569,N_2868);
nand UO_282 (O_282,N_2759,N_2594);
nand UO_283 (O_283,N_2445,N_2100);
xnor UO_284 (O_284,N_2308,N_2164);
nand UO_285 (O_285,N_2584,N_2087);
nor UO_286 (O_286,N_2678,N_2765);
or UO_287 (O_287,N_2902,N_2130);
nand UO_288 (O_288,N_2261,N_2145);
nor UO_289 (O_289,N_2260,N_2081);
or UO_290 (O_290,N_2344,N_2970);
nor UO_291 (O_291,N_2910,N_2263);
nor UO_292 (O_292,N_2465,N_2589);
nand UO_293 (O_293,N_2394,N_2240);
and UO_294 (O_294,N_2663,N_2662);
or UO_295 (O_295,N_2473,N_2601);
nand UO_296 (O_296,N_2819,N_2017);
or UO_297 (O_297,N_2882,N_2659);
nand UO_298 (O_298,N_2670,N_2523);
nand UO_299 (O_299,N_2731,N_2713);
or UO_300 (O_300,N_2303,N_2007);
nor UO_301 (O_301,N_2652,N_2703);
or UO_302 (O_302,N_2720,N_2690);
xor UO_303 (O_303,N_2404,N_2131);
nand UO_304 (O_304,N_2762,N_2862);
nor UO_305 (O_305,N_2398,N_2127);
nand UO_306 (O_306,N_2441,N_2431);
nand UO_307 (O_307,N_2909,N_2012);
xnor UO_308 (O_308,N_2272,N_2502);
xor UO_309 (O_309,N_2185,N_2552);
nand UO_310 (O_310,N_2003,N_2735);
nor UO_311 (O_311,N_2198,N_2612);
or UO_312 (O_312,N_2578,N_2015);
nand UO_313 (O_313,N_2118,N_2851);
xor UO_314 (O_314,N_2739,N_2411);
or UO_315 (O_315,N_2115,N_2402);
nand UO_316 (O_316,N_2399,N_2300);
or UO_317 (O_317,N_2883,N_2234);
and UO_318 (O_318,N_2485,N_2172);
nor UO_319 (O_319,N_2772,N_2456);
or UO_320 (O_320,N_2611,N_2177);
nand UO_321 (O_321,N_2367,N_2573);
xnor UO_322 (O_322,N_2352,N_2549);
nor UO_323 (O_323,N_2841,N_2368);
or UO_324 (O_324,N_2921,N_2435);
xor UO_325 (O_325,N_2356,N_2452);
nand UO_326 (O_326,N_2349,N_2123);
nand UO_327 (O_327,N_2522,N_2354);
or UO_328 (O_328,N_2450,N_2119);
nor UO_329 (O_329,N_2555,N_2725);
or UO_330 (O_330,N_2574,N_2700);
nor UO_331 (O_331,N_2846,N_2782);
nand UO_332 (O_332,N_2781,N_2287);
xnor UO_333 (O_333,N_2037,N_2189);
nor UO_334 (O_334,N_2656,N_2775);
xor UO_335 (O_335,N_2617,N_2068);
nor UO_336 (O_336,N_2872,N_2693);
or UO_337 (O_337,N_2078,N_2488);
or UO_338 (O_338,N_2469,N_2816);
and UO_339 (O_339,N_2838,N_2252);
nor UO_340 (O_340,N_2275,N_2035);
and UO_341 (O_341,N_2581,N_2668);
xor UO_342 (O_342,N_2051,N_2000);
and UO_343 (O_343,N_2034,N_2881);
nor UO_344 (O_344,N_2143,N_2901);
or UO_345 (O_345,N_2632,N_2844);
nand UO_346 (O_346,N_2947,N_2313);
nand UO_347 (O_347,N_2925,N_2646);
and UO_348 (O_348,N_2503,N_2307);
or UO_349 (O_349,N_2318,N_2444);
nor UO_350 (O_350,N_2916,N_2784);
or UO_351 (O_351,N_2550,N_2250);
or UO_352 (O_352,N_2805,N_2544);
or UO_353 (O_353,N_2639,N_2044);
nor UO_354 (O_354,N_2517,N_2060);
nand UO_355 (O_355,N_2305,N_2183);
nor UO_356 (O_356,N_2350,N_2952);
and UO_357 (O_357,N_2673,N_2797);
nand UO_358 (O_358,N_2008,N_2312);
or UO_359 (O_359,N_2038,N_2521);
nand UO_360 (O_360,N_2948,N_2800);
nor UO_361 (O_361,N_2343,N_2254);
nand UO_362 (O_362,N_2325,N_2790);
nor UO_363 (O_363,N_2534,N_2596);
or UO_364 (O_364,N_2181,N_2785);
or UO_365 (O_365,N_2773,N_2988);
nand UO_366 (O_366,N_2945,N_2564);
nand UO_367 (O_367,N_2426,N_2719);
or UO_368 (O_368,N_2634,N_2944);
and UO_369 (O_369,N_2729,N_2530);
or UO_370 (O_370,N_2684,N_2329);
and UO_371 (O_371,N_2084,N_2962);
xor UO_372 (O_372,N_2753,N_2577);
and UO_373 (O_373,N_2913,N_2756);
and UO_374 (O_374,N_2043,N_2718);
or UO_375 (O_375,N_2869,N_2566);
and UO_376 (O_376,N_2649,N_2827);
or UO_377 (O_377,N_2657,N_2406);
and UO_378 (O_378,N_2767,N_2859);
and UO_379 (O_379,N_2464,N_2026);
or UO_380 (O_380,N_2066,N_2849);
xor UO_381 (O_381,N_2090,N_2892);
or UO_382 (O_382,N_2184,N_2205);
nor UO_383 (O_383,N_2637,N_2960);
or UO_384 (O_384,N_2475,N_2073);
nand UO_385 (O_385,N_2710,N_2529);
or UO_386 (O_386,N_2415,N_2395);
and UO_387 (O_387,N_2636,N_2571);
xor UO_388 (O_388,N_2276,N_2461);
nor UO_389 (O_389,N_2192,N_2099);
or UO_390 (O_390,N_2746,N_2380);
nor UO_391 (O_391,N_2787,N_2146);
nand UO_392 (O_392,N_2161,N_2221);
and UO_393 (O_393,N_2745,N_2895);
xnor UO_394 (O_394,N_2393,N_2961);
xor UO_395 (O_395,N_2696,N_2432);
or UO_396 (O_396,N_2245,N_2001);
or UO_397 (O_397,N_2174,N_2167);
xnor UO_398 (O_398,N_2412,N_2247);
and UO_399 (O_399,N_2134,N_2405);
nand UO_400 (O_400,N_2826,N_2677);
and UO_401 (O_401,N_2337,N_2821);
and UO_402 (O_402,N_2176,N_2446);
or UO_403 (O_403,N_2606,N_2227);
nor UO_404 (O_404,N_2116,N_2175);
and UO_405 (O_405,N_2685,N_2187);
or UO_406 (O_406,N_2837,N_2403);
xor UO_407 (O_407,N_2133,N_2538);
nand UO_408 (O_408,N_2080,N_2748);
and UO_409 (O_409,N_2107,N_2360);
and UO_410 (O_410,N_2706,N_2103);
nand UO_411 (O_411,N_2009,N_2644);
xnor UO_412 (O_412,N_2623,N_2466);
or UO_413 (O_413,N_2230,N_2032);
or UO_414 (O_414,N_2239,N_2793);
nor UO_415 (O_415,N_2111,N_2041);
and UO_416 (O_416,N_2832,N_2225);
nor UO_417 (O_417,N_2291,N_2495);
xor UO_418 (O_418,N_2768,N_2158);
or UO_419 (O_419,N_2783,N_2667);
nand UO_420 (O_420,N_2792,N_2311);
xnor UO_421 (O_421,N_2771,N_2182);
or UO_422 (O_422,N_2861,N_2679);
xnor UO_423 (O_423,N_2761,N_2867);
nand UO_424 (O_424,N_2243,N_2018);
nor UO_425 (O_425,N_2077,N_2553);
nor UO_426 (O_426,N_2969,N_2802);
nand UO_427 (O_427,N_2179,N_2510);
or UO_428 (O_428,N_2070,N_2016);
and UO_429 (O_429,N_2381,N_2604);
nand UO_430 (O_430,N_2579,N_2071);
nor UO_431 (O_431,N_2220,N_2126);
nand UO_432 (O_432,N_2973,N_2628);
and UO_433 (O_433,N_2462,N_2336);
nor UO_434 (O_434,N_2125,N_2701);
and UO_435 (O_435,N_2438,N_2141);
and UO_436 (O_436,N_2339,N_2967);
nor UO_437 (O_437,N_2264,N_2941);
nand UO_438 (O_438,N_2328,N_2155);
nand UO_439 (O_439,N_2665,N_2640);
nand UO_440 (O_440,N_2904,N_2024);
or UO_441 (O_441,N_2933,N_2860);
nor UO_442 (O_442,N_2886,N_2592);
xor UO_443 (O_443,N_2327,N_2630);
and UO_444 (O_444,N_2514,N_2420);
nor UO_445 (O_445,N_2568,N_2635);
xor UO_446 (O_446,N_2152,N_2558);
and UO_447 (O_447,N_2113,N_2294);
xnor UO_448 (O_448,N_2457,N_2459);
and UO_449 (O_449,N_2664,N_2235);
xor UO_450 (O_450,N_2213,N_2728);
or UO_451 (O_451,N_2929,N_2917);
or UO_452 (O_452,N_2809,N_2998);
or UO_453 (O_453,N_2856,N_2251);
nand UO_454 (O_454,N_2479,N_2899);
or UO_455 (O_455,N_2215,N_2105);
nand UO_456 (O_456,N_2760,N_2698);
xor UO_457 (O_457,N_2467,N_2120);
and UO_458 (O_458,N_2302,N_2293);
or UO_459 (O_459,N_2614,N_2332);
nand UO_460 (O_460,N_2396,N_2284);
nand UO_461 (O_461,N_2207,N_2980);
or UO_462 (O_462,N_2958,N_2288);
nand UO_463 (O_463,N_2627,N_2897);
xnor UO_464 (O_464,N_2498,N_2833);
xnor UO_465 (O_465,N_2852,N_2201);
and UO_466 (O_466,N_2757,N_2750);
nand UO_467 (O_467,N_2226,N_2915);
or UO_468 (O_468,N_2666,N_2011);
and UO_469 (O_469,N_2075,N_2006);
xor UO_470 (O_470,N_2283,N_2643);
or UO_471 (O_471,N_2362,N_2121);
and UO_472 (O_472,N_2887,N_2858);
and UO_473 (O_473,N_2027,N_2054);
nor UO_474 (O_474,N_2907,N_2128);
nand UO_475 (O_475,N_2583,N_2889);
and UO_476 (O_476,N_2169,N_2689);
xor UO_477 (O_477,N_2877,N_2279);
nor UO_478 (O_478,N_2241,N_2448);
and UO_479 (O_479,N_2585,N_2981);
or UO_480 (O_480,N_2722,N_2180);
and UO_481 (O_481,N_2045,N_2372);
nor UO_482 (O_482,N_2265,N_2208);
nand UO_483 (O_483,N_2067,N_2002);
and UO_484 (O_484,N_2885,N_2013);
or UO_485 (O_485,N_2359,N_2262);
nand UO_486 (O_486,N_2212,N_2545);
and UO_487 (O_487,N_2333,N_2932);
nor UO_488 (O_488,N_2780,N_2520);
nor UO_489 (O_489,N_2610,N_2436);
and UO_490 (O_490,N_2906,N_2655);
nor UO_491 (O_491,N_2624,N_2290);
nor UO_492 (O_492,N_2943,N_2694);
or UO_493 (O_493,N_2661,N_2676);
nand UO_494 (O_494,N_2605,N_2866);
xnor UO_495 (O_495,N_2620,N_2150);
nand UO_496 (O_496,N_2357,N_2516);
xor UO_497 (O_497,N_2255,N_2268);
or UO_498 (O_498,N_2149,N_2749);
and UO_499 (O_499,N_2136,N_2297);
endmodule