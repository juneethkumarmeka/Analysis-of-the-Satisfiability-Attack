module basic_500_3000_500_50_levels_1xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_457,In_369);
nor U1 (N_1,In_23,In_377);
nor U2 (N_2,In_124,In_342);
nand U3 (N_3,In_483,In_33);
nand U4 (N_4,In_452,In_464);
nand U5 (N_5,In_434,In_253);
and U6 (N_6,In_155,In_265);
or U7 (N_7,In_398,In_293);
or U8 (N_8,In_246,In_344);
or U9 (N_9,In_463,In_258);
nor U10 (N_10,In_305,In_169);
or U11 (N_11,In_167,In_96);
and U12 (N_12,In_18,In_481);
or U13 (N_13,In_372,In_394);
or U14 (N_14,In_107,In_373);
and U15 (N_15,In_201,In_172);
and U16 (N_16,In_255,In_269);
nor U17 (N_17,In_208,In_32);
nor U18 (N_18,In_217,In_70);
and U19 (N_19,In_498,In_365);
or U20 (N_20,In_327,In_470);
nand U21 (N_21,In_382,In_163);
and U22 (N_22,In_159,In_476);
nand U23 (N_23,In_26,In_188);
nor U24 (N_24,In_304,In_19);
or U25 (N_25,In_338,In_170);
nor U26 (N_26,In_280,In_77);
nor U27 (N_27,In_162,In_8);
nor U28 (N_28,In_78,In_141);
nand U29 (N_29,In_189,In_419);
or U30 (N_30,In_479,In_408);
nor U31 (N_31,In_227,In_443);
nand U32 (N_32,In_360,In_161);
nand U33 (N_33,In_49,In_12);
nand U34 (N_34,In_199,In_370);
and U35 (N_35,In_371,In_296);
or U36 (N_36,In_390,In_263);
and U37 (N_37,In_134,In_387);
nand U38 (N_38,In_456,In_71);
nand U39 (N_39,In_119,In_55);
nand U40 (N_40,In_166,In_386);
nand U41 (N_41,In_302,In_175);
nand U42 (N_42,In_493,In_95);
and U43 (N_43,In_478,In_142);
nor U44 (N_44,In_30,In_3);
nand U45 (N_45,In_353,In_319);
nand U46 (N_46,In_127,In_31);
nand U47 (N_47,In_471,In_225);
nor U48 (N_48,In_115,In_423);
nand U49 (N_49,In_406,In_299);
nand U50 (N_50,In_67,In_184);
nor U51 (N_51,In_42,In_277);
nand U52 (N_52,In_287,In_278);
nand U53 (N_53,In_58,In_266);
nor U54 (N_54,In_424,In_348);
nor U55 (N_55,In_404,In_47);
nor U56 (N_56,In_139,In_214);
nor U57 (N_57,In_181,In_43);
and U58 (N_58,In_157,In_313);
nand U59 (N_59,In_444,In_484);
nand U60 (N_60,In_100,In_368);
nor U61 (N_61,N_13,In_34);
nor U62 (N_62,N_3,In_216);
and U63 (N_63,In_429,In_282);
or U64 (N_64,In_381,In_194);
and U65 (N_65,In_435,In_272);
nand U66 (N_66,In_379,N_19);
nor U67 (N_67,In_421,In_206);
nand U68 (N_68,N_4,In_25);
or U69 (N_69,In_63,In_494);
or U70 (N_70,N_33,In_416);
nor U71 (N_71,In_37,In_85);
nor U72 (N_72,In_15,N_51);
nor U73 (N_73,In_51,N_32);
nand U74 (N_74,In_279,In_60);
and U75 (N_75,In_200,In_219);
nor U76 (N_76,In_140,In_84);
xnor U77 (N_77,In_380,In_228);
and U78 (N_78,In_105,In_318);
nand U79 (N_79,N_30,In_249);
or U80 (N_80,N_11,N_5);
nand U81 (N_81,In_467,In_146);
and U82 (N_82,In_358,In_164);
nor U83 (N_83,In_461,In_152);
nor U84 (N_84,In_294,In_136);
or U85 (N_85,In_28,In_116);
nand U86 (N_86,In_480,In_359);
nor U87 (N_87,In_221,N_8);
and U88 (N_88,In_462,In_303);
or U89 (N_89,In_357,In_454);
or U90 (N_90,In_430,N_52);
nor U91 (N_91,In_306,In_262);
nor U92 (N_92,In_393,In_286);
and U93 (N_93,In_252,In_364);
and U94 (N_94,In_80,In_234);
nor U95 (N_95,In_106,N_44);
nor U96 (N_96,In_384,In_496);
nor U97 (N_97,In_6,N_47);
nor U98 (N_98,In_367,In_340);
and U99 (N_99,In_300,In_273);
nor U100 (N_100,In_420,In_397);
or U101 (N_101,In_191,In_68);
nor U102 (N_102,N_12,In_195);
and U103 (N_103,In_447,In_190);
xnor U104 (N_104,In_104,In_314);
and U105 (N_105,In_123,In_289);
nor U106 (N_106,In_477,In_7);
nor U107 (N_107,In_57,In_491);
and U108 (N_108,In_165,In_198);
and U109 (N_109,In_325,In_245);
nand U110 (N_110,In_242,In_466);
or U111 (N_111,In_235,In_453);
and U112 (N_112,In_401,In_276);
or U113 (N_113,N_17,N_59);
or U114 (N_114,In_171,N_54);
nor U115 (N_115,In_251,In_324);
and U116 (N_116,In_224,In_10);
and U117 (N_117,N_18,In_337);
or U118 (N_118,In_322,In_499);
or U119 (N_119,In_9,In_237);
nand U120 (N_120,N_92,In_345);
and U121 (N_121,In_418,In_485);
or U122 (N_122,N_85,In_458);
or U123 (N_123,In_138,In_329);
nor U124 (N_124,N_86,In_192);
nand U125 (N_125,In_233,In_145);
or U126 (N_126,In_187,In_413);
and U127 (N_127,In_349,N_79);
nor U128 (N_128,In_450,N_117);
or U129 (N_129,In_405,N_37);
nor U130 (N_130,In_259,N_75);
and U131 (N_131,In_326,In_343);
nand U132 (N_132,In_411,In_341);
nand U133 (N_133,N_118,In_487);
nor U134 (N_134,In_65,In_400);
nand U135 (N_135,In_4,In_182);
and U136 (N_136,In_17,In_90);
and U137 (N_137,In_376,In_308);
and U138 (N_138,In_230,In_218);
nor U139 (N_139,N_29,In_417);
and U140 (N_140,In_250,In_236);
nand U141 (N_141,In_240,In_431);
or U142 (N_142,In_148,In_415);
nand U143 (N_143,In_76,In_283);
or U144 (N_144,N_45,In_366);
nand U145 (N_145,N_73,In_482);
or U146 (N_146,In_399,N_103);
nand U147 (N_147,N_21,In_121);
and U148 (N_148,In_281,N_0);
nor U149 (N_149,In_441,In_363);
or U150 (N_150,N_23,N_71);
nand U151 (N_151,In_53,In_117);
nor U152 (N_152,In_52,In_267);
nand U153 (N_153,In_355,In_465);
and U154 (N_154,In_109,In_73);
nor U155 (N_155,In_254,In_168);
nand U156 (N_156,In_94,In_449);
or U157 (N_157,In_1,In_455);
nor U158 (N_158,N_110,N_10);
or U159 (N_159,In_488,In_178);
nor U160 (N_160,In_425,In_412);
or U161 (N_161,In_437,In_260);
or U162 (N_162,N_112,In_291);
nor U163 (N_163,N_100,In_113);
nor U164 (N_164,In_274,N_77);
nor U165 (N_165,N_50,N_95);
nand U166 (N_166,In_149,In_27);
and U167 (N_167,In_241,In_36);
or U168 (N_168,In_261,In_385);
or U169 (N_169,N_68,N_108);
nand U170 (N_170,N_106,In_183);
or U171 (N_171,In_248,In_323);
and U172 (N_172,In_229,In_432);
nand U173 (N_173,In_247,N_20);
or U174 (N_174,In_137,N_1);
or U175 (N_175,In_203,In_197);
nor U176 (N_176,In_231,In_11);
nor U177 (N_177,N_102,In_122);
nor U178 (N_178,In_213,In_112);
nor U179 (N_179,In_451,N_48);
nand U180 (N_180,N_90,In_285);
and U181 (N_181,N_138,N_46);
and U182 (N_182,In_409,In_298);
nand U183 (N_183,In_48,In_469);
or U184 (N_184,In_103,In_244);
or U185 (N_185,In_495,In_24);
or U186 (N_186,N_127,N_88);
and U187 (N_187,N_69,In_490);
nor U188 (N_188,In_144,In_0);
nand U189 (N_189,In_150,In_375);
or U190 (N_190,In_332,In_440);
nand U191 (N_191,N_111,N_96);
and U192 (N_192,N_145,In_210);
nor U193 (N_193,N_105,N_172);
nand U194 (N_194,N_70,N_169);
or U195 (N_195,In_351,N_178);
and U196 (N_196,N_167,In_226);
or U197 (N_197,In_426,In_174);
nor U198 (N_198,In_328,N_135);
nor U199 (N_199,N_38,In_307);
nor U200 (N_200,In_336,In_207);
or U201 (N_201,In_176,N_109);
nand U202 (N_202,In_114,N_99);
or U203 (N_203,In_75,In_243);
nor U204 (N_204,In_402,In_330);
and U205 (N_205,In_239,N_114);
nor U206 (N_206,N_177,In_442);
or U207 (N_207,In_321,In_131);
nor U208 (N_208,In_158,In_215);
and U209 (N_209,N_131,In_220);
and U210 (N_210,In_29,N_65);
nor U211 (N_211,N_137,N_147);
nor U212 (N_212,In_160,In_331);
and U213 (N_213,In_83,N_58);
or U214 (N_214,In_179,N_173);
nor U215 (N_215,N_63,In_154);
or U216 (N_216,In_128,In_335);
nor U217 (N_217,In_396,In_61);
and U218 (N_218,In_35,In_211);
nor U219 (N_219,N_41,In_41);
nor U220 (N_220,In_354,In_108);
and U221 (N_221,In_40,N_7);
nand U222 (N_222,N_179,N_120);
nand U223 (N_223,In_275,N_15);
or U224 (N_224,N_42,In_392);
or U225 (N_225,In_361,In_407);
nand U226 (N_226,N_89,In_316);
nand U227 (N_227,N_134,N_126);
and U228 (N_228,In_204,N_35);
nand U229 (N_229,In_395,In_232);
and U230 (N_230,N_171,In_414);
nand U231 (N_231,N_28,In_54);
nor U232 (N_232,N_150,N_93);
or U233 (N_233,In_486,In_64);
nor U234 (N_234,N_113,N_148);
nor U235 (N_235,In_315,In_89);
nand U236 (N_236,N_67,N_162);
nor U237 (N_237,In_256,N_123);
nor U238 (N_238,N_43,In_317);
and U239 (N_239,N_161,In_438);
and U240 (N_240,In_301,In_93);
nor U241 (N_241,In_223,In_69);
or U242 (N_242,In_74,N_202);
nor U243 (N_243,N_210,N_154);
nor U244 (N_244,N_222,In_297);
nand U245 (N_245,In_133,In_118);
and U246 (N_246,N_228,In_489);
nor U247 (N_247,N_200,N_144);
nand U248 (N_248,In_292,N_225);
and U249 (N_249,In_92,N_142);
and U250 (N_250,N_24,In_130);
nand U251 (N_251,N_128,N_209);
nand U252 (N_252,N_34,N_116);
nand U253 (N_253,In_311,In_97);
nor U254 (N_254,N_119,N_207);
or U255 (N_255,N_80,N_193);
and U256 (N_256,N_107,In_428);
or U257 (N_257,In_433,N_215);
or U258 (N_258,In_422,In_378);
nor U259 (N_259,N_223,N_229);
and U260 (N_260,In_312,In_16);
and U261 (N_261,In_346,In_13);
nor U262 (N_262,In_72,In_129);
and U263 (N_263,In_448,N_132);
nor U264 (N_264,In_44,N_83);
nor U265 (N_265,N_211,In_62);
and U266 (N_266,N_56,N_194);
nand U267 (N_267,In_101,N_31);
or U268 (N_268,N_78,In_205);
or U269 (N_269,N_183,N_231);
and U270 (N_270,N_6,N_72);
and U271 (N_271,In_5,In_135);
and U272 (N_272,N_197,N_151);
nor U273 (N_273,In_88,N_49);
or U274 (N_274,N_216,In_202);
or U275 (N_275,N_101,N_232);
xnor U276 (N_276,N_36,N_136);
or U277 (N_277,In_2,N_235);
or U278 (N_278,N_226,N_218);
nand U279 (N_279,N_84,In_91);
nand U280 (N_280,N_236,In_59);
nor U281 (N_281,N_2,In_334);
or U282 (N_282,N_149,N_201);
nand U283 (N_283,N_181,In_82);
nand U284 (N_284,In_391,N_190);
nor U285 (N_285,N_220,N_141);
or U286 (N_286,N_186,N_22);
nand U287 (N_287,In_180,N_87);
nand U288 (N_288,N_40,In_50);
and U289 (N_289,In_320,N_156);
or U290 (N_290,In_445,In_147);
and U291 (N_291,In_473,In_99);
nand U292 (N_292,N_94,In_309);
nand U293 (N_293,N_62,In_56);
or U294 (N_294,In_339,In_126);
nand U295 (N_295,N_27,In_222);
and U296 (N_296,N_97,In_111);
or U297 (N_297,In_388,N_180);
nand U298 (N_298,N_16,In_14);
or U299 (N_299,N_191,In_446);
or U300 (N_300,N_240,In_186);
nor U301 (N_301,In_356,N_130);
nor U302 (N_302,In_98,In_153);
and U303 (N_303,In_268,N_196);
or U304 (N_304,In_185,N_271);
nor U305 (N_305,In_459,N_213);
or U306 (N_306,N_163,N_267);
nor U307 (N_307,N_296,N_168);
nor U308 (N_308,N_164,N_104);
nor U309 (N_309,In_350,In_173);
nor U310 (N_310,N_176,N_60);
nand U311 (N_311,In_156,N_166);
and U312 (N_312,N_115,In_22);
and U313 (N_313,N_268,N_295);
and U314 (N_314,N_158,N_82);
or U315 (N_315,N_140,In_492);
nand U316 (N_316,In_132,In_264);
and U317 (N_317,N_286,N_272);
nand U318 (N_318,N_274,N_39);
nand U319 (N_319,N_98,N_241);
nor U320 (N_320,N_91,In_310);
and U321 (N_321,N_254,N_26);
or U322 (N_322,In_38,N_124);
nor U323 (N_323,N_245,N_288);
nand U324 (N_324,N_280,In_389);
nand U325 (N_325,N_227,N_287);
and U326 (N_326,N_159,N_256);
and U327 (N_327,N_293,N_208);
nor U328 (N_328,In_288,N_297);
nor U329 (N_329,N_276,N_221);
and U330 (N_330,In_143,In_79);
or U331 (N_331,N_165,In_21);
nand U332 (N_332,N_214,N_143);
and U333 (N_333,In_333,In_410);
nand U334 (N_334,N_25,N_217);
and U335 (N_335,In_271,N_257);
nor U336 (N_336,N_269,In_110);
or U337 (N_337,N_263,N_282);
nand U338 (N_338,N_244,N_125);
or U339 (N_339,In_81,N_294);
and U340 (N_340,In_295,N_255);
nor U341 (N_341,N_285,N_182);
and U342 (N_342,N_249,In_468);
and U343 (N_343,N_160,N_247);
nor U344 (N_344,In_212,N_262);
nor U345 (N_345,N_248,In_196);
nand U346 (N_346,In_46,N_258);
nor U347 (N_347,N_146,In_427);
nand U348 (N_348,In_290,In_475);
or U349 (N_349,N_290,N_185);
nand U350 (N_350,N_188,In_193);
or U351 (N_351,N_265,N_129);
or U352 (N_352,N_251,N_170);
nor U353 (N_353,N_195,In_352);
or U354 (N_354,N_199,In_472);
or U355 (N_355,In_45,N_204);
nor U356 (N_356,N_14,In_257);
nor U357 (N_357,N_187,In_87);
or U358 (N_358,N_76,In_439);
and U359 (N_359,N_212,N_243);
and U360 (N_360,In_151,N_353);
and U361 (N_361,N_121,In_436);
and U362 (N_362,N_310,N_238);
nor U363 (N_363,N_358,N_329);
and U364 (N_364,N_206,N_316);
and U365 (N_365,N_355,N_189);
or U366 (N_366,N_354,N_299);
nor U367 (N_367,N_234,N_81);
nor U368 (N_368,N_192,N_250);
nand U369 (N_369,N_122,N_326);
or U370 (N_370,N_320,In_66);
nand U371 (N_371,N_270,N_301);
nor U372 (N_372,N_298,N_64);
nand U373 (N_373,N_233,N_334);
nand U374 (N_374,N_335,N_331);
nand U375 (N_375,In_209,N_305);
or U376 (N_376,N_330,In_347);
and U377 (N_377,N_321,N_259);
or U378 (N_378,N_74,N_133);
nor U379 (N_379,N_300,N_289);
and U380 (N_380,In_270,N_239);
or U381 (N_381,In_474,In_177);
or U382 (N_382,N_284,N_337);
nor U383 (N_383,N_317,N_327);
nand U384 (N_384,N_139,N_333);
or U385 (N_385,N_283,N_261);
nand U386 (N_386,N_348,N_260);
nand U387 (N_387,N_157,N_340);
nor U388 (N_388,N_345,N_242);
or U389 (N_389,N_342,N_314);
and U390 (N_390,In_86,N_66);
and U391 (N_391,N_291,In_120);
and U392 (N_392,N_350,In_362);
xor U393 (N_393,In_125,N_152);
and U394 (N_394,N_155,N_344);
or U395 (N_395,N_347,N_328);
nor U396 (N_396,N_252,N_205);
nor U397 (N_397,N_237,N_278);
and U398 (N_398,N_336,N_352);
nand U399 (N_399,N_308,In_403);
nand U400 (N_400,N_307,N_325);
nand U401 (N_401,N_318,In_238);
nor U402 (N_402,N_224,In_374);
or U403 (N_403,N_275,In_102);
nor U404 (N_404,N_322,N_277);
nor U405 (N_405,N_319,N_219);
nand U406 (N_406,N_53,N_273);
nand U407 (N_407,N_306,N_356);
nor U408 (N_408,N_246,N_61);
nand U409 (N_409,N_266,N_203);
nand U410 (N_410,N_230,In_460);
nand U411 (N_411,N_332,N_315);
or U412 (N_412,In_20,N_323);
nand U413 (N_413,N_281,N_343);
nand U414 (N_414,N_302,In_497);
or U415 (N_415,N_304,N_339);
nand U416 (N_416,N_313,N_292);
or U417 (N_417,In_39,N_153);
or U418 (N_418,N_357,N_198);
and U419 (N_419,N_57,N_351);
and U420 (N_420,N_410,N_399);
nand U421 (N_421,N_405,N_376);
or U422 (N_422,N_361,N_383);
nand U423 (N_423,N_174,N_412);
nand U424 (N_424,N_398,N_373);
and U425 (N_425,N_419,N_400);
nand U426 (N_426,N_397,N_380);
and U427 (N_427,N_324,N_382);
or U428 (N_428,N_395,In_383);
nor U429 (N_429,N_392,N_359);
or U430 (N_430,N_417,N_363);
and U431 (N_431,N_396,N_374);
nand U432 (N_432,N_406,N_349);
nor U433 (N_433,N_362,N_408);
nand U434 (N_434,N_381,N_413);
or U435 (N_435,N_311,N_386);
nand U436 (N_436,N_369,N_418);
nor U437 (N_437,N_384,N_370);
nand U438 (N_438,N_372,N_377);
or U439 (N_439,N_341,In_284);
nand U440 (N_440,N_365,N_55);
or U441 (N_441,N_387,N_416);
and U442 (N_442,N_414,N_279);
nand U443 (N_443,N_389,N_385);
nor U444 (N_444,N_402,N_367);
nor U445 (N_445,N_253,N_409);
and U446 (N_446,N_368,N_391);
or U447 (N_447,N_184,N_338);
and U448 (N_448,N_303,N_407);
or U449 (N_449,N_346,N_312);
and U450 (N_450,N_401,N_375);
nand U451 (N_451,N_371,N_378);
and U452 (N_452,N_393,N_309);
nand U453 (N_453,N_415,N_404);
nor U454 (N_454,N_360,N_264);
and U455 (N_455,N_388,N_390);
nand U456 (N_456,N_379,N_403);
nor U457 (N_457,N_411,N_175);
nor U458 (N_458,N_394,N_364);
nor U459 (N_459,N_366,N_9);
nand U460 (N_460,N_397,N_415);
nand U461 (N_461,N_338,N_403);
nor U462 (N_462,N_412,N_395);
and U463 (N_463,N_410,N_395);
or U464 (N_464,N_368,N_410);
nand U465 (N_465,N_303,N_349);
nor U466 (N_466,N_381,N_410);
or U467 (N_467,N_338,N_389);
nand U468 (N_468,N_382,N_366);
nand U469 (N_469,N_338,N_381);
and U470 (N_470,In_284,N_386);
nor U471 (N_471,N_397,N_396);
nand U472 (N_472,N_392,N_367);
or U473 (N_473,N_406,N_375);
nor U474 (N_474,N_363,N_407);
and U475 (N_475,N_409,N_397);
and U476 (N_476,N_349,N_379);
or U477 (N_477,N_414,N_386);
nand U478 (N_478,N_405,N_55);
nand U479 (N_479,N_409,N_311);
nand U480 (N_480,N_450,N_458);
nor U481 (N_481,N_435,N_443);
nand U482 (N_482,N_453,N_447);
or U483 (N_483,N_452,N_436);
or U484 (N_484,N_421,N_459);
nand U485 (N_485,N_475,N_448);
nand U486 (N_486,N_433,N_477);
and U487 (N_487,N_429,N_468);
nand U488 (N_488,N_420,N_455);
nand U489 (N_489,N_469,N_474);
and U490 (N_490,N_457,N_431);
and U491 (N_491,N_444,N_460);
and U492 (N_492,N_476,N_442);
nor U493 (N_493,N_478,N_434);
and U494 (N_494,N_439,N_423);
nand U495 (N_495,N_425,N_430);
and U496 (N_496,N_426,N_428);
nand U497 (N_497,N_451,N_449);
nand U498 (N_498,N_467,N_438);
nand U499 (N_499,N_463,N_427);
or U500 (N_500,N_441,N_473);
nand U501 (N_501,N_446,N_461);
or U502 (N_502,N_470,N_479);
xnor U503 (N_503,N_424,N_445);
nor U504 (N_504,N_422,N_462);
nor U505 (N_505,N_432,N_466);
or U506 (N_506,N_437,N_465);
nor U507 (N_507,N_464,N_440);
nand U508 (N_508,N_471,N_454);
or U509 (N_509,N_472,N_456);
nor U510 (N_510,N_469,N_430);
and U511 (N_511,N_442,N_432);
nand U512 (N_512,N_450,N_479);
or U513 (N_513,N_434,N_438);
nand U514 (N_514,N_430,N_424);
nand U515 (N_515,N_455,N_454);
or U516 (N_516,N_461,N_472);
or U517 (N_517,N_455,N_435);
xor U518 (N_518,N_427,N_458);
nand U519 (N_519,N_432,N_427);
and U520 (N_520,N_455,N_457);
nor U521 (N_521,N_474,N_465);
or U522 (N_522,N_428,N_443);
nor U523 (N_523,N_429,N_469);
nor U524 (N_524,N_452,N_443);
or U525 (N_525,N_430,N_474);
nor U526 (N_526,N_448,N_424);
nor U527 (N_527,N_428,N_448);
nand U528 (N_528,N_454,N_425);
or U529 (N_529,N_420,N_476);
or U530 (N_530,N_426,N_478);
or U531 (N_531,N_433,N_420);
or U532 (N_532,N_423,N_427);
and U533 (N_533,N_470,N_424);
nor U534 (N_534,N_467,N_474);
nor U535 (N_535,N_477,N_424);
or U536 (N_536,N_459,N_422);
nor U537 (N_537,N_443,N_463);
nor U538 (N_538,N_427,N_447);
and U539 (N_539,N_421,N_457);
or U540 (N_540,N_524,N_496);
or U541 (N_541,N_495,N_516);
and U542 (N_542,N_534,N_522);
nand U543 (N_543,N_483,N_539);
nor U544 (N_544,N_525,N_531);
or U545 (N_545,N_500,N_512);
or U546 (N_546,N_503,N_529);
nand U547 (N_547,N_537,N_528);
and U548 (N_548,N_488,N_508);
nand U549 (N_549,N_498,N_499);
nand U550 (N_550,N_504,N_480);
nor U551 (N_551,N_489,N_513);
nand U552 (N_552,N_518,N_519);
nand U553 (N_553,N_538,N_530);
and U554 (N_554,N_514,N_490);
and U555 (N_555,N_492,N_482);
or U556 (N_556,N_497,N_485);
nand U557 (N_557,N_517,N_520);
or U558 (N_558,N_494,N_501);
or U559 (N_559,N_521,N_536);
nor U560 (N_560,N_533,N_502);
nor U561 (N_561,N_506,N_491);
and U562 (N_562,N_487,N_526);
nor U563 (N_563,N_493,N_515);
or U564 (N_564,N_511,N_535);
or U565 (N_565,N_527,N_523);
nand U566 (N_566,N_532,N_509);
nand U567 (N_567,N_484,N_507);
nand U568 (N_568,N_481,N_486);
nor U569 (N_569,N_510,N_505);
nor U570 (N_570,N_539,N_535);
and U571 (N_571,N_516,N_507);
or U572 (N_572,N_528,N_516);
and U573 (N_573,N_496,N_497);
and U574 (N_574,N_488,N_484);
nand U575 (N_575,N_505,N_498);
nand U576 (N_576,N_508,N_516);
nand U577 (N_577,N_502,N_507);
nor U578 (N_578,N_523,N_504);
nor U579 (N_579,N_504,N_506);
nand U580 (N_580,N_506,N_521);
nor U581 (N_581,N_485,N_503);
or U582 (N_582,N_516,N_523);
or U583 (N_583,N_517,N_482);
and U584 (N_584,N_506,N_515);
and U585 (N_585,N_515,N_530);
or U586 (N_586,N_486,N_526);
or U587 (N_587,N_516,N_515);
nor U588 (N_588,N_515,N_505);
nand U589 (N_589,N_495,N_485);
and U590 (N_590,N_524,N_530);
nor U591 (N_591,N_538,N_525);
and U592 (N_592,N_536,N_538);
nor U593 (N_593,N_518,N_505);
nor U594 (N_594,N_490,N_509);
nand U595 (N_595,N_524,N_527);
nor U596 (N_596,N_511,N_507);
or U597 (N_597,N_539,N_517);
or U598 (N_598,N_526,N_537);
or U599 (N_599,N_530,N_526);
nand U600 (N_600,N_563,N_561);
and U601 (N_601,N_565,N_555);
nor U602 (N_602,N_559,N_592);
or U603 (N_603,N_544,N_549);
and U604 (N_604,N_545,N_567);
nand U605 (N_605,N_557,N_540);
and U606 (N_606,N_577,N_598);
or U607 (N_607,N_578,N_576);
nor U608 (N_608,N_582,N_593);
and U609 (N_609,N_568,N_573);
or U610 (N_610,N_597,N_591);
nor U611 (N_611,N_575,N_585);
nor U612 (N_612,N_552,N_580);
nor U613 (N_613,N_572,N_589);
nor U614 (N_614,N_541,N_543);
nand U615 (N_615,N_595,N_566);
nor U616 (N_616,N_586,N_542);
or U617 (N_617,N_550,N_546);
nand U618 (N_618,N_570,N_581);
nand U619 (N_619,N_590,N_569);
nand U620 (N_620,N_547,N_599);
or U621 (N_621,N_574,N_584);
and U622 (N_622,N_551,N_579);
and U623 (N_623,N_588,N_560);
nand U624 (N_624,N_558,N_562);
or U625 (N_625,N_583,N_571);
nor U626 (N_626,N_556,N_553);
nand U627 (N_627,N_587,N_594);
or U628 (N_628,N_596,N_554);
nand U629 (N_629,N_564,N_548);
nand U630 (N_630,N_581,N_542);
and U631 (N_631,N_587,N_591);
nor U632 (N_632,N_552,N_588);
and U633 (N_633,N_592,N_554);
and U634 (N_634,N_592,N_552);
nor U635 (N_635,N_587,N_571);
and U636 (N_636,N_544,N_546);
nor U637 (N_637,N_593,N_544);
and U638 (N_638,N_575,N_599);
nand U639 (N_639,N_554,N_584);
nand U640 (N_640,N_597,N_587);
nand U641 (N_641,N_569,N_586);
nor U642 (N_642,N_598,N_556);
nor U643 (N_643,N_569,N_558);
nand U644 (N_644,N_566,N_596);
nor U645 (N_645,N_564,N_546);
nor U646 (N_646,N_589,N_548);
nor U647 (N_647,N_579,N_554);
and U648 (N_648,N_594,N_589);
or U649 (N_649,N_552,N_570);
xnor U650 (N_650,N_592,N_551);
or U651 (N_651,N_559,N_577);
and U652 (N_652,N_595,N_584);
nor U653 (N_653,N_560,N_556);
or U654 (N_654,N_583,N_559);
or U655 (N_655,N_563,N_567);
nor U656 (N_656,N_598,N_555);
nand U657 (N_657,N_595,N_565);
nand U658 (N_658,N_588,N_563);
nor U659 (N_659,N_593,N_588);
and U660 (N_660,N_642,N_656);
and U661 (N_661,N_657,N_631);
nand U662 (N_662,N_633,N_615);
nor U663 (N_663,N_620,N_607);
and U664 (N_664,N_644,N_641);
nand U665 (N_665,N_622,N_628);
or U666 (N_666,N_611,N_603);
nand U667 (N_667,N_617,N_639);
nor U668 (N_668,N_610,N_646);
nand U669 (N_669,N_613,N_650);
nand U670 (N_670,N_652,N_659);
or U671 (N_671,N_634,N_616);
and U672 (N_672,N_606,N_604);
or U673 (N_673,N_658,N_618);
nand U674 (N_674,N_629,N_637);
nor U675 (N_675,N_653,N_601);
nor U676 (N_676,N_605,N_643);
or U677 (N_677,N_640,N_647);
nor U678 (N_678,N_619,N_636);
and U679 (N_679,N_638,N_632);
nor U680 (N_680,N_649,N_609);
or U681 (N_681,N_600,N_648);
and U682 (N_682,N_602,N_612);
and U683 (N_683,N_655,N_630);
nand U684 (N_684,N_645,N_625);
and U685 (N_685,N_614,N_651);
nor U686 (N_686,N_623,N_635);
nand U687 (N_687,N_608,N_621);
or U688 (N_688,N_627,N_624);
or U689 (N_689,N_654,N_626);
or U690 (N_690,N_606,N_638);
or U691 (N_691,N_615,N_630);
or U692 (N_692,N_608,N_628);
nor U693 (N_693,N_630,N_613);
and U694 (N_694,N_610,N_602);
nor U695 (N_695,N_603,N_635);
and U696 (N_696,N_604,N_645);
nand U697 (N_697,N_622,N_610);
and U698 (N_698,N_613,N_626);
or U699 (N_699,N_643,N_641);
nor U700 (N_700,N_608,N_631);
and U701 (N_701,N_622,N_621);
and U702 (N_702,N_616,N_654);
xnor U703 (N_703,N_623,N_620);
and U704 (N_704,N_640,N_605);
nor U705 (N_705,N_605,N_657);
nand U706 (N_706,N_605,N_603);
xor U707 (N_707,N_659,N_649);
nand U708 (N_708,N_652,N_638);
nand U709 (N_709,N_613,N_614);
and U710 (N_710,N_649,N_603);
nor U711 (N_711,N_641,N_606);
or U712 (N_712,N_647,N_609);
nand U713 (N_713,N_628,N_613);
or U714 (N_714,N_646,N_630);
nand U715 (N_715,N_626,N_656);
nor U716 (N_716,N_617,N_650);
and U717 (N_717,N_651,N_617);
nand U718 (N_718,N_622,N_646);
and U719 (N_719,N_647,N_613);
or U720 (N_720,N_716,N_706);
and U721 (N_721,N_683,N_665);
nor U722 (N_722,N_711,N_708);
or U723 (N_723,N_686,N_674);
or U724 (N_724,N_678,N_663);
nor U725 (N_725,N_673,N_685);
nand U726 (N_726,N_675,N_660);
and U727 (N_727,N_707,N_676);
nand U728 (N_728,N_718,N_669);
nand U729 (N_729,N_679,N_705);
or U730 (N_730,N_687,N_684);
or U731 (N_731,N_661,N_664);
nand U732 (N_732,N_689,N_682);
and U733 (N_733,N_668,N_709);
and U734 (N_734,N_695,N_677);
nor U735 (N_735,N_698,N_681);
nand U736 (N_736,N_712,N_690);
nand U737 (N_737,N_713,N_696);
nor U738 (N_738,N_688,N_691);
and U739 (N_739,N_717,N_697);
or U740 (N_740,N_704,N_693);
or U741 (N_741,N_703,N_700);
nor U742 (N_742,N_672,N_670);
nor U743 (N_743,N_692,N_715);
and U744 (N_744,N_666,N_699);
nor U745 (N_745,N_662,N_702);
and U746 (N_746,N_671,N_701);
nor U747 (N_747,N_714,N_719);
nand U748 (N_748,N_667,N_694);
or U749 (N_749,N_680,N_710);
nor U750 (N_750,N_675,N_674);
nand U751 (N_751,N_687,N_718);
and U752 (N_752,N_683,N_674);
nor U753 (N_753,N_661,N_714);
or U754 (N_754,N_668,N_716);
nand U755 (N_755,N_673,N_708);
and U756 (N_756,N_709,N_715);
nor U757 (N_757,N_690,N_667);
and U758 (N_758,N_705,N_717);
nor U759 (N_759,N_698,N_670);
nand U760 (N_760,N_716,N_698);
nand U761 (N_761,N_706,N_696);
and U762 (N_762,N_705,N_678);
nand U763 (N_763,N_685,N_669);
nand U764 (N_764,N_705,N_709);
and U765 (N_765,N_662,N_684);
nand U766 (N_766,N_696,N_666);
or U767 (N_767,N_674,N_664);
or U768 (N_768,N_680,N_699);
nand U769 (N_769,N_709,N_708);
nor U770 (N_770,N_717,N_700);
nor U771 (N_771,N_660,N_719);
or U772 (N_772,N_704,N_669);
nand U773 (N_773,N_713,N_689);
nand U774 (N_774,N_689,N_706);
nand U775 (N_775,N_718,N_719);
and U776 (N_776,N_714,N_692);
or U777 (N_777,N_704,N_698);
and U778 (N_778,N_718,N_684);
nor U779 (N_779,N_694,N_677);
and U780 (N_780,N_729,N_755);
nand U781 (N_781,N_776,N_771);
or U782 (N_782,N_749,N_745);
or U783 (N_783,N_764,N_746);
and U784 (N_784,N_720,N_735);
nand U785 (N_785,N_747,N_741);
nor U786 (N_786,N_762,N_748);
nand U787 (N_787,N_728,N_721);
or U788 (N_788,N_750,N_736);
or U789 (N_789,N_777,N_772);
and U790 (N_790,N_754,N_737);
nand U791 (N_791,N_739,N_756);
or U792 (N_792,N_765,N_733);
nand U793 (N_793,N_726,N_725);
or U794 (N_794,N_751,N_740);
nor U795 (N_795,N_779,N_724);
nor U796 (N_796,N_727,N_753);
and U797 (N_797,N_723,N_757);
or U798 (N_798,N_738,N_775);
nor U799 (N_799,N_732,N_730);
nand U800 (N_800,N_722,N_773);
nor U801 (N_801,N_731,N_758);
or U802 (N_802,N_742,N_769);
and U803 (N_803,N_778,N_743);
or U804 (N_804,N_770,N_759);
nor U805 (N_805,N_766,N_752);
nand U806 (N_806,N_761,N_734);
and U807 (N_807,N_774,N_744);
and U808 (N_808,N_763,N_767);
and U809 (N_809,N_768,N_760);
or U810 (N_810,N_738,N_732);
nand U811 (N_811,N_748,N_746);
or U812 (N_812,N_751,N_734);
nor U813 (N_813,N_728,N_759);
and U814 (N_814,N_742,N_760);
or U815 (N_815,N_756,N_772);
nand U816 (N_816,N_731,N_740);
nand U817 (N_817,N_749,N_742);
nor U818 (N_818,N_754,N_743);
nand U819 (N_819,N_738,N_768);
nor U820 (N_820,N_777,N_766);
or U821 (N_821,N_775,N_741);
nand U822 (N_822,N_761,N_756);
or U823 (N_823,N_763,N_737);
nor U824 (N_824,N_749,N_733);
nand U825 (N_825,N_762,N_735);
and U826 (N_826,N_728,N_778);
nand U827 (N_827,N_775,N_772);
nor U828 (N_828,N_742,N_754);
nand U829 (N_829,N_752,N_742);
nand U830 (N_830,N_764,N_745);
or U831 (N_831,N_775,N_760);
and U832 (N_832,N_725,N_773);
or U833 (N_833,N_740,N_728);
nand U834 (N_834,N_758,N_773);
nand U835 (N_835,N_720,N_734);
nor U836 (N_836,N_776,N_777);
nand U837 (N_837,N_763,N_765);
nor U838 (N_838,N_775,N_721);
nand U839 (N_839,N_721,N_755);
nand U840 (N_840,N_807,N_827);
nand U841 (N_841,N_836,N_794);
nor U842 (N_842,N_813,N_819);
nor U843 (N_843,N_837,N_793);
and U844 (N_844,N_798,N_828);
or U845 (N_845,N_791,N_839);
or U846 (N_846,N_783,N_832);
and U847 (N_847,N_821,N_809);
or U848 (N_848,N_795,N_784);
nor U849 (N_849,N_834,N_786);
and U850 (N_850,N_790,N_789);
nand U851 (N_851,N_806,N_816);
and U852 (N_852,N_804,N_780);
and U853 (N_853,N_792,N_823);
nand U854 (N_854,N_825,N_785);
and U855 (N_855,N_803,N_824);
nand U856 (N_856,N_812,N_787);
nand U857 (N_857,N_814,N_833);
or U858 (N_858,N_797,N_817);
or U859 (N_859,N_838,N_835);
and U860 (N_860,N_782,N_808);
and U861 (N_861,N_831,N_805);
or U862 (N_862,N_818,N_811);
or U863 (N_863,N_822,N_801);
and U864 (N_864,N_788,N_802);
nand U865 (N_865,N_799,N_800);
nand U866 (N_866,N_830,N_820);
nand U867 (N_867,N_796,N_781);
nor U868 (N_868,N_815,N_810);
or U869 (N_869,N_829,N_826);
nand U870 (N_870,N_831,N_825);
nand U871 (N_871,N_809,N_825);
or U872 (N_872,N_832,N_781);
and U873 (N_873,N_826,N_781);
and U874 (N_874,N_813,N_835);
or U875 (N_875,N_831,N_832);
or U876 (N_876,N_813,N_806);
nand U877 (N_877,N_814,N_819);
and U878 (N_878,N_818,N_822);
nand U879 (N_879,N_796,N_804);
nand U880 (N_880,N_807,N_814);
or U881 (N_881,N_830,N_836);
nor U882 (N_882,N_813,N_834);
nor U883 (N_883,N_792,N_799);
nand U884 (N_884,N_811,N_824);
nor U885 (N_885,N_794,N_833);
or U886 (N_886,N_789,N_784);
or U887 (N_887,N_804,N_839);
or U888 (N_888,N_795,N_820);
and U889 (N_889,N_797,N_799);
and U890 (N_890,N_795,N_821);
or U891 (N_891,N_815,N_804);
and U892 (N_892,N_823,N_819);
or U893 (N_893,N_821,N_801);
nor U894 (N_894,N_821,N_829);
nand U895 (N_895,N_838,N_795);
nor U896 (N_896,N_832,N_819);
and U897 (N_897,N_801,N_818);
xor U898 (N_898,N_806,N_835);
nor U899 (N_899,N_794,N_809);
nand U900 (N_900,N_853,N_886);
or U901 (N_901,N_874,N_848);
or U902 (N_902,N_894,N_860);
nor U903 (N_903,N_840,N_889);
nor U904 (N_904,N_867,N_865);
or U905 (N_905,N_895,N_841);
or U906 (N_906,N_887,N_876);
nor U907 (N_907,N_862,N_890);
and U908 (N_908,N_880,N_854);
and U909 (N_909,N_863,N_879);
and U910 (N_910,N_845,N_870);
and U911 (N_911,N_843,N_851);
nor U912 (N_912,N_892,N_884);
nand U913 (N_913,N_877,N_885);
or U914 (N_914,N_849,N_855);
or U915 (N_915,N_858,N_847);
nor U916 (N_916,N_857,N_872);
or U917 (N_917,N_844,N_846);
and U918 (N_918,N_852,N_842);
or U919 (N_919,N_871,N_899);
nor U920 (N_920,N_864,N_882);
or U921 (N_921,N_869,N_888);
or U922 (N_922,N_898,N_875);
nor U923 (N_923,N_897,N_891);
nor U924 (N_924,N_881,N_856);
or U925 (N_925,N_878,N_868);
nor U926 (N_926,N_873,N_850);
and U927 (N_927,N_893,N_896);
or U928 (N_928,N_883,N_859);
nor U929 (N_929,N_861,N_866);
nand U930 (N_930,N_895,N_882);
nor U931 (N_931,N_878,N_883);
nor U932 (N_932,N_852,N_846);
nand U933 (N_933,N_885,N_895);
or U934 (N_934,N_880,N_881);
or U935 (N_935,N_894,N_881);
and U936 (N_936,N_841,N_871);
nand U937 (N_937,N_872,N_895);
nor U938 (N_938,N_895,N_879);
nor U939 (N_939,N_897,N_876);
and U940 (N_940,N_890,N_865);
or U941 (N_941,N_847,N_896);
and U942 (N_942,N_844,N_853);
nor U943 (N_943,N_840,N_875);
nand U944 (N_944,N_869,N_850);
or U945 (N_945,N_862,N_870);
xnor U946 (N_946,N_851,N_877);
or U947 (N_947,N_851,N_846);
or U948 (N_948,N_878,N_854);
nor U949 (N_949,N_844,N_866);
and U950 (N_950,N_846,N_861);
or U951 (N_951,N_850,N_867);
nor U952 (N_952,N_892,N_847);
and U953 (N_953,N_851,N_896);
or U954 (N_954,N_885,N_845);
or U955 (N_955,N_840,N_871);
or U956 (N_956,N_849,N_881);
or U957 (N_957,N_891,N_844);
or U958 (N_958,N_889,N_845);
nor U959 (N_959,N_899,N_887);
or U960 (N_960,N_915,N_954);
or U961 (N_961,N_948,N_939);
nand U962 (N_962,N_937,N_919);
or U963 (N_963,N_909,N_914);
nor U964 (N_964,N_941,N_924);
nor U965 (N_965,N_947,N_903);
nor U966 (N_966,N_906,N_957);
and U967 (N_967,N_932,N_951);
and U968 (N_968,N_916,N_912);
or U969 (N_969,N_905,N_911);
and U970 (N_970,N_904,N_940);
and U971 (N_971,N_925,N_949);
or U972 (N_972,N_950,N_921);
and U973 (N_973,N_928,N_938);
nand U974 (N_974,N_901,N_959);
nor U975 (N_975,N_929,N_933);
and U976 (N_976,N_955,N_953);
nand U977 (N_977,N_910,N_902);
and U978 (N_978,N_952,N_917);
or U979 (N_979,N_923,N_918);
nand U980 (N_980,N_900,N_931);
nor U981 (N_981,N_945,N_943);
nand U982 (N_982,N_930,N_934);
nand U983 (N_983,N_935,N_956);
or U984 (N_984,N_920,N_907);
nand U985 (N_985,N_908,N_944);
nand U986 (N_986,N_922,N_958);
or U987 (N_987,N_936,N_926);
nor U988 (N_988,N_942,N_927);
or U989 (N_989,N_913,N_946);
nand U990 (N_990,N_951,N_905);
nand U991 (N_991,N_951,N_940);
nor U992 (N_992,N_920,N_940);
and U993 (N_993,N_949,N_905);
and U994 (N_994,N_907,N_919);
or U995 (N_995,N_924,N_933);
nor U996 (N_996,N_948,N_934);
nand U997 (N_997,N_954,N_905);
and U998 (N_998,N_944,N_926);
nand U999 (N_999,N_945,N_941);
or U1000 (N_1000,N_947,N_904);
nor U1001 (N_1001,N_955,N_934);
xor U1002 (N_1002,N_912,N_904);
and U1003 (N_1003,N_916,N_915);
xnor U1004 (N_1004,N_931,N_912);
and U1005 (N_1005,N_903,N_909);
or U1006 (N_1006,N_959,N_922);
nor U1007 (N_1007,N_952,N_918);
nand U1008 (N_1008,N_938,N_904);
nor U1009 (N_1009,N_923,N_942);
xnor U1010 (N_1010,N_944,N_943);
or U1011 (N_1011,N_947,N_910);
nor U1012 (N_1012,N_944,N_905);
and U1013 (N_1013,N_930,N_925);
nor U1014 (N_1014,N_926,N_946);
or U1015 (N_1015,N_950,N_930);
and U1016 (N_1016,N_944,N_911);
nand U1017 (N_1017,N_940,N_918);
nor U1018 (N_1018,N_911,N_937);
nand U1019 (N_1019,N_951,N_925);
or U1020 (N_1020,N_971,N_1016);
nand U1021 (N_1021,N_995,N_980);
and U1022 (N_1022,N_1013,N_1009);
and U1023 (N_1023,N_975,N_1012);
nor U1024 (N_1024,N_973,N_962);
or U1025 (N_1025,N_1014,N_1000);
nor U1026 (N_1026,N_961,N_998);
nor U1027 (N_1027,N_997,N_981);
nand U1028 (N_1028,N_1005,N_1015);
and U1029 (N_1029,N_1017,N_970);
nand U1030 (N_1030,N_977,N_990);
nor U1031 (N_1031,N_984,N_965);
and U1032 (N_1032,N_960,N_982);
or U1033 (N_1033,N_1006,N_974);
or U1034 (N_1034,N_991,N_987);
nand U1035 (N_1035,N_1001,N_993);
nor U1036 (N_1036,N_967,N_969);
and U1037 (N_1037,N_983,N_988);
nor U1038 (N_1038,N_968,N_978);
nor U1039 (N_1039,N_1004,N_999);
xor U1040 (N_1040,N_1011,N_966);
or U1041 (N_1041,N_963,N_979);
xnor U1042 (N_1042,N_989,N_1018);
nor U1043 (N_1043,N_1019,N_1003);
or U1044 (N_1044,N_992,N_1010);
nor U1045 (N_1045,N_985,N_976);
or U1046 (N_1046,N_986,N_1007);
nand U1047 (N_1047,N_996,N_1002);
and U1048 (N_1048,N_994,N_1008);
nand U1049 (N_1049,N_972,N_964);
nor U1050 (N_1050,N_1017,N_1011);
nor U1051 (N_1051,N_965,N_1010);
or U1052 (N_1052,N_1002,N_991);
or U1053 (N_1053,N_983,N_965);
or U1054 (N_1054,N_962,N_991);
and U1055 (N_1055,N_996,N_970);
nor U1056 (N_1056,N_1013,N_1018);
or U1057 (N_1057,N_1008,N_996);
or U1058 (N_1058,N_986,N_961);
nand U1059 (N_1059,N_987,N_1016);
and U1060 (N_1060,N_983,N_996);
nand U1061 (N_1061,N_1002,N_1008);
nand U1062 (N_1062,N_981,N_984);
nor U1063 (N_1063,N_985,N_961);
xnor U1064 (N_1064,N_1016,N_1002);
and U1065 (N_1065,N_987,N_1013);
nor U1066 (N_1066,N_1000,N_989);
nand U1067 (N_1067,N_1005,N_970);
nand U1068 (N_1068,N_960,N_1011);
and U1069 (N_1069,N_969,N_1018);
or U1070 (N_1070,N_1013,N_968);
and U1071 (N_1071,N_987,N_981);
nand U1072 (N_1072,N_1009,N_992);
and U1073 (N_1073,N_973,N_992);
nand U1074 (N_1074,N_996,N_1009);
nand U1075 (N_1075,N_996,N_1006);
or U1076 (N_1076,N_983,N_990);
and U1077 (N_1077,N_1010,N_1003);
nor U1078 (N_1078,N_1002,N_1015);
nor U1079 (N_1079,N_995,N_1005);
or U1080 (N_1080,N_1067,N_1044);
and U1081 (N_1081,N_1060,N_1052);
nand U1082 (N_1082,N_1032,N_1074);
nand U1083 (N_1083,N_1045,N_1072);
nor U1084 (N_1084,N_1049,N_1030);
xor U1085 (N_1085,N_1037,N_1048);
or U1086 (N_1086,N_1068,N_1057);
and U1087 (N_1087,N_1065,N_1054);
and U1088 (N_1088,N_1022,N_1042);
and U1089 (N_1089,N_1028,N_1079);
nor U1090 (N_1090,N_1035,N_1040);
and U1091 (N_1091,N_1043,N_1021);
or U1092 (N_1092,N_1077,N_1033);
nand U1093 (N_1093,N_1073,N_1031);
nand U1094 (N_1094,N_1034,N_1027);
and U1095 (N_1095,N_1023,N_1039);
or U1096 (N_1096,N_1061,N_1020);
nand U1097 (N_1097,N_1041,N_1050);
and U1098 (N_1098,N_1051,N_1063);
nor U1099 (N_1099,N_1059,N_1029);
and U1100 (N_1100,N_1076,N_1078);
or U1101 (N_1101,N_1066,N_1070);
and U1102 (N_1102,N_1055,N_1064);
nand U1103 (N_1103,N_1046,N_1071);
and U1104 (N_1104,N_1026,N_1062);
nor U1105 (N_1105,N_1069,N_1058);
and U1106 (N_1106,N_1056,N_1024);
nand U1107 (N_1107,N_1036,N_1025);
or U1108 (N_1108,N_1047,N_1053);
nor U1109 (N_1109,N_1075,N_1038);
nand U1110 (N_1110,N_1044,N_1056);
nand U1111 (N_1111,N_1029,N_1056);
and U1112 (N_1112,N_1077,N_1064);
and U1113 (N_1113,N_1044,N_1078);
nor U1114 (N_1114,N_1079,N_1056);
or U1115 (N_1115,N_1048,N_1041);
nand U1116 (N_1116,N_1050,N_1070);
and U1117 (N_1117,N_1067,N_1054);
and U1118 (N_1118,N_1033,N_1029);
or U1119 (N_1119,N_1034,N_1054);
or U1120 (N_1120,N_1052,N_1069);
nand U1121 (N_1121,N_1020,N_1024);
xnor U1122 (N_1122,N_1067,N_1073);
and U1123 (N_1123,N_1047,N_1023);
nand U1124 (N_1124,N_1054,N_1070);
nor U1125 (N_1125,N_1031,N_1034);
nand U1126 (N_1126,N_1066,N_1025);
nor U1127 (N_1127,N_1030,N_1051);
nor U1128 (N_1128,N_1033,N_1025);
nor U1129 (N_1129,N_1023,N_1036);
or U1130 (N_1130,N_1074,N_1033);
nand U1131 (N_1131,N_1059,N_1063);
nor U1132 (N_1132,N_1028,N_1040);
or U1133 (N_1133,N_1079,N_1035);
nand U1134 (N_1134,N_1071,N_1077);
nand U1135 (N_1135,N_1049,N_1020);
and U1136 (N_1136,N_1047,N_1069);
nand U1137 (N_1137,N_1050,N_1067);
and U1138 (N_1138,N_1043,N_1027);
nand U1139 (N_1139,N_1039,N_1025);
nor U1140 (N_1140,N_1137,N_1120);
nor U1141 (N_1141,N_1100,N_1135);
nand U1142 (N_1142,N_1133,N_1086);
nand U1143 (N_1143,N_1102,N_1127);
or U1144 (N_1144,N_1091,N_1081);
and U1145 (N_1145,N_1129,N_1109);
and U1146 (N_1146,N_1085,N_1088);
or U1147 (N_1147,N_1096,N_1128);
nor U1148 (N_1148,N_1087,N_1117);
nand U1149 (N_1149,N_1115,N_1095);
nand U1150 (N_1150,N_1094,N_1080);
nand U1151 (N_1151,N_1098,N_1104);
nor U1152 (N_1152,N_1110,N_1125);
nor U1153 (N_1153,N_1103,N_1092);
or U1154 (N_1154,N_1099,N_1093);
nand U1155 (N_1155,N_1134,N_1112);
nor U1156 (N_1156,N_1089,N_1126);
nand U1157 (N_1157,N_1124,N_1131);
nor U1158 (N_1158,N_1105,N_1106);
and U1159 (N_1159,N_1122,N_1123);
or U1160 (N_1160,N_1090,N_1107);
and U1161 (N_1161,N_1083,N_1114);
and U1162 (N_1162,N_1082,N_1111);
or U1163 (N_1163,N_1116,N_1136);
xor U1164 (N_1164,N_1132,N_1119);
nand U1165 (N_1165,N_1084,N_1097);
or U1166 (N_1166,N_1139,N_1138);
nor U1167 (N_1167,N_1108,N_1113);
nor U1168 (N_1168,N_1118,N_1101);
nor U1169 (N_1169,N_1130,N_1121);
or U1170 (N_1170,N_1137,N_1116);
and U1171 (N_1171,N_1139,N_1103);
and U1172 (N_1172,N_1099,N_1121);
and U1173 (N_1173,N_1113,N_1087);
nand U1174 (N_1174,N_1089,N_1094);
and U1175 (N_1175,N_1090,N_1126);
and U1176 (N_1176,N_1086,N_1120);
nor U1177 (N_1177,N_1128,N_1102);
or U1178 (N_1178,N_1087,N_1128);
and U1179 (N_1179,N_1133,N_1084);
nand U1180 (N_1180,N_1125,N_1087);
nand U1181 (N_1181,N_1107,N_1137);
or U1182 (N_1182,N_1087,N_1080);
or U1183 (N_1183,N_1134,N_1132);
or U1184 (N_1184,N_1098,N_1105);
nor U1185 (N_1185,N_1099,N_1133);
or U1186 (N_1186,N_1081,N_1088);
or U1187 (N_1187,N_1131,N_1087);
nand U1188 (N_1188,N_1093,N_1124);
nand U1189 (N_1189,N_1129,N_1115);
nor U1190 (N_1190,N_1090,N_1096);
and U1191 (N_1191,N_1107,N_1098);
and U1192 (N_1192,N_1095,N_1105);
or U1193 (N_1193,N_1096,N_1131);
nor U1194 (N_1194,N_1128,N_1115);
nor U1195 (N_1195,N_1112,N_1080);
nand U1196 (N_1196,N_1110,N_1086);
or U1197 (N_1197,N_1134,N_1084);
nor U1198 (N_1198,N_1109,N_1107);
and U1199 (N_1199,N_1111,N_1098);
and U1200 (N_1200,N_1153,N_1195);
nand U1201 (N_1201,N_1154,N_1156);
nand U1202 (N_1202,N_1143,N_1172);
nand U1203 (N_1203,N_1142,N_1149);
and U1204 (N_1204,N_1176,N_1150);
and U1205 (N_1205,N_1180,N_1191);
or U1206 (N_1206,N_1160,N_1163);
and U1207 (N_1207,N_1173,N_1165);
nor U1208 (N_1208,N_1140,N_1175);
and U1209 (N_1209,N_1187,N_1144);
nand U1210 (N_1210,N_1198,N_1147);
and U1211 (N_1211,N_1157,N_1158);
or U1212 (N_1212,N_1178,N_1188);
nor U1213 (N_1213,N_1171,N_1168);
or U1214 (N_1214,N_1192,N_1152);
or U1215 (N_1215,N_1181,N_1170);
or U1216 (N_1216,N_1196,N_1177);
and U1217 (N_1217,N_1179,N_1161);
and U1218 (N_1218,N_1194,N_1182);
or U1219 (N_1219,N_1184,N_1185);
and U1220 (N_1220,N_1167,N_1166);
nor U1221 (N_1221,N_1145,N_1174);
and U1222 (N_1222,N_1186,N_1183);
nor U1223 (N_1223,N_1164,N_1190);
and U1224 (N_1224,N_1159,N_1193);
nand U1225 (N_1225,N_1141,N_1199);
nand U1226 (N_1226,N_1151,N_1162);
nor U1227 (N_1227,N_1197,N_1148);
nor U1228 (N_1228,N_1146,N_1155);
or U1229 (N_1229,N_1189,N_1169);
nand U1230 (N_1230,N_1140,N_1174);
nand U1231 (N_1231,N_1170,N_1192);
nand U1232 (N_1232,N_1161,N_1142);
or U1233 (N_1233,N_1179,N_1178);
or U1234 (N_1234,N_1146,N_1160);
and U1235 (N_1235,N_1161,N_1169);
nand U1236 (N_1236,N_1173,N_1197);
nor U1237 (N_1237,N_1173,N_1142);
nand U1238 (N_1238,N_1169,N_1190);
or U1239 (N_1239,N_1185,N_1197);
and U1240 (N_1240,N_1144,N_1148);
or U1241 (N_1241,N_1146,N_1164);
nor U1242 (N_1242,N_1175,N_1178);
and U1243 (N_1243,N_1178,N_1148);
nor U1244 (N_1244,N_1153,N_1152);
nor U1245 (N_1245,N_1151,N_1157);
nand U1246 (N_1246,N_1168,N_1183);
and U1247 (N_1247,N_1159,N_1175);
nor U1248 (N_1248,N_1164,N_1169);
or U1249 (N_1249,N_1175,N_1195);
and U1250 (N_1250,N_1179,N_1155);
and U1251 (N_1251,N_1149,N_1141);
nor U1252 (N_1252,N_1182,N_1174);
nor U1253 (N_1253,N_1146,N_1142);
nand U1254 (N_1254,N_1150,N_1190);
nor U1255 (N_1255,N_1175,N_1188);
or U1256 (N_1256,N_1153,N_1194);
and U1257 (N_1257,N_1170,N_1182);
or U1258 (N_1258,N_1198,N_1150);
and U1259 (N_1259,N_1169,N_1182);
or U1260 (N_1260,N_1240,N_1212);
nand U1261 (N_1261,N_1213,N_1252);
or U1262 (N_1262,N_1249,N_1250);
nand U1263 (N_1263,N_1239,N_1218);
or U1264 (N_1264,N_1256,N_1214);
nand U1265 (N_1265,N_1235,N_1246);
nand U1266 (N_1266,N_1200,N_1257);
nand U1267 (N_1267,N_1242,N_1222);
nand U1268 (N_1268,N_1208,N_1238);
or U1269 (N_1269,N_1248,N_1211);
nor U1270 (N_1270,N_1234,N_1226);
or U1271 (N_1271,N_1227,N_1229);
nand U1272 (N_1272,N_1228,N_1232);
xor U1273 (N_1273,N_1258,N_1247);
nand U1274 (N_1274,N_1224,N_1216);
nor U1275 (N_1275,N_1236,N_1206);
nor U1276 (N_1276,N_1201,N_1230);
nor U1277 (N_1277,N_1204,N_1209);
or U1278 (N_1278,N_1245,N_1203);
nand U1279 (N_1279,N_1241,N_1217);
or U1280 (N_1280,N_1205,N_1244);
and U1281 (N_1281,N_1221,N_1255);
nor U1282 (N_1282,N_1237,N_1202);
nor U1283 (N_1283,N_1259,N_1243);
nand U1284 (N_1284,N_1207,N_1215);
and U1285 (N_1285,N_1253,N_1223);
or U1286 (N_1286,N_1220,N_1225);
nor U1287 (N_1287,N_1219,N_1210);
and U1288 (N_1288,N_1231,N_1251);
or U1289 (N_1289,N_1254,N_1233);
or U1290 (N_1290,N_1212,N_1238);
and U1291 (N_1291,N_1245,N_1200);
or U1292 (N_1292,N_1237,N_1215);
or U1293 (N_1293,N_1245,N_1209);
and U1294 (N_1294,N_1240,N_1219);
nor U1295 (N_1295,N_1205,N_1256);
or U1296 (N_1296,N_1231,N_1223);
nand U1297 (N_1297,N_1255,N_1205);
and U1298 (N_1298,N_1228,N_1225);
nor U1299 (N_1299,N_1257,N_1234);
and U1300 (N_1300,N_1207,N_1219);
xor U1301 (N_1301,N_1255,N_1248);
and U1302 (N_1302,N_1220,N_1248);
nand U1303 (N_1303,N_1247,N_1222);
and U1304 (N_1304,N_1213,N_1206);
nor U1305 (N_1305,N_1223,N_1228);
nor U1306 (N_1306,N_1246,N_1242);
or U1307 (N_1307,N_1246,N_1244);
and U1308 (N_1308,N_1236,N_1219);
nand U1309 (N_1309,N_1230,N_1203);
or U1310 (N_1310,N_1252,N_1228);
or U1311 (N_1311,N_1215,N_1209);
or U1312 (N_1312,N_1256,N_1231);
or U1313 (N_1313,N_1216,N_1237);
or U1314 (N_1314,N_1259,N_1210);
or U1315 (N_1315,N_1223,N_1225);
nor U1316 (N_1316,N_1240,N_1257);
or U1317 (N_1317,N_1212,N_1252);
and U1318 (N_1318,N_1246,N_1247);
or U1319 (N_1319,N_1251,N_1219);
nand U1320 (N_1320,N_1307,N_1291);
and U1321 (N_1321,N_1311,N_1292);
nor U1322 (N_1322,N_1270,N_1284);
or U1323 (N_1323,N_1276,N_1308);
nand U1324 (N_1324,N_1314,N_1267);
nand U1325 (N_1325,N_1301,N_1266);
and U1326 (N_1326,N_1319,N_1296);
nand U1327 (N_1327,N_1306,N_1281);
or U1328 (N_1328,N_1300,N_1287);
and U1329 (N_1329,N_1290,N_1268);
nor U1330 (N_1330,N_1318,N_1263);
and U1331 (N_1331,N_1305,N_1278);
nor U1332 (N_1332,N_1262,N_1299);
nor U1333 (N_1333,N_1295,N_1269);
or U1334 (N_1334,N_1273,N_1265);
or U1335 (N_1335,N_1285,N_1275);
and U1336 (N_1336,N_1317,N_1303);
nand U1337 (N_1337,N_1313,N_1260);
or U1338 (N_1338,N_1286,N_1293);
nor U1339 (N_1339,N_1315,N_1316);
or U1340 (N_1340,N_1274,N_1302);
nor U1341 (N_1341,N_1289,N_1261);
or U1342 (N_1342,N_1282,N_1310);
or U1343 (N_1343,N_1304,N_1277);
and U1344 (N_1344,N_1264,N_1280);
xnor U1345 (N_1345,N_1271,N_1297);
or U1346 (N_1346,N_1312,N_1283);
or U1347 (N_1347,N_1272,N_1309);
or U1348 (N_1348,N_1294,N_1298);
and U1349 (N_1349,N_1279,N_1288);
nand U1350 (N_1350,N_1312,N_1285);
and U1351 (N_1351,N_1318,N_1309);
nand U1352 (N_1352,N_1262,N_1286);
and U1353 (N_1353,N_1277,N_1314);
nor U1354 (N_1354,N_1305,N_1292);
or U1355 (N_1355,N_1310,N_1318);
nor U1356 (N_1356,N_1261,N_1288);
nand U1357 (N_1357,N_1303,N_1269);
or U1358 (N_1358,N_1314,N_1291);
nand U1359 (N_1359,N_1311,N_1282);
or U1360 (N_1360,N_1263,N_1317);
nor U1361 (N_1361,N_1267,N_1265);
and U1362 (N_1362,N_1291,N_1305);
or U1363 (N_1363,N_1271,N_1278);
nand U1364 (N_1364,N_1301,N_1283);
and U1365 (N_1365,N_1271,N_1283);
and U1366 (N_1366,N_1307,N_1286);
nor U1367 (N_1367,N_1318,N_1304);
and U1368 (N_1368,N_1309,N_1266);
nand U1369 (N_1369,N_1303,N_1292);
nand U1370 (N_1370,N_1307,N_1279);
and U1371 (N_1371,N_1262,N_1289);
nor U1372 (N_1372,N_1270,N_1294);
and U1373 (N_1373,N_1264,N_1270);
nand U1374 (N_1374,N_1290,N_1280);
nor U1375 (N_1375,N_1262,N_1318);
nor U1376 (N_1376,N_1284,N_1278);
and U1377 (N_1377,N_1299,N_1307);
nor U1378 (N_1378,N_1307,N_1272);
nand U1379 (N_1379,N_1285,N_1300);
nand U1380 (N_1380,N_1324,N_1377);
and U1381 (N_1381,N_1329,N_1357);
or U1382 (N_1382,N_1344,N_1333);
and U1383 (N_1383,N_1355,N_1368);
or U1384 (N_1384,N_1332,N_1367);
and U1385 (N_1385,N_1337,N_1365);
or U1386 (N_1386,N_1334,N_1353);
and U1387 (N_1387,N_1340,N_1335);
nor U1388 (N_1388,N_1328,N_1378);
or U1389 (N_1389,N_1343,N_1366);
or U1390 (N_1390,N_1320,N_1373);
and U1391 (N_1391,N_1360,N_1331);
or U1392 (N_1392,N_1358,N_1356);
nor U1393 (N_1393,N_1327,N_1321);
nor U1394 (N_1394,N_1379,N_1359);
nor U1395 (N_1395,N_1325,N_1372);
nor U1396 (N_1396,N_1323,N_1350);
nor U1397 (N_1397,N_1341,N_1351);
or U1398 (N_1398,N_1336,N_1347);
nand U1399 (N_1399,N_1345,N_1330);
nor U1400 (N_1400,N_1376,N_1338);
nand U1401 (N_1401,N_1369,N_1374);
nor U1402 (N_1402,N_1364,N_1375);
and U1403 (N_1403,N_1339,N_1363);
nand U1404 (N_1404,N_1370,N_1371);
and U1405 (N_1405,N_1354,N_1326);
nand U1406 (N_1406,N_1346,N_1349);
and U1407 (N_1407,N_1352,N_1348);
nor U1408 (N_1408,N_1342,N_1322);
and U1409 (N_1409,N_1362,N_1361);
or U1410 (N_1410,N_1356,N_1339);
and U1411 (N_1411,N_1354,N_1322);
nand U1412 (N_1412,N_1373,N_1363);
and U1413 (N_1413,N_1341,N_1379);
nand U1414 (N_1414,N_1328,N_1367);
nand U1415 (N_1415,N_1352,N_1340);
or U1416 (N_1416,N_1378,N_1340);
and U1417 (N_1417,N_1372,N_1349);
or U1418 (N_1418,N_1320,N_1375);
nand U1419 (N_1419,N_1336,N_1331);
nor U1420 (N_1420,N_1379,N_1353);
nand U1421 (N_1421,N_1340,N_1370);
and U1422 (N_1422,N_1336,N_1329);
or U1423 (N_1423,N_1322,N_1379);
or U1424 (N_1424,N_1351,N_1347);
xnor U1425 (N_1425,N_1347,N_1370);
nor U1426 (N_1426,N_1335,N_1336);
and U1427 (N_1427,N_1360,N_1356);
or U1428 (N_1428,N_1368,N_1376);
nor U1429 (N_1429,N_1369,N_1329);
and U1430 (N_1430,N_1326,N_1357);
and U1431 (N_1431,N_1371,N_1326);
nor U1432 (N_1432,N_1340,N_1325);
and U1433 (N_1433,N_1344,N_1352);
nand U1434 (N_1434,N_1367,N_1355);
nor U1435 (N_1435,N_1374,N_1354);
nand U1436 (N_1436,N_1355,N_1349);
or U1437 (N_1437,N_1372,N_1348);
nor U1438 (N_1438,N_1361,N_1376);
nand U1439 (N_1439,N_1331,N_1342);
and U1440 (N_1440,N_1407,N_1380);
and U1441 (N_1441,N_1394,N_1406);
nand U1442 (N_1442,N_1382,N_1414);
and U1443 (N_1443,N_1392,N_1385);
nor U1444 (N_1444,N_1415,N_1421);
nor U1445 (N_1445,N_1410,N_1426);
nand U1446 (N_1446,N_1416,N_1436);
and U1447 (N_1447,N_1428,N_1393);
or U1448 (N_1448,N_1413,N_1386);
and U1449 (N_1449,N_1391,N_1390);
or U1450 (N_1450,N_1418,N_1425);
nand U1451 (N_1451,N_1429,N_1408);
nand U1452 (N_1452,N_1389,N_1387);
and U1453 (N_1453,N_1422,N_1395);
nand U1454 (N_1454,N_1396,N_1405);
nor U1455 (N_1455,N_1401,N_1397);
nand U1456 (N_1456,N_1432,N_1411);
nand U1457 (N_1457,N_1431,N_1409);
and U1458 (N_1458,N_1381,N_1417);
or U1459 (N_1459,N_1412,N_1402);
or U1460 (N_1460,N_1427,N_1398);
nor U1461 (N_1461,N_1419,N_1435);
or U1462 (N_1462,N_1388,N_1403);
and U1463 (N_1463,N_1433,N_1423);
nand U1464 (N_1464,N_1420,N_1399);
and U1465 (N_1465,N_1434,N_1437);
nor U1466 (N_1466,N_1424,N_1439);
or U1467 (N_1467,N_1384,N_1438);
or U1468 (N_1468,N_1404,N_1400);
nand U1469 (N_1469,N_1430,N_1383);
and U1470 (N_1470,N_1395,N_1392);
nand U1471 (N_1471,N_1394,N_1410);
nand U1472 (N_1472,N_1417,N_1391);
or U1473 (N_1473,N_1413,N_1418);
and U1474 (N_1474,N_1427,N_1418);
nand U1475 (N_1475,N_1429,N_1401);
nand U1476 (N_1476,N_1399,N_1423);
or U1477 (N_1477,N_1406,N_1390);
and U1478 (N_1478,N_1388,N_1387);
or U1479 (N_1479,N_1428,N_1418);
nor U1480 (N_1480,N_1404,N_1382);
or U1481 (N_1481,N_1401,N_1435);
and U1482 (N_1482,N_1410,N_1421);
or U1483 (N_1483,N_1381,N_1389);
nor U1484 (N_1484,N_1432,N_1418);
and U1485 (N_1485,N_1382,N_1397);
nor U1486 (N_1486,N_1389,N_1409);
nor U1487 (N_1487,N_1433,N_1425);
and U1488 (N_1488,N_1389,N_1395);
and U1489 (N_1489,N_1434,N_1430);
nor U1490 (N_1490,N_1381,N_1407);
and U1491 (N_1491,N_1386,N_1418);
and U1492 (N_1492,N_1423,N_1409);
or U1493 (N_1493,N_1385,N_1406);
or U1494 (N_1494,N_1381,N_1422);
xnor U1495 (N_1495,N_1429,N_1415);
and U1496 (N_1496,N_1391,N_1392);
nor U1497 (N_1497,N_1403,N_1412);
nor U1498 (N_1498,N_1386,N_1405);
nand U1499 (N_1499,N_1438,N_1401);
nand U1500 (N_1500,N_1465,N_1485);
nor U1501 (N_1501,N_1443,N_1449);
and U1502 (N_1502,N_1466,N_1458);
and U1503 (N_1503,N_1473,N_1451);
nor U1504 (N_1504,N_1471,N_1462);
nor U1505 (N_1505,N_1487,N_1459);
nor U1506 (N_1506,N_1491,N_1482);
or U1507 (N_1507,N_1444,N_1452);
or U1508 (N_1508,N_1460,N_1484);
and U1509 (N_1509,N_1486,N_1497);
nor U1510 (N_1510,N_1464,N_1499);
nand U1511 (N_1511,N_1468,N_1474);
nand U1512 (N_1512,N_1496,N_1475);
nor U1513 (N_1513,N_1461,N_1489);
nor U1514 (N_1514,N_1472,N_1483);
nand U1515 (N_1515,N_1481,N_1490);
nor U1516 (N_1516,N_1442,N_1453);
nor U1517 (N_1517,N_1492,N_1445);
and U1518 (N_1518,N_1446,N_1457);
or U1519 (N_1519,N_1450,N_1456);
and U1520 (N_1520,N_1447,N_1448);
nor U1521 (N_1521,N_1493,N_1469);
nor U1522 (N_1522,N_1494,N_1498);
nor U1523 (N_1523,N_1477,N_1467);
or U1524 (N_1524,N_1454,N_1479);
nand U1525 (N_1525,N_1478,N_1455);
or U1526 (N_1526,N_1488,N_1463);
nand U1527 (N_1527,N_1440,N_1480);
nor U1528 (N_1528,N_1441,N_1470);
and U1529 (N_1529,N_1495,N_1476);
or U1530 (N_1530,N_1479,N_1490);
and U1531 (N_1531,N_1449,N_1481);
nor U1532 (N_1532,N_1473,N_1481);
or U1533 (N_1533,N_1476,N_1482);
nand U1534 (N_1534,N_1487,N_1451);
and U1535 (N_1535,N_1471,N_1453);
nor U1536 (N_1536,N_1442,N_1491);
and U1537 (N_1537,N_1492,N_1498);
and U1538 (N_1538,N_1443,N_1490);
nor U1539 (N_1539,N_1478,N_1469);
and U1540 (N_1540,N_1453,N_1445);
nand U1541 (N_1541,N_1465,N_1451);
xor U1542 (N_1542,N_1493,N_1452);
nor U1543 (N_1543,N_1462,N_1478);
and U1544 (N_1544,N_1487,N_1475);
xor U1545 (N_1545,N_1453,N_1448);
or U1546 (N_1546,N_1469,N_1468);
nand U1547 (N_1547,N_1471,N_1457);
and U1548 (N_1548,N_1471,N_1467);
nand U1549 (N_1549,N_1470,N_1462);
and U1550 (N_1550,N_1470,N_1447);
or U1551 (N_1551,N_1464,N_1475);
nand U1552 (N_1552,N_1468,N_1487);
and U1553 (N_1553,N_1482,N_1441);
or U1554 (N_1554,N_1455,N_1473);
and U1555 (N_1555,N_1451,N_1472);
nand U1556 (N_1556,N_1456,N_1467);
nor U1557 (N_1557,N_1448,N_1476);
or U1558 (N_1558,N_1479,N_1465);
nand U1559 (N_1559,N_1467,N_1490);
nor U1560 (N_1560,N_1520,N_1541);
nand U1561 (N_1561,N_1546,N_1504);
nand U1562 (N_1562,N_1527,N_1508);
or U1563 (N_1563,N_1531,N_1507);
or U1564 (N_1564,N_1514,N_1551);
or U1565 (N_1565,N_1532,N_1555);
and U1566 (N_1566,N_1529,N_1519);
nand U1567 (N_1567,N_1559,N_1534);
nand U1568 (N_1568,N_1538,N_1525);
or U1569 (N_1569,N_1548,N_1524);
and U1570 (N_1570,N_1509,N_1513);
xor U1571 (N_1571,N_1521,N_1556);
or U1572 (N_1572,N_1539,N_1500);
nand U1573 (N_1573,N_1549,N_1503);
or U1574 (N_1574,N_1516,N_1501);
and U1575 (N_1575,N_1505,N_1550);
or U1576 (N_1576,N_1518,N_1533);
nand U1577 (N_1577,N_1543,N_1552);
nand U1578 (N_1578,N_1547,N_1542);
nor U1579 (N_1579,N_1517,N_1511);
nand U1580 (N_1580,N_1558,N_1540);
or U1581 (N_1581,N_1554,N_1506);
or U1582 (N_1582,N_1545,N_1557);
nor U1583 (N_1583,N_1537,N_1522);
nand U1584 (N_1584,N_1544,N_1510);
nor U1585 (N_1585,N_1515,N_1523);
or U1586 (N_1586,N_1530,N_1536);
nand U1587 (N_1587,N_1502,N_1526);
or U1588 (N_1588,N_1512,N_1535);
and U1589 (N_1589,N_1553,N_1528);
and U1590 (N_1590,N_1526,N_1508);
and U1591 (N_1591,N_1556,N_1502);
nand U1592 (N_1592,N_1513,N_1541);
or U1593 (N_1593,N_1507,N_1519);
nor U1594 (N_1594,N_1557,N_1548);
and U1595 (N_1595,N_1516,N_1557);
nand U1596 (N_1596,N_1527,N_1529);
or U1597 (N_1597,N_1545,N_1506);
nor U1598 (N_1598,N_1550,N_1521);
and U1599 (N_1599,N_1518,N_1538);
nand U1600 (N_1600,N_1541,N_1543);
nor U1601 (N_1601,N_1505,N_1557);
nor U1602 (N_1602,N_1521,N_1524);
nor U1603 (N_1603,N_1517,N_1502);
or U1604 (N_1604,N_1557,N_1520);
or U1605 (N_1605,N_1516,N_1529);
and U1606 (N_1606,N_1502,N_1518);
and U1607 (N_1607,N_1522,N_1517);
nor U1608 (N_1608,N_1507,N_1551);
and U1609 (N_1609,N_1554,N_1524);
nor U1610 (N_1610,N_1516,N_1528);
or U1611 (N_1611,N_1549,N_1554);
nand U1612 (N_1612,N_1547,N_1526);
or U1613 (N_1613,N_1539,N_1553);
nor U1614 (N_1614,N_1520,N_1543);
nor U1615 (N_1615,N_1501,N_1553);
or U1616 (N_1616,N_1515,N_1521);
nand U1617 (N_1617,N_1512,N_1540);
nand U1618 (N_1618,N_1551,N_1503);
or U1619 (N_1619,N_1530,N_1518);
or U1620 (N_1620,N_1575,N_1617);
or U1621 (N_1621,N_1581,N_1582);
nand U1622 (N_1622,N_1588,N_1602);
nand U1623 (N_1623,N_1618,N_1585);
nor U1624 (N_1624,N_1576,N_1597);
or U1625 (N_1625,N_1596,N_1613);
and U1626 (N_1626,N_1563,N_1573);
nor U1627 (N_1627,N_1580,N_1590);
nand U1628 (N_1628,N_1600,N_1574);
nand U1629 (N_1629,N_1609,N_1570);
nor U1630 (N_1630,N_1584,N_1619);
nor U1631 (N_1631,N_1614,N_1566);
and U1632 (N_1632,N_1592,N_1595);
nand U1633 (N_1633,N_1567,N_1565);
nor U1634 (N_1634,N_1583,N_1607);
nand U1635 (N_1635,N_1601,N_1571);
or U1636 (N_1636,N_1605,N_1604);
or U1637 (N_1637,N_1587,N_1562);
or U1638 (N_1638,N_1564,N_1610);
nor U1639 (N_1639,N_1612,N_1560);
nor U1640 (N_1640,N_1569,N_1606);
nand U1641 (N_1641,N_1586,N_1577);
and U1642 (N_1642,N_1579,N_1594);
or U1643 (N_1643,N_1591,N_1603);
nor U1644 (N_1644,N_1599,N_1608);
nor U1645 (N_1645,N_1611,N_1578);
or U1646 (N_1646,N_1568,N_1561);
or U1647 (N_1647,N_1615,N_1598);
or U1648 (N_1648,N_1593,N_1572);
and U1649 (N_1649,N_1616,N_1589);
or U1650 (N_1650,N_1618,N_1567);
and U1651 (N_1651,N_1562,N_1603);
nand U1652 (N_1652,N_1573,N_1596);
nor U1653 (N_1653,N_1571,N_1582);
or U1654 (N_1654,N_1612,N_1617);
nor U1655 (N_1655,N_1561,N_1576);
or U1656 (N_1656,N_1605,N_1560);
and U1657 (N_1657,N_1619,N_1605);
nor U1658 (N_1658,N_1598,N_1612);
or U1659 (N_1659,N_1572,N_1602);
or U1660 (N_1660,N_1610,N_1611);
nand U1661 (N_1661,N_1564,N_1576);
nand U1662 (N_1662,N_1612,N_1562);
or U1663 (N_1663,N_1566,N_1603);
and U1664 (N_1664,N_1564,N_1568);
nand U1665 (N_1665,N_1581,N_1569);
and U1666 (N_1666,N_1607,N_1586);
nand U1667 (N_1667,N_1565,N_1561);
nor U1668 (N_1668,N_1583,N_1585);
or U1669 (N_1669,N_1599,N_1579);
and U1670 (N_1670,N_1584,N_1607);
or U1671 (N_1671,N_1563,N_1600);
nor U1672 (N_1672,N_1609,N_1574);
and U1673 (N_1673,N_1569,N_1578);
and U1674 (N_1674,N_1606,N_1615);
and U1675 (N_1675,N_1588,N_1618);
or U1676 (N_1676,N_1564,N_1597);
nand U1677 (N_1677,N_1616,N_1592);
and U1678 (N_1678,N_1569,N_1580);
and U1679 (N_1679,N_1574,N_1605);
or U1680 (N_1680,N_1670,N_1661);
nand U1681 (N_1681,N_1674,N_1639);
and U1682 (N_1682,N_1651,N_1646);
or U1683 (N_1683,N_1653,N_1655);
nand U1684 (N_1684,N_1627,N_1632);
and U1685 (N_1685,N_1633,N_1623);
nor U1686 (N_1686,N_1673,N_1642);
or U1687 (N_1687,N_1657,N_1667);
nor U1688 (N_1688,N_1641,N_1638);
nor U1689 (N_1689,N_1640,N_1647);
or U1690 (N_1690,N_1672,N_1671);
nand U1691 (N_1691,N_1625,N_1662);
nand U1692 (N_1692,N_1665,N_1676);
nand U1693 (N_1693,N_1666,N_1660);
and U1694 (N_1694,N_1677,N_1658);
nor U1695 (N_1695,N_1668,N_1659);
and U1696 (N_1696,N_1645,N_1679);
nand U1697 (N_1697,N_1669,N_1637);
or U1698 (N_1698,N_1631,N_1630);
nor U1699 (N_1699,N_1626,N_1629);
and U1700 (N_1700,N_1622,N_1650);
nor U1701 (N_1701,N_1636,N_1644);
or U1702 (N_1702,N_1663,N_1649);
nor U1703 (N_1703,N_1656,N_1620);
and U1704 (N_1704,N_1678,N_1675);
nor U1705 (N_1705,N_1652,N_1648);
and U1706 (N_1706,N_1621,N_1635);
nand U1707 (N_1707,N_1654,N_1628);
nor U1708 (N_1708,N_1643,N_1624);
or U1709 (N_1709,N_1634,N_1664);
or U1710 (N_1710,N_1662,N_1663);
or U1711 (N_1711,N_1628,N_1673);
nor U1712 (N_1712,N_1643,N_1631);
and U1713 (N_1713,N_1620,N_1645);
nand U1714 (N_1714,N_1622,N_1678);
and U1715 (N_1715,N_1646,N_1622);
nor U1716 (N_1716,N_1653,N_1630);
nand U1717 (N_1717,N_1649,N_1652);
and U1718 (N_1718,N_1666,N_1648);
nor U1719 (N_1719,N_1665,N_1662);
or U1720 (N_1720,N_1647,N_1656);
and U1721 (N_1721,N_1659,N_1664);
or U1722 (N_1722,N_1674,N_1630);
xnor U1723 (N_1723,N_1634,N_1644);
nand U1724 (N_1724,N_1633,N_1621);
nand U1725 (N_1725,N_1635,N_1629);
and U1726 (N_1726,N_1629,N_1663);
and U1727 (N_1727,N_1652,N_1635);
and U1728 (N_1728,N_1668,N_1642);
nand U1729 (N_1729,N_1655,N_1663);
nand U1730 (N_1730,N_1636,N_1658);
or U1731 (N_1731,N_1626,N_1660);
xnor U1732 (N_1732,N_1626,N_1640);
or U1733 (N_1733,N_1665,N_1638);
nand U1734 (N_1734,N_1648,N_1674);
or U1735 (N_1735,N_1646,N_1653);
or U1736 (N_1736,N_1675,N_1626);
nor U1737 (N_1737,N_1624,N_1645);
nand U1738 (N_1738,N_1638,N_1658);
nor U1739 (N_1739,N_1639,N_1645);
nor U1740 (N_1740,N_1704,N_1688);
nor U1741 (N_1741,N_1739,N_1682);
nand U1742 (N_1742,N_1699,N_1719);
nand U1743 (N_1743,N_1716,N_1702);
nand U1744 (N_1744,N_1712,N_1690);
nor U1745 (N_1745,N_1685,N_1691);
nor U1746 (N_1746,N_1714,N_1709);
or U1747 (N_1747,N_1689,N_1713);
nand U1748 (N_1748,N_1686,N_1723);
nor U1749 (N_1749,N_1684,N_1694);
or U1750 (N_1750,N_1706,N_1700);
nand U1751 (N_1751,N_1728,N_1729);
nand U1752 (N_1752,N_1727,N_1681);
or U1753 (N_1753,N_1687,N_1695);
nand U1754 (N_1754,N_1724,N_1718);
nand U1755 (N_1755,N_1735,N_1737);
and U1756 (N_1756,N_1711,N_1698);
or U1757 (N_1757,N_1736,N_1697);
nand U1758 (N_1758,N_1683,N_1717);
xnor U1759 (N_1759,N_1710,N_1701);
nand U1760 (N_1760,N_1733,N_1692);
and U1761 (N_1761,N_1680,N_1715);
nor U1762 (N_1762,N_1721,N_1730);
or U1763 (N_1763,N_1734,N_1731);
and U1764 (N_1764,N_1705,N_1703);
xor U1765 (N_1765,N_1708,N_1693);
and U1766 (N_1766,N_1720,N_1732);
nand U1767 (N_1767,N_1722,N_1738);
nand U1768 (N_1768,N_1726,N_1725);
nand U1769 (N_1769,N_1696,N_1707);
nor U1770 (N_1770,N_1725,N_1714);
nor U1771 (N_1771,N_1696,N_1717);
and U1772 (N_1772,N_1729,N_1703);
nor U1773 (N_1773,N_1728,N_1725);
and U1774 (N_1774,N_1700,N_1710);
and U1775 (N_1775,N_1682,N_1734);
or U1776 (N_1776,N_1730,N_1737);
and U1777 (N_1777,N_1721,N_1685);
nor U1778 (N_1778,N_1700,N_1705);
nor U1779 (N_1779,N_1693,N_1685);
nor U1780 (N_1780,N_1735,N_1686);
nand U1781 (N_1781,N_1708,N_1710);
nand U1782 (N_1782,N_1690,N_1683);
or U1783 (N_1783,N_1723,N_1714);
and U1784 (N_1784,N_1715,N_1697);
and U1785 (N_1785,N_1699,N_1702);
or U1786 (N_1786,N_1718,N_1693);
or U1787 (N_1787,N_1732,N_1725);
and U1788 (N_1788,N_1719,N_1736);
or U1789 (N_1789,N_1686,N_1700);
or U1790 (N_1790,N_1734,N_1713);
nor U1791 (N_1791,N_1690,N_1686);
and U1792 (N_1792,N_1695,N_1724);
nor U1793 (N_1793,N_1693,N_1704);
or U1794 (N_1794,N_1735,N_1699);
and U1795 (N_1795,N_1708,N_1691);
or U1796 (N_1796,N_1721,N_1709);
nand U1797 (N_1797,N_1681,N_1730);
nand U1798 (N_1798,N_1684,N_1705);
nand U1799 (N_1799,N_1694,N_1703);
nand U1800 (N_1800,N_1748,N_1784);
nor U1801 (N_1801,N_1743,N_1783);
nor U1802 (N_1802,N_1776,N_1791);
and U1803 (N_1803,N_1790,N_1781);
and U1804 (N_1804,N_1767,N_1766);
or U1805 (N_1805,N_1789,N_1792);
nand U1806 (N_1806,N_1764,N_1761);
or U1807 (N_1807,N_1740,N_1796);
nor U1808 (N_1808,N_1768,N_1751);
nand U1809 (N_1809,N_1786,N_1762);
and U1810 (N_1810,N_1788,N_1750);
nand U1811 (N_1811,N_1785,N_1773);
and U1812 (N_1812,N_1779,N_1774);
or U1813 (N_1813,N_1782,N_1775);
or U1814 (N_1814,N_1742,N_1772);
and U1815 (N_1815,N_1754,N_1777);
and U1816 (N_1816,N_1769,N_1771);
and U1817 (N_1817,N_1765,N_1759);
or U1818 (N_1818,N_1799,N_1758);
nor U1819 (N_1819,N_1752,N_1795);
nand U1820 (N_1820,N_1755,N_1746);
and U1821 (N_1821,N_1797,N_1744);
and U1822 (N_1822,N_1793,N_1763);
or U1823 (N_1823,N_1780,N_1787);
nor U1824 (N_1824,N_1778,N_1741);
nor U1825 (N_1825,N_1753,N_1760);
nand U1826 (N_1826,N_1747,N_1770);
nor U1827 (N_1827,N_1749,N_1798);
nand U1828 (N_1828,N_1745,N_1756);
nand U1829 (N_1829,N_1757,N_1794);
and U1830 (N_1830,N_1792,N_1799);
and U1831 (N_1831,N_1782,N_1756);
or U1832 (N_1832,N_1789,N_1790);
nand U1833 (N_1833,N_1748,N_1772);
nand U1834 (N_1834,N_1769,N_1787);
nand U1835 (N_1835,N_1791,N_1769);
nand U1836 (N_1836,N_1755,N_1748);
nor U1837 (N_1837,N_1790,N_1785);
nor U1838 (N_1838,N_1760,N_1762);
or U1839 (N_1839,N_1781,N_1784);
or U1840 (N_1840,N_1752,N_1786);
and U1841 (N_1841,N_1760,N_1759);
nand U1842 (N_1842,N_1767,N_1769);
and U1843 (N_1843,N_1767,N_1772);
and U1844 (N_1844,N_1757,N_1779);
nor U1845 (N_1845,N_1785,N_1792);
nand U1846 (N_1846,N_1757,N_1783);
and U1847 (N_1847,N_1779,N_1767);
and U1848 (N_1848,N_1799,N_1759);
nand U1849 (N_1849,N_1759,N_1750);
or U1850 (N_1850,N_1795,N_1764);
or U1851 (N_1851,N_1743,N_1798);
or U1852 (N_1852,N_1792,N_1775);
and U1853 (N_1853,N_1775,N_1751);
xor U1854 (N_1854,N_1776,N_1766);
nand U1855 (N_1855,N_1775,N_1778);
nor U1856 (N_1856,N_1784,N_1750);
nand U1857 (N_1857,N_1745,N_1741);
and U1858 (N_1858,N_1763,N_1745);
nor U1859 (N_1859,N_1762,N_1747);
nor U1860 (N_1860,N_1827,N_1805);
or U1861 (N_1861,N_1850,N_1817);
nor U1862 (N_1862,N_1859,N_1819);
nor U1863 (N_1863,N_1856,N_1844);
or U1864 (N_1864,N_1854,N_1843);
nand U1865 (N_1865,N_1802,N_1829);
or U1866 (N_1866,N_1822,N_1833);
and U1867 (N_1867,N_1814,N_1834);
nor U1868 (N_1868,N_1858,N_1857);
nand U1869 (N_1869,N_1823,N_1800);
or U1870 (N_1870,N_1821,N_1852);
or U1871 (N_1871,N_1825,N_1841);
nand U1872 (N_1872,N_1809,N_1853);
nor U1873 (N_1873,N_1813,N_1830);
or U1874 (N_1874,N_1801,N_1845);
and U1875 (N_1875,N_1816,N_1804);
or U1876 (N_1876,N_1803,N_1836);
and U1877 (N_1877,N_1824,N_1846);
nand U1878 (N_1878,N_1815,N_1839);
and U1879 (N_1879,N_1828,N_1842);
and U1880 (N_1880,N_1807,N_1837);
and U1881 (N_1881,N_1832,N_1851);
and U1882 (N_1882,N_1826,N_1835);
nand U1883 (N_1883,N_1806,N_1848);
and U1884 (N_1884,N_1849,N_1811);
nand U1885 (N_1885,N_1847,N_1838);
nand U1886 (N_1886,N_1820,N_1840);
nor U1887 (N_1887,N_1810,N_1818);
or U1888 (N_1888,N_1831,N_1812);
nor U1889 (N_1889,N_1855,N_1808);
nor U1890 (N_1890,N_1808,N_1803);
nor U1891 (N_1891,N_1836,N_1849);
nor U1892 (N_1892,N_1812,N_1821);
nor U1893 (N_1893,N_1803,N_1817);
and U1894 (N_1894,N_1832,N_1812);
or U1895 (N_1895,N_1827,N_1816);
and U1896 (N_1896,N_1824,N_1850);
or U1897 (N_1897,N_1840,N_1825);
nor U1898 (N_1898,N_1835,N_1813);
and U1899 (N_1899,N_1816,N_1837);
or U1900 (N_1900,N_1812,N_1853);
or U1901 (N_1901,N_1840,N_1831);
nor U1902 (N_1902,N_1814,N_1818);
or U1903 (N_1903,N_1819,N_1822);
nand U1904 (N_1904,N_1859,N_1808);
nand U1905 (N_1905,N_1811,N_1817);
or U1906 (N_1906,N_1805,N_1839);
and U1907 (N_1907,N_1830,N_1856);
nor U1908 (N_1908,N_1838,N_1828);
nand U1909 (N_1909,N_1820,N_1832);
or U1910 (N_1910,N_1829,N_1840);
nand U1911 (N_1911,N_1835,N_1815);
nand U1912 (N_1912,N_1811,N_1829);
nor U1913 (N_1913,N_1858,N_1802);
nand U1914 (N_1914,N_1823,N_1855);
nor U1915 (N_1915,N_1824,N_1823);
and U1916 (N_1916,N_1829,N_1806);
nor U1917 (N_1917,N_1834,N_1850);
or U1918 (N_1918,N_1849,N_1856);
nor U1919 (N_1919,N_1823,N_1814);
or U1920 (N_1920,N_1919,N_1881);
or U1921 (N_1921,N_1906,N_1875);
nand U1922 (N_1922,N_1895,N_1862);
nand U1923 (N_1923,N_1903,N_1893);
or U1924 (N_1924,N_1897,N_1865);
or U1925 (N_1925,N_1899,N_1873);
or U1926 (N_1926,N_1874,N_1861);
or U1927 (N_1927,N_1907,N_1876);
or U1928 (N_1928,N_1913,N_1889);
nand U1929 (N_1929,N_1910,N_1870);
nand U1930 (N_1930,N_1902,N_1863);
and U1931 (N_1931,N_1884,N_1872);
nor U1932 (N_1932,N_1887,N_1901);
or U1933 (N_1933,N_1864,N_1908);
nor U1934 (N_1934,N_1882,N_1860);
nand U1935 (N_1935,N_1891,N_1914);
or U1936 (N_1936,N_1888,N_1880);
nand U1937 (N_1937,N_1905,N_1909);
nor U1938 (N_1938,N_1900,N_1878);
nor U1939 (N_1939,N_1866,N_1892);
nor U1940 (N_1940,N_1883,N_1916);
nand U1941 (N_1941,N_1911,N_1894);
and U1942 (N_1942,N_1885,N_1886);
or U1943 (N_1943,N_1904,N_1898);
or U1944 (N_1944,N_1915,N_1867);
nand U1945 (N_1945,N_1871,N_1896);
nand U1946 (N_1946,N_1912,N_1877);
nand U1947 (N_1947,N_1879,N_1869);
and U1948 (N_1948,N_1918,N_1890);
or U1949 (N_1949,N_1868,N_1917);
nor U1950 (N_1950,N_1870,N_1901);
nor U1951 (N_1951,N_1872,N_1897);
nand U1952 (N_1952,N_1862,N_1874);
and U1953 (N_1953,N_1900,N_1908);
or U1954 (N_1954,N_1905,N_1899);
or U1955 (N_1955,N_1895,N_1916);
nor U1956 (N_1956,N_1888,N_1860);
and U1957 (N_1957,N_1895,N_1899);
and U1958 (N_1958,N_1910,N_1899);
or U1959 (N_1959,N_1917,N_1919);
xnor U1960 (N_1960,N_1887,N_1898);
nor U1961 (N_1961,N_1862,N_1916);
nand U1962 (N_1962,N_1910,N_1880);
nor U1963 (N_1963,N_1888,N_1905);
nor U1964 (N_1964,N_1869,N_1865);
and U1965 (N_1965,N_1902,N_1894);
and U1966 (N_1966,N_1888,N_1862);
or U1967 (N_1967,N_1894,N_1863);
nor U1968 (N_1968,N_1893,N_1888);
nor U1969 (N_1969,N_1885,N_1899);
or U1970 (N_1970,N_1895,N_1914);
nor U1971 (N_1971,N_1918,N_1912);
nor U1972 (N_1972,N_1864,N_1874);
nor U1973 (N_1973,N_1880,N_1869);
nor U1974 (N_1974,N_1912,N_1862);
or U1975 (N_1975,N_1873,N_1863);
and U1976 (N_1976,N_1901,N_1888);
nor U1977 (N_1977,N_1890,N_1871);
nor U1978 (N_1978,N_1919,N_1882);
nand U1979 (N_1979,N_1915,N_1901);
or U1980 (N_1980,N_1965,N_1939);
and U1981 (N_1981,N_1960,N_1943);
nand U1982 (N_1982,N_1958,N_1972);
nor U1983 (N_1983,N_1922,N_1932);
nand U1984 (N_1984,N_1928,N_1975);
or U1985 (N_1985,N_1920,N_1961);
or U1986 (N_1986,N_1957,N_1924);
nor U1987 (N_1987,N_1976,N_1971);
and U1988 (N_1988,N_1934,N_1968);
nand U1989 (N_1989,N_1973,N_1967);
nand U1990 (N_1990,N_1966,N_1927);
nand U1991 (N_1991,N_1921,N_1969);
nand U1992 (N_1992,N_1940,N_1942);
xnor U1993 (N_1993,N_1936,N_1923);
nor U1994 (N_1994,N_1945,N_1950);
nor U1995 (N_1995,N_1933,N_1931);
nor U1996 (N_1996,N_1978,N_1964);
or U1997 (N_1997,N_1951,N_1930);
and U1998 (N_1998,N_1962,N_1970);
nand U1999 (N_1999,N_1937,N_1954);
or U2000 (N_2000,N_1938,N_1952);
and U2001 (N_2001,N_1949,N_1955);
and U2002 (N_2002,N_1929,N_1959);
nor U2003 (N_2003,N_1974,N_1953);
and U2004 (N_2004,N_1977,N_1935);
and U2005 (N_2005,N_1926,N_1925);
nor U2006 (N_2006,N_1947,N_1963);
nand U2007 (N_2007,N_1956,N_1944);
nand U2008 (N_2008,N_1946,N_1941);
nor U2009 (N_2009,N_1979,N_1948);
nor U2010 (N_2010,N_1970,N_1939);
nand U2011 (N_2011,N_1963,N_1923);
or U2012 (N_2012,N_1977,N_1951);
or U2013 (N_2013,N_1932,N_1943);
nor U2014 (N_2014,N_1953,N_1969);
nor U2015 (N_2015,N_1972,N_1976);
and U2016 (N_2016,N_1924,N_1974);
nand U2017 (N_2017,N_1959,N_1961);
or U2018 (N_2018,N_1949,N_1959);
or U2019 (N_2019,N_1935,N_1944);
nor U2020 (N_2020,N_1945,N_1978);
nand U2021 (N_2021,N_1930,N_1956);
nand U2022 (N_2022,N_1930,N_1958);
nand U2023 (N_2023,N_1964,N_1966);
nor U2024 (N_2024,N_1923,N_1922);
and U2025 (N_2025,N_1966,N_1972);
nand U2026 (N_2026,N_1948,N_1935);
and U2027 (N_2027,N_1948,N_1937);
nor U2028 (N_2028,N_1934,N_1962);
nor U2029 (N_2029,N_1944,N_1925);
or U2030 (N_2030,N_1971,N_1972);
nand U2031 (N_2031,N_1924,N_1971);
nor U2032 (N_2032,N_1933,N_1929);
or U2033 (N_2033,N_1978,N_1941);
or U2034 (N_2034,N_1949,N_1973);
or U2035 (N_2035,N_1976,N_1951);
nor U2036 (N_2036,N_1929,N_1961);
nor U2037 (N_2037,N_1950,N_1936);
nand U2038 (N_2038,N_1977,N_1926);
nor U2039 (N_2039,N_1925,N_1948);
nor U2040 (N_2040,N_1992,N_2017);
and U2041 (N_2041,N_1998,N_1989);
nand U2042 (N_2042,N_2011,N_2029);
or U2043 (N_2043,N_1990,N_2007);
or U2044 (N_2044,N_2009,N_1987);
and U2045 (N_2045,N_2030,N_2006);
or U2046 (N_2046,N_2021,N_2022);
nor U2047 (N_2047,N_2027,N_2036);
and U2048 (N_2048,N_2034,N_2008);
nand U2049 (N_2049,N_2028,N_2012);
and U2050 (N_2050,N_2016,N_2018);
nor U2051 (N_2051,N_1984,N_2003);
or U2052 (N_2052,N_1994,N_2001);
and U2053 (N_2053,N_1983,N_2002);
and U2054 (N_2054,N_2023,N_2026);
nor U2055 (N_2055,N_2014,N_1995);
or U2056 (N_2056,N_2035,N_2005);
and U2057 (N_2057,N_2039,N_1993);
nor U2058 (N_2058,N_1985,N_1980);
and U2059 (N_2059,N_2020,N_2032);
nand U2060 (N_2060,N_2025,N_1997);
nand U2061 (N_2061,N_1991,N_2015);
or U2062 (N_2062,N_1999,N_2031);
nand U2063 (N_2063,N_1981,N_2038);
nor U2064 (N_2064,N_1986,N_2024);
and U2065 (N_2065,N_2010,N_1996);
or U2066 (N_2066,N_2037,N_2013);
xor U2067 (N_2067,N_2000,N_1982);
and U2068 (N_2068,N_2033,N_2019);
nand U2069 (N_2069,N_1988,N_2004);
nand U2070 (N_2070,N_1987,N_1980);
and U2071 (N_2071,N_2020,N_2024);
and U2072 (N_2072,N_1994,N_2025);
nor U2073 (N_2073,N_2016,N_1982);
nand U2074 (N_2074,N_2012,N_2008);
nor U2075 (N_2075,N_2012,N_1987);
and U2076 (N_2076,N_2010,N_2025);
nor U2077 (N_2077,N_2000,N_2033);
nor U2078 (N_2078,N_1989,N_2011);
and U2079 (N_2079,N_2018,N_2014);
nand U2080 (N_2080,N_2032,N_2019);
and U2081 (N_2081,N_2024,N_1997);
nand U2082 (N_2082,N_2027,N_2032);
nand U2083 (N_2083,N_1981,N_2025);
or U2084 (N_2084,N_2036,N_1989);
and U2085 (N_2085,N_1998,N_2035);
nor U2086 (N_2086,N_1992,N_1987);
and U2087 (N_2087,N_2023,N_2028);
and U2088 (N_2088,N_2014,N_2032);
nor U2089 (N_2089,N_2026,N_2010);
nor U2090 (N_2090,N_1988,N_1993);
nor U2091 (N_2091,N_2027,N_2025);
xor U2092 (N_2092,N_2013,N_2001);
or U2093 (N_2093,N_1986,N_1997);
nand U2094 (N_2094,N_2030,N_2008);
xor U2095 (N_2095,N_2039,N_2018);
or U2096 (N_2096,N_2023,N_2032);
nand U2097 (N_2097,N_2029,N_2031);
or U2098 (N_2098,N_1998,N_2022);
nand U2099 (N_2099,N_1983,N_2030);
nor U2100 (N_2100,N_2065,N_2060);
and U2101 (N_2101,N_2056,N_2049);
and U2102 (N_2102,N_2054,N_2051);
nor U2103 (N_2103,N_2057,N_2090);
or U2104 (N_2104,N_2075,N_2083);
nor U2105 (N_2105,N_2070,N_2059);
nor U2106 (N_2106,N_2043,N_2087);
nor U2107 (N_2107,N_2077,N_2096);
nand U2108 (N_2108,N_2078,N_2062);
and U2109 (N_2109,N_2052,N_2058);
and U2110 (N_2110,N_2073,N_2095);
nand U2111 (N_2111,N_2086,N_2046);
or U2112 (N_2112,N_2092,N_2097);
and U2113 (N_2113,N_2048,N_2076);
nor U2114 (N_2114,N_2053,N_2074);
or U2115 (N_2115,N_2099,N_2069);
or U2116 (N_2116,N_2044,N_2047);
and U2117 (N_2117,N_2055,N_2050);
nor U2118 (N_2118,N_2068,N_2045);
nor U2119 (N_2119,N_2091,N_2082);
or U2120 (N_2120,N_2088,N_2042);
nor U2121 (N_2121,N_2093,N_2041);
or U2122 (N_2122,N_2061,N_2072);
and U2123 (N_2123,N_2089,N_2067);
nor U2124 (N_2124,N_2066,N_2063);
nor U2125 (N_2125,N_2084,N_2080);
nor U2126 (N_2126,N_2071,N_2079);
nor U2127 (N_2127,N_2040,N_2085);
and U2128 (N_2128,N_2064,N_2094);
nor U2129 (N_2129,N_2081,N_2098);
xor U2130 (N_2130,N_2055,N_2095);
xnor U2131 (N_2131,N_2082,N_2055);
or U2132 (N_2132,N_2085,N_2058);
nand U2133 (N_2133,N_2087,N_2065);
nand U2134 (N_2134,N_2092,N_2061);
nor U2135 (N_2135,N_2087,N_2076);
or U2136 (N_2136,N_2055,N_2062);
nand U2137 (N_2137,N_2064,N_2040);
nor U2138 (N_2138,N_2047,N_2075);
nor U2139 (N_2139,N_2062,N_2090);
nand U2140 (N_2140,N_2093,N_2083);
nor U2141 (N_2141,N_2054,N_2049);
nand U2142 (N_2142,N_2097,N_2056);
nand U2143 (N_2143,N_2075,N_2056);
nand U2144 (N_2144,N_2071,N_2070);
or U2145 (N_2145,N_2077,N_2074);
or U2146 (N_2146,N_2083,N_2095);
nand U2147 (N_2147,N_2089,N_2080);
nand U2148 (N_2148,N_2048,N_2095);
nor U2149 (N_2149,N_2074,N_2096);
nor U2150 (N_2150,N_2072,N_2064);
nor U2151 (N_2151,N_2076,N_2047);
and U2152 (N_2152,N_2051,N_2092);
and U2153 (N_2153,N_2054,N_2075);
nand U2154 (N_2154,N_2087,N_2059);
and U2155 (N_2155,N_2040,N_2048);
nor U2156 (N_2156,N_2070,N_2093);
nor U2157 (N_2157,N_2053,N_2072);
and U2158 (N_2158,N_2081,N_2091);
or U2159 (N_2159,N_2092,N_2074);
xor U2160 (N_2160,N_2147,N_2133);
and U2161 (N_2161,N_2159,N_2107);
nand U2162 (N_2162,N_2121,N_2100);
and U2163 (N_2163,N_2112,N_2136);
nand U2164 (N_2164,N_2116,N_2144);
or U2165 (N_2165,N_2140,N_2158);
and U2166 (N_2166,N_2148,N_2110);
nor U2167 (N_2167,N_2118,N_2155);
and U2168 (N_2168,N_2117,N_2129);
nor U2169 (N_2169,N_2120,N_2109);
and U2170 (N_2170,N_2123,N_2111);
and U2171 (N_2171,N_2124,N_2138);
and U2172 (N_2172,N_2150,N_2134);
nand U2173 (N_2173,N_2103,N_2122);
and U2174 (N_2174,N_2115,N_2149);
and U2175 (N_2175,N_2113,N_2105);
nand U2176 (N_2176,N_2114,N_2141);
nor U2177 (N_2177,N_2119,N_2145);
or U2178 (N_2178,N_2139,N_2108);
nor U2179 (N_2179,N_2137,N_2106);
nand U2180 (N_2180,N_2126,N_2142);
nor U2181 (N_2181,N_2135,N_2104);
nor U2182 (N_2182,N_2156,N_2127);
or U2183 (N_2183,N_2130,N_2153);
and U2184 (N_2184,N_2132,N_2128);
or U2185 (N_2185,N_2131,N_2152);
nand U2186 (N_2186,N_2151,N_2101);
and U2187 (N_2187,N_2143,N_2146);
nor U2188 (N_2188,N_2125,N_2157);
nor U2189 (N_2189,N_2102,N_2154);
or U2190 (N_2190,N_2122,N_2121);
nand U2191 (N_2191,N_2103,N_2102);
or U2192 (N_2192,N_2154,N_2103);
and U2193 (N_2193,N_2153,N_2132);
and U2194 (N_2194,N_2142,N_2106);
nand U2195 (N_2195,N_2155,N_2115);
nand U2196 (N_2196,N_2129,N_2142);
nand U2197 (N_2197,N_2118,N_2121);
or U2198 (N_2198,N_2117,N_2108);
nor U2199 (N_2199,N_2105,N_2119);
nor U2200 (N_2200,N_2106,N_2143);
and U2201 (N_2201,N_2136,N_2129);
nand U2202 (N_2202,N_2152,N_2110);
or U2203 (N_2203,N_2121,N_2128);
or U2204 (N_2204,N_2126,N_2125);
or U2205 (N_2205,N_2116,N_2150);
nand U2206 (N_2206,N_2138,N_2111);
nand U2207 (N_2207,N_2156,N_2159);
nor U2208 (N_2208,N_2109,N_2157);
and U2209 (N_2209,N_2130,N_2104);
nor U2210 (N_2210,N_2111,N_2114);
nand U2211 (N_2211,N_2100,N_2108);
and U2212 (N_2212,N_2149,N_2134);
nor U2213 (N_2213,N_2114,N_2131);
nor U2214 (N_2214,N_2124,N_2156);
and U2215 (N_2215,N_2149,N_2158);
nor U2216 (N_2216,N_2148,N_2155);
and U2217 (N_2217,N_2149,N_2116);
nand U2218 (N_2218,N_2126,N_2124);
or U2219 (N_2219,N_2143,N_2155);
nor U2220 (N_2220,N_2169,N_2179);
nor U2221 (N_2221,N_2174,N_2164);
or U2222 (N_2222,N_2212,N_2187);
nand U2223 (N_2223,N_2191,N_2168);
or U2224 (N_2224,N_2182,N_2165);
nand U2225 (N_2225,N_2185,N_2184);
nand U2226 (N_2226,N_2207,N_2219);
and U2227 (N_2227,N_2163,N_2217);
and U2228 (N_2228,N_2218,N_2204);
nand U2229 (N_2229,N_2180,N_2190);
and U2230 (N_2230,N_2201,N_2210);
or U2231 (N_2231,N_2178,N_2183);
nor U2232 (N_2232,N_2214,N_2188);
and U2233 (N_2233,N_2197,N_2189);
nand U2234 (N_2234,N_2195,N_2200);
and U2235 (N_2235,N_2175,N_2211);
or U2236 (N_2236,N_2181,N_2203);
nand U2237 (N_2237,N_2194,N_2199);
nand U2238 (N_2238,N_2170,N_2186);
or U2239 (N_2239,N_2173,N_2208);
and U2240 (N_2240,N_2202,N_2166);
nand U2241 (N_2241,N_2206,N_2193);
and U2242 (N_2242,N_2171,N_2172);
nor U2243 (N_2243,N_2177,N_2198);
and U2244 (N_2244,N_2205,N_2160);
nor U2245 (N_2245,N_2167,N_2161);
nor U2246 (N_2246,N_2196,N_2192);
nand U2247 (N_2247,N_2209,N_2213);
or U2248 (N_2248,N_2176,N_2215);
or U2249 (N_2249,N_2216,N_2162);
or U2250 (N_2250,N_2178,N_2175);
nor U2251 (N_2251,N_2179,N_2212);
or U2252 (N_2252,N_2164,N_2200);
nor U2253 (N_2253,N_2169,N_2163);
and U2254 (N_2254,N_2162,N_2172);
and U2255 (N_2255,N_2199,N_2212);
and U2256 (N_2256,N_2190,N_2188);
nand U2257 (N_2257,N_2218,N_2213);
and U2258 (N_2258,N_2210,N_2187);
nor U2259 (N_2259,N_2210,N_2176);
and U2260 (N_2260,N_2166,N_2207);
or U2261 (N_2261,N_2209,N_2163);
and U2262 (N_2262,N_2213,N_2169);
xnor U2263 (N_2263,N_2179,N_2208);
nand U2264 (N_2264,N_2182,N_2213);
or U2265 (N_2265,N_2213,N_2189);
nand U2266 (N_2266,N_2177,N_2188);
or U2267 (N_2267,N_2182,N_2178);
nor U2268 (N_2268,N_2212,N_2168);
nor U2269 (N_2269,N_2171,N_2202);
nand U2270 (N_2270,N_2186,N_2164);
and U2271 (N_2271,N_2186,N_2219);
and U2272 (N_2272,N_2211,N_2212);
nand U2273 (N_2273,N_2192,N_2167);
or U2274 (N_2274,N_2193,N_2192);
or U2275 (N_2275,N_2174,N_2182);
nand U2276 (N_2276,N_2175,N_2194);
nor U2277 (N_2277,N_2219,N_2213);
and U2278 (N_2278,N_2201,N_2178);
nand U2279 (N_2279,N_2162,N_2188);
nand U2280 (N_2280,N_2243,N_2237);
and U2281 (N_2281,N_2272,N_2223);
nand U2282 (N_2282,N_2235,N_2263);
nor U2283 (N_2283,N_2228,N_2246);
or U2284 (N_2284,N_2220,N_2261);
nor U2285 (N_2285,N_2249,N_2221);
or U2286 (N_2286,N_2276,N_2257);
nor U2287 (N_2287,N_2256,N_2260);
and U2288 (N_2288,N_2273,N_2270);
or U2289 (N_2289,N_2265,N_2242);
or U2290 (N_2290,N_2222,N_2262);
and U2291 (N_2291,N_2255,N_2253);
and U2292 (N_2292,N_2236,N_2259);
and U2293 (N_2293,N_2254,N_2230);
and U2294 (N_2294,N_2271,N_2225);
nor U2295 (N_2295,N_2226,N_2240);
nand U2296 (N_2296,N_2234,N_2274);
and U2297 (N_2297,N_2264,N_2229);
and U2298 (N_2298,N_2258,N_2224);
and U2299 (N_2299,N_2268,N_2251);
and U2300 (N_2300,N_2227,N_2239);
xor U2301 (N_2301,N_2269,N_2233);
nand U2302 (N_2302,N_2244,N_2238);
and U2303 (N_2303,N_2232,N_2241);
xnor U2304 (N_2304,N_2245,N_2266);
and U2305 (N_2305,N_2247,N_2248);
nor U2306 (N_2306,N_2252,N_2231);
nand U2307 (N_2307,N_2275,N_2277);
nor U2308 (N_2308,N_2278,N_2250);
or U2309 (N_2309,N_2279,N_2267);
nor U2310 (N_2310,N_2231,N_2257);
nor U2311 (N_2311,N_2242,N_2225);
nand U2312 (N_2312,N_2252,N_2267);
nor U2313 (N_2313,N_2220,N_2254);
or U2314 (N_2314,N_2275,N_2249);
nand U2315 (N_2315,N_2269,N_2232);
nand U2316 (N_2316,N_2266,N_2272);
nand U2317 (N_2317,N_2263,N_2232);
nand U2318 (N_2318,N_2261,N_2276);
or U2319 (N_2319,N_2252,N_2235);
and U2320 (N_2320,N_2275,N_2274);
and U2321 (N_2321,N_2243,N_2272);
nor U2322 (N_2322,N_2275,N_2272);
and U2323 (N_2323,N_2273,N_2264);
and U2324 (N_2324,N_2245,N_2258);
or U2325 (N_2325,N_2279,N_2252);
nand U2326 (N_2326,N_2266,N_2254);
nor U2327 (N_2327,N_2244,N_2262);
nor U2328 (N_2328,N_2252,N_2239);
and U2329 (N_2329,N_2262,N_2232);
nor U2330 (N_2330,N_2262,N_2253);
or U2331 (N_2331,N_2223,N_2248);
and U2332 (N_2332,N_2223,N_2226);
nor U2333 (N_2333,N_2271,N_2251);
or U2334 (N_2334,N_2242,N_2243);
nor U2335 (N_2335,N_2240,N_2267);
nor U2336 (N_2336,N_2251,N_2276);
xor U2337 (N_2337,N_2235,N_2258);
nor U2338 (N_2338,N_2225,N_2267);
nor U2339 (N_2339,N_2277,N_2235);
nand U2340 (N_2340,N_2309,N_2332);
nand U2341 (N_2341,N_2311,N_2310);
or U2342 (N_2342,N_2339,N_2297);
and U2343 (N_2343,N_2301,N_2300);
and U2344 (N_2344,N_2286,N_2285);
and U2345 (N_2345,N_2291,N_2336);
and U2346 (N_2346,N_2293,N_2287);
nand U2347 (N_2347,N_2282,N_2319);
or U2348 (N_2348,N_2315,N_2308);
and U2349 (N_2349,N_2298,N_2320);
nor U2350 (N_2350,N_2304,N_2324);
and U2351 (N_2351,N_2295,N_2314);
or U2352 (N_2352,N_2281,N_2329);
nor U2353 (N_2353,N_2294,N_2321);
nand U2354 (N_2354,N_2305,N_2303);
or U2355 (N_2355,N_2322,N_2283);
nor U2356 (N_2356,N_2318,N_2284);
nand U2357 (N_2357,N_2313,N_2302);
nand U2358 (N_2358,N_2327,N_2338);
nand U2359 (N_2359,N_2330,N_2326);
nand U2360 (N_2360,N_2323,N_2333);
and U2361 (N_2361,N_2325,N_2306);
nand U2362 (N_2362,N_2296,N_2307);
nor U2363 (N_2363,N_2299,N_2280);
nand U2364 (N_2364,N_2288,N_2312);
nand U2365 (N_2365,N_2316,N_2292);
and U2366 (N_2366,N_2328,N_2337);
and U2367 (N_2367,N_2334,N_2317);
nor U2368 (N_2368,N_2331,N_2290);
or U2369 (N_2369,N_2335,N_2289);
or U2370 (N_2370,N_2338,N_2290);
nor U2371 (N_2371,N_2310,N_2293);
nand U2372 (N_2372,N_2290,N_2313);
or U2373 (N_2373,N_2314,N_2322);
or U2374 (N_2374,N_2291,N_2337);
and U2375 (N_2375,N_2288,N_2305);
nand U2376 (N_2376,N_2325,N_2285);
nand U2377 (N_2377,N_2306,N_2281);
xnor U2378 (N_2378,N_2298,N_2284);
or U2379 (N_2379,N_2327,N_2335);
or U2380 (N_2380,N_2324,N_2298);
nor U2381 (N_2381,N_2311,N_2332);
nor U2382 (N_2382,N_2332,N_2327);
nor U2383 (N_2383,N_2318,N_2295);
or U2384 (N_2384,N_2336,N_2298);
nor U2385 (N_2385,N_2293,N_2307);
and U2386 (N_2386,N_2309,N_2326);
and U2387 (N_2387,N_2298,N_2309);
nand U2388 (N_2388,N_2337,N_2289);
and U2389 (N_2389,N_2289,N_2281);
and U2390 (N_2390,N_2285,N_2283);
nor U2391 (N_2391,N_2285,N_2281);
and U2392 (N_2392,N_2287,N_2297);
nand U2393 (N_2393,N_2309,N_2310);
or U2394 (N_2394,N_2300,N_2339);
or U2395 (N_2395,N_2294,N_2302);
nor U2396 (N_2396,N_2318,N_2303);
nand U2397 (N_2397,N_2284,N_2283);
and U2398 (N_2398,N_2328,N_2299);
nand U2399 (N_2399,N_2312,N_2320);
or U2400 (N_2400,N_2366,N_2345);
nor U2401 (N_2401,N_2343,N_2395);
or U2402 (N_2402,N_2372,N_2362);
or U2403 (N_2403,N_2393,N_2392);
nand U2404 (N_2404,N_2379,N_2346);
nor U2405 (N_2405,N_2350,N_2365);
and U2406 (N_2406,N_2368,N_2389);
nor U2407 (N_2407,N_2374,N_2369);
nand U2408 (N_2408,N_2399,N_2384);
and U2409 (N_2409,N_2348,N_2378);
and U2410 (N_2410,N_2347,N_2386);
nor U2411 (N_2411,N_2371,N_2357);
or U2412 (N_2412,N_2364,N_2341);
and U2413 (N_2413,N_2381,N_2340);
and U2414 (N_2414,N_2359,N_2342);
or U2415 (N_2415,N_2380,N_2383);
or U2416 (N_2416,N_2385,N_2375);
or U2417 (N_2417,N_2344,N_2349);
nand U2418 (N_2418,N_2353,N_2358);
and U2419 (N_2419,N_2376,N_2387);
nor U2420 (N_2420,N_2354,N_2373);
and U2421 (N_2421,N_2377,N_2397);
nand U2422 (N_2422,N_2367,N_2356);
or U2423 (N_2423,N_2352,N_2360);
and U2424 (N_2424,N_2351,N_2396);
and U2425 (N_2425,N_2388,N_2355);
and U2426 (N_2426,N_2390,N_2398);
nor U2427 (N_2427,N_2382,N_2363);
nor U2428 (N_2428,N_2391,N_2361);
or U2429 (N_2429,N_2394,N_2370);
or U2430 (N_2430,N_2354,N_2375);
nor U2431 (N_2431,N_2379,N_2397);
nor U2432 (N_2432,N_2362,N_2392);
and U2433 (N_2433,N_2372,N_2354);
and U2434 (N_2434,N_2384,N_2358);
nor U2435 (N_2435,N_2395,N_2354);
or U2436 (N_2436,N_2361,N_2358);
nor U2437 (N_2437,N_2341,N_2387);
or U2438 (N_2438,N_2398,N_2393);
nor U2439 (N_2439,N_2382,N_2387);
nand U2440 (N_2440,N_2373,N_2364);
and U2441 (N_2441,N_2368,N_2395);
and U2442 (N_2442,N_2347,N_2358);
or U2443 (N_2443,N_2365,N_2381);
and U2444 (N_2444,N_2356,N_2341);
and U2445 (N_2445,N_2390,N_2378);
or U2446 (N_2446,N_2355,N_2395);
nand U2447 (N_2447,N_2353,N_2359);
or U2448 (N_2448,N_2363,N_2356);
nor U2449 (N_2449,N_2386,N_2361);
nand U2450 (N_2450,N_2352,N_2342);
nor U2451 (N_2451,N_2383,N_2370);
nor U2452 (N_2452,N_2366,N_2341);
nor U2453 (N_2453,N_2393,N_2391);
or U2454 (N_2454,N_2344,N_2366);
nor U2455 (N_2455,N_2354,N_2390);
and U2456 (N_2456,N_2341,N_2346);
nand U2457 (N_2457,N_2399,N_2364);
and U2458 (N_2458,N_2387,N_2381);
or U2459 (N_2459,N_2361,N_2375);
nand U2460 (N_2460,N_2418,N_2413);
nand U2461 (N_2461,N_2427,N_2401);
nand U2462 (N_2462,N_2440,N_2435);
and U2463 (N_2463,N_2430,N_2448);
nor U2464 (N_2464,N_2423,N_2416);
nand U2465 (N_2465,N_2438,N_2417);
nor U2466 (N_2466,N_2451,N_2403);
nand U2467 (N_2467,N_2449,N_2434);
nor U2468 (N_2468,N_2429,N_2437);
and U2469 (N_2469,N_2455,N_2411);
nor U2470 (N_2470,N_2405,N_2443);
nor U2471 (N_2471,N_2452,N_2456);
nor U2472 (N_2472,N_2424,N_2408);
or U2473 (N_2473,N_2436,N_2453);
nand U2474 (N_2474,N_2409,N_2410);
nand U2475 (N_2475,N_2450,N_2419);
nand U2476 (N_2476,N_2447,N_2445);
and U2477 (N_2477,N_2415,N_2414);
and U2478 (N_2478,N_2431,N_2439);
nor U2479 (N_2479,N_2406,N_2432);
nor U2480 (N_2480,N_2428,N_2444);
or U2481 (N_2481,N_2459,N_2400);
and U2482 (N_2482,N_2458,N_2404);
nand U2483 (N_2483,N_2412,N_2446);
and U2484 (N_2484,N_2442,N_2426);
nand U2485 (N_2485,N_2402,N_2421);
and U2486 (N_2486,N_2425,N_2457);
nand U2487 (N_2487,N_2441,N_2433);
and U2488 (N_2488,N_2420,N_2454);
or U2489 (N_2489,N_2422,N_2407);
and U2490 (N_2490,N_2456,N_2441);
and U2491 (N_2491,N_2423,N_2432);
nor U2492 (N_2492,N_2422,N_2445);
nand U2493 (N_2493,N_2443,N_2447);
nand U2494 (N_2494,N_2434,N_2416);
nor U2495 (N_2495,N_2456,N_2417);
nor U2496 (N_2496,N_2437,N_2456);
or U2497 (N_2497,N_2456,N_2444);
or U2498 (N_2498,N_2417,N_2449);
and U2499 (N_2499,N_2421,N_2413);
nor U2500 (N_2500,N_2455,N_2421);
nor U2501 (N_2501,N_2400,N_2402);
or U2502 (N_2502,N_2409,N_2434);
or U2503 (N_2503,N_2415,N_2408);
nand U2504 (N_2504,N_2418,N_2406);
nor U2505 (N_2505,N_2426,N_2414);
or U2506 (N_2506,N_2405,N_2427);
and U2507 (N_2507,N_2438,N_2429);
and U2508 (N_2508,N_2431,N_2445);
nor U2509 (N_2509,N_2441,N_2431);
or U2510 (N_2510,N_2430,N_2441);
nand U2511 (N_2511,N_2437,N_2408);
nor U2512 (N_2512,N_2411,N_2405);
or U2513 (N_2513,N_2418,N_2423);
nand U2514 (N_2514,N_2407,N_2404);
or U2515 (N_2515,N_2416,N_2433);
or U2516 (N_2516,N_2401,N_2416);
nor U2517 (N_2517,N_2402,N_2440);
nand U2518 (N_2518,N_2454,N_2400);
or U2519 (N_2519,N_2414,N_2403);
nand U2520 (N_2520,N_2464,N_2501);
and U2521 (N_2521,N_2474,N_2484);
and U2522 (N_2522,N_2508,N_2489);
and U2523 (N_2523,N_2485,N_2514);
nand U2524 (N_2524,N_2481,N_2505);
nand U2525 (N_2525,N_2482,N_2471);
or U2526 (N_2526,N_2495,N_2494);
nand U2527 (N_2527,N_2462,N_2478);
nor U2528 (N_2528,N_2504,N_2463);
and U2529 (N_2529,N_2517,N_2487);
nor U2530 (N_2530,N_2519,N_2512);
nor U2531 (N_2531,N_2461,N_2509);
nor U2532 (N_2532,N_2476,N_2499);
and U2533 (N_2533,N_2493,N_2472);
or U2534 (N_2534,N_2510,N_2475);
nand U2535 (N_2535,N_2513,N_2502);
xor U2536 (N_2536,N_2488,N_2469);
and U2537 (N_2537,N_2491,N_2506);
or U2538 (N_2538,N_2518,N_2486);
nand U2539 (N_2539,N_2490,N_2479);
or U2540 (N_2540,N_2497,N_2498);
and U2541 (N_2541,N_2467,N_2503);
nor U2542 (N_2542,N_2500,N_2465);
or U2543 (N_2543,N_2515,N_2468);
and U2544 (N_2544,N_2470,N_2492);
or U2545 (N_2545,N_2507,N_2477);
nand U2546 (N_2546,N_2511,N_2483);
or U2547 (N_2547,N_2516,N_2466);
nor U2548 (N_2548,N_2473,N_2496);
or U2549 (N_2549,N_2460,N_2480);
nand U2550 (N_2550,N_2512,N_2463);
and U2551 (N_2551,N_2505,N_2478);
nor U2552 (N_2552,N_2479,N_2474);
or U2553 (N_2553,N_2512,N_2496);
and U2554 (N_2554,N_2480,N_2479);
or U2555 (N_2555,N_2500,N_2478);
xnor U2556 (N_2556,N_2494,N_2512);
nor U2557 (N_2557,N_2515,N_2518);
or U2558 (N_2558,N_2467,N_2518);
or U2559 (N_2559,N_2486,N_2460);
or U2560 (N_2560,N_2489,N_2473);
or U2561 (N_2561,N_2494,N_2489);
nor U2562 (N_2562,N_2474,N_2493);
xor U2563 (N_2563,N_2498,N_2510);
nand U2564 (N_2564,N_2493,N_2480);
and U2565 (N_2565,N_2466,N_2488);
and U2566 (N_2566,N_2488,N_2491);
nand U2567 (N_2567,N_2505,N_2466);
nor U2568 (N_2568,N_2503,N_2509);
nand U2569 (N_2569,N_2469,N_2498);
nor U2570 (N_2570,N_2490,N_2472);
nor U2571 (N_2571,N_2502,N_2464);
nand U2572 (N_2572,N_2485,N_2463);
and U2573 (N_2573,N_2470,N_2506);
and U2574 (N_2574,N_2486,N_2497);
or U2575 (N_2575,N_2466,N_2485);
and U2576 (N_2576,N_2478,N_2495);
and U2577 (N_2577,N_2490,N_2471);
or U2578 (N_2578,N_2500,N_2486);
xor U2579 (N_2579,N_2494,N_2474);
and U2580 (N_2580,N_2534,N_2557);
nor U2581 (N_2581,N_2555,N_2569);
or U2582 (N_2582,N_2530,N_2522);
and U2583 (N_2583,N_2537,N_2551);
and U2584 (N_2584,N_2546,N_2570);
nand U2585 (N_2585,N_2575,N_2566);
or U2586 (N_2586,N_2542,N_2558);
nor U2587 (N_2587,N_2552,N_2538);
and U2588 (N_2588,N_2526,N_2579);
nand U2589 (N_2589,N_2573,N_2520);
nor U2590 (N_2590,N_2547,N_2565);
nand U2591 (N_2591,N_2525,N_2536);
or U2592 (N_2592,N_2567,N_2564);
nand U2593 (N_2593,N_2529,N_2523);
or U2594 (N_2594,N_2560,N_2550);
nor U2595 (N_2595,N_2521,N_2554);
or U2596 (N_2596,N_2563,N_2541);
nand U2597 (N_2597,N_2577,N_2548);
nor U2598 (N_2598,N_2561,N_2574);
nand U2599 (N_2599,N_2556,N_2539);
nor U2600 (N_2600,N_2535,N_2553);
or U2601 (N_2601,N_2528,N_2544);
nand U2602 (N_2602,N_2568,N_2576);
or U2603 (N_2603,N_2572,N_2532);
nor U2604 (N_2604,N_2549,N_2562);
nand U2605 (N_2605,N_2571,N_2540);
and U2606 (N_2606,N_2543,N_2533);
or U2607 (N_2607,N_2578,N_2527);
and U2608 (N_2608,N_2545,N_2524);
nor U2609 (N_2609,N_2559,N_2531);
nand U2610 (N_2610,N_2533,N_2523);
nor U2611 (N_2611,N_2579,N_2536);
nor U2612 (N_2612,N_2547,N_2533);
or U2613 (N_2613,N_2523,N_2562);
nand U2614 (N_2614,N_2536,N_2562);
nor U2615 (N_2615,N_2534,N_2532);
or U2616 (N_2616,N_2578,N_2550);
nand U2617 (N_2617,N_2539,N_2567);
or U2618 (N_2618,N_2529,N_2565);
nor U2619 (N_2619,N_2538,N_2521);
nand U2620 (N_2620,N_2533,N_2536);
nor U2621 (N_2621,N_2530,N_2531);
and U2622 (N_2622,N_2537,N_2569);
nand U2623 (N_2623,N_2568,N_2546);
and U2624 (N_2624,N_2530,N_2544);
and U2625 (N_2625,N_2525,N_2534);
and U2626 (N_2626,N_2550,N_2542);
nor U2627 (N_2627,N_2566,N_2570);
nor U2628 (N_2628,N_2532,N_2560);
or U2629 (N_2629,N_2532,N_2553);
nand U2630 (N_2630,N_2523,N_2539);
nor U2631 (N_2631,N_2575,N_2528);
nand U2632 (N_2632,N_2554,N_2579);
nand U2633 (N_2633,N_2529,N_2531);
and U2634 (N_2634,N_2532,N_2530);
nor U2635 (N_2635,N_2562,N_2554);
nor U2636 (N_2636,N_2569,N_2548);
nand U2637 (N_2637,N_2527,N_2571);
and U2638 (N_2638,N_2572,N_2533);
nor U2639 (N_2639,N_2552,N_2544);
or U2640 (N_2640,N_2589,N_2599);
nor U2641 (N_2641,N_2584,N_2616);
nor U2642 (N_2642,N_2613,N_2638);
nand U2643 (N_2643,N_2609,N_2593);
nand U2644 (N_2644,N_2582,N_2581);
nand U2645 (N_2645,N_2592,N_2639);
and U2646 (N_2646,N_2627,N_2605);
nor U2647 (N_2647,N_2617,N_2600);
xnor U2648 (N_2648,N_2632,N_2628);
nor U2649 (N_2649,N_2635,N_2619);
nor U2650 (N_2650,N_2634,N_2621);
nand U2651 (N_2651,N_2586,N_2596);
nand U2652 (N_2652,N_2604,N_2629);
nor U2653 (N_2653,N_2618,N_2580);
or U2654 (N_2654,N_2611,N_2612);
nor U2655 (N_2655,N_2633,N_2583);
and U2656 (N_2656,N_2597,N_2595);
or U2657 (N_2657,N_2637,N_2601);
or U2658 (N_2658,N_2620,N_2594);
and U2659 (N_2659,N_2606,N_2615);
nand U2660 (N_2660,N_2585,N_2631);
nor U2661 (N_2661,N_2607,N_2598);
and U2662 (N_2662,N_2630,N_2588);
nand U2663 (N_2663,N_2610,N_2591);
nand U2664 (N_2664,N_2625,N_2626);
and U2665 (N_2665,N_2602,N_2624);
nand U2666 (N_2666,N_2608,N_2603);
nand U2667 (N_2667,N_2636,N_2623);
and U2668 (N_2668,N_2587,N_2590);
nor U2669 (N_2669,N_2614,N_2622);
nand U2670 (N_2670,N_2632,N_2614);
and U2671 (N_2671,N_2601,N_2608);
and U2672 (N_2672,N_2586,N_2623);
nor U2673 (N_2673,N_2634,N_2615);
nor U2674 (N_2674,N_2602,N_2617);
nand U2675 (N_2675,N_2609,N_2600);
nor U2676 (N_2676,N_2607,N_2605);
and U2677 (N_2677,N_2608,N_2619);
nor U2678 (N_2678,N_2628,N_2602);
xor U2679 (N_2679,N_2610,N_2613);
or U2680 (N_2680,N_2610,N_2606);
nor U2681 (N_2681,N_2618,N_2638);
nand U2682 (N_2682,N_2625,N_2603);
and U2683 (N_2683,N_2618,N_2592);
nand U2684 (N_2684,N_2637,N_2587);
or U2685 (N_2685,N_2587,N_2618);
nor U2686 (N_2686,N_2613,N_2601);
and U2687 (N_2687,N_2616,N_2588);
nor U2688 (N_2688,N_2639,N_2605);
or U2689 (N_2689,N_2612,N_2631);
or U2690 (N_2690,N_2604,N_2609);
or U2691 (N_2691,N_2593,N_2633);
or U2692 (N_2692,N_2580,N_2631);
and U2693 (N_2693,N_2589,N_2617);
nand U2694 (N_2694,N_2589,N_2595);
nor U2695 (N_2695,N_2605,N_2616);
nor U2696 (N_2696,N_2581,N_2633);
nor U2697 (N_2697,N_2622,N_2591);
nand U2698 (N_2698,N_2610,N_2611);
and U2699 (N_2699,N_2585,N_2616);
or U2700 (N_2700,N_2642,N_2682);
nand U2701 (N_2701,N_2663,N_2664);
nand U2702 (N_2702,N_2695,N_2681);
or U2703 (N_2703,N_2692,N_2693);
or U2704 (N_2704,N_2640,N_2680);
nand U2705 (N_2705,N_2648,N_2644);
nand U2706 (N_2706,N_2670,N_2691);
and U2707 (N_2707,N_2684,N_2671);
or U2708 (N_2708,N_2659,N_2689);
nand U2709 (N_2709,N_2688,N_2650);
and U2710 (N_2710,N_2687,N_2672);
nand U2711 (N_2711,N_2655,N_2665);
nand U2712 (N_2712,N_2658,N_2679);
nand U2713 (N_2713,N_2643,N_2647);
and U2714 (N_2714,N_2675,N_2690);
or U2715 (N_2715,N_2668,N_2657);
nor U2716 (N_2716,N_2660,N_2698);
nand U2717 (N_2717,N_2641,N_2649);
nand U2718 (N_2718,N_2697,N_2651);
nand U2719 (N_2719,N_2661,N_2646);
and U2720 (N_2720,N_2676,N_2696);
or U2721 (N_2721,N_2677,N_2685);
nand U2722 (N_2722,N_2666,N_2686);
nor U2723 (N_2723,N_2645,N_2662);
and U2724 (N_2724,N_2669,N_2673);
or U2725 (N_2725,N_2694,N_2654);
nor U2726 (N_2726,N_2653,N_2674);
nand U2727 (N_2727,N_2678,N_2683);
and U2728 (N_2728,N_2667,N_2699);
and U2729 (N_2729,N_2656,N_2652);
nand U2730 (N_2730,N_2654,N_2674);
xnor U2731 (N_2731,N_2673,N_2661);
and U2732 (N_2732,N_2688,N_2644);
nor U2733 (N_2733,N_2661,N_2664);
nand U2734 (N_2734,N_2646,N_2658);
and U2735 (N_2735,N_2654,N_2682);
or U2736 (N_2736,N_2696,N_2675);
or U2737 (N_2737,N_2690,N_2670);
and U2738 (N_2738,N_2649,N_2672);
nor U2739 (N_2739,N_2658,N_2673);
nor U2740 (N_2740,N_2679,N_2657);
nor U2741 (N_2741,N_2676,N_2654);
nor U2742 (N_2742,N_2697,N_2654);
or U2743 (N_2743,N_2661,N_2652);
nor U2744 (N_2744,N_2655,N_2689);
nand U2745 (N_2745,N_2649,N_2661);
xnor U2746 (N_2746,N_2663,N_2692);
nor U2747 (N_2747,N_2675,N_2685);
nand U2748 (N_2748,N_2696,N_2657);
nand U2749 (N_2749,N_2696,N_2669);
nor U2750 (N_2750,N_2673,N_2678);
or U2751 (N_2751,N_2692,N_2696);
xor U2752 (N_2752,N_2645,N_2684);
and U2753 (N_2753,N_2678,N_2679);
nor U2754 (N_2754,N_2689,N_2690);
nand U2755 (N_2755,N_2696,N_2664);
nor U2756 (N_2756,N_2645,N_2697);
and U2757 (N_2757,N_2652,N_2659);
nor U2758 (N_2758,N_2658,N_2653);
or U2759 (N_2759,N_2643,N_2667);
and U2760 (N_2760,N_2712,N_2727);
and U2761 (N_2761,N_2738,N_2725);
nor U2762 (N_2762,N_2741,N_2757);
or U2763 (N_2763,N_2732,N_2728);
nor U2764 (N_2764,N_2735,N_2724);
or U2765 (N_2765,N_2756,N_2720);
nand U2766 (N_2766,N_2734,N_2711);
nor U2767 (N_2767,N_2750,N_2721);
nor U2768 (N_2768,N_2751,N_2744);
or U2769 (N_2769,N_2737,N_2703);
and U2770 (N_2770,N_2705,N_2746);
nand U2771 (N_2771,N_2719,N_2715);
and U2772 (N_2772,N_2736,N_2723);
nor U2773 (N_2773,N_2730,N_2707);
and U2774 (N_2774,N_2733,N_2729);
nor U2775 (N_2775,N_2714,N_2743);
nor U2776 (N_2776,N_2709,N_2700);
and U2777 (N_2777,N_2748,N_2742);
nand U2778 (N_2778,N_2753,N_2754);
or U2779 (N_2779,N_2745,N_2739);
or U2780 (N_2780,N_2717,N_2702);
nand U2781 (N_2781,N_2718,N_2713);
nor U2782 (N_2782,N_2740,N_2749);
or U2783 (N_2783,N_2701,N_2726);
nor U2784 (N_2784,N_2752,N_2708);
nand U2785 (N_2785,N_2716,N_2722);
or U2786 (N_2786,N_2747,N_2706);
nor U2787 (N_2787,N_2710,N_2755);
nand U2788 (N_2788,N_2704,N_2758);
or U2789 (N_2789,N_2759,N_2731);
and U2790 (N_2790,N_2753,N_2732);
and U2791 (N_2791,N_2705,N_2708);
nor U2792 (N_2792,N_2748,N_2741);
and U2793 (N_2793,N_2752,N_2734);
and U2794 (N_2794,N_2741,N_2758);
nand U2795 (N_2795,N_2728,N_2740);
and U2796 (N_2796,N_2758,N_2751);
and U2797 (N_2797,N_2725,N_2732);
nor U2798 (N_2798,N_2738,N_2749);
nor U2799 (N_2799,N_2725,N_2739);
nor U2800 (N_2800,N_2701,N_2750);
nand U2801 (N_2801,N_2759,N_2717);
or U2802 (N_2802,N_2747,N_2712);
nand U2803 (N_2803,N_2759,N_2755);
or U2804 (N_2804,N_2748,N_2703);
and U2805 (N_2805,N_2724,N_2707);
nand U2806 (N_2806,N_2727,N_2749);
nor U2807 (N_2807,N_2713,N_2710);
nor U2808 (N_2808,N_2727,N_2719);
or U2809 (N_2809,N_2718,N_2748);
nor U2810 (N_2810,N_2744,N_2719);
or U2811 (N_2811,N_2727,N_2713);
or U2812 (N_2812,N_2727,N_2715);
or U2813 (N_2813,N_2702,N_2712);
or U2814 (N_2814,N_2705,N_2721);
nor U2815 (N_2815,N_2722,N_2726);
nand U2816 (N_2816,N_2744,N_2713);
and U2817 (N_2817,N_2721,N_2703);
nor U2818 (N_2818,N_2758,N_2706);
and U2819 (N_2819,N_2737,N_2738);
nand U2820 (N_2820,N_2779,N_2793);
nand U2821 (N_2821,N_2775,N_2772);
xnor U2822 (N_2822,N_2774,N_2814);
xnor U2823 (N_2823,N_2765,N_2813);
or U2824 (N_2824,N_2796,N_2787);
nor U2825 (N_2825,N_2781,N_2762);
nor U2826 (N_2826,N_2769,N_2782);
and U2827 (N_2827,N_2806,N_2805);
nor U2828 (N_2828,N_2770,N_2780);
nor U2829 (N_2829,N_2777,N_2815);
nand U2830 (N_2830,N_2800,N_2791);
or U2831 (N_2831,N_2812,N_2790);
or U2832 (N_2832,N_2817,N_2766);
and U2833 (N_2833,N_2792,N_2807);
nor U2834 (N_2834,N_2761,N_2767);
nor U2835 (N_2835,N_2768,N_2803);
nand U2836 (N_2836,N_2771,N_2764);
nor U2837 (N_2837,N_2799,N_2818);
or U2838 (N_2838,N_2788,N_2811);
or U2839 (N_2839,N_2789,N_2797);
and U2840 (N_2840,N_2810,N_2808);
or U2841 (N_2841,N_2798,N_2776);
and U2842 (N_2842,N_2785,N_2783);
and U2843 (N_2843,N_2773,N_2778);
nor U2844 (N_2844,N_2819,N_2795);
or U2845 (N_2845,N_2786,N_2784);
nand U2846 (N_2846,N_2802,N_2809);
or U2847 (N_2847,N_2804,N_2763);
nand U2848 (N_2848,N_2760,N_2801);
nand U2849 (N_2849,N_2816,N_2794);
or U2850 (N_2850,N_2790,N_2766);
nor U2851 (N_2851,N_2770,N_2812);
or U2852 (N_2852,N_2779,N_2774);
or U2853 (N_2853,N_2814,N_2770);
nand U2854 (N_2854,N_2766,N_2789);
nor U2855 (N_2855,N_2793,N_2766);
nor U2856 (N_2856,N_2772,N_2760);
nand U2857 (N_2857,N_2796,N_2760);
nand U2858 (N_2858,N_2801,N_2778);
or U2859 (N_2859,N_2798,N_2773);
nand U2860 (N_2860,N_2790,N_2762);
and U2861 (N_2861,N_2811,N_2815);
nand U2862 (N_2862,N_2810,N_2798);
nor U2863 (N_2863,N_2767,N_2783);
nor U2864 (N_2864,N_2803,N_2813);
nand U2865 (N_2865,N_2787,N_2792);
or U2866 (N_2866,N_2810,N_2814);
nor U2867 (N_2867,N_2765,N_2761);
and U2868 (N_2868,N_2769,N_2784);
nand U2869 (N_2869,N_2787,N_2818);
or U2870 (N_2870,N_2760,N_2816);
nor U2871 (N_2871,N_2800,N_2795);
and U2872 (N_2872,N_2764,N_2818);
nand U2873 (N_2873,N_2819,N_2814);
nand U2874 (N_2874,N_2779,N_2764);
or U2875 (N_2875,N_2774,N_2803);
or U2876 (N_2876,N_2774,N_2788);
or U2877 (N_2877,N_2805,N_2797);
or U2878 (N_2878,N_2809,N_2813);
nor U2879 (N_2879,N_2786,N_2807);
nor U2880 (N_2880,N_2820,N_2870);
nand U2881 (N_2881,N_2879,N_2873);
nor U2882 (N_2882,N_2876,N_2868);
nand U2883 (N_2883,N_2836,N_2838);
xnor U2884 (N_2884,N_2844,N_2878);
nor U2885 (N_2885,N_2863,N_2875);
or U2886 (N_2886,N_2824,N_2841);
nor U2887 (N_2887,N_2861,N_2867);
or U2888 (N_2888,N_2835,N_2862);
and U2889 (N_2889,N_2860,N_2831);
nand U2890 (N_2890,N_2833,N_2874);
and U2891 (N_2891,N_2837,N_2854);
nor U2892 (N_2892,N_2859,N_2832);
nand U2893 (N_2893,N_2855,N_2846);
nor U2894 (N_2894,N_2853,N_2858);
and U2895 (N_2895,N_2840,N_2865);
and U2896 (N_2896,N_2848,N_2857);
nand U2897 (N_2897,N_2847,N_2851);
or U2898 (N_2898,N_2839,N_2823);
xor U2899 (N_2899,N_2866,N_2849);
and U2900 (N_2900,N_2871,N_2845);
nor U2901 (N_2901,N_2869,N_2830);
and U2902 (N_2902,N_2827,N_2864);
nand U2903 (N_2903,N_2821,N_2828);
and U2904 (N_2904,N_2826,N_2822);
nor U2905 (N_2905,N_2843,N_2856);
and U2906 (N_2906,N_2852,N_2842);
and U2907 (N_2907,N_2877,N_2829);
or U2908 (N_2908,N_2872,N_2834);
or U2909 (N_2909,N_2850,N_2825);
or U2910 (N_2910,N_2846,N_2866);
and U2911 (N_2911,N_2837,N_2872);
nor U2912 (N_2912,N_2848,N_2866);
or U2913 (N_2913,N_2840,N_2848);
and U2914 (N_2914,N_2830,N_2844);
and U2915 (N_2915,N_2856,N_2827);
nor U2916 (N_2916,N_2828,N_2864);
nand U2917 (N_2917,N_2822,N_2830);
and U2918 (N_2918,N_2860,N_2841);
nand U2919 (N_2919,N_2840,N_2842);
nor U2920 (N_2920,N_2873,N_2822);
nand U2921 (N_2921,N_2832,N_2846);
or U2922 (N_2922,N_2851,N_2864);
nor U2923 (N_2923,N_2823,N_2820);
or U2924 (N_2924,N_2837,N_2840);
and U2925 (N_2925,N_2856,N_2832);
and U2926 (N_2926,N_2835,N_2828);
nand U2927 (N_2927,N_2825,N_2849);
nand U2928 (N_2928,N_2861,N_2856);
and U2929 (N_2929,N_2839,N_2873);
nand U2930 (N_2930,N_2821,N_2866);
nor U2931 (N_2931,N_2847,N_2833);
nand U2932 (N_2932,N_2826,N_2862);
nand U2933 (N_2933,N_2875,N_2853);
nand U2934 (N_2934,N_2861,N_2872);
or U2935 (N_2935,N_2861,N_2865);
nand U2936 (N_2936,N_2826,N_2875);
nand U2937 (N_2937,N_2864,N_2850);
or U2938 (N_2938,N_2866,N_2865);
nor U2939 (N_2939,N_2834,N_2866);
or U2940 (N_2940,N_2908,N_2926);
or U2941 (N_2941,N_2883,N_2937);
or U2942 (N_2942,N_2917,N_2938);
or U2943 (N_2943,N_2911,N_2882);
or U2944 (N_2944,N_2922,N_2903);
nor U2945 (N_2945,N_2929,N_2925);
nor U2946 (N_2946,N_2918,N_2899);
nand U2947 (N_2947,N_2910,N_2914);
or U2948 (N_2948,N_2885,N_2894);
nand U2949 (N_2949,N_2924,N_2912);
or U2950 (N_2950,N_2921,N_2905);
nor U2951 (N_2951,N_2900,N_2931);
and U2952 (N_2952,N_2881,N_2904);
and U2953 (N_2953,N_2928,N_2884);
and U2954 (N_2954,N_2880,N_2923);
nand U2955 (N_2955,N_2886,N_2895);
nand U2956 (N_2956,N_2891,N_2890);
nor U2957 (N_2957,N_2933,N_2913);
nand U2958 (N_2958,N_2930,N_2892);
nor U2959 (N_2959,N_2934,N_2932);
nand U2960 (N_2960,N_2935,N_2920);
or U2961 (N_2961,N_2898,N_2897);
or U2962 (N_2962,N_2919,N_2939);
and U2963 (N_2963,N_2887,N_2889);
and U2964 (N_2964,N_2936,N_2916);
nor U2965 (N_2965,N_2907,N_2896);
and U2966 (N_2966,N_2915,N_2927);
and U2967 (N_2967,N_2902,N_2906);
or U2968 (N_2968,N_2909,N_2893);
or U2969 (N_2969,N_2888,N_2901);
or U2970 (N_2970,N_2934,N_2897);
nand U2971 (N_2971,N_2916,N_2926);
nor U2972 (N_2972,N_2880,N_2883);
or U2973 (N_2973,N_2902,N_2927);
and U2974 (N_2974,N_2882,N_2937);
and U2975 (N_2975,N_2901,N_2916);
nor U2976 (N_2976,N_2932,N_2906);
and U2977 (N_2977,N_2908,N_2880);
nor U2978 (N_2978,N_2914,N_2935);
or U2979 (N_2979,N_2923,N_2932);
or U2980 (N_2980,N_2899,N_2886);
and U2981 (N_2981,N_2896,N_2913);
nand U2982 (N_2982,N_2891,N_2907);
nand U2983 (N_2983,N_2885,N_2892);
nor U2984 (N_2984,N_2890,N_2900);
and U2985 (N_2985,N_2936,N_2885);
nand U2986 (N_2986,N_2887,N_2939);
nor U2987 (N_2987,N_2930,N_2897);
nor U2988 (N_2988,N_2880,N_2905);
or U2989 (N_2989,N_2936,N_2903);
and U2990 (N_2990,N_2886,N_2918);
or U2991 (N_2991,N_2908,N_2906);
and U2992 (N_2992,N_2938,N_2889);
nand U2993 (N_2993,N_2893,N_2934);
nor U2994 (N_2994,N_2934,N_2886);
nand U2995 (N_2995,N_2908,N_2911);
nand U2996 (N_2996,N_2917,N_2894);
nor U2997 (N_2997,N_2891,N_2920);
and U2998 (N_2998,N_2904,N_2895);
nor U2999 (N_2999,N_2917,N_2882);
and UO_0 (O_0,N_2987,N_2998);
nand UO_1 (O_1,N_2975,N_2979);
nor UO_2 (O_2,N_2959,N_2976);
nand UO_3 (O_3,N_2946,N_2944);
nor UO_4 (O_4,N_2985,N_2948);
and UO_5 (O_5,N_2977,N_2964);
or UO_6 (O_6,N_2949,N_2957);
nor UO_7 (O_7,N_2974,N_2954);
and UO_8 (O_8,N_2988,N_2972);
nand UO_9 (O_9,N_2993,N_2994);
and UO_10 (O_10,N_2986,N_2984);
and UO_11 (O_11,N_2999,N_2956);
or UO_12 (O_12,N_2951,N_2983);
and UO_13 (O_13,N_2981,N_2990);
nand UO_14 (O_14,N_2978,N_2953);
nor UO_15 (O_15,N_2971,N_2962);
nor UO_16 (O_16,N_2950,N_2966);
and UO_17 (O_17,N_2989,N_2952);
and UO_18 (O_18,N_2960,N_2968);
or UO_19 (O_19,N_2963,N_2973);
or UO_20 (O_20,N_2942,N_2955);
nor UO_21 (O_21,N_2961,N_2997);
nor UO_22 (O_22,N_2940,N_2947);
nand UO_23 (O_23,N_2982,N_2996);
nor UO_24 (O_24,N_2943,N_2965);
or UO_25 (O_25,N_2970,N_2945);
nor UO_26 (O_26,N_2995,N_2969);
or UO_27 (O_27,N_2980,N_2991);
nand UO_28 (O_28,N_2992,N_2958);
or UO_29 (O_29,N_2967,N_2941);
or UO_30 (O_30,N_2986,N_2975);
or UO_31 (O_31,N_2972,N_2982);
nor UO_32 (O_32,N_2982,N_2976);
nor UO_33 (O_33,N_2975,N_2954);
nor UO_34 (O_34,N_2992,N_2953);
nor UO_35 (O_35,N_2986,N_2993);
and UO_36 (O_36,N_2953,N_2959);
nand UO_37 (O_37,N_2952,N_2963);
and UO_38 (O_38,N_2945,N_2983);
or UO_39 (O_39,N_2970,N_2993);
and UO_40 (O_40,N_2973,N_2964);
and UO_41 (O_41,N_2987,N_2947);
nand UO_42 (O_42,N_2966,N_2965);
nand UO_43 (O_43,N_2995,N_2989);
or UO_44 (O_44,N_2958,N_2988);
or UO_45 (O_45,N_2944,N_2955);
or UO_46 (O_46,N_2944,N_2963);
nand UO_47 (O_47,N_2984,N_2953);
nand UO_48 (O_48,N_2990,N_2975);
and UO_49 (O_49,N_2940,N_2984);
nand UO_50 (O_50,N_2991,N_2999);
and UO_51 (O_51,N_2958,N_2940);
or UO_52 (O_52,N_2944,N_2985);
and UO_53 (O_53,N_2989,N_2945);
nand UO_54 (O_54,N_2951,N_2957);
and UO_55 (O_55,N_2949,N_2998);
nand UO_56 (O_56,N_2981,N_2995);
and UO_57 (O_57,N_2969,N_2955);
nand UO_58 (O_58,N_2979,N_2940);
and UO_59 (O_59,N_2942,N_2987);
and UO_60 (O_60,N_2991,N_2981);
or UO_61 (O_61,N_2956,N_2977);
and UO_62 (O_62,N_2961,N_2957);
nand UO_63 (O_63,N_2949,N_2970);
nor UO_64 (O_64,N_2948,N_2992);
xor UO_65 (O_65,N_2988,N_2960);
nor UO_66 (O_66,N_2991,N_2960);
or UO_67 (O_67,N_2997,N_2992);
or UO_68 (O_68,N_2976,N_2989);
nand UO_69 (O_69,N_2982,N_2970);
xnor UO_70 (O_70,N_2967,N_2950);
and UO_71 (O_71,N_2949,N_2971);
or UO_72 (O_72,N_2941,N_2945);
nand UO_73 (O_73,N_2992,N_2975);
or UO_74 (O_74,N_2951,N_2962);
and UO_75 (O_75,N_2997,N_2968);
nor UO_76 (O_76,N_2981,N_2954);
nor UO_77 (O_77,N_2960,N_2969);
or UO_78 (O_78,N_2980,N_2970);
nor UO_79 (O_79,N_2959,N_2979);
nor UO_80 (O_80,N_2952,N_2942);
nand UO_81 (O_81,N_2950,N_2976);
nand UO_82 (O_82,N_2962,N_2967);
or UO_83 (O_83,N_2951,N_2948);
or UO_84 (O_84,N_2952,N_2948);
and UO_85 (O_85,N_2982,N_2984);
nor UO_86 (O_86,N_2972,N_2956);
and UO_87 (O_87,N_2942,N_2994);
and UO_88 (O_88,N_2960,N_2976);
and UO_89 (O_89,N_2940,N_2974);
and UO_90 (O_90,N_2940,N_2952);
nor UO_91 (O_91,N_2994,N_2941);
nor UO_92 (O_92,N_2941,N_2959);
nand UO_93 (O_93,N_2980,N_2947);
nand UO_94 (O_94,N_2972,N_2987);
nor UO_95 (O_95,N_2954,N_2942);
and UO_96 (O_96,N_2949,N_2975);
nand UO_97 (O_97,N_2948,N_2942);
or UO_98 (O_98,N_2976,N_2949);
nor UO_99 (O_99,N_2981,N_2947);
nand UO_100 (O_100,N_2983,N_2953);
nor UO_101 (O_101,N_2982,N_2960);
nand UO_102 (O_102,N_2973,N_2972);
and UO_103 (O_103,N_2990,N_2984);
nor UO_104 (O_104,N_2990,N_2964);
nor UO_105 (O_105,N_2965,N_2963);
nor UO_106 (O_106,N_2959,N_2997);
nor UO_107 (O_107,N_2980,N_2986);
nor UO_108 (O_108,N_2950,N_2972);
nor UO_109 (O_109,N_2953,N_2997);
and UO_110 (O_110,N_2966,N_2986);
and UO_111 (O_111,N_2989,N_2956);
nand UO_112 (O_112,N_2993,N_2979);
and UO_113 (O_113,N_2988,N_2965);
nand UO_114 (O_114,N_2994,N_2955);
and UO_115 (O_115,N_2985,N_2970);
and UO_116 (O_116,N_2984,N_2988);
or UO_117 (O_117,N_2966,N_2949);
and UO_118 (O_118,N_2994,N_2959);
and UO_119 (O_119,N_2964,N_2963);
nor UO_120 (O_120,N_2991,N_2959);
nor UO_121 (O_121,N_2959,N_2969);
and UO_122 (O_122,N_2949,N_2951);
and UO_123 (O_123,N_2945,N_2963);
nor UO_124 (O_124,N_2975,N_2966);
and UO_125 (O_125,N_2963,N_2998);
nand UO_126 (O_126,N_2995,N_2963);
and UO_127 (O_127,N_2985,N_2952);
nor UO_128 (O_128,N_2978,N_2950);
and UO_129 (O_129,N_2948,N_2978);
nand UO_130 (O_130,N_2964,N_2989);
or UO_131 (O_131,N_2970,N_2992);
or UO_132 (O_132,N_2951,N_2984);
or UO_133 (O_133,N_2945,N_2947);
and UO_134 (O_134,N_2977,N_2951);
nand UO_135 (O_135,N_2962,N_2989);
and UO_136 (O_136,N_2987,N_2944);
nand UO_137 (O_137,N_2953,N_2945);
or UO_138 (O_138,N_2999,N_2961);
nor UO_139 (O_139,N_2974,N_2959);
nand UO_140 (O_140,N_2974,N_2982);
nand UO_141 (O_141,N_2996,N_2995);
nor UO_142 (O_142,N_2958,N_2971);
or UO_143 (O_143,N_2960,N_2966);
or UO_144 (O_144,N_2960,N_2992);
and UO_145 (O_145,N_2941,N_2963);
xor UO_146 (O_146,N_2979,N_2945);
and UO_147 (O_147,N_2997,N_2975);
nor UO_148 (O_148,N_2942,N_2975);
xnor UO_149 (O_149,N_2990,N_2941);
and UO_150 (O_150,N_2991,N_2975);
nor UO_151 (O_151,N_2971,N_2955);
and UO_152 (O_152,N_2977,N_2979);
or UO_153 (O_153,N_2970,N_2974);
nand UO_154 (O_154,N_2967,N_2960);
and UO_155 (O_155,N_2950,N_2940);
nand UO_156 (O_156,N_2998,N_2950);
nand UO_157 (O_157,N_2951,N_2970);
or UO_158 (O_158,N_2958,N_2984);
or UO_159 (O_159,N_2978,N_2968);
nor UO_160 (O_160,N_2961,N_2998);
nor UO_161 (O_161,N_2960,N_2957);
nor UO_162 (O_162,N_2940,N_2956);
and UO_163 (O_163,N_2981,N_2970);
nor UO_164 (O_164,N_2976,N_2984);
and UO_165 (O_165,N_2950,N_2959);
or UO_166 (O_166,N_2982,N_2968);
nand UO_167 (O_167,N_2951,N_2950);
or UO_168 (O_168,N_2945,N_2993);
nand UO_169 (O_169,N_2969,N_2986);
nor UO_170 (O_170,N_2962,N_2984);
nor UO_171 (O_171,N_2945,N_2985);
or UO_172 (O_172,N_2941,N_2972);
nand UO_173 (O_173,N_2997,N_2966);
and UO_174 (O_174,N_2955,N_2963);
and UO_175 (O_175,N_2952,N_2955);
and UO_176 (O_176,N_2971,N_2950);
nor UO_177 (O_177,N_2974,N_2977);
nand UO_178 (O_178,N_2942,N_2950);
nand UO_179 (O_179,N_2968,N_2988);
nand UO_180 (O_180,N_2991,N_2978);
or UO_181 (O_181,N_2949,N_2984);
nand UO_182 (O_182,N_2946,N_2998);
and UO_183 (O_183,N_2999,N_2958);
nor UO_184 (O_184,N_2986,N_2948);
and UO_185 (O_185,N_2965,N_2947);
nor UO_186 (O_186,N_2996,N_2948);
and UO_187 (O_187,N_2987,N_2967);
nand UO_188 (O_188,N_2972,N_2948);
nor UO_189 (O_189,N_2963,N_2948);
and UO_190 (O_190,N_2954,N_2955);
nand UO_191 (O_191,N_2965,N_2982);
or UO_192 (O_192,N_2956,N_2987);
and UO_193 (O_193,N_2980,N_2994);
and UO_194 (O_194,N_2950,N_2979);
nor UO_195 (O_195,N_2992,N_2972);
and UO_196 (O_196,N_2980,N_2943);
and UO_197 (O_197,N_2954,N_2951);
and UO_198 (O_198,N_2982,N_2985);
nand UO_199 (O_199,N_2971,N_2996);
or UO_200 (O_200,N_2996,N_2987);
or UO_201 (O_201,N_2966,N_2977);
nand UO_202 (O_202,N_2960,N_2956);
and UO_203 (O_203,N_2940,N_2945);
nor UO_204 (O_204,N_2945,N_2968);
nor UO_205 (O_205,N_2964,N_2945);
and UO_206 (O_206,N_2947,N_2974);
or UO_207 (O_207,N_2971,N_2975);
nand UO_208 (O_208,N_2992,N_2976);
nor UO_209 (O_209,N_2966,N_2948);
nand UO_210 (O_210,N_2980,N_2977);
and UO_211 (O_211,N_2959,N_2945);
or UO_212 (O_212,N_2953,N_2948);
nand UO_213 (O_213,N_2959,N_2996);
xor UO_214 (O_214,N_2997,N_2999);
and UO_215 (O_215,N_2985,N_2993);
and UO_216 (O_216,N_2971,N_2999);
or UO_217 (O_217,N_2965,N_2994);
nor UO_218 (O_218,N_2997,N_2947);
and UO_219 (O_219,N_2953,N_2949);
nand UO_220 (O_220,N_2958,N_2950);
or UO_221 (O_221,N_2942,N_2957);
and UO_222 (O_222,N_2992,N_2945);
and UO_223 (O_223,N_2957,N_2968);
nor UO_224 (O_224,N_2947,N_2971);
and UO_225 (O_225,N_2940,N_2948);
nor UO_226 (O_226,N_2989,N_2959);
and UO_227 (O_227,N_2989,N_2975);
and UO_228 (O_228,N_2963,N_2974);
and UO_229 (O_229,N_2974,N_2995);
and UO_230 (O_230,N_2991,N_2964);
and UO_231 (O_231,N_2971,N_2957);
or UO_232 (O_232,N_2947,N_2942);
or UO_233 (O_233,N_2974,N_2988);
or UO_234 (O_234,N_2969,N_2976);
nor UO_235 (O_235,N_2963,N_2971);
or UO_236 (O_236,N_2993,N_2965);
or UO_237 (O_237,N_2987,N_2995);
or UO_238 (O_238,N_2985,N_2978);
nand UO_239 (O_239,N_2983,N_2988);
nand UO_240 (O_240,N_2941,N_2975);
nand UO_241 (O_241,N_2971,N_2965);
or UO_242 (O_242,N_2971,N_2985);
or UO_243 (O_243,N_2973,N_2970);
nand UO_244 (O_244,N_2967,N_2983);
or UO_245 (O_245,N_2978,N_2979);
nor UO_246 (O_246,N_2981,N_2977);
and UO_247 (O_247,N_2988,N_2944);
nor UO_248 (O_248,N_2959,N_2942);
and UO_249 (O_249,N_2957,N_2958);
nand UO_250 (O_250,N_2965,N_2981);
and UO_251 (O_251,N_2975,N_2976);
and UO_252 (O_252,N_2991,N_2949);
nand UO_253 (O_253,N_2985,N_2946);
nor UO_254 (O_254,N_2981,N_2982);
and UO_255 (O_255,N_2982,N_2990);
and UO_256 (O_256,N_2993,N_2950);
nor UO_257 (O_257,N_2970,N_2975);
or UO_258 (O_258,N_2971,N_2969);
nand UO_259 (O_259,N_2973,N_2940);
nand UO_260 (O_260,N_2954,N_2947);
and UO_261 (O_261,N_2959,N_2975);
nand UO_262 (O_262,N_2997,N_2972);
nor UO_263 (O_263,N_2991,N_2947);
nand UO_264 (O_264,N_2975,N_2977);
nand UO_265 (O_265,N_2950,N_2994);
and UO_266 (O_266,N_2996,N_2953);
or UO_267 (O_267,N_2998,N_2947);
or UO_268 (O_268,N_2948,N_2998);
nor UO_269 (O_269,N_2951,N_2987);
nand UO_270 (O_270,N_2955,N_2949);
nor UO_271 (O_271,N_2991,N_2962);
nor UO_272 (O_272,N_2943,N_2967);
nand UO_273 (O_273,N_2941,N_2971);
nand UO_274 (O_274,N_2993,N_2999);
or UO_275 (O_275,N_2968,N_2942);
nand UO_276 (O_276,N_2940,N_2954);
nand UO_277 (O_277,N_2986,N_2945);
nand UO_278 (O_278,N_2942,N_2999);
and UO_279 (O_279,N_2994,N_2987);
or UO_280 (O_280,N_2949,N_2987);
or UO_281 (O_281,N_2980,N_2983);
nand UO_282 (O_282,N_2988,N_2952);
or UO_283 (O_283,N_2974,N_2951);
nand UO_284 (O_284,N_2975,N_2967);
nand UO_285 (O_285,N_2991,N_2966);
or UO_286 (O_286,N_2979,N_2951);
nor UO_287 (O_287,N_2981,N_2980);
and UO_288 (O_288,N_2964,N_2999);
or UO_289 (O_289,N_2997,N_2982);
and UO_290 (O_290,N_2980,N_2961);
nor UO_291 (O_291,N_2947,N_2952);
nand UO_292 (O_292,N_2953,N_2940);
or UO_293 (O_293,N_2969,N_2999);
or UO_294 (O_294,N_2944,N_2974);
nor UO_295 (O_295,N_2954,N_2977);
and UO_296 (O_296,N_2980,N_2993);
and UO_297 (O_297,N_2947,N_2946);
or UO_298 (O_298,N_2999,N_2968);
nor UO_299 (O_299,N_2952,N_2981);
or UO_300 (O_300,N_2980,N_2992);
nand UO_301 (O_301,N_2974,N_2996);
nand UO_302 (O_302,N_2971,N_2991);
or UO_303 (O_303,N_2970,N_2967);
nand UO_304 (O_304,N_2977,N_2988);
or UO_305 (O_305,N_2949,N_2986);
and UO_306 (O_306,N_2963,N_2985);
and UO_307 (O_307,N_2948,N_2984);
or UO_308 (O_308,N_2964,N_2974);
nor UO_309 (O_309,N_2942,N_2977);
or UO_310 (O_310,N_2985,N_2975);
or UO_311 (O_311,N_2963,N_2950);
and UO_312 (O_312,N_2986,N_2985);
nor UO_313 (O_313,N_2961,N_2949);
nor UO_314 (O_314,N_2977,N_2963);
or UO_315 (O_315,N_2979,N_2942);
nand UO_316 (O_316,N_2945,N_2944);
or UO_317 (O_317,N_2978,N_2977);
nand UO_318 (O_318,N_2958,N_2979);
xnor UO_319 (O_319,N_2968,N_2977);
nor UO_320 (O_320,N_2980,N_2941);
and UO_321 (O_321,N_2967,N_2959);
nand UO_322 (O_322,N_2950,N_2990);
nor UO_323 (O_323,N_2969,N_2966);
and UO_324 (O_324,N_2985,N_2942);
nand UO_325 (O_325,N_2971,N_2973);
nor UO_326 (O_326,N_2962,N_2985);
nand UO_327 (O_327,N_2997,N_2994);
or UO_328 (O_328,N_2957,N_2992);
and UO_329 (O_329,N_2951,N_2976);
nor UO_330 (O_330,N_2945,N_2950);
or UO_331 (O_331,N_2988,N_2987);
nor UO_332 (O_332,N_2979,N_2991);
and UO_333 (O_333,N_2974,N_2973);
and UO_334 (O_334,N_2969,N_2953);
or UO_335 (O_335,N_2940,N_2960);
or UO_336 (O_336,N_2985,N_2977);
and UO_337 (O_337,N_2978,N_2969);
nand UO_338 (O_338,N_2985,N_2998);
or UO_339 (O_339,N_2948,N_2973);
nor UO_340 (O_340,N_2995,N_2978);
nor UO_341 (O_341,N_2984,N_2994);
and UO_342 (O_342,N_2996,N_2962);
or UO_343 (O_343,N_2995,N_2988);
or UO_344 (O_344,N_2996,N_2958);
or UO_345 (O_345,N_2998,N_2976);
and UO_346 (O_346,N_2956,N_2963);
and UO_347 (O_347,N_2966,N_2961);
nand UO_348 (O_348,N_2989,N_2984);
nand UO_349 (O_349,N_2945,N_2971);
nor UO_350 (O_350,N_2962,N_2949);
nand UO_351 (O_351,N_2966,N_2976);
nor UO_352 (O_352,N_2974,N_2966);
nor UO_353 (O_353,N_2988,N_2970);
and UO_354 (O_354,N_2977,N_2972);
nor UO_355 (O_355,N_2978,N_2988);
and UO_356 (O_356,N_2974,N_2958);
nor UO_357 (O_357,N_2981,N_2979);
and UO_358 (O_358,N_2980,N_2965);
and UO_359 (O_359,N_2993,N_2949);
or UO_360 (O_360,N_2981,N_2948);
and UO_361 (O_361,N_2990,N_2946);
nand UO_362 (O_362,N_2980,N_2995);
or UO_363 (O_363,N_2953,N_2976);
and UO_364 (O_364,N_2964,N_2984);
and UO_365 (O_365,N_2943,N_2978);
and UO_366 (O_366,N_2962,N_2969);
or UO_367 (O_367,N_2982,N_2989);
nand UO_368 (O_368,N_2984,N_2963);
nand UO_369 (O_369,N_2941,N_2955);
nor UO_370 (O_370,N_2947,N_2969);
and UO_371 (O_371,N_2989,N_2981);
nor UO_372 (O_372,N_2962,N_2963);
and UO_373 (O_373,N_2947,N_2993);
nand UO_374 (O_374,N_2966,N_2999);
and UO_375 (O_375,N_2950,N_2944);
nand UO_376 (O_376,N_2965,N_2949);
and UO_377 (O_377,N_2966,N_2964);
nor UO_378 (O_378,N_2975,N_2968);
and UO_379 (O_379,N_2963,N_2981);
or UO_380 (O_380,N_2968,N_2970);
nor UO_381 (O_381,N_2995,N_2994);
nor UO_382 (O_382,N_2944,N_2977);
or UO_383 (O_383,N_2997,N_2973);
and UO_384 (O_384,N_2983,N_2974);
nand UO_385 (O_385,N_2956,N_2957);
nor UO_386 (O_386,N_2959,N_2980);
and UO_387 (O_387,N_2955,N_2976);
and UO_388 (O_388,N_2965,N_2989);
nor UO_389 (O_389,N_2945,N_2974);
and UO_390 (O_390,N_2940,N_2992);
and UO_391 (O_391,N_2949,N_2999);
nor UO_392 (O_392,N_2980,N_2985);
nor UO_393 (O_393,N_2948,N_2955);
nand UO_394 (O_394,N_2964,N_2957);
nand UO_395 (O_395,N_2997,N_2970);
and UO_396 (O_396,N_2996,N_2966);
nand UO_397 (O_397,N_2990,N_2954);
nor UO_398 (O_398,N_2942,N_2993);
nor UO_399 (O_399,N_2969,N_2977);
nand UO_400 (O_400,N_2974,N_2946);
nand UO_401 (O_401,N_2999,N_2953);
and UO_402 (O_402,N_2998,N_2940);
nand UO_403 (O_403,N_2988,N_2957);
nand UO_404 (O_404,N_2956,N_2975);
and UO_405 (O_405,N_2959,N_2947);
or UO_406 (O_406,N_2945,N_2942);
and UO_407 (O_407,N_2993,N_2998);
nand UO_408 (O_408,N_2981,N_2988);
and UO_409 (O_409,N_2943,N_2994);
nor UO_410 (O_410,N_2968,N_2973);
nor UO_411 (O_411,N_2971,N_2972);
or UO_412 (O_412,N_2971,N_2987);
nand UO_413 (O_413,N_2958,N_2942);
nor UO_414 (O_414,N_2942,N_2974);
nand UO_415 (O_415,N_2951,N_2966);
nand UO_416 (O_416,N_2961,N_2941);
nand UO_417 (O_417,N_2999,N_2977);
nand UO_418 (O_418,N_2964,N_2975);
and UO_419 (O_419,N_2961,N_2983);
and UO_420 (O_420,N_2940,N_2987);
nor UO_421 (O_421,N_2944,N_2942);
nand UO_422 (O_422,N_2953,N_2956);
nand UO_423 (O_423,N_2987,N_2997);
or UO_424 (O_424,N_2979,N_2987);
and UO_425 (O_425,N_2955,N_2998);
and UO_426 (O_426,N_2980,N_2963);
nand UO_427 (O_427,N_2965,N_2998);
nand UO_428 (O_428,N_2983,N_2959);
nor UO_429 (O_429,N_2968,N_2949);
nand UO_430 (O_430,N_2971,N_2952);
or UO_431 (O_431,N_2997,N_2948);
nor UO_432 (O_432,N_2959,N_2949);
nand UO_433 (O_433,N_2977,N_2961);
or UO_434 (O_434,N_2952,N_2956);
nor UO_435 (O_435,N_2945,N_2977);
and UO_436 (O_436,N_2974,N_2986);
nand UO_437 (O_437,N_2982,N_2992);
or UO_438 (O_438,N_2982,N_2945);
nand UO_439 (O_439,N_2998,N_2966);
nor UO_440 (O_440,N_2968,N_2940);
nor UO_441 (O_441,N_2947,N_2964);
or UO_442 (O_442,N_2991,N_2972);
and UO_443 (O_443,N_2996,N_2983);
or UO_444 (O_444,N_2941,N_2965);
or UO_445 (O_445,N_2983,N_2975);
and UO_446 (O_446,N_2962,N_2998);
nand UO_447 (O_447,N_2966,N_2941);
nor UO_448 (O_448,N_2942,N_2967);
nor UO_449 (O_449,N_2943,N_2966);
or UO_450 (O_450,N_2944,N_2969);
or UO_451 (O_451,N_2977,N_2976);
nand UO_452 (O_452,N_2994,N_2964);
nand UO_453 (O_453,N_2972,N_2957);
or UO_454 (O_454,N_2976,N_2965);
and UO_455 (O_455,N_2955,N_2972);
or UO_456 (O_456,N_2983,N_2973);
or UO_457 (O_457,N_2957,N_2959);
or UO_458 (O_458,N_2953,N_2991);
or UO_459 (O_459,N_2950,N_2992);
nor UO_460 (O_460,N_2966,N_2940);
and UO_461 (O_461,N_2972,N_2974);
or UO_462 (O_462,N_2953,N_2941);
or UO_463 (O_463,N_2969,N_2973);
nor UO_464 (O_464,N_2956,N_2943);
and UO_465 (O_465,N_2993,N_2954);
nand UO_466 (O_466,N_2990,N_2966);
nand UO_467 (O_467,N_2987,N_2975);
and UO_468 (O_468,N_2962,N_2997);
and UO_469 (O_469,N_2968,N_2966);
nand UO_470 (O_470,N_2961,N_2967);
nand UO_471 (O_471,N_2941,N_2944);
or UO_472 (O_472,N_2978,N_2989);
or UO_473 (O_473,N_2952,N_2943);
nand UO_474 (O_474,N_2967,N_2991);
xnor UO_475 (O_475,N_2978,N_2984);
nor UO_476 (O_476,N_2982,N_2962);
or UO_477 (O_477,N_2954,N_2978);
and UO_478 (O_478,N_2943,N_2954);
nand UO_479 (O_479,N_2981,N_2983);
nor UO_480 (O_480,N_2952,N_2946);
or UO_481 (O_481,N_2949,N_2985);
or UO_482 (O_482,N_2958,N_2966);
or UO_483 (O_483,N_2947,N_2990);
and UO_484 (O_484,N_2949,N_2948);
nand UO_485 (O_485,N_2973,N_2994);
and UO_486 (O_486,N_2954,N_2949);
nand UO_487 (O_487,N_2975,N_2995);
nor UO_488 (O_488,N_2993,N_2952);
and UO_489 (O_489,N_2985,N_2992);
or UO_490 (O_490,N_2985,N_2947);
and UO_491 (O_491,N_2957,N_2943);
or UO_492 (O_492,N_2971,N_2948);
nor UO_493 (O_493,N_2967,N_2988);
nand UO_494 (O_494,N_2946,N_2999);
and UO_495 (O_495,N_2957,N_2941);
nor UO_496 (O_496,N_2944,N_2991);
or UO_497 (O_497,N_2998,N_2953);
or UO_498 (O_498,N_2955,N_2975);
or UO_499 (O_499,N_2983,N_2966);
endmodule