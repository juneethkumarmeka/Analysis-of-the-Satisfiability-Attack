module basic_750_5000_1000_5_levels_1xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_459,In_353);
and U1 (N_1,In_150,In_337);
and U2 (N_2,In_69,In_267);
nand U3 (N_3,In_406,In_471);
nor U4 (N_4,In_190,In_559);
and U5 (N_5,In_143,In_141);
or U6 (N_6,In_264,In_438);
or U7 (N_7,In_107,In_218);
nand U8 (N_8,In_594,In_330);
and U9 (N_9,In_42,In_126);
or U10 (N_10,In_339,In_85);
nor U11 (N_11,In_213,In_159);
or U12 (N_12,In_268,In_611);
or U13 (N_13,In_333,In_451);
and U14 (N_14,In_442,In_184);
or U15 (N_15,In_281,In_696);
or U16 (N_16,In_313,In_655);
or U17 (N_17,In_157,In_191);
nor U18 (N_18,In_635,In_530);
or U19 (N_19,In_448,In_284);
nor U20 (N_20,In_325,In_675);
and U21 (N_21,In_163,In_223);
and U22 (N_22,In_60,In_362);
nor U23 (N_23,In_619,In_248);
or U24 (N_24,In_430,In_260);
nor U25 (N_25,In_685,In_639);
or U26 (N_26,In_713,In_81);
nand U27 (N_27,In_52,In_158);
nor U28 (N_28,In_324,In_634);
nand U29 (N_29,In_343,In_543);
nor U30 (N_30,In_691,In_389);
nand U31 (N_31,In_22,In_243);
nor U32 (N_32,In_562,In_228);
nand U33 (N_33,In_628,In_73);
and U34 (N_34,In_27,In_583);
nand U35 (N_35,In_689,In_54);
or U36 (N_36,In_261,In_289);
or U37 (N_37,In_1,In_422);
nor U38 (N_38,In_677,In_478);
nor U39 (N_39,In_116,In_624);
and U40 (N_40,In_443,In_332);
or U41 (N_41,In_597,In_433);
nor U42 (N_42,In_255,In_467);
nand U43 (N_43,In_545,In_263);
or U44 (N_44,In_650,In_674);
and U45 (N_45,In_210,In_600);
and U46 (N_46,In_70,In_652);
nor U47 (N_47,In_623,In_269);
nand U48 (N_48,In_607,In_79);
or U49 (N_49,In_534,In_32);
nor U50 (N_50,In_167,In_490);
and U51 (N_51,In_728,In_250);
or U52 (N_52,In_693,In_294);
or U53 (N_53,In_475,In_214);
nor U54 (N_54,In_512,In_51);
and U55 (N_55,In_36,In_444);
nor U56 (N_56,In_435,In_97);
and U57 (N_57,In_564,In_217);
nor U58 (N_58,In_449,In_346);
and U59 (N_59,In_702,In_578);
and U60 (N_60,In_252,In_119);
or U61 (N_61,In_549,In_50);
nand U62 (N_62,In_651,In_112);
nor U63 (N_63,In_441,In_349);
nand U64 (N_64,In_114,In_481);
or U65 (N_65,In_288,In_102);
and U66 (N_66,In_173,In_323);
nor U67 (N_67,In_698,In_482);
nor U68 (N_68,In_727,In_37);
or U69 (N_69,In_560,In_47);
nor U70 (N_70,In_335,In_11);
or U71 (N_71,In_357,In_747);
or U72 (N_72,In_569,In_476);
nor U73 (N_73,In_66,In_486);
and U74 (N_74,In_188,In_164);
and U75 (N_75,In_436,In_732);
nand U76 (N_76,In_285,In_371);
or U77 (N_77,In_359,In_579);
and U78 (N_78,In_596,In_493);
and U79 (N_79,In_402,In_720);
nor U80 (N_80,In_301,In_429);
and U81 (N_81,In_226,In_322);
or U82 (N_82,In_717,In_312);
nor U83 (N_83,In_340,In_584);
and U84 (N_84,In_369,In_55);
and U85 (N_85,In_453,In_5);
and U86 (N_86,In_718,In_273);
or U87 (N_87,In_484,In_193);
nor U88 (N_88,In_351,In_94);
or U89 (N_89,In_197,In_591);
or U90 (N_90,In_204,In_707);
or U91 (N_91,In_44,In_544);
nand U92 (N_92,In_287,In_598);
nand U93 (N_93,In_195,In_219);
nand U94 (N_94,In_663,In_404);
and U95 (N_95,In_588,In_24);
or U96 (N_96,In_474,In_140);
and U97 (N_97,In_242,In_649);
or U98 (N_98,In_413,In_676);
nand U99 (N_99,In_412,In_88);
nor U100 (N_100,In_233,In_692);
nor U101 (N_101,In_9,In_71);
or U102 (N_102,In_145,In_385);
or U103 (N_103,In_298,In_177);
or U104 (N_104,In_19,In_26);
nor U105 (N_105,In_20,In_122);
nand U106 (N_106,In_83,In_643);
and U107 (N_107,In_407,In_179);
nand U108 (N_108,In_33,In_237);
nor U109 (N_109,In_504,In_507);
or U110 (N_110,In_524,In_270);
nand U111 (N_111,In_182,In_419);
and U112 (N_112,In_721,In_581);
and U113 (N_113,In_347,In_314);
and U114 (N_114,In_169,In_35);
nor U115 (N_115,In_679,In_168);
xnor U116 (N_116,In_230,In_129);
and U117 (N_117,In_440,In_25);
nand U118 (N_118,In_132,In_708);
and U119 (N_119,In_489,In_151);
nor U120 (N_120,In_16,In_606);
nand U121 (N_121,In_421,In_98);
or U122 (N_122,In_405,In_201);
nor U123 (N_123,In_654,In_501);
nor U124 (N_124,In_90,In_236);
and U125 (N_125,In_662,In_196);
nand U126 (N_126,In_161,In_719);
or U127 (N_127,In_497,In_286);
nor U128 (N_128,In_743,In_77);
nor U129 (N_129,In_673,In_626);
and U130 (N_130,In_587,In_472);
nor U131 (N_131,In_423,In_556);
nand U132 (N_132,In_235,In_576);
and U133 (N_133,In_45,In_603);
and U134 (N_134,In_118,In_317);
and U135 (N_135,In_306,In_334);
and U136 (N_136,In_61,In_483);
nand U137 (N_137,In_160,In_388);
xnor U138 (N_138,In_245,In_608);
or U139 (N_139,In_181,In_239);
nand U140 (N_140,In_15,In_365);
or U141 (N_141,In_176,In_657);
nand U142 (N_142,In_625,In_455);
or U143 (N_143,In_152,In_106);
nor U144 (N_144,In_741,In_113);
or U145 (N_145,In_590,In_445);
nand U146 (N_146,In_612,In_394);
nor U147 (N_147,In_307,In_180);
nor U148 (N_148,In_465,In_640);
nor U149 (N_149,In_671,In_234);
nor U150 (N_150,In_200,In_171);
nand U151 (N_151,In_621,In_418);
nor U152 (N_152,In_420,In_454);
or U153 (N_153,In_220,In_296);
and U154 (N_154,In_730,In_710);
nor U155 (N_155,In_58,In_715);
and U156 (N_156,In_616,In_428);
nand U157 (N_157,In_28,In_316);
or U158 (N_158,In_291,In_589);
nor U159 (N_159,In_686,In_704);
and U160 (N_160,In_238,In_739);
nor U161 (N_161,In_211,In_279);
or U162 (N_162,In_117,In_745);
nor U163 (N_163,In_68,In_345);
or U164 (N_164,In_658,In_417);
nand U165 (N_165,In_552,In_225);
nor U166 (N_166,In_733,In_31);
nand U167 (N_167,In_508,In_30);
nor U168 (N_168,In_310,In_63);
nand U169 (N_169,In_580,In_84);
nor U170 (N_170,In_723,In_229);
or U171 (N_171,In_108,In_403);
and U172 (N_172,In_397,In_280);
and U173 (N_173,In_396,In_638);
nand U174 (N_174,In_198,In_485);
nand U175 (N_175,In_415,In_139);
or U176 (N_176,In_183,In_372);
or U177 (N_177,In_586,In_749);
nor U178 (N_178,In_10,In_684);
or U179 (N_179,In_672,In_192);
nor U180 (N_180,In_149,In_427);
xor U181 (N_181,In_328,In_683);
nor U182 (N_182,In_480,In_105);
nand U183 (N_183,In_463,In_391);
nand U184 (N_184,In_87,In_91);
or U185 (N_185,In_618,In_709);
and U186 (N_186,In_514,In_277);
and U187 (N_187,In_155,In_297);
nor U188 (N_188,In_207,In_437);
and U189 (N_189,In_75,In_82);
and U190 (N_190,In_3,In_110);
nor U191 (N_191,In_633,In_678);
or U192 (N_192,In_144,In_642);
nand U193 (N_193,In_746,In_615);
and U194 (N_194,In_411,In_452);
xnor U195 (N_195,In_240,In_115);
or U196 (N_196,In_130,In_386);
and U197 (N_197,In_203,In_740);
or U198 (N_198,In_215,In_535);
or U199 (N_199,In_670,In_521);
or U200 (N_200,In_522,In_729);
or U201 (N_201,In_80,In_199);
or U202 (N_202,In_266,In_665);
nor U203 (N_203,In_393,In_206);
nand U204 (N_204,In_599,In_309);
or U205 (N_205,In_148,In_450);
xor U206 (N_206,In_488,In_613);
and U207 (N_207,In_464,In_282);
nand U208 (N_208,In_505,In_376);
and U209 (N_209,In_373,In_124);
and U210 (N_210,In_342,In_392);
nand U211 (N_211,In_636,In_614);
nor U212 (N_212,In_256,In_278);
and U213 (N_213,In_632,In_523);
and U214 (N_214,In_516,In_142);
and U215 (N_215,In_567,In_382);
nor U216 (N_216,In_64,In_517);
and U217 (N_217,In_468,In_528);
nand U218 (N_218,In_541,In_185);
or U219 (N_219,In_553,In_377);
nand U220 (N_220,In_360,In_222);
nor U221 (N_221,In_664,In_518);
nand U222 (N_222,In_401,In_62);
or U223 (N_223,In_131,In_4);
or U224 (N_224,In_384,In_470);
or U225 (N_225,In_326,In_414);
or U226 (N_226,In_716,In_364);
or U227 (N_227,In_631,In_509);
or U228 (N_228,In_526,In_249);
nand U229 (N_229,In_460,In_358);
and U230 (N_230,In_456,In_272);
or U231 (N_231,In_540,In_712);
or U232 (N_232,In_154,In_156);
nand U233 (N_233,In_604,In_416);
or U234 (N_234,In_93,In_17);
nor U235 (N_235,In_295,In_629);
nor U236 (N_236,In_500,In_172);
and U237 (N_237,In_561,In_566);
nand U238 (N_238,In_38,In_506);
and U239 (N_239,In_439,In_147);
nor U240 (N_240,In_532,In_166);
and U241 (N_241,In_536,In_627);
nand U242 (N_242,In_92,In_12);
or U243 (N_243,In_216,In_734);
and U244 (N_244,In_300,In_645);
nand U245 (N_245,In_378,In_356);
and U246 (N_246,In_99,In_711);
nor U247 (N_247,In_14,In_424);
nor U248 (N_248,In_315,In_434);
or U249 (N_249,In_660,In_361);
nand U250 (N_250,In_533,In_100);
and U251 (N_251,In_375,In_65);
nand U252 (N_252,In_542,In_537);
nor U253 (N_253,In_341,In_290);
nor U254 (N_254,In_321,In_368);
nor U255 (N_255,In_104,In_18);
nor U256 (N_256,In_189,In_299);
or U257 (N_257,In_563,In_381);
nor U258 (N_258,In_23,In_682);
nand U259 (N_259,In_178,In_725);
or U260 (N_260,In_276,In_0);
nor U261 (N_261,In_601,In_477);
nor U262 (N_262,In_558,In_555);
nand U263 (N_263,In_426,In_29);
nor U264 (N_264,In_74,In_123);
nand U265 (N_265,In_554,In_661);
or U266 (N_266,In_374,In_136);
and U267 (N_267,In_492,In_609);
and U268 (N_268,In_303,In_7);
nor U269 (N_269,In_259,In_53);
and U270 (N_270,In_432,In_46);
nor U271 (N_271,In_165,In_302);
and U272 (N_272,In_305,In_251);
nor U273 (N_273,In_247,In_694);
nor U274 (N_274,In_146,In_699);
and U275 (N_275,In_78,In_703);
nand U276 (N_276,In_348,In_510);
nor U277 (N_277,In_293,In_101);
nand U278 (N_278,In_700,In_695);
nand U279 (N_279,In_308,In_408);
and U280 (N_280,In_637,In_331);
or U281 (N_281,In_574,In_446);
nand U282 (N_282,In_503,In_205);
nor U283 (N_283,In_6,In_669);
and U284 (N_284,In_76,In_380);
and U285 (N_285,In_539,In_546);
or U286 (N_286,In_447,In_551);
and U287 (N_287,In_121,In_494);
nand U288 (N_288,In_726,In_227);
nand U289 (N_289,In_257,In_570);
and U290 (N_290,In_244,In_519);
nor U291 (N_291,In_466,In_224);
nor U292 (N_292,In_212,In_547);
and U293 (N_293,In_647,In_43);
nor U294 (N_294,In_274,In_431);
or U295 (N_295,In_258,In_398);
nor U296 (N_296,In_722,In_593);
nor U297 (N_297,In_620,In_292);
and U298 (N_298,In_137,In_262);
nand U299 (N_299,In_511,In_125);
or U300 (N_300,In_363,In_605);
and U301 (N_301,In_736,In_458);
nor U302 (N_302,In_602,In_688);
nor U303 (N_303,In_573,In_59);
nor U304 (N_304,In_496,In_352);
nor U305 (N_305,In_469,In_656);
nand U306 (N_306,In_648,In_86);
nor U307 (N_307,In_221,In_592);
nor U308 (N_308,In_706,In_187);
and U309 (N_309,In_209,In_350);
or U310 (N_310,In_21,In_367);
nor U311 (N_311,In_557,In_383);
or U312 (N_312,In_338,In_742);
or U313 (N_313,In_246,In_194);
nor U314 (N_314,In_525,In_538);
nor U315 (N_315,In_491,In_120);
nor U316 (N_316,In_646,In_253);
nand U317 (N_317,In_13,In_399);
nor U318 (N_318,In_320,In_103);
nor U319 (N_319,In_495,In_271);
or U320 (N_320,In_659,In_701);
and U321 (N_321,In_153,In_8);
nor U322 (N_322,In_666,In_697);
nand U323 (N_323,In_134,In_41);
nor U324 (N_324,In_111,In_135);
nor U325 (N_325,In_366,In_327);
nor U326 (N_326,In_109,In_232);
or U327 (N_327,In_138,In_653);
nor U328 (N_328,In_175,In_329);
or U329 (N_329,In_577,In_610);
or U330 (N_330,In_127,In_748);
nand U331 (N_331,In_585,In_668);
and U332 (N_332,In_714,In_479);
nand U333 (N_333,In_487,In_410);
nor U334 (N_334,In_738,In_575);
or U335 (N_335,In_318,In_265);
nor U336 (N_336,In_617,In_622);
or U337 (N_337,In_641,In_40);
and U338 (N_338,In_170,In_49);
or U339 (N_339,In_667,In_344);
nor U340 (N_340,In_128,In_680);
or U341 (N_341,In_531,In_34);
and U342 (N_342,In_457,In_56);
nor U343 (N_343,In_336,In_400);
nand U344 (N_344,In_548,In_744);
nor U345 (N_345,In_387,In_644);
nor U346 (N_346,In_690,In_513);
nor U347 (N_347,In_731,In_395);
and U348 (N_348,In_498,In_425);
or U349 (N_349,In_254,In_582);
nor U350 (N_350,In_568,In_595);
nor U351 (N_351,In_96,In_737);
and U352 (N_352,In_571,In_572);
and U353 (N_353,In_550,In_202);
nor U354 (N_354,In_89,In_354);
nand U355 (N_355,In_527,In_390);
and U356 (N_356,In_319,In_275);
or U357 (N_357,In_208,In_355);
or U358 (N_358,In_630,In_473);
or U359 (N_359,In_461,In_39);
and U360 (N_360,In_499,In_72);
nand U361 (N_361,In_735,In_57);
or U362 (N_362,In_133,In_311);
or U363 (N_363,In_565,In_515);
nor U364 (N_364,In_520,In_174);
or U365 (N_365,In_370,In_95);
nand U366 (N_366,In_462,In_687);
nand U367 (N_367,In_283,In_502);
and U368 (N_368,In_2,In_48);
nor U369 (N_369,In_724,In_186);
nor U370 (N_370,In_379,In_241);
or U371 (N_371,In_67,In_529);
and U372 (N_372,In_409,In_304);
or U373 (N_373,In_162,In_705);
nor U374 (N_374,In_231,In_681);
nor U375 (N_375,In_271,In_410);
nand U376 (N_376,In_173,In_199);
nor U377 (N_377,In_190,In_206);
nand U378 (N_378,In_620,In_509);
nor U379 (N_379,In_418,In_548);
nand U380 (N_380,In_475,In_311);
nor U381 (N_381,In_717,In_299);
nand U382 (N_382,In_202,In_365);
or U383 (N_383,In_726,In_409);
nand U384 (N_384,In_98,In_469);
nand U385 (N_385,In_429,In_586);
or U386 (N_386,In_356,In_507);
nand U387 (N_387,In_524,In_680);
or U388 (N_388,In_112,In_321);
or U389 (N_389,In_261,In_190);
or U390 (N_390,In_56,In_221);
nand U391 (N_391,In_497,In_532);
nand U392 (N_392,In_77,In_665);
or U393 (N_393,In_7,In_338);
or U394 (N_394,In_590,In_584);
or U395 (N_395,In_51,In_516);
nor U396 (N_396,In_340,In_278);
or U397 (N_397,In_571,In_51);
and U398 (N_398,In_85,In_628);
nand U399 (N_399,In_203,In_133);
and U400 (N_400,In_157,In_379);
nor U401 (N_401,In_379,In_522);
nand U402 (N_402,In_110,In_630);
nand U403 (N_403,In_557,In_25);
nor U404 (N_404,In_439,In_598);
or U405 (N_405,In_616,In_460);
nand U406 (N_406,In_130,In_307);
xnor U407 (N_407,In_375,In_243);
nand U408 (N_408,In_0,In_532);
or U409 (N_409,In_209,In_378);
nand U410 (N_410,In_512,In_523);
or U411 (N_411,In_199,In_153);
nand U412 (N_412,In_42,In_409);
or U413 (N_413,In_462,In_258);
and U414 (N_414,In_125,In_218);
nor U415 (N_415,In_367,In_717);
nor U416 (N_416,In_48,In_212);
and U417 (N_417,In_24,In_131);
nand U418 (N_418,In_550,In_430);
or U419 (N_419,In_222,In_115);
nand U420 (N_420,In_430,In_434);
or U421 (N_421,In_631,In_571);
and U422 (N_422,In_415,In_379);
and U423 (N_423,In_275,In_504);
or U424 (N_424,In_321,In_247);
or U425 (N_425,In_377,In_441);
or U426 (N_426,In_205,In_125);
or U427 (N_427,In_469,In_570);
or U428 (N_428,In_651,In_94);
or U429 (N_429,In_473,In_348);
or U430 (N_430,In_605,In_622);
nand U431 (N_431,In_79,In_193);
and U432 (N_432,In_13,In_46);
nand U433 (N_433,In_425,In_225);
nor U434 (N_434,In_384,In_497);
nor U435 (N_435,In_196,In_246);
or U436 (N_436,In_374,In_596);
nor U437 (N_437,In_479,In_274);
nand U438 (N_438,In_276,In_495);
nand U439 (N_439,In_589,In_522);
nand U440 (N_440,In_709,In_120);
nor U441 (N_441,In_225,In_11);
or U442 (N_442,In_147,In_155);
or U443 (N_443,In_147,In_429);
or U444 (N_444,In_294,In_85);
and U445 (N_445,In_143,In_412);
and U446 (N_446,In_587,In_160);
and U447 (N_447,In_685,In_681);
and U448 (N_448,In_664,In_287);
and U449 (N_449,In_60,In_409);
or U450 (N_450,In_334,In_251);
and U451 (N_451,In_192,In_60);
and U452 (N_452,In_563,In_232);
nor U453 (N_453,In_53,In_347);
or U454 (N_454,In_533,In_745);
nand U455 (N_455,In_260,In_4);
or U456 (N_456,In_257,In_736);
or U457 (N_457,In_513,In_714);
xnor U458 (N_458,In_366,In_496);
nand U459 (N_459,In_526,In_144);
xor U460 (N_460,In_307,In_275);
nand U461 (N_461,In_382,In_37);
nor U462 (N_462,In_54,In_123);
or U463 (N_463,In_699,In_729);
and U464 (N_464,In_65,In_663);
or U465 (N_465,In_271,In_524);
and U466 (N_466,In_294,In_729);
nand U467 (N_467,In_420,In_457);
nor U468 (N_468,In_58,In_92);
nor U469 (N_469,In_273,In_382);
or U470 (N_470,In_148,In_688);
nand U471 (N_471,In_650,In_659);
nor U472 (N_472,In_150,In_671);
nor U473 (N_473,In_270,In_443);
or U474 (N_474,In_40,In_461);
nor U475 (N_475,In_347,In_693);
and U476 (N_476,In_243,In_136);
nand U477 (N_477,In_287,In_201);
or U478 (N_478,In_611,In_640);
and U479 (N_479,In_527,In_428);
and U480 (N_480,In_622,In_524);
nor U481 (N_481,In_502,In_629);
and U482 (N_482,In_194,In_243);
or U483 (N_483,In_270,In_361);
and U484 (N_484,In_35,In_669);
and U485 (N_485,In_453,In_600);
or U486 (N_486,In_306,In_43);
or U487 (N_487,In_331,In_622);
nand U488 (N_488,In_165,In_160);
or U489 (N_489,In_684,In_433);
or U490 (N_490,In_715,In_538);
and U491 (N_491,In_429,In_584);
nor U492 (N_492,In_79,In_309);
nand U493 (N_493,In_302,In_138);
or U494 (N_494,In_585,In_611);
nor U495 (N_495,In_383,In_734);
nor U496 (N_496,In_566,In_75);
or U497 (N_497,In_508,In_23);
nand U498 (N_498,In_189,In_240);
and U499 (N_499,In_683,In_342);
or U500 (N_500,In_684,In_466);
nor U501 (N_501,In_295,In_235);
and U502 (N_502,In_515,In_288);
nor U503 (N_503,In_577,In_92);
and U504 (N_504,In_67,In_730);
nand U505 (N_505,In_310,In_550);
or U506 (N_506,In_714,In_717);
nor U507 (N_507,In_715,In_431);
or U508 (N_508,In_518,In_586);
and U509 (N_509,In_680,In_513);
nand U510 (N_510,In_288,In_155);
nor U511 (N_511,In_591,In_171);
nand U512 (N_512,In_49,In_161);
nor U513 (N_513,In_41,In_606);
or U514 (N_514,In_498,In_108);
or U515 (N_515,In_110,In_363);
or U516 (N_516,In_91,In_288);
and U517 (N_517,In_629,In_424);
nand U518 (N_518,In_292,In_655);
or U519 (N_519,In_556,In_267);
nand U520 (N_520,In_505,In_437);
nor U521 (N_521,In_588,In_441);
or U522 (N_522,In_380,In_325);
nor U523 (N_523,In_559,In_539);
nor U524 (N_524,In_195,In_606);
and U525 (N_525,In_278,In_129);
and U526 (N_526,In_55,In_277);
and U527 (N_527,In_708,In_705);
or U528 (N_528,In_428,In_133);
nand U529 (N_529,In_593,In_423);
nand U530 (N_530,In_110,In_230);
nand U531 (N_531,In_102,In_257);
or U532 (N_532,In_304,In_111);
nor U533 (N_533,In_498,In_214);
nand U534 (N_534,In_109,In_510);
nor U535 (N_535,In_38,In_281);
and U536 (N_536,In_464,In_264);
nand U537 (N_537,In_278,In_12);
nand U538 (N_538,In_208,In_5);
nor U539 (N_539,In_280,In_650);
and U540 (N_540,In_673,In_141);
or U541 (N_541,In_570,In_739);
nor U542 (N_542,In_257,In_465);
or U543 (N_543,In_559,In_653);
or U544 (N_544,In_441,In_683);
and U545 (N_545,In_585,In_16);
nand U546 (N_546,In_173,In_381);
and U547 (N_547,In_285,In_739);
or U548 (N_548,In_566,In_568);
and U549 (N_549,In_56,In_124);
nor U550 (N_550,In_709,In_574);
nor U551 (N_551,In_543,In_40);
nor U552 (N_552,In_73,In_20);
nand U553 (N_553,In_331,In_311);
nor U554 (N_554,In_460,In_510);
nand U555 (N_555,In_473,In_432);
nor U556 (N_556,In_97,In_35);
nor U557 (N_557,In_674,In_61);
nor U558 (N_558,In_512,In_519);
xor U559 (N_559,In_333,In_41);
nand U560 (N_560,In_432,In_3);
or U561 (N_561,In_709,In_539);
or U562 (N_562,In_169,In_424);
or U563 (N_563,In_201,In_369);
and U564 (N_564,In_94,In_178);
or U565 (N_565,In_289,In_499);
nand U566 (N_566,In_354,In_448);
and U567 (N_567,In_375,In_251);
or U568 (N_568,In_375,In_577);
nand U569 (N_569,In_702,In_589);
or U570 (N_570,In_357,In_416);
xnor U571 (N_571,In_464,In_447);
nor U572 (N_572,In_179,In_353);
nor U573 (N_573,In_363,In_440);
nand U574 (N_574,In_720,In_212);
nor U575 (N_575,In_256,In_627);
nand U576 (N_576,In_484,In_269);
nand U577 (N_577,In_60,In_373);
nor U578 (N_578,In_671,In_407);
or U579 (N_579,In_562,In_149);
nand U580 (N_580,In_653,In_71);
or U581 (N_581,In_59,In_566);
nand U582 (N_582,In_55,In_605);
nand U583 (N_583,In_238,In_40);
or U584 (N_584,In_540,In_189);
nor U585 (N_585,In_329,In_378);
nand U586 (N_586,In_643,In_450);
nor U587 (N_587,In_316,In_541);
nand U588 (N_588,In_633,In_515);
nand U589 (N_589,In_46,In_366);
nor U590 (N_590,In_268,In_67);
nand U591 (N_591,In_137,In_307);
nor U592 (N_592,In_425,In_379);
nor U593 (N_593,In_597,In_465);
nand U594 (N_594,In_678,In_445);
or U595 (N_595,In_27,In_416);
and U596 (N_596,In_262,In_239);
and U597 (N_597,In_277,In_271);
and U598 (N_598,In_301,In_189);
or U599 (N_599,In_91,In_682);
nand U600 (N_600,In_687,In_302);
nor U601 (N_601,In_63,In_255);
or U602 (N_602,In_37,In_678);
nand U603 (N_603,In_192,In_53);
and U604 (N_604,In_72,In_96);
and U605 (N_605,In_609,In_529);
nand U606 (N_606,In_497,In_113);
nor U607 (N_607,In_399,In_60);
or U608 (N_608,In_351,In_618);
nand U609 (N_609,In_657,In_66);
nor U610 (N_610,In_519,In_207);
and U611 (N_611,In_736,In_107);
and U612 (N_612,In_51,In_63);
nor U613 (N_613,In_374,In_129);
or U614 (N_614,In_502,In_660);
nor U615 (N_615,In_611,In_59);
nand U616 (N_616,In_605,In_325);
or U617 (N_617,In_36,In_547);
or U618 (N_618,In_271,In_191);
or U619 (N_619,In_322,In_213);
and U620 (N_620,In_624,In_427);
nor U621 (N_621,In_253,In_644);
or U622 (N_622,In_263,In_504);
nand U623 (N_623,In_57,In_668);
or U624 (N_624,In_39,In_127);
and U625 (N_625,In_499,In_316);
and U626 (N_626,In_540,In_38);
or U627 (N_627,In_280,In_71);
and U628 (N_628,In_64,In_458);
and U629 (N_629,In_488,In_151);
or U630 (N_630,In_99,In_524);
nand U631 (N_631,In_745,In_262);
nand U632 (N_632,In_310,In_746);
nor U633 (N_633,In_246,In_10);
nand U634 (N_634,In_502,In_688);
or U635 (N_635,In_580,In_15);
nand U636 (N_636,In_659,In_510);
nand U637 (N_637,In_200,In_732);
nand U638 (N_638,In_606,In_654);
nand U639 (N_639,In_112,In_94);
nor U640 (N_640,In_341,In_567);
nand U641 (N_641,In_450,In_448);
nand U642 (N_642,In_518,In_169);
nand U643 (N_643,In_464,In_119);
nand U644 (N_644,In_274,In_67);
nor U645 (N_645,In_416,In_748);
and U646 (N_646,In_17,In_44);
and U647 (N_647,In_479,In_71);
nand U648 (N_648,In_698,In_101);
nor U649 (N_649,In_249,In_230);
nand U650 (N_650,In_719,In_747);
or U651 (N_651,In_271,In_654);
nand U652 (N_652,In_747,In_741);
nor U653 (N_653,In_185,In_408);
and U654 (N_654,In_81,In_306);
nand U655 (N_655,In_588,In_502);
nor U656 (N_656,In_366,In_514);
nand U657 (N_657,In_543,In_723);
nand U658 (N_658,In_626,In_583);
nand U659 (N_659,In_608,In_47);
or U660 (N_660,In_531,In_677);
or U661 (N_661,In_578,In_382);
and U662 (N_662,In_433,In_197);
nor U663 (N_663,In_678,In_68);
and U664 (N_664,In_446,In_406);
or U665 (N_665,In_177,In_369);
nor U666 (N_666,In_678,In_453);
nor U667 (N_667,In_506,In_543);
and U668 (N_668,In_154,In_273);
or U669 (N_669,In_474,In_87);
and U670 (N_670,In_155,In_274);
nand U671 (N_671,In_96,In_714);
nand U672 (N_672,In_37,In_295);
nand U673 (N_673,In_316,In_83);
nor U674 (N_674,In_75,In_359);
and U675 (N_675,In_137,In_654);
nand U676 (N_676,In_78,In_398);
nand U677 (N_677,In_320,In_434);
nor U678 (N_678,In_30,In_119);
nand U679 (N_679,In_77,In_99);
xor U680 (N_680,In_735,In_487);
and U681 (N_681,In_119,In_183);
or U682 (N_682,In_545,In_35);
nor U683 (N_683,In_380,In_280);
nand U684 (N_684,In_323,In_391);
nand U685 (N_685,In_718,In_18);
or U686 (N_686,In_223,In_387);
and U687 (N_687,In_393,In_439);
nor U688 (N_688,In_189,In_17);
and U689 (N_689,In_377,In_296);
nand U690 (N_690,In_374,In_280);
nor U691 (N_691,In_465,In_272);
nand U692 (N_692,In_301,In_613);
and U693 (N_693,In_255,In_102);
nand U694 (N_694,In_677,In_301);
nand U695 (N_695,In_48,In_277);
and U696 (N_696,In_426,In_154);
nor U697 (N_697,In_107,In_515);
nor U698 (N_698,In_3,In_276);
nand U699 (N_699,In_33,In_54);
nor U700 (N_700,In_749,In_206);
nor U701 (N_701,In_271,In_103);
nor U702 (N_702,In_560,In_156);
nand U703 (N_703,In_203,In_426);
nor U704 (N_704,In_219,In_201);
and U705 (N_705,In_302,In_516);
or U706 (N_706,In_484,In_343);
nand U707 (N_707,In_627,In_112);
nor U708 (N_708,In_239,In_681);
nor U709 (N_709,In_714,In_466);
and U710 (N_710,In_21,In_130);
nand U711 (N_711,In_673,In_147);
and U712 (N_712,In_72,In_55);
nor U713 (N_713,In_433,In_159);
nand U714 (N_714,In_232,In_733);
or U715 (N_715,In_307,In_685);
or U716 (N_716,In_146,In_227);
nor U717 (N_717,In_381,In_74);
or U718 (N_718,In_162,In_421);
nor U719 (N_719,In_459,In_486);
nand U720 (N_720,In_357,In_600);
nor U721 (N_721,In_626,In_142);
or U722 (N_722,In_66,In_560);
nand U723 (N_723,In_98,In_407);
and U724 (N_724,In_128,In_165);
and U725 (N_725,In_749,In_418);
nor U726 (N_726,In_240,In_328);
and U727 (N_727,In_96,In_419);
and U728 (N_728,In_270,In_414);
or U729 (N_729,In_238,In_309);
or U730 (N_730,In_271,In_60);
or U731 (N_731,In_312,In_490);
nor U732 (N_732,In_333,In_579);
and U733 (N_733,In_604,In_122);
and U734 (N_734,In_27,In_132);
and U735 (N_735,In_269,In_605);
or U736 (N_736,In_480,In_27);
or U737 (N_737,In_100,In_40);
nor U738 (N_738,In_488,In_348);
nor U739 (N_739,In_18,In_44);
nand U740 (N_740,In_667,In_218);
nor U741 (N_741,In_0,In_292);
or U742 (N_742,In_105,In_637);
nand U743 (N_743,In_132,In_582);
or U744 (N_744,In_428,In_243);
nor U745 (N_745,In_677,In_378);
nor U746 (N_746,In_254,In_612);
and U747 (N_747,In_563,In_379);
nand U748 (N_748,In_582,In_569);
or U749 (N_749,In_566,In_359);
or U750 (N_750,In_442,In_498);
and U751 (N_751,In_399,In_259);
nor U752 (N_752,In_292,In_622);
nor U753 (N_753,In_235,In_525);
or U754 (N_754,In_354,In_680);
nand U755 (N_755,In_511,In_324);
nor U756 (N_756,In_147,In_519);
and U757 (N_757,In_321,In_84);
and U758 (N_758,In_362,In_326);
and U759 (N_759,In_155,In_594);
nand U760 (N_760,In_131,In_706);
nor U761 (N_761,In_661,In_377);
or U762 (N_762,In_138,In_316);
and U763 (N_763,In_444,In_527);
nand U764 (N_764,In_735,In_610);
and U765 (N_765,In_662,In_426);
nor U766 (N_766,In_20,In_154);
nor U767 (N_767,In_606,In_512);
nor U768 (N_768,In_507,In_263);
nand U769 (N_769,In_392,In_45);
nor U770 (N_770,In_465,In_231);
or U771 (N_771,In_296,In_686);
nor U772 (N_772,In_522,In_658);
or U773 (N_773,In_104,In_368);
or U774 (N_774,In_379,In_385);
nor U775 (N_775,In_535,In_394);
or U776 (N_776,In_85,In_651);
and U777 (N_777,In_226,In_25);
nor U778 (N_778,In_692,In_330);
xor U779 (N_779,In_282,In_664);
nand U780 (N_780,In_433,In_122);
and U781 (N_781,In_226,In_671);
and U782 (N_782,In_687,In_89);
or U783 (N_783,In_502,In_108);
nand U784 (N_784,In_654,In_656);
or U785 (N_785,In_153,In_70);
nor U786 (N_786,In_736,In_294);
nor U787 (N_787,In_540,In_490);
nand U788 (N_788,In_492,In_524);
nor U789 (N_789,In_599,In_590);
or U790 (N_790,In_28,In_362);
nor U791 (N_791,In_223,In_173);
xnor U792 (N_792,In_286,In_548);
nor U793 (N_793,In_92,In_594);
nor U794 (N_794,In_573,In_63);
or U795 (N_795,In_96,In_666);
nor U796 (N_796,In_421,In_489);
nand U797 (N_797,In_25,In_301);
nor U798 (N_798,In_706,In_663);
and U799 (N_799,In_203,In_70);
and U800 (N_800,In_522,In_394);
nor U801 (N_801,In_9,In_686);
and U802 (N_802,In_728,In_541);
nor U803 (N_803,In_468,In_44);
and U804 (N_804,In_545,In_443);
nor U805 (N_805,In_262,In_450);
nor U806 (N_806,In_80,In_166);
nor U807 (N_807,In_451,In_362);
or U808 (N_808,In_525,In_313);
nor U809 (N_809,In_6,In_670);
or U810 (N_810,In_29,In_220);
or U811 (N_811,In_303,In_184);
and U812 (N_812,In_438,In_283);
or U813 (N_813,In_580,In_496);
nand U814 (N_814,In_258,In_287);
nor U815 (N_815,In_694,In_180);
nor U816 (N_816,In_734,In_153);
nor U817 (N_817,In_200,In_228);
nor U818 (N_818,In_196,In_695);
or U819 (N_819,In_479,In_403);
or U820 (N_820,In_697,In_354);
or U821 (N_821,In_657,In_682);
nand U822 (N_822,In_300,In_537);
nand U823 (N_823,In_400,In_690);
or U824 (N_824,In_431,In_286);
nor U825 (N_825,In_46,In_365);
nand U826 (N_826,In_9,In_17);
and U827 (N_827,In_670,In_664);
and U828 (N_828,In_379,In_470);
or U829 (N_829,In_628,In_707);
or U830 (N_830,In_650,In_191);
or U831 (N_831,In_524,In_490);
nor U832 (N_832,In_415,In_700);
nor U833 (N_833,In_747,In_376);
nor U834 (N_834,In_110,In_241);
and U835 (N_835,In_33,In_297);
nor U836 (N_836,In_176,In_70);
or U837 (N_837,In_713,In_296);
or U838 (N_838,In_628,In_625);
and U839 (N_839,In_523,In_743);
nor U840 (N_840,In_663,In_700);
nor U841 (N_841,In_337,In_379);
and U842 (N_842,In_398,In_193);
or U843 (N_843,In_515,In_563);
nor U844 (N_844,In_482,In_631);
or U845 (N_845,In_135,In_203);
or U846 (N_846,In_483,In_504);
nor U847 (N_847,In_704,In_578);
nand U848 (N_848,In_315,In_242);
nand U849 (N_849,In_277,In_675);
or U850 (N_850,In_692,In_596);
and U851 (N_851,In_126,In_709);
nor U852 (N_852,In_241,In_733);
or U853 (N_853,In_385,In_527);
nand U854 (N_854,In_164,In_33);
or U855 (N_855,In_386,In_54);
or U856 (N_856,In_6,In_279);
and U857 (N_857,In_157,In_210);
or U858 (N_858,In_636,In_391);
nand U859 (N_859,In_107,In_723);
or U860 (N_860,In_664,In_248);
nor U861 (N_861,In_345,In_577);
xnor U862 (N_862,In_120,In_113);
or U863 (N_863,In_286,In_295);
nand U864 (N_864,In_460,In_169);
nand U865 (N_865,In_55,In_398);
or U866 (N_866,In_587,In_131);
or U867 (N_867,In_284,In_556);
nand U868 (N_868,In_18,In_713);
nor U869 (N_869,In_74,In_473);
and U870 (N_870,In_708,In_115);
or U871 (N_871,In_216,In_112);
nand U872 (N_872,In_430,In_19);
nor U873 (N_873,In_243,In_463);
nand U874 (N_874,In_157,In_594);
nor U875 (N_875,In_266,In_718);
nand U876 (N_876,In_66,In_719);
nand U877 (N_877,In_500,In_77);
nor U878 (N_878,In_359,In_397);
nor U879 (N_879,In_179,In_56);
nand U880 (N_880,In_172,In_105);
and U881 (N_881,In_555,In_464);
or U882 (N_882,In_173,In_26);
nor U883 (N_883,In_58,In_582);
or U884 (N_884,In_114,In_595);
and U885 (N_885,In_288,In_632);
or U886 (N_886,In_491,In_253);
and U887 (N_887,In_536,In_216);
nor U888 (N_888,In_285,In_549);
or U889 (N_889,In_37,In_340);
nor U890 (N_890,In_344,In_307);
or U891 (N_891,In_373,In_391);
or U892 (N_892,In_276,In_325);
nor U893 (N_893,In_181,In_377);
or U894 (N_894,In_548,In_111);
or U895 (N_895,In_254,In_482);
nor U896 (N_896,In_105,In_129);
nand U897 (N_897,In_537,In_650);
or U898 (N_898,In_491,In_683);
or U899 (N_899,In_494,In_419);
nor U900 (N_900,In_353,In_650);
and U901 (N_901,In_632,In_560);
or U902 (N_902,In_351,In_229);
nand U903 (N_903,In_388,In_595);
or U904 (N_904,In_633,In_599);
and U905 (N_905,In_306,In_473);
or U906 (N_906,In_702,In_63);
nand U907 (N_907,In_236,In_290);
nor U908 (N_908,In_470,In_308);
nand U909 (N_909,In_579,In_563);
or U910 (N_910,In_627,In_531);
and U911 (N_911,In_416,In_234);
nand U912 (N_912,In_608,In_708);
nor U913 (N_913,In_169,In_39);
and U914 (N_914,In_664,In_607);
and U915 (N_915,In_6,In_126);
or U916 (N_916,In_474,In_466);
or U917 (N_917,In_89,In_680);
nand U918 (N_918,In_364,In_92);
nor U919 (N_919,In_85,In_525);
nand U920 (N_920,In_735,In_551);
nor U921 (N_921,In_604,In_167);
and U922 (N_922,In_97,In_260);
and U923 (N_923,In_220,In_557);
nand U924 (N_924,In_580,In_238);
or U925 (N_925,In_124,In_352);
nand U926 (N_926,In_34,In_18);
nor U927 (N_927,In_536,In_156);
nand U928 (N_928,In_672,In_600);
nand U929 (N_929,In_28,In_45);
xor U930 (N_930,In_586,In_285);
and U931 (N_931,In_746,In_112);
and U932 (N_932,In_110,In_488);
nor U933 (N_933,In_386,In_421);
or U934 (N_934,In_524,In_151);
nand U935 (N_935,In_601,In_541);
or U936 (N_936,In_352,In_335);
or U937 (N_937,In_159,In_77);
or U938 (N_938,In_25,In_171);
and U939 (N_939,In_33,In_171);
or U940 (N_940,In_322,In_460);
or U941 (N_941,In_331,In_230);
or U942 (N_942,In_564,In_344);
and U943 (N_943,In_351,In_257);
nor U944 (N_944,In_565,In_696);
nor U945 (N_945,In_613,In_726);
nor U946 (N_946,In_93,In_692);
and U947 (N_947,In_335,In_482);
nand U948 (N_948,In_23,In_634);
and U949 (N_949,In_438,In_732);
nand U950 (N_950,In_224,In_222);
or U951 (N_951,In_716,In_115);
nand U952 (N_952,In_554,In_66);
nor U953 (N_953,In_125,In_204);
nand U954 (N_954,In_128,In_557);
and U955 (N_955,In_617,In_695);
xnor U956 (N_956,In_66,In_145);
and U957 (N_957,In_341,In_456);
and U958 (N_958,In_667,In_440);
nor U959 (N_959,In_650,In_113);
or U960 (N_960,In_232,In_35);
and U961 (N_961,In_500,In_515);
nand U962 (N_962,In_558,In_544);
and U963 (N_963,In_18,In_379);
nor U964 (N_964,In_586,In_461);
nor U965 (N_965,In_80,In_468);
and U966 (N_966,In_2,In_50);
nand U967 (N_967,In_73,In_37);
nor U968 (N_968,In_444,In_616);
and U969 (N_969,In_408,In_34);
nor U970 (N_970,In_514,In_4);
nand U971 (N_971,In_445,In_21);
or U972 (N_972,In_72,In_34);
or U973 (N_973,In_316,In_14);
nor U974 (N_974,In_599,In_686);
nand U975 (N_975,In_129,In_456);
nand U976 (N_976,In_70,In_433);
nand U977 (N_977,In_642,In_258);
or U978 (N_978,In_544,In_74);
or U979 (N_979,In_46,In_507);
nand U980 (N_980,In_58,In_142);
or U981 (N_981,In_76,In_132);
nor U982 (N_982,In_441,In_749);
nor U983 (N_983,In_633,In_705);
nand U984 (N_984,In_301,In_331);
nand U985 (N_985,In_723,In_708);
nor U986 (N_986,In_158,In_428);
and U987 (N_987,In_572,In_585);
and U988 (N_988,In_699,In_588);
nand U989 (N_989,In_114,In_100);
nor U990 (N_990,In_166,In_55);
nor U991 (N_991,In_472,In_357);
nor U992 (N_992,In_404,In_507);
nor U993 (N_993,In_578,In_554);
or U994 (N_994,In_372,In_310);
or U995 (N_995,In_345,In_65);
nand U996 (N_996,In_526,In_242);
nor U997 (N_997,In_198,In_100);
nor U998 (N_998,In_634,In_165);
nor U999 (N_999,In_664,In_526);
nor U1000 (N_1000,N_184,N_996);
nand U1001 (N_1001,N_244,N_160);
or U1002 (N_1002,N_751,N_580);
and U1003 (N_1003,N_743,N_274);
or U1004 (N_1004,N_871,N_865);
or U1005 (N_1005,N_651,N_703);
nor U1006 (N_1006,N_632,N_532);
and U1007 (N_1007,N_605,N_959);
or U1008 (N_1008,N_335,N_812);
nor U1009 (N_1009,N_132,N_89);
nand U1010 (N_1010,N_297,N_406);
and U1011 (N_1011,N_26,N_428);
nand U1012 (N_1012,N_737,N_255);
nor U1013 (N_1013,N_117,N_223);
nor U1014 (N_1014,N_181,N_732);
or U1015 (N_1015,N_834,N_457);
nand U1016 (N_1016,N_424,N_962);
nor U1017 (N_1017,N_275,N_427);
or U1018 (N_1018,N_788,N_515);
nand U1019 (N_1019,N_248,N_250);
or U1020 (N_1020,N_866,N_260);
and U1021 (N_1021,N_446,N_876);
nand U1022 (N_1022,N_572,N_571);
nand U1023 (N_1023,N_574,N_257);
nor U1024 (N_1024,N_169,N_887);
nand U1025 (N_1025,N_444,N_816);
nor U1026 (N_1026,N_28,N_644);
and U1027 (N_1027,N_649,N_553);
or U1028 (N_1028,N_736,N_848);
nand U1029 (N_1029,N_771,N_977);
or U1030 (N_1030,N_221,N_964);
nand U1031 (N_1031,N_186,N_304);
nor U1032 (N_1032,N_606,N_12);
nor U1033 (N_1033,N_863,N_104);
nand U1034 (N_1034,N_382,N_960);
and U1035 (N_1035,N_313,N_661);
nor U1036 (N_1036,N_49,N_711);
nand U1037 (N_1037,N_264,N_203);
or U1038 (N_1038,N_623,N_589);
nand U1039 (N_1039,N_10,N_123);
and U1040 (N_1040,N_608,N_95);
and U1041 (N_1041,N_521,N_722);
and U1042 (N_1042,N_449,N_84);
or U1043 (N_1043,N_170,N_481);
and U1044 (N_1044,N_310,N_761);
nand U1045 (N_1045,N_319,N_460);
xor U1046 (N_1046,N_942,N_293);
nor U1047 (N_1047,N_835,N_631);
nor U1048 (N_1048,N_204,N_693);
and U1049 (N_1049,N_641,N_781);
nand U1050 (N_1050,N_719,N_557);
nor U1051 (N_1051,N_998,N_196);
or U1052 (N_1052,N_206,N_913);
nor U1053 (N_1053,N_487,N_576);
nor U1054 (N_1054,N_137,N_5);
nand U1055 (N_1055,N_584,N_462);
and U1056 (N_1056,N_493,N_873);
nand U1057 (N_1057,N_272,N_30);
or U1058 (N_1058,N_935,N_669);
and U1059 (N_1059,N_763,N_941);
nand U1060 (N_1060,N_337,N_854);
nand U1061 (N_1061,N_650,N_594);
and U1062 (N_1062,N_65,N_24);
nor U1063 (N_1063,N_249,N_586);
nand U1064 (N_1064,N_738,N_520);
and U1065 (N_1065,N_473,N_536);
and U1066 (N_1066,N_119,N_106);
and U1067 (N_1067,N_896,N_225);
xor U1068 (N_1068,N_948,N_979);
nor U1069 (N_1069,N_893,N_683);
nor U1070 (N_1070,N_407,N_862);
nand U1071 (N_1071,N_360,N_373);
nor U1072 (N_1072,N_602,N_830);
xnor U1073 (N_1073,N_115,N_949);
and U1074 (N_1074,N_980,N_734);
nand U1075 (N_1075,N_789,N_383);
and U1076 (N_1076,N_695,N_111);
and U1077 (N_1077,N_534,N_885);
or U1078 (N_1078,N_279,N_421);
and U1079 (N_1079,N_923,N_684);
nand U1080 (N_1080,N_653,N_218);
or U1081 (N_1081,N_320,N_826);
nand U1082 (N_1082,N_450,N_409);
nand U1083 (N_1083,N_555,N_135);
or U1084 (N_1084,N_116,N_51);
nor U1085 (N_1085,N_400,N_901);
and U1086 (N_1086,N_397,N_418);
and U1087 (N_1087,N_814,N_891);
or U1088 (N_1088,N_262,N_61);
or U1089 (N_1089,N_479,N_668);
or U1090 (N_1090,N_491,N_802);
nor U1091 (N_1091,N_29,N_114);
and U1092 (N_1092,N_844,N_105);
and U1093 (N_1093,N_806,N_251);
nand U1094 (N_1094,N_920,N_285);
and U1095 (N_1095,N_537,N_73);
nor U1096 (N_1096,N_646,N_359);
nand U1097 (N_1097,N_765,N_573);
nor U1098 (N_1098,N_903,N_499);
xor U1099 (N_1099,N_549,N_961);
and U1100 (N_1100,N_577,N_224);
nand U1101 (N_1101,N_987,N_514);
and U1102 (N_1102,N_603,N_899);
nor U1103 (N_1103,N_367,N_944);
nor U1104 (N_1104,N_875,N_66);
nor U1105 (N_1105,N_759,N_859);
nor U1106 (N_1106,N_627,N_940);
and U1107 (N_1107,N_388,N_474);
or U1108 (N_1108,N_813,N_365);
xor U1109 (N_1109,N_152,N_209);
nand U1110 (N_1110,N_452,N_617);
nand U1111 (N_1111,N_656,N_202);
nor U1112 (N_1112,N_775,N_681);
or U1113 (N_1113,N_680,N_380);
nor U1114 (N_1114,N_276,N_195);
or U1115 (N_1115,N_648,N_246);
or U1116 (N_1116,N_433,N_587);
or U1117 (N_1117,N_707,N_420);
or U1118 (N_1118,N_83,N_416);
and U1119 (N_1119,N_639,N_983);
nor U1120 (N_1120,N_674,N_194);
xor U1121 (N_1121,N_370,N_91);
and U1122 (N_1122,N_945,N_3);
or U1123 (N_1123,N_544,N_868);
nor U1124 (N_1124,N_861,N_58);
and U1125 (N_1125,N_592,N_328);
or U1126 (N_1126,N_689,N_773);
or U1127 (N_1127,N_134,N_405);
and U1128 (N_1128,N_102,N_989);
and U1129 (N_1129,N_927,N_966);
nor U1130 (N_1130,N_618,N_166);
or U1131 (N_1131,N_20,N_305);
nand U1132 (N_1132,N_289,N_124);
nor U1133 (N_1133,N_197,N_227);
or U1134 (N_1134,N_506,N_583);
and U1135 (N_1135,N_192,N_528);
nand U1136 (N_1136,N_235,N_870);
and U1137 (N_1137,N_769,N_512);
nand U1138 (N_1138,N_56,N_149);
nor U1139 (N_1139,N_500,N_317);
nand U1140 (N_1140,N_448,N_794);
nor U1141 (N_1141,N_570,N_645);
nor U1142 (N_1142,N_688,N_995);
nor U1143 (N_1143,N_894,N_292);
and U1144 (N_1144,N_157,N_183);
nand U1145 (N_1145,N_867,N_748);
and U1146 (N_1146,N_598,N_219);
or U1147 (N_1147,N_847,N_706);
xor U1148 (N_1148,N_762,N_322);
nand U1149 (N_1149,N_154,N_174);
nand U1150 (N_1150,N_821,N_916);
or U1151 (N_1151,N_151,N_810);
and U1152 (N_1152,N_526,N_671);
or U1153 (N_1153,N_226,N_142);
or U1154 (N_1154,N_538,N_569);
nand U1155 (N_1155,N_364,N_931);
or U1156 (N_1156,N_801,N_430);
or U1157 (N_1157,N_956,N_677);
or U1158 (N_1158,N_120,N_616);
nor U1159 (N_1159,N_890,N_662);
nor U1160 (N_1160,N_687,N_864);
nor U1161 (N_1161,N_978,N_634);
nand U1162 (N_1162,N_558,N_659);
nor U1163 (N_1163,N_808,N_377);
or U1164 (N_1164,N_145,N_193);
and U1165 (N_1165,N_126,N_451);
nor U1166 (N_1166,N_971,N_82);
and U1167 (N_1167,N_331,N_23);
nor U1168 (N_1168,N_880,N_216);
and U1169 (N_1169,N_198,N_22);
or U1170 (N_1170,N_108,N_306);
and U1171 (N_1171,N_746,N_552);
and U1172 (N_1172,N_234,N_981);
nor U1173 (N_1173,N_750,N_175);
nand U1174 (N_1174,N_437,N_256);
and U1175 (N_1175,N_754,N_879);
and U1176 (N_1176,N_352,N_76);
or U1177 (N_1177,N_469,N_682);
or U1178 (N_1178,N_640,N_431);
nand U1179 (N_1179,N_60,N_540);
nor U1180 (N_1180,N_494,N_906);
or U1181 (N_1181,N_829,N_485);
or U1182 (N_1182,N_349,N_395);
or U1183 (N_1183,N_130,N_519);
and U1184 (N_1184,N_658,N_701);
or U1185 (N_1185,N_182,N_888);
nor U1186 (N_1186,N_579,N_811);
and U1187 (N_1187,N_670,N_79);
or U1188 (N_1188,N_220,N_163);
nor U1189 (N_1189,N_34,N_283);
and U1190 (N_1190,N_265,N_509);
nor U1191 (N_1191,N_399,N_635);
or U1192 (N_1192,N_27,N_15);
nand U1193 (N_1193,N_356,N_363);
nand U1194 (N_1194,N_714,N_807);
or U1195 (N_1195,N_368,N_231);
nand U1196 (N_1196,N_189,N_838);
xor U1197 (N_1197,N_443,N_325);
or U1198 (N_1198,N_140,N_261);
or U1199 (N_1199,N_575,N_560);
or U1200 (N_1200,N_269,N_168);
nand U1201 (N_1201,N_884,N_905);
nor U1202 (N_1202,N_94,N_475);
xor U1203 (N_1203,N_975,N_343);
or U1204 (N_1204,N_533,N_8);
nor U1205 (N_1205,N_822,N_836);
nor U1206 (N_1206,N_40,N_378);
nand U1207 (N_1207,N_59,N_904);
and U1208 (N_1208,N_318,N_128);
and U1209 (N_1209,N_665,N_303);
nand U1210 (N_1210,N_122,N_778);
and U1211 (N_1211,N_486,N_882);
and U1212 (N_1212,N_776,N_963);
or U1213 (N_1213,N_311,N_9);
and U1214 (N_1214,N_92,N_717);
or U1215 (N_1215,N_1,N_718);
nand U1216 (N_1216,N_898,N_456);
or U1217 (N_1217,N_624,N_245);
nand U1218 (N_1218,N_419,N_567);
or U1219 (N_1219,N_770,N_477);
nand U1220 (N_1220,N_562,N_466);
nor U1221 (N_1221,N_14,N_372);
and U1222 (N_1222,N_915,N_839);
nor U1223 (N_1223,N_889,N_101);
and U1224 (N_1224,N_259,N_429);
and U1225 (N_1225,N_414,N_369);
nand U1226 (N_1226,N_381,N_910);
nor U1227 (N_1227,N_455,N_277);
nand U1228 (N_1228,N_852,N_955);
nor U1229 (N_1229,N_78,N_582);
nand U1230 (N_1230,N_615,N_842);
nor U1231 (N_1231,N_478,N_967);
nor U1232 (N_1232,N_921,N_841);
or U1233 (N_1233,N_131,N_180);
or U1234 (N_1234,N_673,N_440);
or U1235 (N_1235,N_326,N_11);
and U1236 (N_1236,N_112,N_45);
or U1237 (N_1237,N_926,N_869);
and U1238 (N_1238,N_797,N_502);
and U1239 (N_1239,N_721,N_601);
and U1240 (N_1240,N_323,N_404);
and U1241 (N_1241,N_764,N_127);
and U1242 (N_1242,N_158,N_675);
or U1243 (N_1243,N_663,N_666);
nand U1244 (N_1244,N_18,N_969);
and U1245 (N_1245,N_425,N_612);
nor U1246 (N_1246,N_547,N_976);
nor U1247 (N_1247,N_691,N_556);
nand U1248 (N_1248,N_753,N_697);
nand U1249 (N_1249,N_804,N_148);
nand U1250 (N_1250,N_109,N_236);
or U1251 (N_1251,N_434,N_986);
and U1252 (N_1252,N_713,N_88);
and U1253 (N_1253,N_464,N_539);
nand U1254 (N_1254,N_883,N_386);
nor U1255 (N_1255,N_951,N_930);
and U1256 (N_1256,N_741,N_952);
nor U1257 (N_1257,N_595,N_749);
or U1258 (N_1258,N_690,N_190);
and U1259 (N_1259,N_215,N_176);
nor U1260 (N_1260,N_912,N_340);
nor U1261 (N_1261,N_374,N_630);
and U1262 (N_1262,N_417,N_413);
or U1263 (N_1263,N_622,N_777);
and U1264 (N_1264,N_832,N_379);
nor U1265 (N_1265,N_796,N_53);
or U1266 (N_1266,N_321,N_917);
nor U1267 (N_1267,N_954,N_818);
nand U1268 (N_1268,N_679,N_161);
xnor U1269 (N_1269,N_513,N_990);
and U1270 (N_1270,N_667,N_68);
nor U1271 (N_1271,N_708,N_55);
nor U1272 (N_1272,N_389,N_858);
nor U1273 (N_1273,N_191,N_786);
and U1274 (N_1274,N_657,N_286);
or U1275 (N_1275,N_438,N_568);
nand U1276 (N_1276,N_733,N_943);
nand U1277 (N_1277,N_241,N_445);
or U1278 (N_1278,N_32,N_398);
and U1279 (N_1279,N_729,N_924);
nand U1280 (N_1280,N_72,N_441);
nor U1281 (N_1281,N_302,N_900);
and U1282 (N_1282,N_877,N_823);
nand U1283 (N_1283,N_600,N_212);
nor U1284 (N_1284,N_345,N_93);
or U1285 (N_1285,N_242,N_342);
and U1286 (N_1286,N_881,N_239);
nand U1287 (N_1287,N_287,N_774);
and U1288 (N_1288,N_745,N_790);
or U1289 (N_1289,N_87,N_200);
and U1290 (N_1290,N_237,N_886);
nand U1291 (N_1291,N_937,N_758);
nand U1292 (N_1292,N_655,N_596);
and U1293 (N_1293,N_636,N_613);
nor U1294 (N_1294,N_50,N_38);
and U1295 (N_1295,N_394,N_71);
and U1296 (N_1296,N_290,N_435);
or U1297 (N_1297,N_704,N_97);
or U1298 (N_1298,N_36,N_178);
and U1299 (N_1299,N_610,N_965);
or U1300 (N_1300,N_334,N_564);
nor U1301 (N_1301,N_21,N_447);
and U1302 (N_1302,N_205,N_48);
nand U1303 (N_1303,N_874,N_548);
and U1304 (N_1304,N_840,N_715);
nor U1305 (N_1305,N_831,N_25);
and U1306 (N_1306,N_288,N_207);
nand U1307 (N_1307,N_222,N_86);
or U1308 (N_1308,N_525,N_353);
or U1309 (N_1309,N_43,N_411);
nor U1310 (N_1310,N_495,N_100);
and U1311 (N_1311,N_52,N_785);
or U1312 (N_1312,N_173,N_860);
nand U1313 (N_1313,N_467,N_354);
or U1314 (N_1314,N_415,N_517);
nand U1315 (N_1315,N_107,N_339);
nand U1316 (N_1316,N_757,N_361);
nand U1317 (N_1317,N_57,N_187);
and U1318 (N_1318,N_110,N_599);
or U1319 (N_1319,N_6,N_483);
nand U1320 (N_1320,N_270,N_39);
nor U1321 (N_1321,N_928,N_850);
nor U1322 (N_1322,N_314,N_280);
nand U1323 (N_1323,N_98,N_702);
nand U1324 (N_1324,N_694,N_845);
nand U1325 (N_1325,N_795,N_254);
or U1326 (N_1326,N_725,N_676);
and U1327 (N_1327,N_344,N_803);
or U1328 (N_1328,N_988,N_113);
nand U1329 (N_1329,N_308,N_63);
and U1330 (N_1330,N_902,N_554);
nor U1331 (N_1331,N_74,N_946);
nor U1332 (N_1332,N_267,N_699);
nor U1333 (N_1333,N_492,N_188);
nor U1334 (N_1334,N_984,N_565);
nand U1335 (N_1335,N_217,N_484);
nor U1336 (N_1336,N_504,N_42);
and U1337 (N_1337,N_301,N_471);
and U1338 (N_1338,N_614,N_739);
or U1339 (N_1339,N_578,N_141);
nor U1340 (N_1340,N_507,N_77);
or U1341 (N_1341,N_179,N_208);
nor U1342 (N_1342,N_185,N_633);
nand U1343 (N_1343,N_609,N_709);
and U1344 (N_1344,N_793,N_597);
or U1345 (N_1345,N_299,N_240);
or U1346 (N_1346,N_31,N_637);
and U1347 (N_1347,N_19,N_468);
and U1348 (N_1348,N_607,N_619);
nor U1349 (N_1349,N_787,N_164);
nand U1350 (N_1350,N_529,N_230);
and U1351 (N_1351,N_201,N_970);
nor U1352 (N_1352,N_638,N_792);
or U1353 (N_1353,N_139,N_266);
nand U1354 (N_1354,N_351,N_720);
and U1355 (N_1355,N_233,N_329);
and U1356 (N_1356,N_727,N_156);
nor U1357 (N_1357,N_103,N_531);
or U1358 (N_1358,N_779,N_390);
nand U1359 (N_1359,N_70,N_550);
nand U1360 (N_1360,N_401,N_523);
and U1361 (N_1361,N_543,N_90);
nand U1362 (N_1362,N_933,N_341);
or U1363 (N_1363,N_291,N_843);
nor U1364 (N_1364,N_125,N_642);
and U1365 (N_1365,N_159,N_54);
nand U1366 (N_1366,N_593,N_273);
and U1367 (N_1367,N_731,N_392);
or U1368 (N_1368,N_664,N_505);
or U1369 (N_1369,N_535,N_756);
and U1370 (N_1370,N_999,N_150);
or U1371 (N_1371,N_740,N_710);
or U1372 (N_1372,N_80,N_643);
nand U1373 (N_1373,N_138,N_284);
or U1374 (N_1374,N_992,N_621);
nor U1375 (N_1375,N_647,N_974);
and U1376 (N_1376,N_700,N_393);
nor U1377 (N_1377,N_96,N_895);
nor U1378 (N_1378,N_33,N_735);
and U1379 (N_1379,N_805,N_872);
nor U1380 (N_1380,N_892,N_358);
and U1381 (N_1381,N_426,N_371);
and U1382 (N_1382,N_403,N_561);
and U1383 (N_1383,N_17,N_375);
or U1384 (N_1384,N_263,N_324);
and U1385 (N_1385,N_897,N_968);
nand U1386 (N_1386,N_947,N_37);
and U1387 (N_1387,N_489,N_972);
and U1388 (N_1388,N_307,N_837);
and U1389 (N_1389,N_162,N_387);
nor U1390 (N_1390,N_490,N_384);
nor U1391 (N_1391,N_228,N_133);
nand U1392 (N_1392,N_985,N_851);
nor U1393 (N_1393,N_522,N_2);
or U1394 (N_1394,N_332,N_652);
and U1395 (N_1395,N_716,N_857);
xor U1396 (N_1396,N_747,N_585);
nor U1397 (N_1397,N_376,N_783);
nand U1398 (N_1398,N_497,N_780);
or U1399 (N_1399,N_482,N_496);
nor U1400 (N_1400,N_121,N_672);
or U1401 (N_1401,N_213,N_846);
nand U1402 (N_1402,N_827,N_476);
nor U1403 (N_1403,N_67,N_768);
or U1404 (N_1404,N_336,N_692);
and U1405 (N_1405,N_503,N_686);
nand U1406 (N_1406,N_147,N_993);
or U1407 (N_1407,N_542,N_620);
nor U1408 (N_1408,N_799,N_791);
or U1409 (N_1409,N_118,N_129);
or U1410 (N_1410,N_412,N_13);
nor U1411 (N_1411,N_938,N_590);
and U1412 (N_1412,N_546,N_423);
nor U1413 (N_1413,N_755,N_472);
or U1414 (N_1414,N_516,N_357);
and U1415 (N_1415,N_611,N_396);
xnor U1416 (N_1416,N_934,N_0);
xor U1417 (N_1417,N_766,N_391);
nor U1418 (N_1418,N_171,N_698);
xor U1419 (N_1419,N_909,N_199);
or U1420 (N_1420,N_918,N_69);
and U1421 (N_1421,N_309,N_510);
nor U1422 (N_1422,N_654,N_410);
nand U1423 (N_1423,N_282,N_271);
or U1424 (N_1424,N_524,N_936);
or U1425 (N_1425,N_723,N_824);
nand U1426 (N_1426,N_432,N_258);
nor U1427 (N_1427,N_950,N_685);
nand U1428 (N_1428,N_458,N_712);
nand U1429 (N_1429,N_581,N_143);
and U1430 (N_1430,N_346,N_402);
nor U1431 (N_1431,N_350,N_165);
or U1432 (N_1432,N_465,N_243);
nor U1433 (N_1433,N_825,N_167);
or U1434 (N_1434,N_800,N_878);
nand U1435 (N_1435,N_752,N_767);
or U1436 (N_1436,N_817,N_238);
and U1437 (N_1437,N_366,N_563);
and U1438 (N_1438,N_742,N_146);
nand U1439 (N_1439,N_44,N_760);
or U1440 (N_1440,N_75,N_62);
nor U1441 (N_1441,N_628,N_488);
nand U1442 (N_1442,N_136,N_300);
or U1443 (N_1443,N_922,N_347);
nand U1444 (N_1444,N_296,N_798);
nor U1445 (N_1445,N_728,N_81);
or U1446 (N_1446,N_408,N_991);
nor U1447 (N_1447,N_518,N_994);
and U1448 (N_1448,N_16,N_315);
and U1449 (N_1449,N_177,N_281);
nand U1450 (N_1450,N_362,N_155);
and U1451 (N_1451,N_541,N_232);
or U1452 (N_1452,N_253,N_588);
and U1453 (N_1453,N_41,N_982);
xor U1454 (N_1454,N_463,N_439);
xnor U1455 (N_1455,N_153,N_298);
nand U1456 (N_1456,N_591,N_907);
or U1457 (N_1457,N_330,N_385);
or U1458 (N_1458,N_784,N_470);
or U1459 (N_1459,N_453,N_958);
or U1460 (N_1460,N_932,N_46);
or U1461 (N_1461,N_459,N_229);
nor U1462 (N_1462,N_730,N_530);
and U1463 (N_1463,N_422,N_626);
nor U1464 (N_1464,N_696,N_294);
nand U1465 (N_1465,N_772,N_47);
nand U1466 (N_1466,N_604,N_501);
or U1467 (N_1467,N_625,N_348);
nor U1468 (N_1468,N_461,N_726);
and U1469 (N_1469,N_144,N_247);
nand U1470 (N_1470,N_914,N_480);
nand U1471 (N_1471,N_782,N_559);
and U1472 (N_1472,N_856,N_833);
and U1473 (N_1473,N_849,N_925);
and U1474 (N_1474,N_511,N_828);
or U1475 (N_1475,N_953,N_7);
nor U1476 (N_1476,N_99,N_35);
nor U1477 (N_1477,N_678,N_508);
xor U1478 (N_1478,N_744,N_327);
or U1479 (N_1479,N_929,N_815);
or U1480 (N_1480,N_172,N_333);
or U1481 (N_1481,N_312,N_660);
or U1482 (N_1482,N_629,N_295);
nor U1483 (N_1483,N_64,N_498);
nor U1484 (N_1484,N_214,N_705);
nor U1485 (N_1485,N_939,N_997);
or U1486 (N_1486,N_355,N_853);
nand U1487 (N_1487,N_454,N_566);
nand U1488 (N_1488,N_436,N_252);
and U1489 (N_1489,N_957,N_527);
nand U1490 (N_1490,N_908,N_211);
or U1491 (N_1491,N_338,N_919);
or U1492 (N_1492,N_545,N_268);
or U1493 (N_1493,N_973,N_855);
nor U1494 (N_1494,N_278,N_819);
nand U1495 (N_1495,N_911,N_316);
nand U1496 (N_1496,N_442,N_809);
or U1497 (N_1497,N_4,N_210);
and U1498 (N_1498,N_724,N_551);
nand U1499 (N_1499,N_820,N_85);
nor U1500 (N_1500,N_156,N_235);
nand U1501 (N_1501,N_809,N_374);
or U1502 (N_1502,N_23,N_536);
nor U1503 (N_1503,N_629,N_452);
or U1504 (N_1504,N_860,N_730);
or U1505 (N_1505,N_662,N_458);
nor U1506 (N_1506,N_402,N_589);
nor U1507 (N_1507,N_554,N_445);
nand U1508 (N_1508,N_81,N_358);
and U1509 (N_1509,N_0,N_528);
nand U1510 (N_1510,N_51,N_114);
and U1511 (N_1511,N_187,N_984);
and U1512 (N_1512,N_874,N_748);
and U1513 (N_1513,N_814,N_336);
nor U1514 (N_1514,N_429,N_789);
nand U1515 (N_1515,N_656,N_653);
and U1516 (N_1516,N_68,N_381);
and U1517 (N_1517,N_434,N_13);
and U1518 (N_1518,N_337,N_52);
or U1519 (N_1519,N_57,N_33);
and U1520 (N_1520,N_945,N_288);
nor U1521 (N_1521,N_889,N_867);
or U1522 (N_1522,N_52,N_245);
nor U1523 (N_1523,N_691,N_495);
and U1524 (N_1524,N_56,N_524);
or U1525 (N_1525,N_67,N_128);
or U1526 (N_1526,N_736,N_165);
and U1527 (N_1527,N_356,N_698);
or U1528 (N_1528,N_418,N_826);
nand U1529 (N_1529,N_917,N_293);
or U1530 (N_1530,N_780,N_80);
nor U1531 (N_1531,N_76,N_70);
and U1532 (N_1532,N_83,N_391);
nor U1533 (N_1533,N_177,N_504);
nand U1534 (N_1534,N_908,N_677);
and U1535 (N_1535,N_856,N_806);
nor U1536 (N_1536,N_402,N_29);
nor U1537 (N_1537,N_737,N_462);
and U1538 (N_1538,N_111,N_719);
or U1539 (N_1539,N_902,N_270);
nor U1540 (N_1540,N_326,N_219);
or U1541 (N_1541,N_480,N_63);
nand U1542 (N_1542,N_109,N_420);
or U1543 (N_1543,N_563,N_586);
nor U1544 (N_1544,N_380,N_162);
and U1545 (N_1545,N_897,N_713);
or U1546 (N_1546,N_384,N_904);
or U1547 (N_1547,N_260,N_919);
or U1548 (N_1548,N_426,N_14);
and U1549 (N_1549,N_962,N_217);
or U1550 (N_1550,N_809,N_329);
nor U1551 (N_1551,N_444,N_878);
nor U1552 (N_1552,N_856,N_587);
or U1553 (N_1553,N_126,N_464);
nor U1554 (N_1554,N_496,N_931);
or U1555 (N_1555,N_921,N_544);
nor U1556 (N_1556,N_919,N_777);
nand U1557 (N_1557,N_34,N_637);
and U1558 (N_1558,N_814,N_980);
and U1559 (N_1559,N_52,N_325);
nor U1560 (N_1560,N_860,N_791);
and U1561 (N_1561,N_705,N_638);
and U1562 (N_1562,N_893,N_911);
nand U1563 (N_1563,N_322,N_658);
and U1564 (N_1564,N_692,N_358);
nand U1565 (N_1565,N_313,N_237);
or U1566 (N_1566,N_125,N_431);
nor U1567 (N_1567,N_889,N_167);
and U1568 (N_1568,N_841,N_258);
or U1569 (N_1569,N_162,N_920);
nand U1570 (N_1570,N_135,N_413);
nand U1571 (N_1571,N_33,N_370);
and U1572 (N_1572,N_658,N_759);
or U1573 (N_1573,N_226,N_73);
nand U1574 (N_1574,N_410,N_613);
or U1575 (N_1575,N_768,N_869);
or U1576 (N_1576,N_304,N_913);
or U1577 (N_1577,N_519,N_568);
and U1578 (N_1578,N_191,N_225);
and U1579 (N_1579,N_926,N_809);
and U1580 (N_1580,N_187,N_620);
and U1581 (N_1581,N_240,N_180);
nor U1582 (N_1582,N_964,N_445);
nor U1583 (N_1583,N_840,N_965);
nor U1584 (N_1584,N_567,N_863);
and U1585 (N_1585,N_628,N_2);
xnor U1586 (N_1586,N_591,N_818);
and U1587 (N_1587,N_110,N_68);
and U1588 (N_1588,N_84,N_20);
or U1589 (N_1589,N_460,N_57);
and U1590 (N_1590,N_411,N_926);
or U1591 (N_1591,N_425,N_67);
or U1592 (N_1592,N_414,N_647);
and U1593 (N_1593,N_909,N_818);
nand U1594 (N_1594,N_506,N_845);
or U1595 (N_1595,N_447,N_51);
or U1596 (N_1596,N_433,N_462);
nor U1597 (N_1597,N_816,N_401);
nand U1598 (N_1598,N_142,N_992);
or U1599 (N_1599,N_288,N_630);
nand U1600 (N_1600,N_911,N_214);
and U1601 (N_1601,N_46,N_63);
xor U1602 (N_1602,N_360,N_574);
nor U1603 (N_1603,N_461,N_693);
and U1604 (N_1604,N_527,N_307);
nor U1605 (N_1605,N_389,N_387);
nand U1606 (N_1606,N_631,N_682);
nand U1607 (N_1607,N_758,N_933);
or U1608 (N_1608,N_181,N_628);
or U1609 (N_1609,N_251,N_814);
nor U1610 (N_1610,N_169,N_751);
or U1611 (N_1611,N_447,N_722);
and U1612 (N_1612,N_603,N_937);
and U1613 (N_1613,N_632,N_812);
nor U1614 (N_1614,N_979,N_189);
and U1615 (N_1615,N_645,N_64);
nor U1616 (N_1616,N_472,N_346);
nand U1617 (N_1617,N_576,N_326);
or U1618 (N_1618,N_655,N_980);
and U1619 (N_1619,N_213,N_272);
and U1620 (N_1620,N_305,N_739);
and U1621 (N_1621,N_605,N_242);
nor U1622 (N_1622,N_644,N_94);
or U1623 (N_1623,N_127,N_316);
nor U1624 (N_1624,N_909,N_118);
nor U1625 (N_1625,N_142,N_274);
nand U1626 (N_1626,N_830,N_304);
nand U1627 (N_1627,N_225,N_498);
nor U1628 (N_1628,N_968,N_315);
nor U1629 (N_1629,N_784,N_301);
and U1630 (N_1630,N_12,N_73);
or U1631 (N_1631,N_110,N_299);
nor U1632 (N_1632,N_743,N_413);
nor U1633 (N_1633,N_880,N_155);
and U1634 (N_1634,N_990,N_311);
nand U1635 (N_1635,N_122,N_645);
nor U1636 (N_1636,N_192,N_850);
or U1637 (N_1637,N_802,N_48);
or U1638 (N_1638,N_757,N_373);
nand U1639 (N_1639,N_266,N_489);
nand U1640 (N_1640,N_106,N_323);
and U1641 (N_1641,N_654,N_439);
and U1642 (N_1642,N_393,N_200);
nand U1643 (N_1643,N_966,N_877);
and U1644 (N_1644,N_711,N_130);
nand U1645 (N_1645,N_44,N_780);
and U1646 (N_1646,N_354,N_482);
or U1647 (N_1647,N_385,N_858);
nand U1648 (N_1648,N_520,N_998);
nand U1649 (N_1649,N_565,N_136);
nor U1650 (N_1650,N_406,N_99);
and U1651 (N_1651,N_668,N_932);
nand U1652 (N_1652,N_614,N_886);
nand U1653 (N_1653,N_525,N_396);
and U1654 (N_1654,N_807,N_18);
nand U1655 (N_1655,N_744,N_422);
and U1656 (N_1656,N_947,N_237);
nand U1657 (N_1657,N_734,N_264);
nand U1658 (N_1658,N_604,N_656);
nor U1659 (N_1659,N_657,N_504);
nand U1660 (N_1660,N_585,N_151);
nor U1661 (N_1661,N_491,N_742);
or U1662 (N_1662,N_996,N_225);
nand U1663 (N_1663,N_8,N_574);
nand U1664 (N_1664,N_692,N_932);
or U1665 (N_1665,N_799,N_807);
nor U1666 (N_1666,N_239,N_49);
or U1667 (N_1667,N_148,N_742);
or U1668 (N_1668,N_368,N_482);
and U1669 (N_1669,N_904,N_640);
and U1670 (N_1670,N_556,N_174);
nor U1671 (N_1671,N_730,N_188);
nor U1672 (N_1672,N_101,N_305);
nor U1673 (N_1673,N_119,N_772);
and U1674 (N_1674,N_295,N_99);
nand U1675 (N_1675,N_577,N_442);
nor U1676 (N_1676,N_792,N_817);
nand U1677 (N_1677,N_437,N_961);
and U1678 (N_1678,N_644,N_513);
and U1679 (N_1679,N_358,N_876);
or U1680 (N_1680,N_873,N_381);
and U1681 (N_1681,N_822,N_472);
nand U1682 (N_1682,N_411,N_953);
and U1683 (N_1683,N_334,N_135);
and U1684 (N_1684,N_516,N_205);
or U1685 (N_1685,N_415,N_768);
nor U1686 (N_1686,N_883,N_503);
or U1687 (N_1687,N_866,N_722);
nand U1688 (N_1688,N_630,N_487);
nor U1689 (N_1689,N_217,N_216);
nor U1690 (N_1690,N_902,N_644);
and U1691 (N_1691,N_403,N_4);
nand U1692 (N_1692,N_118,N_226);
nor U1693 (N_1693,N_650,N_630);
nand U1694 (N_1694,N_789,N_330);
nand U1695 (N_1695,N_708,N_73);
nand U1696 (N_1696,N_726,N_30);
and U1697 (N_1697,N_888,N_473);
or U1698 (N_1698,N_783,N_102);
nor U1699 (N_1699,N_839,N_934);
and U1700 (N_1700,N_57,N_79);
nor U1701 (N_1701,N_684,N_635);
nand U1702 (N_1702,N_359,N_436);
or U1703 (N_1703,N_224,N_839);
and U1704 (N_1704,N_966,N_190);
and U1705 (N_1705,N_750,N_986);
nor U1706 (N_1706,N_861,N_230);
nor U1707 (N_1707,N_984,N_390);
or U1708 (N_1708,N_716,N_312);
nor U1709 (N_1709,N_51,N_326);
or U1710 (N_1710,N_532,N_806);
or U1711 (N_1711,N_507,N_236);
and U1712 (N_1712,N_29,N_770);
or U1713 (N_1713,N_890,N_11);
or U1714 (N_1714,N_971,N_55);
and U1715 (N_1715,N_482,N_453);
and U1716 (N_1716,N_978,N_18);
and U1717 (N_1717,N_803,N_411);
or U1718 (N_1718,N_753,N_7);
or U1719 (N_1719,N_611,N_883);
or U1720 (N_1720,N_788,N_592);
or U1721 (N_1721,N_365,N_388);
nand U1722 (N_1722,N_787,N_675);
nand U1723 (N_1723,N_175,N_669);
nor U1724 (N_1724,N_796,N_605);
nand U1725 (N_1725,N_588,N_331);
nand U1726 (N_1726,N_37,N_450);
nand U1727 (N_1727,N_367,N_324);
nand U1728 (N_1728,N_486,N_558);
nor U1729 (N_1729,N_185,N_175);
nor U1730 (N_1730,N_200,N_449);
and U1731 (N_1731,N_213,N_333);
or U1732 (N_1732,N_19,N_717);
or U1733 (N_1733,N_796,N_748);
or U1734 (N_1734,N_528,N_129);
nor U1735 (N_1735,N_201,N_827);
nand U1736 (N_1736,N_455,N_902);
nand U1737 (N_1737,N_54,N_205);
and U1738 (N_1738,N_503,N_484);
nand U1739 (N_1739,N_669,N_902);
nand U1740 (N_1740,N_310,N_815);
nor U1741 (N_1741,N_157,N_138);
nor U1742 (N_1742,N_636,N_729);
nor U1743 (N_1743,N_619,N_144);
nand U1744 (N_1744,N_41,N_549);
or U1745 (N_1745,N_498,N_748);
and U1746 (N_1746,N_309,N_370);
nor U1747 (N_1747,N_244,N_420);
and U1748 (N_1748,N_47,N_357);
and U1749 (N_1749,N_990,N_645);
and U1750 (N_1750,N_353,N_826);
nor U1751 (N_1751,N_833,N_14);
or U1752 (N_1752,N_462,N_569);
or U1753 (N_1753,N_878,N_959);
nor U1754 (N_1754,N_344,N_582);
nor U1755 (N_1755,N_81,N_473);
nor U1756 (N_1756,N_971,N_711);
and U1757 (N_1757,N_781,N_523);
nor U1758 (N_1758,N_708,N_19);
nand U1759 (N_1759,N_975,N_492);
nor U1760 (N_1760,N_662,N_348);
nand U1761 (N_1761,N_811,N_822);
nor U1762 (N_1762,N_355,N_162);
nor U1763 (N_1763,N_756,N_653);
and U1764 (N_1764,N_405,N_706);
nor U1765 (N_1765,N_883,N_705);
or U1766 (N_1766,N_763,N_639);
nor U1767 (N_1767,N_183,N_42);
and U1768 (N_1768,N_627,N_387);
xor U1769 (N_1769,N_422,N_215);
and U1770 (N_1770,N_458,N_152);
and U1771 (N_1771,N_194,N_850);
nor U1772 (N_1772,N_378,N_796);
and U1773 (N_1773,N_347,N_120);
and U1774 (N_1774,N_529,N_724);
nand U1775 (N_1775,N_247,N_159);
and U1776 (N_1776,N_945,N_30);
nor U1777 (N_1777,N_478,N_783);
or U1778 (N_1778,N_772,N_33);
nor U1779 (N_1779,N_319,N_431);
or U1780 (N_1780,N_700,N_370);
nand U1781 (N_1781,N_803,N_71);
nand U1782 (N_1782,N_502,N_665);
nor U1783 (N_1783,N_735,N_703);
and U1784 (N_1784,N_390,N_410);
nor U1785 (N_1785,N_978,N_208);
nand U1786 (N_1786,N_177,N_575);
nor U1787 (N_1787,N_91,N_151);
and U1788 (N_1788,N_351,N_108);
nand U1789 (N_1789,N_667,N_777);
nor U1790 (N_1790,N_68,N_254);
nor U1791 (N_1791,N_980,N_795);
and U1792 (N_1792,N_420,N_111);
nand U1793 (N_1793,N_449,N_824);
or U1794 (N_1794,N_984,N_518);
and U1795 (N_1795,N_753,N_931);
nor U1796 (N_1796,N_980,N_480);
or U1797 (N_1797,N_749,N_29);
nand U1798 (N_1798,N_464,N_578);
nor U1799 (N_1799,N_392,N_185);
nor U1800 (N_1800,N_995,N_201);
or U1801 (N_1801,N_99,N_109);
and U1802 (N_1802,N_642,N_923);
nand U1803 (N_1803,N_904,N_606);
and U1804 (N_1804,N_25,N_842);
nor U1805 (N_1805,N_235,N_200);
nor U1806 (N_1806,N_128,N_627);
and U1807 (N_1807,N_891,N_225);
nor U1808 (N_1808,N_850,N_943);
nor U1809 (N_1809,N_205,N_943);
nor U1810 (N_1810,N_760,N_22);
nand U1811 (N_1811,N_74,N_782);
and U1812 (N_1812,N_23,N_294);
nand U1813 (N_1813,N_807,N_585);
nor U1814 (N_1814,N_784,N_617);
nor U1815 (N_1815,N_270,N_896);
and U1816 (N_1816,N_230,N_266);
and U1817 (N_1817,N_494,N_873);
or U1818 (N_1818,N_699,N_373);
and U1819 (N_1819,N_270,N_825);
and U1820 (N_1820,N_910,N_312);
nand U1821 (N_1821,N_979,N_267);
xnor U1822 (N_1822,N_554,N_608);
or U1823 (N_1823,N_316,N_190);
nor U1824 (N_1824,N_448,N_309);
or U1825 (N_1825,N_991,N_111);
and U1826 (N_1826,N_768,N_270);
and U1827 (N_1827,N_323,N_623);
and U1828 (N_1828,N_953,N_901);
nand U1829 (N_1829,N_440,N_749);
and U1830 (N_1830,N_805,N_118);
nor U1831 (N_1831,N_781,N_319);
nand U1832 (N_1832,N_818,N_254);
or U1833 (N_1833,N_837,N_862);
or U1834 (N_1834,N_422,N_903);
nor U1835 (N_1835,N_699,N_766);
and U1836 (N_1836,N_319,N_749);
and U1837 (N_1837,N_645,N_968);
nor U1838 (N_1838,N_112,N_360);
and U1839 (N_1839,N_20,N_619);
nor U1840 (N_1840,N_424,N_712);
or U1841 (N_1841,N_821,N_654);
nand U1842 (N_1842,N_367,N_729);
and U1843 (N_1843,N_933,N_32);
or U1844 (N_1844,N_362,N_326);
nand U1845 (N_1845,N_798,N_839);
nor U1846 (N_1846,N_245,N_418);
or U1847 (N_1847,N_436,N_922);
nand U1848 (N_1848,N_237,N_646);
xor U1849 (N_1849,N_276,N_485);
and U1850 (N_1850,N_634,N_665);
and U1851 (N_1851,N_539,N_643);
and U1852 (N_1852,N_851,N_96);
nor U1853 (N_1853,N_514,N_819);
or U1854 (N_1854,N_87,N_775);
nor U1855 (N_1855,N_306,N_866);
and U1856 (N_1856,N_662,N_397);
or U1857 (N_1857,N_327,N_454);
nor U1858 (N_1858,N_320,N_59);
nand U1859 (N_1859,N_405,N_951);
or U1860 (N_1860,N_560,N_709);
nor U1861 (N_1861,N_911,N_851);
nand U1862 (N_1862,N_383,N_321);
nand U1863 (N_1863,N_240,N_597);
nand U1864 (N_1864,N_372,N_20);
nor U1865 (N_1865,N_894,N_785);
and U1866 (N_1866,N_474,N_30);
or U1867 (N_1867,N_1,N_518);
nor U1868 (N_1868,N_209,N_501);
or U1869 (N_1869,N_813,N_604);
nand U1870 (N_1870,N_120,N_911);
nand U1871 (N_1871,N_889,N_675);
nor U1872 (N_1872,N_540,N_847);
nand U1873 (N_1873,N_900,N_511);
or U1874 (N_1874,N_507,N_301);
and U1875 (N_1875,N_605,N_899);
nand U1876 (N_1876,N_143,N_759);
or U1877 (N_1877,N_221,N_637);
nand U1878 (N_1878,N_34,N_645);
and U1879 (N_1879,N_627,N_838);
or U1880 (N_1880,N_950,N_911);
nand U1881 (N_1881,N_229,N_442);
nand U1882 (N_1882,N_729,N_354);
nor U1883 (N_1883,N_296,N_956);
nor U1884 (N_1884,N_576,N_205);
or U1885 (N_1885,N_139,N_648);
and U1886 (N_1886,N_208,N_562);
nor U1887 (N_1887,N_374,N_415);
nand U1888 (N_1888,N_901,N_845);
nand U1889 (N_1889,N_926,N_678);
or U1890 (N_1890,N_204,N_598);
nor U1891 (N_1891,N_912,N_792);
and U1892 (N_1892,N_711,N_308);
and U1893 (N_1893,N_355,N_826);
nor U1894 (N_1894,N_428,N_278);
and U1895 (N_1895,N_78,N_403);
and U1896 (N_1896,N_184,N_713);
and U1897 (N_1897,N_568,N_552);
nand U1898 (N_1898,N_788,N_212);
and U1899 (N_1899,N_252,N_805);
nor U1900 (N_1900,N_130,N_241);
nand U1901 (N_1901,N_690,N_625);
and U1902 (N_1902,N_572,N_518);
nor U1903 (N_1903,N_94,N_270);
nor U1904 (N_1904,N_956,N_550);
nor U1905 (N_1905,N_43,N_338);
and U1906 (N_1906,N_128,N_233);
nand U1907 (N_1907,N_973,N_145);
or U1908 (N_1908,N_841,N_520);
nand U1909 (N_1909,N_299,N_656);
nand U1910 (N_1910,N_379,N_133);
and U1911 (N_1911,N_819,N_776);
nor U1912 (N_1912,N_653,N_697);
or U1913 (N_1913,N_100,N_75);
nor U1914 (N_1914,N_98,N_189);
nor U1915 (N_1915,N_413,N_955);
nor U1916 (N_1916,N_29,N_324);
and U1917 (N_1917,N_233,N_537);
or U1918 (N_1918,N_514,N_551);
nand U1919 (N_1919,N_176,N_292);
nor U1920 (N_1920,N_992,N_445);
nor U1921 (N_1921,N_210,N_796);
nor U1922 (N_1922,N_90,N_695);
or U1923 (N_1923,N_486,N_343);
nand U1924 (N_1924,N_724,N_917);
or U1925 (N_1925,N_822,N_337);
nor U1926 (N_1926,N_740,N_37);
and U1927 (N_1927,N_278,N_578);
or U1928 (N_1928,N_452,N_450);
nand U1929 (N_1929,N_218,N_682);
nand U1930 (N_1930,N_682,N_651);
or U1931 (N_1931,N_299,N_406);
nor U1932 (N_1932,N_391,N_309);
and U1933 (N_1933,N_579,N_839);
nor U1934 (N_1934,N_791,N_493);
nor U1935 (N_1935,N_807,N_880);
or U1936 (N_1936,N_450,N_814);
nor U1937 (N_1937,N_279,N_67);
nand U1938 (N_1938,N_946,N_540);
nor U1939 (N_1939,N_97,N_562);
and U1940 (N_1940,N_261,N_902);
nor U1941 (N_1941,N_51,N_635);
nor U1942 (N_1942,N_789,N_871);
or U1943 (N_1943,N_604,N_52);
and U1944 (N_1944,N_155,N_372);
nand U1945 (N_1945,N_933,N_92);
nand U1946 (N_1946,N_180,N_37);
nand U1947 (N_1947,N_626,N_837);
or U1948 (N_1948,N_587,N_689);
or U1949 (N_1949,N_589,N_75);
and U1950 (N_1950,N_527,N_574);
and U1951 (N_1951,N_382,N_334);
nor U1952 (N_1952,N_343,N_13);
nor U1953 (N_1953,N_310,N_628);
or U1954 (N_1954,N_913,N_217);
or U1955 (N_1955,N_471,N_642);
nor U1956 (N_1956,N_953,N_246);
or U1957 (N_1957,N_50,N_381);
or U1958 (N_1958,N_313,N_140);
and U1959 (N_1959,N_105,N_937);
or U1960 (N_1960,N_61,N_499);
or U1961 (N_1961,N_822,N_264);
or U1962 (N_1962,N_841,N_621);
or U1963 (N_1963,N_340,N_671);
or U1964 (N_1964,N_969,N_70);
nand U1965 (N_1965,N_120,N_4);
and U1966 (N_1966,N_46,N_665);
nor U1967 (N_1967,N_415,N_649);
nand U1968 (N_1968,N_544,N_613);
or U1969 (N_1969,N_771,N_685);
nand U1970 (N_1970,N_87,N_964);
nand U1971 (N_1971,N_88,N_436);
nor U1972 (N_1972,N_611,N_422);
and U1973 (N_1973,N_812,N_571);
or U1974 (N_1974,N_334,N_592);
nor U1975 (N_1975,N_637,N_344);
nor U1976 (N_1976,N_335,N_257);
nand U1977 (N_1977,N_101,N_842);
nor U1978 (N_1978,N_321,N_238);
and U1979 (N_1979,N_569,N_306);
or U1980 (N_1980,N_507,N_398);
nor U1981 (N_1981,N_197,N_646);
and U1982 (N_1982,N_306,N_36);
and U1983 (N_1983,N_511,N_158);
or U1984 (N_1984,N_922,N_447);
nor U1985 (N_1985,N_751,N_482);
or U1986 (N_1986,N_838,N_786);
nor U1987 (N_1987,N_683,N_133);
nand U1988 (N_1988,N_357,N_402);
or U1989 (N_1989,N_10,N_116);
nor U1990 (N_1990,N_590,N_870);
nand U1991 (N_1991,N_228,N_399);
nand U1992 (N_1992,N_949,N_92);
nor U1993 (N_1993,N_290,N_336);
nand U1994 (N_1994,N_210,N_386);
nand U1995 (N_1995,N_70,N_348);
nand U1996 (N_1996,N_286,N_973);
and U1997 (N_1997,N_237,N_508);
or U1998 (N_1998,N_326,N_767);
nor U1999 (N_1999,N_831,N_11);
nor U2000 (N_2000,N_1733,N_1217);
and U2001 (N_2001,N_1761,N_1920);
or U2002 (N_2002,N_1596,N_1014);
nor U2003 (N_2003,N_1111,N_1650);
nand U2004 (N_2004,N_1592,N_1712);
or U2005 (N_2005,N_1750,N_1113);
and U2006 (N_2006,N_1143,N_1969);
nand U2007 (N_2007,N_1424,N_1739);
and U2008 (N_2008,N_1495,N_1049);
or U2009 (N_2009,N_1986,N_1076);
and U2010 (N_2010,N_1188,N_1843);
nand U2011 (N_2011,N_1058,N_1308);
or U2012 (N_2012,N_1720,N_1734);
or U2013 (N_2013,N_1430,N_1862);
or U2014 (N_2014,N_1698,N_1857);
and U2015 (N_2015,N_1150,N_1011);
or U2016 (N_2016,N_1778,N_1919);
and U2017 (N_2017,N_1764,N_1556);
nand U2018 (N_2018,N_1293,N_1263);
or U2019 (N_2019,N_1410,N_1906);
nor U2020 (N_2020,N_1114,N_1674);
or U2021 (N_2021,N_1020,N_1291);
nand U2022 (N_2022,N_1854,N_1528);
nand U2023 (N_2023,N_1483,N_1184);
and U2024 (N_2024,N_1790,N_1061);
nor U2025 (N_2025,N_1318,N_1851);
nand U2026 (N_2026,N_1891,N_1865);
nor U2027 (N_2027,N_1322,N_1497);
or U2028 (N_2028,N_1725,N_1962);
nand U2029 (N_2029,N_1486,N_1446);
nand U2030 (N_2030,N_1794,N_1785);
nand U2031 (N_2031,N_1043,N_1417);
nand U2032 (N_2032,N_1988,N_1493);
nor U2033 (N_2033,N_1035,N_1386);
nand U2034 (N_2034,N_1861,N_1628);
and U2035 (N_2035,N_1543,N_1363);
and U2036 (N_2036,N_1411,N_1910);
or U2037 (N_2037,N_1859,N_1335);
or U2038 (N_2038,N_1309,N_1983);
or U2039 (N_2039,N_1173,N_1894);
and U2040 (N_2040,N_1618,N_1566);
nand U2041 (N_2041,N_1075,N_1577);
nor U2042 (N_2042,N_1632,N_1029);
nor U2043 (N_2043,N_1202,N_1547);
nor U2044 (N_2044,N_1824,N_1998);
and U2045 (N_2045,N_1179,N_1615);
nor U2046 (N_2046,N_1956,N_1228);
nor U2047 (N_2047,N_1849,N_1685);
nor U2048 (N_2048,N_1837,N_1203);
nand U2049 (N_2049,N_1270,N_1071);
nand U2050 (N_2050,N_1719,N_1783);
nand U2051 (N_2051,N_1044,N_1256);
nor U2052 (N_2052,N_1868,N_1244);
nand U2053 (N_2053,N_1468,N_1091);
nor U2054 (N_2054,N_1673,N_1893);
and U2055 (N_2055,N_1409,N_1925);
and U2056 (N_2056,N_1737,N_1062);
and U2057 (N_2057,N_1554,N_1816);
nand U2058 (N_2058,N_1182,N_1999);
nand U2059 (N_2059,N_1141,N_1505);
nand U2060 (N_2060,N_1457,N_1985);
or U2061 (N_2061,N_1022,N_1162);
and U2062 (N_2062,N_1569,N_1520);
nand U2063 (N_2063,N_1531,N_1881);
and U2064 (N_2064,N_1214,N_1169);
and U2065 (N_2065,N_1391,N_1670);
nor U2066 (N_2066,N_1819,N_1453);
nand U2067 (N_2067,N_1423,N_1436);
and U2068 (N_2068,N_1589,N_1081);
nor U2069 (N_2069,N_1835,N_1025);
or U2070 (N_2070,N_1361,N_1137);
and U2071 (N_2071,N_1357,N_1401);
and U2072 (N_2072,N_1311,N_1106);
nand U2073 (N_2073,N_1458,N_1475);
nor U2074 (N_2074,N_1372,N_1266);
and U2075 (N_2075,N_1504,N_1017);
nand U2076 (N_2076,N_1271,N_1492);
nand U2077 (N_2077,N_1220,N_1665);
nand U2078 (N_2078,N_1482,N_1333);
nand U2079 (N_2079,N_1353,N_1287);
or U2080 (N_2080,N_1642,N_1339);
or U2081 (N_2081,N_1388,N_1187);
or U2082 (N_2082,N_1845,N_1542);
and U2083 (N_2083,N_1275,N_1779);
or U2084 (N_2084,N_1261,N_1591);
nor U2085 (N_2085,N_1935,N_1623);
nand U2086 (N_2086,N_1129,N_1756);
nand U2087 (N_2087,N_1957,N_1107);
nor U2088 (N_2088,N_1503,N_1329);
and U2089 (N_2089,N_1358,N_1747);
nor U2090 (N_2090,N_1929,N_1715);
or U2091 (N_2091,N_1234,N_1200);
or U2092 (N_2092,N_1099,N_1751);
nand U2093 (N_2093,N_1343,N_1989);
and U2094 (N_2094,N_1472,N_1175);
nor U2095 (N_2095,N_1146,N_1965);
and U2096 (N_2096,N_1347,N_1498);
nand U2097 (N_2097,N_1240,N_1827);
and U2098 (N_2098,N_1947,N_1094);
nor U2099 (N_2099,N_1594,N_1237);
nor U2100 (N_2100,N_1330,N_1127);
and U2101 (N_2101,N_1158,N_1197);
and U2102 (N_2102,N_1770,N_1995);
nor U2103 (N_2103,N_1860,N_1112);
or U2104 (N_2104,N_1675,N_1908);
nand U2105 (N_2105,N_1494,N_1006);
nand U2106 (N_2106,N_1808,N_1300);
nand U2107 (N_2107,N_1428,N_1139);
or U2108 (N_2108,N_1433,N_1342);
and U2109 (N_2109,N_1344,N_1422);
and U2110 (N_2110,N_1312,N_1806);
or U2111 (N_2111,N_1366,N_1839);
nor U2112 (N_2112,N_1306,N_1717);
nor U2113 (N_2113,N_1087,N_1277);
and U2114 (N_2114,N_1211,N_1905);
nor U2115 (N_2115,N_1926,N_1641);
or U2116 (N_2116,N_1939,N_1879);
or U2117 (N_2117,N_1648,N_1192);
nor U2118 (N_2118,N_1359,N_1053);
nor U2119 (N_2119,N_1400,N_1721);
nand U2120 (N_2120,N_1616,N_1658);
nor U2121 (N_2121,N_1239,N_1491);
or U2122 (N_2122,N_1105,N_1195);
nor U2123 (N_2123,N_1584,N_1888);
nor U2124 (N_2124,N_1606,N_1752);
and U2125 (N_2125,N_1223,N_1264);
nand U2126 (N_2126,N_1221,N_1257);
and U2127 (N_2127,N_1360,N_1152);
nor U2128 (N_2128,N_1915,N_1406);
and U2129 (N_2129,N_1274,N_1567);
nand U2130 (N_2130,N_1464,N_1031);
nand U2131 (N_2131,N_1654,N_1976);
and U2132 (N_2132,N_1512,N_1762);
or U2133 (N_2133,N_1145,N_1617);
nand U2134 (N_2134,N_1365,N_1607);
nor U2135 (N_2135,N_1033,N_1758);
or U2136 (N_2136,N_1686,N_1927);
and U2137 (N_2137,N_1896,N_1130);
and U2138 (N_2138,N_1117,N_1307);
nand U2139 (N_2139,N_1624,N_1368);
and U2140 (N_2140,N_1198,N_1518);
nor U2141 (N_2141,N_1352,N_1074);
or U2142 (N_2142,N_1979,N_1413);
or U2143 (N_2143,N_1523,N_1399);
nor U2144 (N_2144,N_1877,N_1496);
and U2145 (N_2145,N_1278,N_1276);
nand U2146 (N_2146,N_1236,N_1166);
nand U2147 (N_2147,N_1181,N_1160);
or U2148 (N_2148,N_1867,N_1077);
nand U2149 (N_2149,N_1010,N_1883);
nor U2150 (N_2150,N_1814,N_1807);
nand U2151 (N_2151,N_1793,N_1533);
or U2152 (N_2152,N_1298,N_1627);
nand U2153 (N_2153,N_1799,N_1955);
nor U2154 (N_2154,N_1305,N_1323);
or U2155 (N_2155,N_1073,N_1706);
and U2156 (N_2156,N_1208,N_1887);
nor U2157 (N_2157,N_1163,N_1059);
and U2158 (N_2158,N_1229,N_1697);
or U2159 (N_2159,N_1735,N_1599);
and U2160 (N_2160,N_1850,N_1171);
nor U2161 (N_2161,N_1602,N_1301);
or U2162 (N_2162,N_1026,N_1870);
nand U2163 (N_2163,N_1959,N_1948);
or U2164 (N_2164,N_1924,N_1765);
and U2165 (N_2165,N_1684,N_1703);
nor U2166 (N_2166,N_1502,N_1499);
and U2167 (N_2167,N_1831,N_1371);
and U2168 (N_2168,N_1763,N_1346);
and U2169 (N_2169,N_1572,N_1190);
nor U2170 (N_2170,N_1093,N_1377);
and U2171 (N_2171,N_1633,N_1787);
nand U2172 (N_2172,N_1248,N_1488);
and U2173 (N_2173,N_1289,N_1644);
or U2174 (N_2174,N_1296,N_1967);
or U2175 (N_2175,N_1390,N_1479);
nor U2176 (N_2176,N_1527,N_1431);
nor U2177 (N_2177,N_1821,N_1243);
or U2178 (N_2178,N_1434,N_1191);
nor U2179 (N_2179,N_1951,N_1509);
and U2180 (N_2180,N_1226,N_1748);
or U2181 (N_2181,N_1313,N_1683);
and U2182 (N_2182,N_1448,N_1830);
and U2183 (N_2183,N_1462,N_1530);
nand U2184 (N_2184,N_1384,N_1964);
nor U2185 (N_2185,N_1515,N_1696);
and U2186 (N_2186,N_1978,N_1836);
and U2187 (N_2187,N_1555,N_1545);
nor U2188 (N_2188,N_1484,N_1984);
or U2189 (N_2189,N_1176,N_1536);
and U2190 (N_2190,N_1437,N_1945);
nor U2191 (N_2191,N_1420,N_1662);
or U2192 (N_2192,N_1705,N_1439);
or U2193 (N_2193,N_1884,N_1841);
nand U2194 (N_2194,N_1710,N_1397);
and U2195 (N_2195,N_1728,N_1631);
and U2196 (N_2196,N_1522,N_1302);
nand U2197 (N_2197,N_1678,N_1156);
nand U2198 (N_2198,N_1564,N_1711);
nor U2199 (N_2199,N_1600,N_1265);
and U2200 (N_2200,N_1900,N_1822);
nor U2201 (N_2201,N_1269,N_1326);
or U2202 (N_2202,N_1856,N_1246);
and U2203 (N_2203,N_1350,N_1120);
or U2204 (N_2204,N_1252,N_1089);
and U2205 (N_2205,N_1051,N_1019);
and U2206 (N_2206,N_1514,N_1147);
or U2207 (N_2207,N_1354,N_1723);
nor U2208 (N_2208,N_1281,N_1932);
nor U2209 (N_2209,N_1385,N_1619);
nand U2210 (N_2210,N_1279,N_1272);
or U2211 (N_2211,N_1471,N_1916);
and U2212 (N_2212,N_1213,N_1940);
or U2213 (N_2213,N_1110,N_1730);
nor U2214 (N_2214,N_1918,N_1048);
or U2215 (N_2215,N_1622,N_1138);
or U2216 (N_2216,N_1885,N_1818);
nor U2217 (N_2217,N_1174,N_1122);
nand U2218 (N_2218,N_1241,N_1108);
nor U2219 (N_2219,N_1579,N_1946);
nor U2220 (N_2220,N_1655,N_1395);
nand U2221 (N_2221,N_1500,N_1524);
and U2222 (N_2222,N_1485,N_1115);
nor U2223 (N_2223,N_1320,N_1574);
nor U2224 (N_2224,N_1370,N_1224);
or U2225 (N_2225,N_1557,N_1376);
nor U2226 (N_2226,N_1991,N_1027);
and U2227 (N_2227,N_1303,N_1651);
nor U2228 (N_2228,N_1427,N_1899);
nand U2229 (N_2229,N_1452,N_1669);
nand U2230 (N_2230,N_1796,N_1653);
and U2231 (N_2231,N_1407,N_1218);
and U2232 (N_2232,N_1656,N_1381);
and U2233 (N_2233,N_1561,N_1327);
nand U2234 (N_2234,N_1538,N_1404);
nor U2235 (N_2235,N_1421,N_1069);
and U2236 (N_2236,N_1032,N_1992);
or U2237 (N_2237,N_1078,N_1054);
nor U2238 (N_2238,N_1040,N_1671);
and U2239 (N_2239,N_1016,N_1340);
nand U2240 (N_2240,N_1249,N_1348);
nand U2241 (N_2241,N_1771,N_1310);
and U2242 (N_2242,N_1903,N_1255);
nor U2243 (N_2243,N_1866,N_1052);
nor U2244 (N_2244,N_1487,N_1933);
nor U2245 (N_2245,N_1980,N_1328);
nand U2246 (N_2246,N_1098,N_1212);
and U2247 (N_2247,N_1461,N_1247);
nor U2248 (N_2248,N_1950,N_1429);
or U2249 (N_2249,N_1425,N_1781);
nor U2250 (N_2250,N_1511,N_1636);
and U2251 (N_2251,N_1949,N_1295);
nor U2252 (N_2252,N_1858,N_1444);
nand U2253 (N_2253,N_1104,N_1936);
or U2254 (N_2254,N_1463,N_1873);
or U2255 (N_2255,N_1699,N_1609);
or U2256 (N_2256,N_1018,N_1125);
nand U2257 (N_2257,N_1123,N_1451);
and U2258 (N_2258,N_1874,N_1418);
nor U2259 (N_2259,N_1096,N_1971);
nand U2260 (N_2260,N_1757,N_1285);
or U2261 (N_2261,N_1772,N_1317);
and U2262 (N_2262,N_1718,N_1826);
or U2263 (N_2263,N_1086,N_1447);
nor U2264 (N_2264,N_1299,N_1741);
and U2265 (N_2265,N_1337,N_1913);
or U2266 (N_2266,N_1440,N_1205);
or U2267 (N_2267,N_1535,N_1562);
nand U2268 (N_2268,N_1100,N_1852);
and U2269 (N_2269,N_1657,N_1977);
nor U2270 (N_2270,N_1405,N_1912);
and U2271 (N_2271,N_1768,N_1907);
nor U2272 (N_2272,N_1460,N_1412);
nand U2273 (N_2273,N_1286,N_1990);
or U2274 (N_2274,N_1063,N_1701);
or U2275 (N_2275,N_1154,N_1612);
or U2276 (N_2276,N_1469,N_1004);
or U2277 (N_2277,N_1441,N_1754);
or U2278 (N_2278,N_1369,N_1639);
nand U2279 (N_2279,N_1151,N_1708);
or U2280 (N_2280,N_1349,N_1880);
nor U2281 (N_2281,N_1805,N_1064);
nor U2282 (N_2282,N_1972,N_1966);
or U2283 (N_2283,N_1941,N_1811);
nor U2284 (N_2284,N_1290,N_1103);
and U2285 (N_2285,N_1914,N_1646);
and U2286 (N_2286,N_1975,N_1953);
or U2287 (N_2287,N_1829,N_1393);
and U2288 (N_2288,N_1598,N_1416);
and U2289 (N_2289,N_1034,N_1732);
and U2290 (N_2290,N_1872,N_1414);
nand U2291 (N_2291,N_1119,N_1593);
or U2292 (N_2292,N_1801,N_1563);
nor U2293 (N_2293,N_1336,N_1537);
nor U2294 (N_2294,N_1996,N_1573);
nand U2295 (N_2295,N_1645,N_1519);
and U2296 (N_2296,N_1245,N_1126);
or U2297 (N_2297,N_1148,N_1315);
or U2298 (N_2298,N_1997,N_1042);
nand U2299 (N_2299,N_1201,N_1659);
or U2300 (N_2300,N_1525,N_1743);
and U2301 (N_2301,N_1605,N_1037);
nor U2302 (N_2302,N_1209,N_1324);
nand U2303 (N_2303,N_1570,N_1426);
and U2304 (N_2304,N_1634,N_1118);
or U2305 (N_2305,N_1812,N_1892);
nor U2306 (N_2306,N_1140,N_1024);
or U2307 (N_2307,N_1398,N_1338);
and U2308 (N_2308,N_1611,N_1193);
nor U2309 (N_2309,N_1109,N_1581);
nor U2310 (N_2310,N_1041,N_1981);
nand U2311 (N_2311,N_1454,N_1047);
and U2312 (N_2312,N_1745,N_1846);
nor U2313 (N_2313,N_1954,N_1432);
and U2314 (N_2314,N_1601,N_1679);
and U2315 (N_2315,N_1157,N_1876);
or U2316 (N_2316,N_1832,N_1539);
nor U2317 (N_2317,N_1481,N_1007);
nor U2318 (N_2318,N_1797,N_1789);
nor U2319 (N_2319,N_1005,N_1435);
nor U2320 (N_2320,N_1056,N_1825);
nor U2321 (N_2321,N_1838,N_1736);
or U2322 (N_2322,N_1604,N_1911);
and U2323 (N_2323,N_1470,N_1844);
and U2324 (N_2324,N_1786,N_1379);
or U2325 (N_2325,N_1647,N_1389);
nand U2326 (N_2326,N_1944,N_1459);
and U2327 (N_2327,N_1516,N_1544);
nand U2328 (N_2328,N_1552,N_1691);
nand U2329 (N_2329,N_1476,N_1687);
nor U2330 (N_2330,N_1132,N_1116);
and U2331 (N_2331,N_1057,N_1963);
and U2332 (N_2332,N_1586,N_1629);
nor U2333 (N_2333,N_1853,N_1630);
and U2334 (N_2334,N_1689,N_1834);
or U2335 (N_2335,N_1036,N_1288);
and U2336 (N_2336,N_1961,N_1766);
and U2337 (N_2337,N_1597,N_1474);
nor U2338 (N_2338,N_1273,N_1080);
or U2339 (N_2339,N_1682,N_1066);
nand U2340 (N_2340,N_1415,N_1373);
nand U2341 (N_2341,N_1886,N_1704);
nor U2342 (N_2342,N_1942,N_1693);
and U2343 (N_2343,N_1250,N_1380);
nand U2344 (N_2344,N_1777,N_1331);
or U2345 (N_2345,N_1590,N_1578);
and U2346 (N_2346,N_1185,N_1922);
nand U2347 (N_2347,N_1661,N_1660);
nand U2348 (N_2348,N_1131,N_1702);
nor U2349 (N_2349,N_1206,N_1232);
or U2350 (N_2350,N_1183,N_1782);
or U2351 (N_2351,N_1928,N_1321);
and U2352 (N_2352,N_1165,N_1039);
nor U2353 (N_2353,N_1958,N_1694);
or U2354 (N_2354,N_1828,N_1013);
and U2355 (N_2355,N_1161,N_1960);
or U2356 (N_2356,N_1260,N_1550);
nand U2357 (N_2357,N_1374,N_1155);
nor U2358 (N_2358,N_1784,N_1517);
nor U2359 (N_2359,N_1970,N_1795);
and U2360 (N_2360,N_1878,N_1023);
and U2361 (N_2361,N_1378,N_1178);
nor U2362 (N_2362,N_1635,N_1196);
and U2363 (N_2363,N_1677,N_1144);
and U2364 (N_2364,N_1199,N_1553);
or U2365 (N_2365,N_1466,N_1334);
nor U2366 (N_2366,N_1890,N_1097);
nand U2367 (N_2367,N_1521,N_1583);
nor U2368 (N_2368,N_1297,N_1219);
nor U2369 (N_2369,N_1803,N_1455);
or U2370 (N_2370,N_1325,N_1529);
nand U2371 (N_2371,N_1314,N_1242);
nand U2372 (N_2372,N_1136,N_1753);
and U2373 (N_2373,N_1727,N_1847);
and U2374 (N_2374,N_1864,N_1707);
nor U2375 (N_2375,N_1442,N_1480);
or U2376 (N_2376,N_1001,N_1383);
and U2377 (N_2377,N_1180,N_1294);
nor U2378 (N_2378,N_1225,N_1608);
nor U2379 (N_2379,N_1142,N_1084);
nand U2380 (N_2380,N_1501,N_1382);
nand U2381 (N_2381,N_1668,N_1800);
nor U2382 (N_2382,N_1930,N_1603);
and U2383 (N_2383,N_1724,N_1931);
or U2384 (N_2384,N_1092,N_1050);
nor U2385 (N_2385,N_1450,N_1804);
nand U2386 (N_2386,N_1489,N_1210);
nor U2387 (N_2387,N_1810,N_1823);
and U2388 (N_2388,N_1403,N_1251);
nor U2389 (N_2389,N_1082,N_1934);
or U2390 (N_2390,N_1419,N_1587);
nor U2391 (N_2391,N_1367,N_1438);
and U2392 (N_2392,N_1028,N_1576);
nor U2393 (N_2393,N_1000,N_1588);
nand U2394 (N_2394,N_1769,N_1280);
and U2395 (N_2395,N_1731,N_1134);
nand U2396 (N_2396,N_1170,N_1559);
and U2397 (N_2397,N_1952,N_1575);
nand U2398 (N_2398,N_1060,N_1571);
nor U2399 (N_2399,N_1012,N_1667);
nor U2400 (N_2400,N_1095,N_1284);
or U2401 (N_2401,N_1540,N_1254);
nor U2402 (N_2402,N_1124,N_1402);
nand U2403 (N_2403,N_1714,N_1643);
and U2404 (N_2404,N_1003,N_1316);
nand U2405 (N_2405,N_1065,N_1937);
nand U2406 (N_2406,N_1083,N_1351);
nor U2407 (N_2407,N_1921,N_1534);
and U2408 (N_2408,N_1030,N_1585);
and U2409 (N_2409,N_1046,N_1672);
nor U2410 (N_2410,N_1688,N_1809);
or U2411 (N_2411,N_1613,N_1759);
or U2412 (N_2412,N_1760,N_1207);
or U2413 (N_2413,N_1938,N_1002);
and U2414 (N_2414,N_1833,N_1128);
nand U2415 (N_2415,N_1982,N_1773);
nand U2416 (N_2416,N_1079,N_1445);
xnor U2417 (N_2417,N_1638,N_1135);
or U2418 (N_2418,N_1716,N_1780);
and U2419 (N_2419,N_1738,N_1478);
and U2420 (N_2420,N_1072,N_1133);
nand U2421 (N_2421,N_1580,N_1709);
nand U2422 (N_2422,N_1652,N_1626);
or U2423 (N_2423,N_1943,N_1820);
nor U2424 (N_2424,N_1067,N_1258);
and U2425 (N_2425,N_1394,N_1994);
nor U2426 (N_2426,N_1490,N_1513);
or U2427 (N_2427,N_1233,N_1749);
or U2428 (N_2428,N_1121,N_1364);
xnor U2429 (N_2429,N_1088,N_1568);
nor U2430 (N_2430,N_1477,N_1798);
or U2431 (N_2431,N_1898,N_1015);
nand U2432 (N_2432,N_1869,N_1595);
and U2433 (N_2433,N_1726,N_1055);
or U2434 (N_2434,N_1506,N_1238);
and U2435 (N_2435,N_1341,N_1268);
nor U2436 (N_2436,N_1038,N_1871);
nor U2437 (N_2437,N_1507,N_1102);
and U2438 (N_2438,N_1901,N_1902);
nor U2439 (N_2439,N_1253,N_1889);
and U2440 (N_2440,N_1755,N_1532);
nor U2441 (N_2441,N_1740,N_1802);
nor U2442 (N_2442,N_1560,N_1090);
nor U2443 (N_2443,N_1546,N_1548);
nor U2444 (N_2444,N_1663,N_1167);
and U2445 (N_2445,N_1582,N_1909);
and U2446 (N_2446,N_1625,N_1637);
or U2447 (N_2447,N_1021,N_1356);
and U2448 (N_2448,N_1332,N_1692);
nor U2449 (N_2449,N_1283,N_1775);
nor U2450 (N_2450,N_1456,N_1551);
or U2451 (N_2451,N_1680,N_1558);
and U2452 (N_2452,N_1204,N_1904);
nand U2453 (N_2453,N_1443,N_1070);
nor U2454 (N_2454,N_1304,N_1863);
nand U2455 (N_2455,N_1345,N_1355);
nor U2456 (N_2456,N_1235,N_1614);
nor U2457 (N_2457,N_1974,N_1159);
and U2458 (N_2458,N_1815,N_1713);
or U2459 (N_2459,N_1729,N_1259);
nand U2460 (N_2460,N_1101,N_1923);
or U2461 (N_2461,N_1009,N_1875);
or U2462 (N_2462,N_1895,N_1695);
nor U2463 (N_2463,N_1817,N_1473);
or U2464 (N_2464,N_1855,N_1774);
nor U2465 (N_2465,N_1362,N_1282);
and U2466 (N_2466,N_1186,N_1465);
or U2467 (N_2467,N_1168,N_1776);
and U2468 (N_2468,N_1664,N_1177);
nor U2469 (N_2469,N_1227,N_1164);
or U2470 (N_2470,N_1149,N_1788);
nand U2471 (N_2471,N_1230,N_1526);
nor U2472 (N_2472,N_1319,N_1987);
and U2473 (N_2473,N_1744,N_1392);
or U2474 (N_2474,N_1840,N_1508);
nor U2475 (N_2475,N_1541,N_1897);
xnor U2476 (N_2476,N_1681,N_1216);
nor U2477 (N_2477,N_1387,N_1375);
xor U2478 (N_2478,N_1467,N_1742);
nand U2479 (N_2479,N_1882,N_1215);
nand U2480 (N_2480,N_1791,N_1666);
and U2481 (N_2481,N_1813,N_1231);
nand U2482 (N_2482,N_1792,N_1700);
nor U2483 (N_2483,N_1620,N_1153);
nor U2484 (N_2484,N_1993,N_1045);
or U2485 (N_2485,N_1722,N_1172);
nor U2486 (N_2486,N_1917,N_1008);
or U2487 (N_2487,N_1746,N_1973);
and U2488 (N_2488,N_1510,N_1085);
and U2489 (N_2489,N_1767,N_1690);
nand U2490 (N_2490,N_1267,N_1610);
and U2491 (N_2491,N_1292,N_1222);
or U2492 (N_2492,N_1194,N_1262);
nor U2493 (N_2493,N_1968,N_1449);
nand U2494 (N_2494,N_1640,N_1842);
xnor U2495 (N_2495,N_1408,N_1565);
nor U2496 (N_2496,N_1621,N_1848);
nand U2497 (N_2497,N_1396,N_1189);
and U2498 (N_2498,N_1549,N_1649);
and U2499 (N_2499,N_1676,N_1068);
or U2500 (N_2500,N_1888,N_1841);
and U2501 (N_2501,N_1285,N_1491);
and U2502 (N_2502,N_1397,N_1823);
nor U2503 (N_2503,N_1316,N_1033);
nand U2504 (N_2504,N_1675,N_1258);
and U2505 (N_2505,N_1158,N_1331);
and U2506 (N_2506,N_1895,N_1643);
or U2507 (N_2507,N_1871,N_1730);
and U2508 (N_2508,N_1657,N_1444);
or U2509 (N_2509,N_1100,N_1455);
nor U2510 (N_2510,N_1388,N_1545);
nor U2511 (N_2511,N_1642,N_1567);
nand U2512 (N_2512,N_1616,N_1432);
or U2513 (N_2513,N_1057,N_1815);
nor U2514 (N_2514,N_1667,N_1399);
and U2515 (N_2515,N_1352,N_1525);
nand U2516 (N_2516,N_1207,N_1753);
and U2517 (N_2517,N_1502,N_1665);
or U2518 (N_2518,N_1309,N_1988);
and U2519 (N_2519,N_1109,N_1640);
nand U2520 (N_2520,N_1320,N_1820);
nand U2521 (N_2521,N_1749,N_1444);
nor U2522 (N_2522,N_1953,N_1764);
or U2523 (N_2523,N_1870,N_1655);
or U2524 (N_2524,N_1550,N_1027);
or U2525 (N_2525,N_1724,N_1506);
or U2526 (N_2526,N_1407,N_1705);
nor U2527 (N_2527,N_1589,N_1935);
nor U2528 (N_2528,N_1299,N_1996);
or U2529 (N_2529,N_1661,N_1134);
nor U2530 (N_2530,N_1904,N_1745);
or U2531 (N_2531,N_1635,N_1413);
and U2532 (N_2532,N_1539,N_1621);
nor U2533 (N_2533,N_1190,N_1012);
nor U2534 (N_2534,N_1049,N_1769);
or U2535 (N_2535,N_1427,N_1215);
nand U2536 (N_2536,N_1446,N_1030);
nand U2537 (N_2537,N_1391,N_1722);
nor U2538 (N_2538,N_1793,N_1491);
nor U2539 (N_2539,N_1967,N_1911);
or U2540 (N_2540,N_1161,N_1269);
and U2541 (N_2541,N_1141,N_1905);
or U2542 (N_2542,N_1253,N_1849);
and U2543 (N_2543,N_1480,N_1758);
nand U2544 (N_2544,N_1414,N_1549);
nor U2545 (N_2545,N_1967,N_1620);
nor U2546 (N_2546,N_1421,N_1256);
and U2547 (N_2547,N_1593,N_1385);
and U2548 (N_2548,N_1265,N_1931);
or U2549 (N_2549,N_1609,N_1114);
or U2550 (N_2550,N_1073,N_1113);
nor U2551 (N_2551,N_1252,N_1372);
and U2552 (N_2552,N_1570,N_1060);
and U2553 (N_2553,N_1202,N_1606);
and U2554 (N_2554,N_1754,N_1230);
or U2555 (N_2555,N_1879,N_1022);
nand U2556 (N_2556,N_1438,N_1574);
nor U2557 (N_2557,N_1296,N_1748);
or U2558 (N_2558,N_1934,N_1749);
and U2559 (N_2559,N_1397,N_1514);
and U2560 (N_2560,N_1178,N_1552);
nor U2561 (N_2561,N_1674,N_1539);
or U2562 (N_2562,N_1644,N_1123);
nand U2563 (N_2563,N_1587,N_1141);
nor U2564 (N_2564,N_1602,N_1903);
nand U2565 (N_2565,N_1121,N_1329);
and U2566 (N_2566,N_1952,N_1934);
and U2567 (N_2567,N_1344,N_1268);
and U2568 (N_2568,N_1005,N_1825);
xnor U2569 (N_2569,N_1936,N_1989);
nor U2570 (N_2570,N_1469,N_1250);
nor U2571 (N_2571,N_1308,N_1296);
or U2572 (N_2572,N_1986,N_1607);
and U2573 (N_2573,N_1180,N_1604);
and U2574 (N_2574,N_1634,N_1307);
and U2575 (N_2575,N_1515,N_1103);
nand U2576 (N_2576,N_1572,N_1387);
and U2577 (N_2577,N_1689,N_1831);
nand U2578 (N_2578,N_1432,N_1738);
nand U2579 (N_2579,N_1743,N_1238);
and U2580 (N_2580,N_1805,N_1418);
and U2581 (N_2581,N_1661,N_1962);
nor U2582 (N_2582,N_1612,N_1409);
and U2583 (N_2583,N_1674,N_1054);
nand U2584 (N_2584,N_1355,N_1425);
nand U2585 (N_2585,N_1685,N_1611);
and U2586 (N_2586,N_1673,N_1916);
nand U2587 (N_2587,N_1084,N_1259);
or U2588 (N_2588,N_1953,N_1205);
nand U2589 (N_2589,N_1371,N_1080);
nor U2590 (N_2590,N_1472,N_1781);
and U2591 (N_2591,N_1622,N_1943);
nor U2592 (N_2592,N_1521,N_1168);
nor U2593 (N_2593,N_1650,N_1838);
nand U2594 (N_2594,N_1579,N_1803);
or U2595 (N_2595,N_1657,N_1260);
or U2596 (N_2596,N_1602,N_1630);
nand U2597 (N_2597,N_1530,N_1629);
and U2598 (N_2598,N_1548,N_1542);
nand U2599 (N_2599,N_1476,N_1784);
or U2600 (N_2600,N_1016,N_1045);
nor U2601 (N_2601,N_1826,N_1873);
nor U2602 (N_2602,N_1156,N_1762);
or U2603 (N_2603,N_1055,N_1638);
nor U2604 (N_2604,N_1312,N_1076);
nor U2605 (N_2605,N_1904,N_1886);
and U2606 (N_2606,N_1926,N_1081);
and U2607 (N_2607,N_1276,N_1168);
nand U2608 (N_2608,N_1560,N_1786);
and U2609 (N_2609,N_1337,N_1129);
or U2610 (N_2610,N_1533,N_1943);
nor U2611 (N_2611,N_1945,N_1266);
or U2612 (N_2612,N_1232,N_1333);
and U2613 (N_2613,N_1953,N_1000);
and U2614 (N_2614,N_1844,N_1375);
and U2615 (N_2615,N_1235,N_1582);
nand U2616 (N_2616,N_1311,N_1231);
or U2617 (N_2617,N_1175,N_1442);
nor U2618 (N_2618,N_1594,N_1850);
nand U2619 (N_2619,N_1658,N_1721);
nor U2620 (N_2620,N_1834,N_1526);
nor U2621 (N_2621,N_1668,N_1976);
nor U2622 (N_2622,N_1181,N_1210);
nor U2623 (N_2623,N_1816,N_1957);
nand U2624 (N_2624,N_1063,N_1058);
or U2625 (N_2625,N_1389,N_1083);
nor U2626 (N_2626,N_1131,N_1217);
nor U2627 (N_2627,N_1046,N_1632);
and U2628 (N_2628,N_1356,N_1726);
nand U2629 (N_2629,N_1008,N_1936);
and U2630 (N_2630,N_1023,N_1108);
nor U2631 (N_2631,N_1180,N_1319);
nand U2632 (N_2632,N_1486,N_1749);
or U2633 (N_2633,N_1790,N_1709);
nor U2634 (N_2634,N_1205,N_1319);
and U2635 (N_2635,N_1481,N_1347);
nand U2636 (N_2636,N_1362,N_1327);
nor U2637 (N_2637,N_1016,N_1697);
nor U2638 (N_2638,N_1524,N_1650);
nand U2639 (N_2639,N_1217,N_1469);
nor U2640 (N_2640,N_1548,N_1678);
or U2641 (N_2641,N_1440,N_1907);
nand U2642 (N_2642,N_1575,N_1383);
nand U2643 (N_2643,N_1543,N_1072);
nand U2644 (N_2644,N_1541,N_1543);
and U2645 (N_2645,N_1669,N_1874);
and U2646 (N_2646,N_1445,N_1898);
nand U2647 (N_2647,N_1836,N_1983);
and U2648 (N_2648,N_1948,N_1760);
and U2649 (N_2649,N_1758,N_1986);
nor U2650 (N_2650,N_1556,N_1988);
and U2651 (N_2651,N_1477,N_1422);
and U2652 (N_2652,N_1017,N_1000);
or U2653 (N_2653,N_1873,N_1899);
nand U2654 (N_2654,N_1710,N_1602);
nor U2655 (N_2655,N_1709,N_1886);
and U2656 (N_2656,N_1372,N_1812);
nor U2657 (N_2657,N_1960,N_1030);
or U2658 (N_2658,N_1597,N_1049);
nand U2659 (N_2659,N_1000,N_1492);
or U2660 (N_2660,N_1553,N_1890);
nand U2661 (N_2661,N_1843,N_1397);
or U2662 (N_2662,N_1556,N_1827);
or U2663 (N_2663,N_1318,N_1324);
and U2664 (N_2664,N_1730,N_1193);
and U2665 (N_2665,N_1002,N_1350);
and U2666 (N_2666,N_1454,N_1282);
or U2667 (N_2667,N_1468,N_1989);
or U2668 (N_2668,N_1323,N_1746);
or U2669 (N_2669,N_1182,N_1337);
or U2670 (N_2670,N_1877,N_1586);
and U2671 (N_2671,N_1189,N_1432);
or U2672 (N_2672,N_1853,N_1305);
and U2673 (N_2673,N_1331,N_1748);
nand U2674 (N_2674,N_1399,N_1175);
nand U2675 (N_2675,N_1322,N_1144);
xnor U2676 (N_2676,N_1050,N_1559);
and U2677 (N_2677,N_1357,N_1651);
or U2678 (N_2678,N_1409,N_1450);
nand U2679 (N_2679,N_1579,N_1045);
or U2680 (N_2680,N_1742,N_1356);
and U2681 (N_2681,N_1416,N_1126);
nor U2682 (N_2682,N_1070,N_1544);
and U2683 (N_2683,N_1610,N_1133);
and U2684 (N_2684,N_1249,N_1170);
nor U2685 (N_2685,N_1513,N_1758);
nand U2686 (N_2686,N_1133,N_1792);
nor U2687 (N_2687,N_1504,N_1818);
nor U2688 (N_2688,N_1168,N_1200);
and U2689 (N_2689,N_1748,N_1676);
or U2690 (N_2690,N_1163,N_1402);
or U2691 (N_2691,N_1631,N_1579);
or U2692 (N_2692,N_1045,N_1138);
nand U2693 (N_2693,N_1318,N_1770);
or U2694 (N_2694,N_1222,N_1892);
or U2695 (N_2695,N_1279,N_1772);
nand U2696 (N_2696,N_1920,N_1819);
nor U2697 (N_2697,N_1041,N_1016);
nor U2698 (N_2698,N_1589,N_1948);
and U2699 (N_2699,N_1059,N_1501);
nor U2700 (N_2700,N_1129,N_1924);
and U2701 (N_2701,N_1571,N_1801);
or U2702 (N_2702,N_1560,N_1101);
or U2703 (N_2703,N_1688,N_1661);
nor U2704 (N_2704,N_1416,N_1714);
nor U2705 (N_2705,N_1890,N_1625);
nor U2706 (N_2706,N_1548,N_1283);
nor U2707 (N_2707,N_1927,N_1285);
nor U2708 (N_2708,N_1441,N_1473);
and U2709 (N_2709,N_1217,N_1788);
nand U2710 (N_2710,N_1205,N_1968);
nor U2711 (N_2711,N_1646,N_1426);
nand U2712 (N_2712,N_1315,N_1170);
nand U2713 (N_2713,N_1731,N_1090);
nand U2714 (N_2714,N_1599,N_1474);
nor U2715 (N_2715,N_1621,N_1323);
nor U2716 (N_2716,N_1586,N_1262);
nand U2717 (N_2717,N_1985,N_1261);
nand U2718 (N_2718,N_1200,N_1512);
nand U2719 (N_2719,N_1064,N_1479);
and U2720 (N_2720,N_1564,N_1175);
nor U2721 (N_2721,N_1904,N_1939);
nor U2722 (N_2722,N_1209,N_1957);
or U2723 (N_2723,N_1732,N_1737);
nor U2724 (N_2724,N_1718,N_1603);
or U2725 (N_2725,N_1256,N_1156);
or U2726 (N_2726,N_1490,N_1001);
or U2727 (N_2727,N_1277,N_1565);
nor U2728 (N_2728,N_1585,N_1839);
nand U2729 (N_2729,N_1999,N_1388);
nand U2730 (N_2730,N_1475,N_1281);
and U2731 (N_2731,N_1805,N_1200);
nand U2732 (N_2732,N_1957,N_1807);
nor U2733 (N_2733,N_1824,N_1916);
nor U2734 (N_2734,N_1263,N_1267);
or U2735 (N_2735,N_1659,N_1047);
and U2736 (N_2736,N_1050,N_1492);
or U2737 (N_2737,N_1612,N_1796);
and U2738 (N_2738,N_1015,N_1312);
and U2739 (N_2739,N_1415,N_1571);
and U2740 (N_2740,N_1347,N_1920);
or U2741 (N_2741,N_1835,N_1470);
nand U2742 (N_2742,N_1137,N_1738);
and U2743 (N_2743,N_1670,N_1393);
nand U2744 (N_2744,N_1584,N_1901);
or U2745 (N_2745,N_1176,N_1608);
nor U2746 (N_2746,N_1439,N_1005);
or U2747 (N_2747,N_1854,N_1979);
and U2748 (N_2748,N_1444,N_1693);
or U2749 (N_2749,N_1222,N_1761);
or U2750 (N_2750,N_1267,N_1327);
or U2751 (N_2751,N_1617,N_1858);
nand U2752 (N_2752,N_1453,N_1204);
nand U2753 (N_2753,N_1245,N_1317);
nand U2754 (N_2754,N_1447,N_1688);
nand U2755 (N_2755,N_1760,N_1975);
nand U2756 (N_2756,N_1255,N_1091);
nand U2757 (N_2757,N_1538,N_1374);
nor U2758 (N_2758,N_1783,N_1905);
and U2759 (N_2759,N_1087,N_1359);
or U2760 (N_2760,N_1900,N_1605);
nand U2761 (N_2761,N_1422,N_1122);
nand U2762 (N_2762,N_1914,N_1884);
and U2763 (N_2763,N_1441,N_1997);
nor U2764 (N_2764,N_1625,N_1316);
or U2765 (N_2765,N_1547,N_1339);
and U2766 (N_2766,N_1022,N_1394);
nand U2767 (N_2767,N_1822,N_1865);
nor U2768 (N_2768,N_1189,N_1904);
or U2769 (N_2769,N_1072,N_1793);
nand U2770 (N_2770,N_1696,N_1265);
xor U2771 (N_2771,N_1791,N_1423);
nor U2772 (N_2772,N_1526,N_1414);
or U2773 (N_2773,N_1048,N_1720);
or U2774 (N_2774,N_1307,N_1493);
nor U2775 (N_2775,N_1916,N_1935);
and U2776 (N_2776,N_1046,N_1584);
nor U2777 (N_2777,N_1175,N_1071);
and U2778 (N_2778,N_1176,N_1123);
or U2779 (N_2779,N_1348,N_1375);
and U2780 (N_2780,N_1132,N_1060);
nand U2781 (N_2781,N_1549,N_1535);
and U2782 (N_2782,N_1550,N_1540);
xnor U2783 (N_2783,N_1100,N_1388);
or U2784 (N_2784,N_1486,N_1038);
nor U2785 (N_2785,N_1009,N_1076);
nand U2786 (N_2786,N_1358,N_1204);
or U2787 (N_2787,N_1828,N_1880);
and U2788 (N_2788,N_1281,N_1433);
and U2789 (N_2789,N_1193,N_1871);
nor U2790 (N_2790,N_1727,N_1528);
nor U2791 (N_2791,N_1267,N_1289);
nand U2792 (N_2792,N_1085,N_1011);
or U2793 (N_2793,N_1611,N_1726);
and U2794 (N_2794,N_1788,N_1873);
nand U2795 (N_2795,N_1945,N_1436);
nor U2796 (N_2796,N_1569,N_1492);
and U2797 (N_2797,N_1460,N_1856);
nand U2798 (N_2798,N_1545,N_1548);
and U2799 (N_2799,N_1363,N_1213);
or U2800 (N_2800,N_1668,N_1682);
nand U2801 (N_2801,N_1108,N_1608);
nand U2802 (N_2802,N_1659,N_1861);
nand U2803 (N_2803,N_1144,N_1365);
nand U2804 (N_2804,N_1185,N_1773);
and U2805 (N_2805,N_1189,N_1699);
nand U2806 (N_2806,N_1389,N_1064);
or U2807 (N_2807,N_1435,N_1618);
or U2808 (N_2808,N_1638,N_1870);
nor U2809 (N_2809,N_1343,N_1168);
and U2810 (N_2810,N_1361,N_1700);
nor U2811 (N_2811,N_1493,N_1886);
nand U2812 (N_2812,N_1852,N_1340);
or U2813 (N_2813,N_1099,N_1867);
or U2814 (N_2814,N_1346,N_1544);
nor U2815 (N_2815,N_1373,N_1475);
and U2816 (N_2816,N_1628,N_1407);
nor U2817 (N_2817,N_1119,N_1026);
nand U2818 (N_2818,N_1571,N_1881);
nand U2819 (N_2819,N_1438,N_1460);
nor U2820 (N_2820,N_1681,N_1352);
xnor U2821 (N_2821,N_1781,N_1111);
nand U2822 (N_2822,N_1531,N_1424);
nand U2823 (N_2823,N_1059,N_1096);
xnor U2824 (N_2824,N_1136,N_1287);
nand U2825 (N_2825,N_1969,N_1193);
nand U2826 (N_2826,N_1323,N_1716);
nand U2827 (N_2827,N_1205,N_1713);
and U2828 (N_2828,N_1892,N_1786);
nor U2829 (N_2829,N_1936,N_1244);
and U2830 (N_2830,N_1199,N_1613);
nor U2831 (N_2831,N_1085,N_1017);
nand U2832 (N_2832,N_1622,N_1853);
or U2833 (N_2833,N_1763,N_1143);
nor U2834 (N_2834,N_1053,N_1796);
and U2835 (N_2835,N_1789,N_1428);
xnor U2836 (N_2836,N_1580,N_1734);
nand U2837 (N_2837,N_1033,N_1859);
nor U2838 (N_2838,N_1998,N_1889);
or U2839 (N_2839,N_1994,N_1697);
and U2840 (N_2840,N_1827,N_1114);
or U2841 (N_2841,N_1858,N_1140);
and U2842 (N_2842,N_1760,N_1199);
and U2843 (N_2843,N_1732,N_1166);
and U2844 (N_2844,N_1848,N_1953);
nor U2845 (N_2845,N_1339,N_1174);
nor U2846 (N_2846,N_1192,N_1128);
and U2847 (N_2847,N_1140,N_1715);
nand U2848 (N_2848,N_1409,N_1974);
and U2849 (N_2849,N_1186,N_1904);
or U2850 (N_2850,N_1987,N_1012);
nand U2851 (N_2851,N_1128,N_1079);
nand U2852 (N_2852,N_1654,N_1358);
nor U2853 (N_2853,N_1607,N_1430);
and U2854 (N_2854,N_1520,N_1248);
or U2855 (N_2855,N_1306,N_1883);
nor U2856 (N_2856,N_1280,N_1294);
nand U2857 (N_2857,N_1247,N_1469);
or U2858 (N_2858,N_1019,N_1979);
nor U2859 (N_2859,N_1924,N_1998);
nor U2860 (N_2860,N_1313,N_1831);
nor U2861 (N_2861,N_1594,N_1557);
nand U2862 (N_2862,N_1816,N_1901);
nor U2863 (N_2863,N_1760,N_1444);
nand U2864 (N_2864,N_1955,N_1998);
nor U2865 (N_2865,N_1439,N_1642);
nand U2866 (N_2866,N_1222,N_1661);
and U2867 (N_2867,N_1797,N_1574);
nor U2868 (N_2868,N_1566,N_1004);
nand U2869 (N_2869,N_1306,N_1305);
nor U2870 (N_2870,N_1098,N_1203);
or U2871 (N_2871,N_1469,N_1483);
or U2872 (N_2872,N_1667,N_1756);
or U2873 (N_2873,N_1195,N_1890);
and U2874 (N_2874,N_1737,N_1052);
nand U2875 (N_2875,N_1458,N_1025);
and U2876 (N_2876,N_1393,N_1231);
nand U2877 (N_2877,N_1104,N_1021);
nor U2878 (N_2878,N_1213,N_1199);
nand U2879 (N_2879,N_1571,N_1763);
nor U2880 (N_2880,N_1129,N_1486);
or U2881 (N_2881,N_1577,N_1831);
or U2882 (N_2882,N_1824,N_1208);
and U2883 (N_2883,N_1317,N_1876);
or U2884 (N_2884,N_1489,N_1442);
or U2885 (N_2885,N_1846,N_1603);
nor U2886 (N_2886,N_1582,N_1257);
and U2887 (N_2887,N_1499,N_1071);
nand U2888 (N_2888,N_1735,N_1381);
xnor U2889 (N_2889,N_1181,N_1859);
and U2890 (N_2890,N_1202,N_1330);
nor U2891 (N_2891,N_1375,N_1228);
nand U2892 (N_2892,N_1010,N_1861);
nand U2893 (N_2893,N_1659,N_1944);
xor U2894 (N_2894,N_1387,N_1784);
nor U2895 (N_2895,N_1459,N_1434);
or U2896 (N_2896,N_1325,N_1629);
or U2897 (N_2897,N_1925,N_1090);
and U2898 (N_2898,N_1696,N_1560);
or U2899 (N_2899,N_1985,N_1621);
nand U2900 (N_2900,N_1038,N_1071);
nand U2901 (N_2901,N_1894,N_1988);
nand U2902 (N_2902,N_1610,N_1782);
nand U2903 (N_2903,N_1902,N_1265);
nor U2904 (N_2904,N_1874,N_1622);
nor U2905 (N_2905,N_1992,N_1887);
and U2906 (N_2906,N_1113,N_1287);
nand U2907 (N_2907,N_1149,N_1303);
nor U2908 (N_2908,N_1044,N_1527);
and U2909 (N_2909,N_1142,N_1324);
or U2910 (N_2910,N_1349,N_1163);
or U2911 (N_2911,N_1267,N_1342);
and U2912 (N_2912,N_1406,N_1936);
or U2913 (N_2913,N_1896,N_1355);
nor U2914 (N_2914,N_1297,N_1893);
nor U2915 (N_2915,N_1770,N_1507);
nor U2916 (N_2916,N_1643,N_1629);
and U2917 (N_2917,N_1534,N_1004);
or U2918 (N_2918,N_1413,N_1010);
nor U2919 (N_2919,N_1498,N_1977);
and U2920 (N_2920,N_1325,N_1802);
or U2921 (N_2921,N_1490,N_1882);
nand U2922 (N_2922,N_1972,N_1786);
or U2923 (N_2923,N_1826,N_1844);
nand U2924 (N_2924,N_1217,N_1477);
nor U2925 (N_2925,N_1747,N_1563);
and U2926 (N_2926,N_1831,N_1743);
nor U2927 (N_2927,N_1291,N_1615);
nand U2928 (N_2928,N_1324,N_1366);
nor U2929 (N_2929,N_1584,N_1763);
nand U2930 (N_2930,N_1625,N_1779);
nor U2931 (N_2931,N_1184,N_1987);
nor U2932 (N_2932,N_1071,N_1502);
or U2933 (N_2933,N_1987,N_1336);
or U2934 (N_2934,N_1985,N_1054);
and U2935 (N_2935,N_1756,N_1243);
nand U2936 (N_2936,N_1985,N_1473);
nand U2937 (N_2937,N_1989,N_1417);
nand U2938 (N_2938,N_1716,N_1993);
xnor U2939 (N_2939,N_1609,N_1749);
or U2940 (N_2940,N_1582,N_1507);
and U2941 (N_2941,N_1583,N_1750);
nand U2942 (N_2942,N_1498,N_1552);
or U2943 (N_2943,N_1707,N_1516);
nand U2944 (N_2944,N_1840,N_1965);
or U2945 (N_2945,N_1284,N_1031);
and U2946 (N_2946,N_1852,N_1327);
or U2947 (N_2947,N_1019,N_1720);
nand U2948 (N_2948,N_1630,N_1060);
xnor U2949 (N_2949,N_1739,N_1458);
nand U2950 (N_2950,N_1102,N_1823);
or U2951 (N_2951,N_1571,N_1437);
xnor U2952 (N_2952,N_1702,N_1629);
and U2953 (N_2953,N_1007,N_1614);
nor U2954 (N_2954,N_1665,N_1944);
and U2955 (N_2955,N_1849,N_1132);
and U2956 (N_2956,N_1338,N_1826);
and U2957 (N_2957,N_1106,N_1749);
nor U2958 (N_2958,N_1955,N_1440);
nor U2959 (N_2959,N_1279,N_1830);
nor U2960 (N_2960,N_1046,N_1124);
nor U2961 (N_2961,N_1928,N_1440);
or U2962 (N_2962,N_1172,N_1278);
nor U2963 (N_2963,N_1797,N_1069);
nor U2964 (N_2964,N_1075,N_1260);
or U2965 (N_2965,N_1775,N_1205);
and U2966 (N_2966,N_1527,N_1530);
nor U2967 (N_2967,N_1947,N_1245);
nor U2968 (N_2968,N_1754,N_1665);
or U2969 (N_2969,N_1019,N_1065);
and U2970 (N_2970,N_1098,N_1375);
nand U2971 (N_2971,N_1896,N_1372);
nand U2972 (N_2972,N_1225,N_1000);
nor U2973 (N_2973,N_1744,N_1784);
and U2974 (N_2974,N_1970,N_1008);
nor U2975 (N_2975,N_1824,N_1628);
and U2976 (N_2976,N_1860,N_1116);
nor U2977 (N_2977,N_1802,N_1756);
or U2978 (N_2978,N_1324,N_1971);
nor U2979 (N_2979,N_1971,N_1726);
and U2980 (N_2980,N_1916,N_1367);
and U2981 (N_2981,N_1510,N_1872);
and U2982 (N_2982,N_1844,N_1179);
and U2983 (N_2983,N_1066,N_1377);
nor U2984 (N_2984,N_1747,N_1044);
nor U2985 (N_2985,N_1836,N_1182);
and U2986 (N_2986,N_1308,N_1614);
and U2987 (N_2987,N_1226,N_1689);
and U2988 (N_2988,N_1879,N_1018);
and U2989 (N_2989,N_1595,N_1322);
nand U2990 (N_2990,N_1559,N_1036);
nand U2991 (N_2991,N_1627,N_1292);
or U2992 (N_2992,N_1683,N_1888);
nor U2993 (N_2993,N_1278,N_1832);
or U2994 (N_2994,N_1230,N_1847);
and U2995 (N_2995,N_1391,N_1473);
nand U2996 (N_2996,N_1165,N_1865);
xnor U2997 (N_2997,N_1001,N_1412);
nand U2998 (N_2998,N_1824,N_1668);
nor U2999 (N_2999,N_1166,N_1743);
nand U3000 (N_3000,N_2523,N_2316);
or U3001 (N_3001,N_2929,N_2518);
or U3002 (N_3002,N_2222,N_2897);
and U3003 (N_3003,N_2394,N_2680);
or U3004 (N_3004,N_2564,N_2577);
nand U3005 (N_3005,N_2857,N_2977);
or U3006 (N_3006,N_2024,N_2665);
and U3007 (N_3007,N_2639,N_2839);
and U3008 (N_3008,N_2908,N_2931);
nand U3009 (N_3009,N_2158,N_2776);
or U3010 (N_3010,N_2837,N_2195);
nor U3011 (N_3011,N_2666,N_2988);
nand U3012 (N_3012,N_2039,N_2312);
and U3013 (N_3013,N_2346,N_2229);
nand U3014 (N_3014,N_2924,N_2128);
nor U3015 (N_3015,N_2901,N_2983);
nor U3016 (N_3016,N_2487,N_2053);
nor U3017 (N_3017,N_2359,N_2586);
or U3018 (N_3018,N_2253,N_2736);
or U3019 (N_3019,N_2446,N_2542);
or U3020 (N_3020,N_2937,N_2696);
nor U3021 (N_3021,N_2580,N_2871);
nand U3022 (N_3022,N_2991,N_2131);
nor U3023 (N_3023,N_2828,N_2519);
and U3024 (N_3024,N_2202,N_2961);
and U3025 (N_3025,N_2042,N_2959);
and U3026 (N_3026,N_2513,N_2812);
nor U3027 (N_3027,N_2074,N_2159);
or U3028 (N_3028,N_2259,N_2488);
and U3029 (N_3029,N_2390,N_2714);
nand U3030 (N_3030,N_2778,N_2300);
and U3031 (N_3031,N_2473,N_2620);
and U3032 (N_3032,N_2900,N_2150);
nand U3033 (N_3033,N_2412,N_2560);
or U3034 (N_3034,N_2921,N_2726);
nand U3035 (N_3035,N_2647,N_2392);
and U3036 (N_3036,N_2790,N_2920);
nor U3037 (N_3037,N_2362,N_2214);
or U3038 (N_3038,N_2122,N_2444);
nor U3039 (N_3039,N_2808,N_2764);
nor U3040 (N_3040,N_2766,N_2065);
and U3041 (N_3041,N_2759,N_2092);
and U3042 (N_3042,N_2958,N_2091);
nor U3043 (N_3043,N_2052,N_2252);
nand U3044 (N_3044,N_2372,N_2025);
nor U3045 (N_3045,N_2136,N_2045);
nor U3046 (N_3046,N_2238,N_2060);
and U3047 (N_3047,N_2781,N_2701);
nand U3048 (N_3048,N_2532,N_2850);
and U3049 (N_3049,N_2330,N_2244);
and U3050 (N_3050,N_2310,N_2894);
nand U3051 (N_3051,N_2228,N_2435);
nand U3052 (N_3052,N_2964,N_2420);
or U3053 (N_3053,N_2332,N_2942);
and U3054 (N_3054,N_2290,N_2996);
nand U3055 (N_3055,N_2307,N_2479);
nand U3056 (N_3056,N_2489,N_2910);
or U3057 (N_3057,N_2711,N_2089);
nor U3058 (N_3058,N_2561,N_2892);
and U3059 (N_3059,N_2719,N_2268);
nor U3060 (N_3060,N_2006,N_2410);
or U3061 (N_3061,N_2795,N_2842);
and U3062 (N_3062,N_2474,N_2124);
and U3063 (N_3063,N_2567,N_2890);
or U3064 (N_3064,N_2118,N_2787);
nand U3065 (N_3065,N_2831,N_2686);
or U3066 (N_3066,N_2297,N_2695);
or U3067 (N_3067,N_2585,N_2744);
nand U3068 (N_3068,N_2514,N_2311);
and U3069 (N_3069,N_2792,N_2434);
or U3070 (N_3070,N_2399,N_2725);
and U3071 (N_3071,N_2611,N_2555);
nor U3072 (N_3072,N_2997,N_2544);
and U3073 (N_3073,N_2369,N_2236);
and U3074 (N_3074,N_2440,N_2504);
or U3075 (N_3075,N_2438,N_2437);
nor U3076 (N_3076,N_2391,N_2044);
nand U3077 (N_3077,N_2037,N_2738);
or U3078 (N_3078,N_2535,N_2050);
nor U3079 (N_3079,N_2660,N_2218);
nor U3080 (N_3080,N_2094,N_2872);
nor U3081 (N_3081,N_2062,N_2129);
nor U3082 (N_3082,N_2589,N_2067);
xnor U3083 (N_3083,N_2141,N_2189);
or U3084 (N_3084,N_2130,N_2486);
or U3085 (N_3085,N_2888,N_2713);
and U3086 (N_3086,N_2728,N_2454);
and U3087 (N_3087,N_2134,N_2273);
nand U3088 (N_3088,N_2969,N_2351);
and U3089 (N_3089,N_2098,N_2603);
or U3090 (N_3090,N_2791,N_2557);
and U3091 (N_3091,N_2581,N_2638);
nor U3092 (N_3092,N_2706,N_2995);
or U3093 (N_3093,N_2682,N_2190);
nand U3094 (N_3094,N_2017,N_2135);
nor U3095 (N_3095,N_2971,N_2395);
nand U3096 (N_3096,N_2380,N_2972);
nand U3097 (N_3097,N_2676,N_2856);
nor U3098 (N_3098,N_2646,N_2443);
nand U3099 (N_3099,N_2840,N_2112);
and U3100 (N_3100,N_2344,N_2260);
nor U3101 (N_3101,N_2215,N_2397);
and U3102 (N_3102,N_2785,N_2626);
nand U3103 (N_3103,N_2002,N_2863);
nor U3104 (N_3104,N_2595,N_2153);
nand U3105 (N_3105,N_2334,N_2191);
nand U3106 (N_3106,N_2175,N_2993);
nand U3107 (N_3107,N_2800,N_2343);
or U3108 (N_3108,N_2278,N_2406);
nor U3109 (N_3109,N_2623,N_2289);
and U3110 (N_3110,N_2464,N_2957);
or U3111 (N_3111,N_2370,N_2182);
or U3112 (N_3112,N_2318,N_2569);
or U3113 (N_3113,N_2678,N_2777);
nand U3114 (N_3114,N_2949,N_2799);
or U3115 (N_3115,N_2246,N_2865);
or U3116 (N_3116,N_2771,N_2484);
or U3117 (N_3117,N_2427,N_2408);
and U3118 (N_3118,N_2166,N_2357);
nor U3119 (N_3119,N_2866,N_2822);
and U3120 (N_3120,N_2447,N_2819);
or U3121 (N_3121,N_2176,N_2256);
or U3122 (N_3122,N_2756,N_2715);
nand U3123 (N_3123,N_2783,N_2152);
nor U3124 (N_3124,N_2192,N_2164);
nand U3125 (N_3125,N_2951,N_2525);
and U3126 (N_3126,N_2517,N_2775);
or U3127 (N_3127,N_2163,N_2201);
xor U3128 (N_3128,N_2693,N_2597);
or U3129 (N_3129,N_2876,N_2617);
and U3130 (N_3130,N_2106,N_2655);
or U3131 (N_3131,N_2896,N_2178);
nor U3132 (N_3132,N_2482,N_2944);
and U3133 (N_3133,N_2827,N_2078);
or U3134 (N_3134,N_2559,N_2952);
or U3135 (N_3135,N_2541,N_2833);
or U3136 (N_3136,N_2388,N_2076);
or U3137 (N_3137,N_2345,N_2494);
or U3138 (N_3138,N_2223,N_2167);
or U3139 (N_3139,N_2085,N_2441);
nor U3140 (N_3140,N_2099,N_2954);
and U3141 (N_3141,N_2948,N_2095);
nor U3142 (N_3142,N_2267,N_2142);
nor U3143 (N_3143,N_2398,N_2433);
nor U3144 (N_3144,N_2859,N_2043);
nor U3145 (N_3145,N_2020,N_2613);
nor U3146 (N_3146,N_2788,N_2409);
nand U3147 (N_3147,N_2622,N_2374);
nor U3148 (N_3148,N_2279,N_2763);
and U3149 (N_3149,N_2070,N_2625);
xor U3150 (N_3150,N_2832,N_2291);
or U3151 (N_3151,N_2926,N_2331);
nor U3152 (N_3152,N_2459,N_2976);
nor U3153 (N_3153,N_2478,N_2919);
or U3154 (N_3154,N_2619,N_2093);
and U3155 (N_3155,N_2361,N_2377);
and U3156 (N_3156,N_2923,N_2907);
and U3157 (N_3157,N_2905,N_2855);
and U3158 (N_3158,N_2879,N_2063);
nand U3159 (N_3159,N_2220,N_2698);
and U3160 (N_3160,N_2064,N_2242);
or U3161 (N_3161,N_2430,N_2366);
or U3162 (N_3162,N_2174,N_2087);
nor U3163 (N_3163,N_2426,N_2990);
nor U3164 (N_3164,N_2315,N_2632);
nand U3165 (N_3165,N_2480,N_2934);
or U3166 (N_3166,N_2165,N_2097);
xor U3167 (N_3167,N_2739,N_2904);
nand U3168 (N_3168,N_2211,N_2858);
or U3169 (N_3169,N_2936,N_2336);
nor U3170 (N_3170,N_2825,N_2008);
and U3171 (N_3171,N_2265,N_2975);
xnor U3172 (N_3172,N_2533,N_2393);
xnor U3173 (N_3173,N_2594,N_2467);
and U3174 (N_3174,N_2452,N_2335);
nor U3175 (N_3175,N_2009,N_2047);
or U3176 (N_3176,N_2111,N_2630);
nand U3177 (N_3177,N_2477,N_2015);
and U3178 (N_3178,N_2621,N_2154);
nand U3179 (N_3179,N_2531,N_2319);
nand U3180 (N_3180,N_2151,N_2575);
nand U3181 (N_3181,N_2610,N_2574);
nor U3182 (N_3182,N_2168,N_2662);
nor U3183 (N_3183,N_2329,N_2700);
nor U3184 (N_3184,N_2180,N_2127);
or U3185 (N_3185,N_2768,N_2930);
nor U3186 (N_3186,N_2634,N_2707);
or U3187 (N_3187,N_2925,N_2173);
nand U3188 (N_3188,N_2249,N_2558);
nor U3189 (N_3189,N_2472,N_2605);
or U3190 (N_3190,N_2225,N_2465);
nand U3191 (N_3191,N_2084,N_2549);
nand U3192 (N_3192,N_2028,N_2294);
and U3193 (N_3193,N_2498,N_2295);
nor U3194 (N_3194,N_2852,N_2512);
or U3195 (N_3195,N_2079,N_2609);
nor U3196 (N_3196,N_2687,N_2608);
or U3197 (N_3197,N_2684,N_2432);
nor U3198 (N_3198,N_2301,N_2679);
and U3199 (N_3199,N_2341,N_2974);
and U3200 (N_3200,N_2068,N_2889);
and U3201 (N_3201,N_2618,N_2939);
or U3202 (N_3202,N_2891,N_2875);
nand U3203 (N_3203,N_2524,N_2199);
xnor U3204 (N_3204,N_2817,N_2132);
and U3205 (N_3205,N_2641,N_2116);
nor U3206 (N_3206,N_2963,N_2635);
or U3207 (N_3207,N_2515,N_2456);
nand U3208 (N_3208,N_2054,N_2539);
or U3209 (N_3209,N_2970,N_2554);
or U3210 (N_3210,N_2709,N_2100);
nand U3211 (N_3211,N_2149,N_2522);
nand U3212 (N_3212,N_2500,N_2540);
or U3213 (N_3213,N_2598,N_2418);
or U3214 (N_3214,N_2965,N_2227);
nand U3215 (N_3215,N_2762,N_2461);
nand U3216 (N_3216,N_2004,N_2770);
or U3217 (N_3217,N_2333,N_2258);
nand U3218 (N_3218,N_2587,N_2731);
or U3219 (N_3219,N_2439,N_2945);
nand U3220 (N_3220,N_2013,N_2146);
and U3221 (N_3221,N_2906,N_2987);
nand U3222 (N_3222,N_2046,N_2108);
and U3223 (N_3223,N_2668,N_2276);
nor U3224 (N_3224,N_2749,N_2740);
nor U3225 (N_3225,N_2296,N_2272);
or U3226 (N_3226,N_2022,N_2962);
and U3227 (N_3227,N_2019,N_2520);
nand U3228 (N_3228,N_2615,N_2212);
nor U3229 (N_3229,N_2162,N_2860);
or U3230 (N_3230,N_2526,N_2255);
nor U3231 (N_3231,N_2348,N_2119);
or U3232 (N_3232,N_2502,N_2287);
nand U3233 (N_3233,N_2221,N_2462);
nor U3234 (N_3234,N_2172,N_2233);
nand U3235 (N_3235,N_2798,N_2985);
or U3236 (N_3236,N_2917,N_2773);
or U3237 (N_3237,N_2234,N_2803);
nand U3238 (N_3238,N_2056,N_2080);
nand U3239 (N_3239,N_2177,N_2838);
and U3240 (N_3240,N_2813,N_2968);
nand U3241 (N_3241,N_2774,N_2210);
nand U3242 (N_3242,N_2356,N_2612);
and U3243 (N_3243,N_2846,N_2818);
nand U3244 (N_3244,N_2724,N_2292);
or U3245 (N_3245,N_2789,N_2378);
nand U3246 (N_3246,N_2844,N_2385);
or U3247 (N_3247,N_2805,N_2286);
and U3248 (N_3248,N_2281,N_2881);
nor U3249 (N_3249,N_2932,N_2353);
and U3250 (N_3250,N_2324,N_2072);
or U3251 (N_3251,N_2349,N_2027);
nand U3252 (N_3252,N_2001,N_2882);
nor U3253 (N_3253,N_2120,N_2508);
or U3254 (N_3254,N_2873,N_2947);
nand U3255 (N_3255,N_2697,N_2148);
nor U3256 (N_3256,N_2614,N_2752);
and U3257 (N_3257,N_2185,N_2760);
nor U3258 (N_3258,N_2110,N_2326);
nand U3259 (N_3259,N_2735,N_2381);
nor U3260 (N_3260,N_2509,N_2683);
or U3261 (N_3261,N_2553,N_2946);
nand U3262 (N_3262,N_2811,N_2914);
nor U3263 (N_3263,N_2648,N_2835);
or U3264 (N_3264,N_2782,N_2563);
nor U3265 (N_3265,N_2673,N_2217);
and U3266 (N_3266,N_2967,N_2848);
and U3267 (N_3267,N_2516,N_2672);
nand U3268 (N_3268,N_2371,N_2083);
nor U3269 (N_3269,N_2007,N_2911);
nand U3270 (N_3270,N_2703,N_2566);
xor U3271 (N_3271,N_2144,N_2354);
and U3272 (N_3272,N_2841,N_2137);
nand U3273 (N_3273,N_2821,N_2186);
or U3274 (N_3274,N_2237,N_2868);
and U3275 (N_3275,N_2145,N_2556);
nor U3276 (N_3276,N_2796,N_2355);
or U3277 (N_3277,N_2075,N_2179);
or U3278 (N_3278,N_2373,N_2205);
and U3279 (N_3279,N_2547,N_2629);
and U3280 (N_3280,N_2893,N_2845);
or U3281 (N_3281,N_2637,N_2160);
or U3282 (N_3282,N_2950,N_2196);
or U3283 (N_3283,N_2723,N_2854);
nor U3284 (N_3284,N_2704,N_2722);
and U3285 (N_3285,N_2506,N_2309);
or U3286 (N_3286,N_2123,N_2867);
nor U3287 (N_3287,N_2208,N_2669);
nor U3288 (N_3288,N_2633,N_2030);
nand U3289 (N_3289,N_2384,N_2694);
or U3290 (N_3290,N_2671,N_2584);
and U3291 (N_3291,N_2747,N_2973);
and U3292 (N_3292,N_2011,N_2627);
nand U3293 (N_3293,N_2884,N_2853);
nand U3294 (N_3294,N_2449,N_2018);
nand U3295 (N_3295,N_2862,N_2143);
nor U3296 (N_3296,N_2654,N_2457);
nand U3297 (N_3297,N_2601,N_2263);
nor U3298 (N_3298,N_2029,N_2328);
nor U3299 (N_3299,N_2960,N_2741);
or U3300 (N_3300,N_2302,N_2299);
or U3301 (N_3301,N_2732,N_2401);
nand U3302 (N_3302,N_2224,N_2986);
nand U3303 (N_3303,N_2170,N_2802);
and U3304 (N_3304,N_2667,N_2303);
nand U3305 (N_3305,N_2448,N_2801);
nand U3306 (N_3306,N_2424,N_2415);
nand U3307 (N_3307,N_2103,N_2927);
nand U3308 (N_3308,N_2023,N_2583);
and U3309 (N_3309,N_2748,N_2998);
or U3310 (N_3310,N_2016,N_2365);
and U3311 (N_3311,N_2293,N_2308);
or U3312 (N_3312,N_2270,N_2797);
nor U3313 (N_3313,N_2849,N_2313);
nand U3314 (N_3314,N_2471,N_2705);
nand U3315 (N_3315,N_2400,N_2994);
and U3316 (N_3316,N_2499,N_2643);
or U3317 (N_3317,N_2602,N_2870);
or U3318 (N_3318,N_2898,N_2031);
and U3319 (N_3319,N_2721,N_2049);
nand U3320 (N_3320,N_2829,N_2830);
nor U3321 (N_3321,N_2109,N_2710);
and U3322 (N_3322,N_2032,N_2451);
and U3323 (N_3323,N_2413,N_2277);
nor U3324 (N_3324,N_2073,N_2599);
or U3325 (N_3325,N_2941,N_2729);
or U3326 (N_3326,N_2284,N_2491);
or U3327 (N_3327,N_2593,N_2241);
or U3328 (N_3328,N_2712,N_2262);
nor U3329 (N_3329,N_2507,N_2423);
or U3330 (N_3330,N_2922,N_2984);
nand U3331 (N_3331,N_2530,N_2915);
nor U3332 (N_3332,N_2588,N_2363);
and U3333 (N_3333,N_2003,N_2576);
or U3334 (N_3334,N_2306,N_2982);
and U3335 (N_3335,N_2989,N_2652);
nor U3336 (N_3336,N_2836,N_2733);
nor U3337 (N_3337,N_2198,N_2183);
nand U3338 (N_3338,N_2887,N_2264);
or U3339 (N_3339,N_2463,N_2940);
xnor U3340 (N_3340,N_2543,N_2718);
and U3341 (N_3341,N_2193,N_2081);
nand U3342 (N_3342,N_2360,N_2383);
and U3343 (N_3343,N_2240,N_2226);
and U3344 (N_3344,N_2628,N_2653);
or U3345 (N_3345,N_2405,N_2537);
or U3346 (N_3346,N_2981,N_2470);
nand U3347 (N_3347,N_2490,N_2903);
nor U3348 (N_3348,N_2751,N_2431);
or U3349 (N_3349,N_2592,N_2661);
nand U3350 (N_3350,N_2352,N_2235);
or U3351 (N_3351,N_2935,N_2493);
nand U3352 (N_3352,N_2161,N_2114);
or U3353 (N_3353,N_2057,N_2036);
nor U3354 (N_3354,N_2650,N_2271);
and U3355 (N_3355,N_2035,N_2786);
or U3356 (N_3356,N_2815,N_2659);
or U3357 (N_3357,N_2651,N_2206);
or U3358 (N_3358,N_2913,N_2861);
or U3359 (N_3359,N_2347,N_2780);
nor U3360 (N_3360,N_2288,N_2458);
nand U3361 (N_3361,N_2690,N_2501);
and U3362 (N_3362,N_2794,N_2282);
or U3363 (N_3363,N_2505,N_2834);
nand U3364 (N_3364,N_2232,N_2304);
and U3365 (N_3365,N_2536,N_2061);
and U3366 (N_3366,N_2257,N_2285);
nor U3367 (N_3367,N_2342,N_2527);
or U3368 (N_3368,N_2104,N_2869);
nor U3369 (N_3369,N_2283,N_2274);
nor U3370 (N_3370,N_2953,N_2386);
nand U3371 (N_3371,N_2207,N_2026);
nand U3372 (N_3372,N_2758,N_2495);
nand U3373 (N_3373,N_2743,N_2455);
or U3374 (N_3374,N_2885,N_2475);
or U3375 (N_3375,N_2139,N_2496);
or U3376 (N_3376,N_2538,N_2445);
nand U3377 (N_3377,N_2197,N_2082);
or U3378 (N_3378,N_2823,N_2396);
and U3379 (N_3379,N_2529,N_2243);
or U3380 (N_3380,N_2928,N_2674);
nor U3381 (N_3381,N_2250,N_2375);
or U3382 (N_3382,N_2916,N_2720);
and U3383 (N_3383,N_2090,N_2247);
nand U3384 (N_3384,N_2269,N_2442);
or U3385 (N_3385,N_2086,N_2573);
nor U3386 (N_3386,N_2428,N_2322);
and U3387 (N_3387,N_2677,N_2568);
nor U3388 (N_3388,N_2992,N_2938);
nand U3389 (N_3389,N_2784,N_2670);
and U3390 (N_3390,N_2364,N_2403);
or U3391 (N_3391,N_2570,N_2656);
or U3392 (N_3392,N_2126,N_2000);
nor U3393 (N_3393,N_2231,N_2699);
or U3394 (N_3394,N_2716,N_2809);
or U3395 (N_3395,N_2816,N_2772);
xor U3396 (N_3396,N_2181,N_2010);
and U3397 (N_3397,N_2203,N_2600);
nor U3398 (N_3398,N_2209,N_2414);
and U3399 (N_3399,N_2460,N_2708);
nand U3400 (N_3400,N_2298,N_2769);
nor U3401 (N_3401,N_2978,N_2305);
and U3402 (N_3402,N_2266,N_2320);
and U3403 (N_3403,N_2909,N_2402);
nor U3404 (N_3404,N_2497,N_2545);
nor U3405 (N_3405,N_2810,N_2757);
or U3406 (N_3406,N_2806,N_2765);
nand U3407 (N_3407,N_2675,N_2096);
or U3408 (N_3408,N_2562,N_2337);
nand U3409 (N_3409,N_2636,N_2481);
or U3410 (N_3410,N_2847,N_2469);
nand U3411 (N_3411,N_2552,N_2419);
nand U3412 (N_3412,N_2883,N_2327);
nand U3413 (N_3413,N_2033,N_2933);
xor U3414 (N_3414,N_2314,N_2350);
or U3415 (N_3415,N_2737,N_2807);
and U3416 (N_3416,N_2604,N_2213);
and U3417 (N_3417,N_2980,N_2804);
and U3418 (N_3418,N_2691,N_2843);
nand U3419 (N_3419,N_2321,N_2730);
or U3420 (N_3420,N_2358,N_2658);
nand U3421 (N_3421,N_2546,N_2387);
nor U3422 (N_3422,N_2105,N_2503);
or U3423 (N_3423,N_2579,N_2548);
nor U3424 (N_3424,N_2066,N_2793);
nor U3425 (N_3425,N_2761,N_2820);
xnor U3426 (N_3426,N_2014,N_2956);
and U3427 (N_3427,N_2416,N_2999);
nand U3428 (N_3428,N_2171,N_2453);
nor U3429 (N_3429,N_2102,N_2874);
nand U3430 (N_3430,N_2902,N_2204);
and U3431 (N_3431,N_2323,N_2059);
and U3432 (N_3432,N_2382,N_2966);
or U3433 (N_3433,N_2631,N_2685);
nor U3434 (N_3434,N_2239,N_2492);
nor U3435 (N_3435,N_2169,N_2483);
or U3436 (N_3436,N_2367,N_2750);
and U3437 (N_3437,N_2943,N_2734);
nor U3438 (N_3438,N_2245,N_2389);
and U3439 (N_3439,N_2663,N_2582);
and U3440 (N_3440,N_2779,N_2038);
nand U3441 (N_3441,N_2254,N_2664);
or U3442 (N_3442,N_2754,N_2755);
or U3443 (N_3443,N_2899,N_2551);
or U3444 (N_3444,N_2912,N_2115);
nand U3445 (N_3445,N_2688,N_2878);
nand U3446 (N_3446,N_2261,N_2826);
nand U3447 (N_3447,N_2534,N_2689);
nor U3448 (N_3448,N_2101,N_2717);
and U3449 (N_3449,N_2051,N_2644);
or U3450 (N_3450,N_2468,N_2550);
or U3451 (N_3451,N_2125,N_2476);
nand U3452 (N_3452,N_2767,N_2745);
nor U3453 (N_3453,N_2048,N_2607);
and U3454 (N_3454,N_2591,N_2578);
and U3455 (N_3455,N_2280,N_2147);
and U3456 (N_3456,N_2230,N_2877);
nor U3457 (N_3457,N_2034,N_2521);
and U3458 (N_3458,N_2485,N_2590);
nand U3459 (N_3459,N_2157,N_2979);
nor U3460 (N_3460,N_2184,N_2742);
and U3461 (N_3461,N_2746,N_2624);
nand U3462 (N_3462,N_2572,N_2155);
nand U3463 (N_3463,N_2436,N_2851);
nor U3464 (N_3464,N_2021,N_2317);
or U3465 (N_3465,N_2058,N_2117);
and U3466 (N_3466,N_2140,N_2133);
nor U3467 (N_3467,N_2379,N_2156);
or U3468 (N_3468,N_2368,N_2088);
and U3469 (N_3469,N_2640,N_2753);
or U3470 (N_3470,N_2325,N_2421);
nand U3471 (N_3471,N_2187,N_2616);
or U3472 (N_3472,N_2113,N_2692);
and U3473 (N_3473,N_2571,N_2404);
nand U3474 (N_3474,N_2077,N_2340);
nor U3475 (N_3475,N_2138,N_2248);
nor U3476 (N_3476,N_2727,N_2814);
or U3477 (N_3477,N_2642,N_2606);
nor U3478 (N_3478,N_2376,N_2895);
or U3479 (N_3479,N_2251,N_2012);
and U3480 (N_3480,N_2216,N_2041);
nand U3481 (N_3481,N_2411,N_2275);
nand U3482 (N_3482,N_2955,N_2466);
nand U3483 (N_3483,N_2511,N_2510);
nor U3484 (N_3484,N_2055,N_2824);
nand U3485 (N_3485,N_2219,N_2194);
nand U3486 (N_3486,N_2339,N_2918);
nand U3487 (N_3487,N_2040,N_2681);
nor U3488 (N_3488,N_2528,N_2645);
nor U3489 (N_3489,N_2657,N_2702);
or U3490 (N_3490,N_2649,N_2407);
or U3491 (N_3491,N_2425,N_2338);
nor U3492 (N_3492,N_2596,N_2880);
and U3493 (N_3493,N_2417,N_2121);
nand U3494 (N_3494,N_2429,N_2069);
nor U3495 (N_3495,N_2188,N_2864);
nor U3496 (N_3496,N_2422,N_2200);
and U3497 (N_3497,N_2005,N_2565);
nor U3498 (N_3498,N_2107,N_2071);
nor U3499 (N_3499,N_2450,N_2886);
nor U3500 (N_3500,N_2781,N_2727);
nand U3501 (N_3501,N_2623,N_2581);
and U3502 (N_3502,N_2333,N_2274);
nand U3503 (N_3503,N_2076,N_2213);
nand U3504 (N_3504,N_2446,N_2086);
nand U3505 (N_3505,N_2470,N_2186);
or U3506 (N_3506,N_2573,N_2789);
nor U3507 (N_3507,N_2725,N_2632);
nor U3508 (N_3508,N_2190,N_2019);
xnor U3509 (N_3509,N_2075,N_2034);
and U3510 (N_3510,N_2492,N_2142);
and U3511 (N_3511,N_2236,N_2918);
nor U3512 (N_3512,N_2605,N_2597);
or U3513 (N_3513,N_2579,N_2689);
nor U3514 (N_3514,N_2119,N_2150);
and U3515 (N_3515,N_2625,N_2504);
or U3516 (N_3516,N_2980,N_2628);
nand U3517 (N_3517,N_2091,N_2189);
nor U3518 (N_3518,N_2667,N_2774);
nor U3519 (N_3519,N_2692,N_2179);
nand U3520 (N_3520,N_2535,N_2738);
nor U3521 (N_3521,N_2927,N_2338);
and U3522 (N_3522,N_2630,N_2497);
and U3523 (N_3523,N_2579,N_2482);
and U3524 (N_3524,N_2976,N_2590);
or U3525 (N_3525,N_2790,N_2713);
or U3526 (N_3526,N_2703,N_2539);
and U3527 (N_3527,N_2136,N_2002);
and U3528 (N_3528,N_2811,N_2047);
and U3529 (N_3529,N_2628,N_2486);
and U3530 (N_3530,N_2400,N_2536);
nand U3531 (N_3531,N_2164,N_2138);
or U3532 (N_3532,N_2893,N_2215);
or U3533 (N_3533,N_2649,N_2625);
nor U3534 (N_3534,N_2227,N_2252);
nand U3535 (N_3535,N_2925,N_2903);
or U3536 (N_3536,N_2210,N_2329);
and U3537 (N_3537,N_2833,N_2198);
or U3538 (N_3538,N_2821,N_2861);
and U3539 (N_3539,N_2717,N_2728);
and U3540 (N_3540,N_2508,N_2666);
and U3541 (N_3541,N_2005,N_2490);
and U3542 (N_3542,N_2066,N_2146);
nand U3543 (N_3543,N_2241,N_2524);
and U3544 (N_3544,N_2187,N_2568);
nor U3545 (N_3545,N_2225,N_2046);
nor U3546 (N_3546,N_2047,N_2074);
nor U3547 (N_3547,N_2090,N_2107);
or U3548 (N_3548,N_2844,N_2348);
or U3549 (N_3549,N_2451,N_2410);
and U3550 (N_3550,N_2613,N_2707);
or U3551 (N_3551,N_2800,N_2895);
or U3552 (N_3552,N_2866,N_2821);
and U3553 (N_3553,N_2395,N_2933);
nor U3554 (N_3554,N_2749,N_2348);
and U3555 (N_3555,N_2259,N_2749);
and U3556 (N_3556,N_2467,N_2578);
nand U3557 (N_3557,N_2033,N_2544);
nand U3558 (N_3558,N_2226,N_2219);
and U3559 (N_3559,N_2124,N_2878);
nand U3560 (N_3560,N_2864,N_2220);
and U3561 (N_3561,N_2355,N_2467);
nor U3562 (N_3562,N_2487,N_2758);
and U3563 (N_3563,N_2319,N_2729);
and U3564 (N_3564,N_2707,N_2653);
nor U3565 (N_3565,N_2792,N_2800);
or U3566 (N_3566,N_2068,N_2215);
nand U3567 (N_3567,N_2706,N_2890);
nand U3568 (N_3568,N_2787,N_2294);
nand U3569 (N_3569,N_2173,N_2641);
and U3570 (N_3570,N_2000,N_2836);
and U3571 (N_3571,N_2766,N_2823);
or U3572 (N_3572,N_2594,N_2795);
and U3573 (N_3573,N_2650,N_2227);
or U3574 (N_3574,N_2472,N_2771);
nand U3575 (N_3575,N_2186,N_2777);
or U3576 (N_3576,N_2127,N_2251);
and U3577 (N_3577,N_2670,N_2923);
nor U3578 (N_3578,N_2622,N_2117);
nor U3579 (N_3579,N_2152,N_2658);
and U3580 (N_3580,N_2933,N_2273);
and U3581 (N_3581,N_2238,N_2186);
nor U3582 (N_3582,N_2153,N_2258);
nor U3583 (N_3583,N_2652,N_2570);
nand U3584 (N_3584,N_2220,N_2348);
nor U3585 (N_3585,N_2559,N_2010);
or U3586 (N_3586,N_2445,N_2015);
or U3587 (N_3587,N_2737,N_2843);
and U3588 (N_3588,N_2783,N_2577);
and U3589 (N_3589,N_2570,N_2045);
and U3590 (N_3590,N_2032,N_2757);
or U3591 (N_3591,N_2772,N_2178);
nor U3592 (N_3592,N_2091,N_2315);
or U3593 (N_3593,N_2907,N_2950);
nand U3594 (N_3594,N_2212,N_2096);
nor U3595 (N_3595,N_2465,N_2714);
nor U3596 (N_3596,N_2489,N_2731);
nor U3597 (N_3597,N_2453,N_2656);
and U3598 (N_3598,N_2690,N_2596);
nand U3599 (N_3599,N_2989,N_2862);
and U3600 (N_3600,N_2648,N_2866);
nand U3601 (N_3601,N_2664,N_2507);
and U3602 (N_3602,N_2307,N_2997);
nand U3603 (N_3603,N_2275,N_2527);
or U3604 (N_3604,N_2302,N_2152);
or U3605 (N_3605,N_2089,N_2785);
nand U3606 (N_3606,N_2948,N_2870);
or U3607 (N_3607,N_2291,N_2740);
and U3608 (N_3608,N_2000,N_2633);
and U3609 (N_3609,N_2014,N_2928);
nand U3610 (N_3610,N_2957,N_2382);
or U3611 (N_3611,N_2490,N_2830);
or U3612 (N_3612,N_2117,N_2185);
nor U3613 (N_3613,N_2343,N_2413);
nand U3614 (N_3614,N_2185,N_2093);
nor U3615 (N_3615,N_2860,N_2550);
nor U3616 (N_3616,N_2100,N_2385);
and U3617 (N_3617,N_2983,N_2170);
or U3618 (N_3618,N_2117,N_2440);
nor U3619 (N_3619,N_2619,N_2416);
and U3620 (N_3620,N_2214,N_2960);
nand U3621 (N_3621,N_2971,N_2176);
and U3622 (N_3622,N_2540,N_2782);
and U3623 (N_3623,N_2524,N_2550);
nor U3624 (N_3624,N_2022,N_2806);
or U3625 (N_3625,N_2695,N_2236);
and U3626 (N_3626,N_2492,N_2882);
and U3627 (N_3627,N_2083,N_2550);
nand U3628 (N_3628,N_2527,N_2635);
nand U3629 (N_3629,N_2031,N_2980);
nor U3630 (N_3630,N_2746,N_2535);
or U3631 (N_3631,N_2744,N_2458);
nand U3632 (N_3632,N_2481,N_2203);
or U3633 (N_3633,N_2324,N_2103);
nor U3634 (N_3634,N_2300,N_2009);
and U3635 (N_3635,N_2375,N_2622);
or U3636 (N_3636,N_2654,N_2862);
and U3637 (N_3637,N_2384,N_2689);
and U3638 (N_3638,N_2357,N_2304);
nor U3639 (N_3639,N_2369,N_2484);
or U3640 (N_3640,N_2318,N_2927);
or U3641 (N_3641,N_2931,N_2481);
and U3642 (N_3642,N_2740,N_2981);
nor U3643 (N_3643,N_2933,N_2635);
or U3644 (N_3644,N_2835,N_2421);
nor U3645 (N_3645,N_2339,N_2510);
nor U3646 (N_3646,N_2865,N_2216);
or U3647 (N_3647,N_2858,N_2314);
nor U3648 (N_3648,N_2243,N_2747);
nand U3649 (N_3649,N_2989,N_2857);
nor U3650 (N_3650,N_2607,N_2452);
nand U3651 (N_3651,N_2079,N_2598);
nor U3652 (N_3652,N_2053,N_2036);
nand U3653 (N_3653,N_2657,N_2045);
nor U3654 (N_3654,N_2196,N_2481);
and U3655 (N_3655,N_2889,N_2158);
nand U3656 (N_3656,N_2698,N_2565);
or U3657 (N_3657,N_2024,N_2212);
nor U3658 (N_3658,N_2367,N_2170);
or U3659 (N_3659,N_2905,N_2580);
and U3660 (N_3660,N_2348,N_2123);
nand U3661 (N_3661,N_2685,N_2591);
nor U3662 (N_3662,N_2048,N_2080);
or U3663 (N_3663,N_2825,N_2129);
or U3664 (N_3664,N_2658,N_2385);
nor U3665 (N_3665,N_2938,N_2797);
nand U3666 (N_3666,N_2307,N_2747);
nor U3667 (N_3667,N_2734,N_2588);
or U3668 (N_3668,N_2209,N_2767);
and U3669 (N_3669,N_2003,N_2332);
nand U3670 (N_3670,N_2335,N_2142);
or U3671 (N_3671,N_2019,N_2777);
nand U3672 (N_3672,N_2486,N_2938);
nor U3673 (N_3673,N_2544,N_2743);
and U3674 (N_3674,N_2649,N_2338);
nand U3675 (N_3675,N_2846,N_2479);
nand U3676 (N_3676,N_2718,N_2546);
nand U3677 (N_3677,N_2929,N_2311);
or U3678 (N_3678,N_2946,N_2983);
nand U3679 (N_3679,N_2844,N_2418);
nor U3680 (N_3680,N_2706,N_2050);
nand U3681 (N_3681,N_2695,N_2471);
and U3682 (N_3682,N_2312,N_2292);
nor U3683 (N_3683,N_2489,N_2821);
nand U3684 (N_3684,N_2278,N_2322);
or U3685 (N_3685,N_2394,N_2498);
nand U3686 (N_3686,N_2545,N_2781);
nor U3687 (N_3687,N_2692,N_2292);
nor U3688 (N_3688,N_2539,N_2394);
nor U3689 (N_3689,N_2440,N_2629);
and U3690 (N_3690,N_2686,N_2402);
nand U3691 (N_3691,N_2549,N_2327);
nand U3692 (N_3692,N_2922,N_2355);
and U3693 (N_3693,N_2513,N_2391);
nand U3694 (N_3694,N_2115,N_2708);
nand U3695 (N_3695,N_2722,N_2452);
or U3696 (N_3696,N_2147,N_2029);
and U3697 (N_3697,N_2085,N_2956);
and U3698 (N_3698,N_2723,N_2910);
nor U3699 (N_3699,N_2279,N_2229);
or U3700 (N_3700,N_2162,N_2055);
nor U3701 (N_3701,N_2418,N_2038);
or U3702 (N_3702,N_2341,N_2124);
nand U3703 (N_3703,N_2757,N_2748);
nand U3704 (N_3704,N_2200,N_2571);
and U3705 (N_3705,N_2701,N_2850);
or U3706 (N_3706,N_2503,N_2090);
nor U3707 (N_3707,N_2057,N_2228);
and U3708 (N_3708,N_2596,N_2689);
nand U3709 (N_3709,N_2616,N_2371);
and U3710 (N_3710,N_2289,N_2636);
and U3711 (N_3711,N_2374,N_2299);
xnor U3712 (N_3712,N_2881,N_2825);
nand U3713 (N_3713,N_2638,N_2831);
or U3714 (N_3714,N_2931,N_2699);
nand U3715 (N_3715,N_2352,N_2171);
nand U3716 (N_3716,N_2383,N_2664);
nand U3717 (N_3717,N_2304,N_2634);
or U3718 (N_3718,N_2390,N_2360);
nand U3719 (N_3719,N_2002,N_2116);
and U3720 (N_3720,N_2813,N_2374);
nor U3721 (N_3721,N_2954,N_2542);
or U3722 (N_3722,N_2074,N_2443);
nor U3723 (N_3723,N_2032,N_2201);
or U3724 (N_3724,N_2070,N_2097);
nor U3725 (N_3725,N_2478,N_2244);
and U3726 (N_3726,N_2171,N_2841);
or U3727 (N_3727,N_2606,N_2662);
or U3728 (N_3728,N_2150,N_2928);
and U3729 (N_3729,N_2318,N_2459);
nand U3730 (N_3730,N_2016,N_2547);
or U3731 (N_3731,N_2362,N_2468);
and U3732 (N_3732,N_2010,N_2527);
nand U3733 (N_3733,N_2969,N_2458);
or U3734 (N_3734,N_2161,N_2890);
or U3735 (N_3735,N_2805,N_2791);
and U3736 (N_3736,N_2055,N_2146);
nand U3737 (N_3737,N_2544,N_2291);
xor U3738 (N_3738,N_2887,N_2102);
or U3739 (N_3739,N_2138,N_2882);
or U3740 (N_3740,N_2663,N_2422);
nand U3741 (N_3741,N_2018,N_2159);
nor U3742 (N_3742,N_2159,N_2337);
nand U3743 (N_3743,N_2566,N_2753);
or U3744 (N_3744,N_2938,N_2131);
xor U3745 (N_3745,N_2903,N_2058);
nor U3746 (N_3746,N_2336,N_2175);
or U3747 (N_3747,N_2351,N_2204);
nor U3748 (N_3748,N_2690,N_2533);
nor U3749 (N_3749,N_2975,N_2569);
nand U3750 (N_3750,N_2829,N_2673);
or U3751 (N_3751,N_2100,N_2915);
or U3752 (N_3752,N_2941,N_2611);
xnor U3753 (N_3753,N_2997,N_2071);
nand U3754 (N_3754,N_2209,N_2956);
and U3755 (N_3755,N_2103,N_2819);
nor U3756 (N_3756,N_2076,N_2934);
and U3757 (N_3757,N_2617,N_2330);
nand U3758 (N_3758,N_2492,N_2553);
nand U3759 (N_3759,N_2022,N_2278);
nand U3760 (N_3760,N_2907,N_2679);
or U3761 (N_3761,N_2553,N_2179);
or U3762 (N_3762,N_2485,N_2006);
or U3763 (N_3763,N_2734,N_2369);
and U3764 (N_3764,N_2627,N_2791);
nor U3765 (N_3765,N_2167,N_2249);
nand U3766 (N_3766,N_2090,N_2217);
nand U3767 (N_3767,N_2738,N_2945);
or U3768 (N_3768,N_2482,N_2053);
or U3769 (N_3769,N_2493,N_2587);
and U3770 (N_3770,N_2713,N_2621);
or U3771 (N_3771,N_2625,N_2600);
nor U3772 (N_3772,N_2048,N_2753);
nor U3773 (N_3773,N_2296,N_2489);
and U3774 (N_3774,N_2559,N_2763);
or U3775 (N_3775,N_2568,N_2844);
nand U3776 (N_3776,N_2611,N_2164);
nor U3777 (N_3777,N_2845,N_2943);
nand U3778 (N_3778,N_2064,N_2216);
nand U3779 (N_3779,N_2396,N_2813);
or U3780 (N_3780,N_2654,N_2406);
nand U3781 (N_3781,N_2564,N_2299);
or U3782 (N_3782,N_2630,N_2347);
and U3783 (N_3783,N_2442,N_2851);
or U3784 (N_3784,N_2949,N_2377);
nand U3785 (N_3785,N_2849,N_2787);
nor U3786 (N_3786,N_2614,N_2279);
or U3787 (N_3787,N_2311,N_2528);
and U3788 (N_3788,N_2022,N_2291);
nand U3789 (N_3789,N_2169,N_2815);
nor U3790 (N_3790,N_2026,N_2093);
nor U3791 (N_3791,N_2334,N_2301);
nor U3792 (N_3792,N_2672,N_2830);
or U3793 (N_3793,N_2468,N_2711);
and U3794 (N_3794,N_2790,N_2575);
and U3795 (N_3795,N_2171,N_2296);
and U3796 (N_3796,N_2365,N_2610);
and U3797 (N_3797,N_2437,N_2256);
and U3798 (N_3798,N_2972,N_2185);
nor U3799 (N_3799,N_2326,N_2081);
nor U3800 (N_3800,N_2177,N_2370);
and U3801 (N_3801,N_2615,N_2296);
or U3802 (N_3802,N_2013,N_2478);
nor U3803 (N_3803,N_2410,N_2321);
and U3804 (N_3804,N_2821,N_2362);
or U3805 (N_3805,N_2712,N_2633);
or U3806 (N_3806,N_2478,N_2703);
or U3807 (N_3807,N_2487,N_2888);
and U3808 (N_3808,N_2998,N_2868);
or U3809 (N_3809,N_2169,N_2239);
nand U3810 (N_3810,N_2539,N_2420);
or U3811 (N_3811,N_2858,N_2013);
and U3812 (N_3812,N_2218,N_2127);
nand U3813 (N_3813,N_2098,N_2866);
and U3814 (N_3814,N_2316,N_2890);
nor U3815 (N_3815,N_2677,N_2581);
and U3816 (N_3816,N_2710,N_2399);
nor U3817 (N_3817,N_2643,N_2541);
nor U3818 (N_3818,N_2288,N_2360);
nor U3819 (N_3819,N_2266,N_2154);
nor U3820 (N_3820,N_2469,N_2157);
xor U3821 (N_3821,N_2732,N_2190);
nand U3822 (N_3822,N_2453,N_2978);
nor U3823 (N_3823,N_2973,N_2362);
and U3824 (N_3824,N_2888,N_2250);
or U3825 (N_3825,N_2856,N_2570);
or U3826 (N_3826,N_2282,N_2621);
or U3827 (N_3827,N_2788,N_2523);
or U3828 (N_3828,N_2843,N_2424);
nand U3829 (N_3829,N_2390,N_2008);
nand U3830 (N_3830,N_2492,N_2630);
nand U3831 (N_3831,N_2522,N_2503);
nor U3832 (N_3832,N_2774,N_2074);
nor U3833 (N_3833,N_2195,N_2896);
or U3834 (N_3834,N_2585,N_2308);
or U3835 (N_3835,N_2554,N_2936);
nand U3836 (N_3836,N_2002,N_2819);
and U3837 (N_3837,N_2634,N_2528);
nor U3838 (N_3838,N_2082,N_2011);
and U3839 (N_3839,N_2212,N_2281);
nor U3840 (N_3840,N_2213,N_2820);
or U3841 (N_3841,N_2870,N_2372);
or U3842 (N_3842,N_2602,N_2712);
and U3843 (N_3843,N_2942,N_2868);
nor U3844 (N_3844,N_2243,N_2213);
or U3845 (N_3845,N_2216,N_2989);
nor U3846 (N_3846,N_2630,N_2780);
and U3847 (N_3847,N_2477,N_2376);
nand U3848 (N_3848,N_2311,N_2913);
or U3849 (N_3849,N_2210,N_2977);
and U3850 (N_3850,N_2560,N_2064);
nor U3851 (N_3851,N_2343,N_2341);
or U3852 (N_3852,N_2897,N_2842);
and U3853 (N_3853,N_2814,N_2389);
nor U3854 (N_3854,N_2510,N_2983);
and U3855 (N_3855,N_2928,N_2943);
or U3856 (N_3856,N_2219,N_2987);
nand U3857 (N_3857,N_2016,N_2900);
nor U3858 (N_3858,N_2561,N_2817);
nor U3859 (N_3859,N_2752,N_2720);
and U3860 (N_3860,N_2367,N_2454);
nor U3861 (N_3861,N_2103,N_2297);
nand U3862 (N_3862,N_2498,N_2464);
nor U3863 (N_3863,N_2921,N_2883);
and U3864 (N_3864,N_2163,N_2564);
or U3865 (N_3865,N_2942,N_2106);
and U3866 (N_3866,N_2906,N_2569);
nor U3867 (N_3867,N_2695,N_2268);
nor U3868 (N_3868,N_2407,N_2759);
or U3869 (N_3869,N_2874,N_2859);
nand U3870 (N_3870,N_2076,N_2826);
and U3871 (N_3871,N_2133,N_2790);
nand U3872 (N_3872,N_2541,N_2302);
nor U3873 (N_3873,N_2570,N_2403);
nand U3874 (N_3874,N_2424,N_2458);
or U3875 (N_3875,N_2209,N_2311);
nor U3876 (N_3876,N_2112,N_2511);
or U3877 (N_3877,N_2633,N_2838);
or U3878 (N_3878,N_2066,N_2679);
xor U3879 (N_3879,N_2884,N_2455);
and U3880 (N_3880,N_2730,N_2536);
nand U3881 (N_3881,N_2990,N_2327);
nor U3882 (N_3882,N_2690,N_2495);
or U3883 (N_3883,N_2221,N_2363);
or U3884 (N_3884,N_2531,N_2888);
nand U3885 (N_3885,N_2877,N_2807);
nor U3886 (N_3886,N_2684,N_2036);
nand U3887 (N_3887,N_2846,N_2447);
and U3888 (N_3888,N_2878,N_2708);
or U3889 (N_3889,N_2574,N_2967);
nor U3890 (N_3890,N_2576,N_2794);
nand U3891 (N_3891,N_2161,N_2846);
nand U3892 (N_3892,N_2701,N_2237);
and U3893 (N_3893,N_2628,N_2777);
nand U3894 (N_3894,N_2589,N_2040);
nand U3895 (N_3895,N_2902,N_2256);
and U3896 (N_3896,N_2269,N_2835);
and U3897 (N_3897,N_2660,N_2343);
nand U3898 (N_3898,N_2326,N_2257);
and U3899 (N_3899,N_2534,N_2031);
nand U3900 (N_3900,N_2979,N_2101);
and U3901 (N_3901,N_2443,N_2634);
nor U3902 (N_3902,N_2480,N_2985);
nand U3903 (N_3903,N_2031,N_2392);
nand U3904 (N_3904,N_2179,N_2893);
or U3905 (N_3905,N_2475,N_2903);
and U3906 (N_3906,N_2447,N_2315);
or U3907 (N_3907,N_2037,N_2236);
nor U3908 (N_3908,N_2206,N_2016);
nor U3909 (N_3909,N_2184,N_2710);
and U3910 (N_3910,N_2751,N_2405);
or U3911 (N_3911,N_2846,N_2511);
or U3912 (N_3912,N_2281,N_2248);
nor U3913 (N_3913,N_2541,N_2462);
nor U3914 (N_3914,N_2886,N_2892);
and U3915 (N_3915,N_2260,N_2925);
nor U3916 (N_3916,N_2106,N_2475);
or U3917 (N_3917,N_2590,N_2455);
nand U3918 (N_3918,N_2467,N_2322);
and U3919 (N_3919,N_2288,N_2340);
and U3920 (N_3920,N_2812,N_2808);
or U3921 (N_3921,N_2696,N_2286);
and U3922 (N_3922,N_2431,N_2612);
and U3923 (N_3923,N_2583,N_2610);
nand U3924 (N_3924,N_2671,N_2810);
nand U3925 (N_3925,N_2541,N_2175);
nand U3926 (N_3926,N_2337,N_2584);
nor U3927 (N_3927,N_2621,N_2307);
or U3928 (N_3928,N_2385,N_2756);
nor U3929 (N_3929,N_2133,N_2924);
nor U3930 (N_3930,N_2873,N_2695);
and U3931 (N_3931,N_2429,N_2893);
or U3932 (N_3932,N_2405,N_2255);
or U3933 (N_3933,N_2556,N_2732);
or U3934 (N_3934,N_2214,N_2038);
nand U3935 (N_3935,N_2196,N_2275);
nand U3936 (N_3936,N_2324,N_2642);
nand U3937 (N_3937,N_2756,N_2365);
nand U3938 (N_3938,N_2848,N_2499);
nand U3939 (N_3939,N_2484,N_2695);
or U3940 (N_3940,N_2649,N_2852);
or U3941 (N_3941,N_2629,N_2334);
or U3942 (N_3942,N_2813,N_2281);
or U3943 (N_3943,N_2862,N_2982);
nand U3944 (N_3944,N_2819,N_2211);
nand U3945 (N_3945,N_2486,N_2587);
nor U3946 (N_3946,N_2888,N_2937);
and U3947 (N_3947,N_2052,N_2849);
nor U3948 (N_3948,N_2300,N_2285);
nand U3949 (N_3949,N_2202,N_2409);
and U3950 (N_3950,N_2965,N_2897);
nor U3951 (N_3951,N_2675,N_2462);
and U3952 (N_3952,N_2706,N_2155);
nand U3953 (N_3953,N_2425,N_2672);
nor U3954 (N_3954,N_2602,N_2601);
or U3955 (N_3955,N_2367,N_2356);
nor U3956 (N_3956,N_2684,N_2873);
and U3957 (N_3957,N_2442,N_2914);
nand U3958 (N_3958,N_2540,N_2213);
or U3959 (N_3959,N_2172,N_2096);
nor U3960 (N_3960,N_2715,N_2731);
nor U3961 (N_3961,N_2124,N_2741);
nor U3962 (N_3962,N_2519,N_2565);
nor U3963 (N_3963,N_2556,N_2553);
and U3964 (N_3964,N_2246,N_2986);
xnor U3965 (N_3965,N_2247,N_2851);
nor U3966 (N_3966,N_2292,N_2605);
nor U3967 (N_3967,N_2894,N_2276);
nand U3968 (N_3968,N_2426,N_2411);
or U3969 (N_3969,N_2513,N_2610);
or U3970 (N_3970,N_2047,N_2618);
nand U3971 (N_3971,N_2129,N_2966);
and U3972 (N_3972,N_2185,N_2715);
nand U3973 (N_3973,N_2624,N_2509);
nand U3974 (N_3974,N_2282,N_2769);
or U3975 (N_3975,N_2999,N_2225);
nor U3976 (N_3976,N_2746,N_2588);
nand U3977 (N_3977,N_2604,N_2608);
or U3978 (N_3978,N_2472,N_2731);
or U3979 (N_3979,N_2432,N_2299);
nor U3980 (N_3980,N_2340,N_2801);
or U3981 (N_3981,N_2164,N_2251);
and U3982 (N_3982,N_2465,N_2455);
nand U3983 (N_3983,N_2465,N_2081);
nor U3984 (N_3984,N_2769,N_2186);
nor U3985 (N_3985,N_2896,N_2342);
nor U3986 (N_3986,N_2243,N_2498);
nand U3987 (N_3987,N_2798,N_2138);
and U3988 (N_3988,N_2543,N_2863);
or U3989 (N_3989,N_2735,N_2897);
or U3990 (N_3990,N_2046,N_2410);
or U3991 (N_3991,N_2553,N_2905);
nor U3992 (N_3992,N_2590,N_2793);
and U3993 (N_3993,N_2015,N_2360);
nand U3994 (N_3994,N_2310,N_2778);
or U3995 (N_3995,N_2733,N_2492);
and U3996 (N_3996,N_2611,N_2452);
or U3997 (N_3997,N_2585,N_2121);
nor U3998 (N_3998,N_2744,N_2981);
and U3999 (N_3999,N_2629,N_2357);
and U4000 (N_4000,N_3339,N_3341);
or U4001 (N_4001,N_3338,N_3721);
nand U4002 (N_4002,N_3719,N_3847);
and U4003 (N_4003,N_3095,N_3350);
nor U4004 (N_4004,N_3749,N_3865);
nor U4005 (N_4005,N_3432,N_3690);
and U4006 (N_4006,N_3337,N_3305);
nand U4007 (N_4007,N_3767,N_3023);
or U4008 (N_4008,N_3279,N_3075);
nand U4009 (N_4009,N_3886,N_3144);
nor U4010 (N_4010,N_3856,N_3435);
nor U4011 (N_4011,N_3716,N_3622);
or U4012 (N_4012,N_3970,N_3146);
nor U4013 (N_4013,N_3581,N_3608);
nor U4014 (N_4014,N_3322,N_3898);
nand U4015 (N_4015,N_3018,N_3654);
or U4016 (N_4016,N_3377,N_3897);
or U4017 (N_4017,N_3065,N_3820);
nor U4018 (N_4018,N_3159,N_3662);
or U4019 (N_4019,N_3702,N_3974);
or U4020 (N_4020,N_3384,N_3262);
or U4021 (N_4021,N_3227,N_3631);
nand U4022 (N_4022,N_3200,N_3110);
or U4023 (N_4023,N_3866,N_3940);
nand U4024 (N_4024,N_3442,N_3805);
nor U4025 (N_4025,N_3443,N_3671);
or U4026 (N_4026,N_3240,N_3924);
nand U4027 (N_4027,N_3187,N_3819);
and U4028 (N_4028,N_3378,N_3046);
nand U4029 (N_4029,N_3786,N_3737);
and U4030 (N_4030,N_3685,N_3076);
or U4031 (N_4031,N_3619,N_3463);
nor U4032 (N_4032,N_3366,N_3155);
or U4033 (N_4033,N_3609,N_3951);
nor U4034 (N_4034,N_3299,N_3400);
or U4035 (N_4035,N_3540,N_3170);
nor U4036 (N_4036,N_3004,N_3682);
or U4037 (N_4037,N_3461,N_3000);
nand U4038 (N_4038,N_3616,N_3293);
nor U4039 (N_4039,N_3750,N_3912);
or U4040 (N_4040,N_3879,N_3978);
nand U4041 (N_4041,N_3610,N_3298);
or U4042 (N_4042,N_3954,N_3321);
and U4043 (N_4043,N_3862,N_3165);
nor U4044 (N_4044,N_3241,N_3100);
nand U4045 (N_4045,N_3278,N_3704);
nor U4046 (N_4046,N_3618,N_3256);
or U4047 (N_4047,N_3031,N_3013);
nand U4048 (N_4048,N_3854,N_3390);
or U4049 (N_4049,N_3128,N_3996);
nor U4050 (N_4050,N_3414,N_3948);
and U4051 (N_4051,N_3109,N_3320);
and U4052 (N_4052,N_3229,N_3746);
nor U4053 (N_4053,N_3641,N_3203);
nor U4054 (N_4054,N_3106,N_3927);
nand U4055 (N_4055,N_3519,N_3582);
and U4056 (N_4056,N_3172,N_3994);
and U4057 (N_4057,N_3041,N_3148);
or U4058 (N_4058,N_3349,N_3402);
or U4059 (N_4059,N_3953,N_3909);
nand U4060 (N_4060,N_3498,N_3571);
nand U4061 (N_4061,N_3637,N_3930);
nor U4062 (N_4062,N_3989,N_3529);
nor U4063 (N_4063,N_3964,N_3792);
or U4064 (N_4064,N_3732,N_3931);
or U4065 (N_4065,N_3422,N_3538);
nand U4066 (N_4066,N_3361,N_3491);
xor U4067 (N_4067,N_3925,N_3425);
and U4068 (N_4068,N_3555,N_3703);
or U4069 (N_4069,N_3272,N_3525);
and U4070 (N_4070,N_3212,N_3330);
and U4071 (N_4071,N_3372,N_3517);
nor U4072 (N_4072,N_3890,N_3143);
or U4073 (N_4073,N_3777,N_3899);
nor U4074 (N_4074,N_3120,N_3135);
nand U4075 (N_4075,N_3199,N_3762);
or U4076 (N_4076,N_3530,N_3583);
nand U4077 (N_4077,N_3250,N_3874);
or U4078 (N_4078,N_3754,N_3068);
or U4079 (N_4079,N_3543,N_3449);
nor U4080 (N_4080,N_3015,N_3674);
nand U4081 (N_4081,N_3916,N_3423);
or U4082 (N_4082,N_3304,N_3444);
or U4083 (N_4083,N_3539,N_3171);
nor U4084 (N_4084,N_3426,N_3271);
nand U4085 (N_4085,N_3326,N_3313);
or U4086 (N_4086,N_3531,N_3441);
nor U4087 (N_4087,N_3549,N_3607);
nor U4088 (N_4088,N_3815,N_3052);
nor U4089 (N_4089,N_3301,N_3118);
nor U4090 (N_4090,N_3055,N_3037);
nor U4091 (N_4091,N_3096,N_3197);
nand U4092 (N_4092,N_3870,N_3929);
or U4093 (N_4093,N_3542,N_3917);
and U4094 (N_4094,N_3606,N_3800);
nor U4095 (N_4095,N_3009,N_3764);
and U4096 (N_4096,N_3504,N_3079);
and U4097 (N_4097,N_3741,N_3962);
nand U4098 (N_4098,N_3413,N_3454);
nand U4099 (N_4099,N_3557,N_3437);
or U4100 (N_4100,N_3353,N_3231);
or U4101 (N_4101,N_3154,N_3869);
nor U4102 (N_4102,N_3357,N_3518);
nand U4103 (N_4103,N_3692,N_3230);
and U4104 (N_4104,N_3730,N_3082);
and U4105 (N_4105,N_3334,N_3968);
nand U4106 (N_4106,N_3876,N_3035);
nand U4107 (N_4107,N_3615,N_3290);
nand U4108 (N_4108,N_3864,N_3238);
nand U4109 (N_4109,N_3484,N_3104);
and U4110 (N_4110,N_3034,N_3412);
nor U4111 (N_4111,N_3826,N_3488);
or U4112 (N_4112,N_3878,N_3103);
nand U4113 (N_4113,N_3825,N_3896);
nor U4114 (N_4114,N_3291,N_3772);
or U4115 (N_4115,N_3708,N_3051);
nor U4116 (N_4116,N_3505,N_3177);
nand U4117 (N_4117,N_3681,N_3027);
and U4118 (N_4118,N_3205,N_3132);
or U4119 (N_4119,N_3248,N_3783);
nand U4120 (N_4120,N_3111,N_3045);
nand U4121 (N_4121,N_3768,N_3431);
or U4122 (N_4122,N_3880,N_3336);
nor U4123 (N_4123,N_3537,N_3220);
nand U4124 (N_4124,N_3476,N_3507);
and U4125 (N_4125,N_3329,N_3006);
nand U4126 (N_4126,N_3528,N_3625);
nand U4127 (N_4127,N_3875,N_3687);
nand U4128 (N_4128,N_3280,N_3058);
nor U4129 (N_4129,N_3577,N_3101);
xnor U4130 (N_4130,N_3714,N_3913);
nand U4131 (N_4131,N_3789,N_3829);
nor U4132 (N_4132,N_3603,N_3446);
and U4133 (N_4133,N_3524,N_3142);
and U4134 (N_4134,N_3558,N_3904);
nand U4135 (N_4135,N_3419,N_3102);
or U4136 (N_4136,N_3806,N_3655);
nand U4137 (N_4137,N_3673,N_3914);
nand U4138 (N_4138,N_3393,N_3209);
or U4139 (N_4139,N_3753,N_3892);
nor U4140 (N_4140,N_3121,N_3678);
nand U4141 (N_4141,N_3947,N_3675);
nand U4142 (N_4142,N_3303,N_3564);
and U4143 (N_4143,N_3300,N_3570);
or U4144 (N_4144,N_3253,N_3776);
nor U4145 (N_4145,N_3744,N_3287);
or U4146 (N_4146,N_3668,N_3218);
or U4147 (N_4147,N_3054,N_3801);
and U4148 (N_4148,N_3010,N_3080);
or U4149 (N_4149,N_3883,N_3575);
and U4150 (N_4150,N_3345,N_3473);
or U4151 (N_4151,N_3623,N_3288);
nand U4152 (N_4152,N_3434,N_3286);
nand U4153 (N_4153,N_3952,N_3511);
xor U4154 (N_4154,N_3684,N_3281);
nor U4155 (N_4155,N_3460,N_3889);
nand U4156 (N_4156,N_3153,N_3276);
and U4157 (N_4157,N_3131,N_3285);
nor U4158 (N_4158,N_3822,N_3723);
and U4159 (N_4159,N_3823,N_3039);
nor U4160 (N_4160,N_3314,N_3302);
nand U4161 (N_4161,N_3204,N_3907);
nand U4162 (N_4162,N_3945,N_3375);
nor U4163 (N_4163,N_3228,N_3691);
and U4164 (N_4164,N_3072,N_3657);
or U4165 (N_4165,N_3568,N_3332);
and U4166 (N_4166,N_3644,N_3267);
nand U4167 (N_4167,N_3595,N_3355);
nor U4168 (N_4168,N_3791,N_3427);
nand U4169 (N_4169,N_3922,N_3482);
nor U4170 (N_4170,N_3032,N_3191);
and U4171 (N_4171,N_3048,N_3918);
nor U4172 (N_4172,N_3294,N_3310);
and U4173 (N_4173,N_3560,N_3474);
nor U4174 (N_4174,N_3991,N_3589);
and U4175 (N_4175,N_3067,N_3411);
and U4176 (N_4176,N_3450,N_3022);
nor U4177 (N_4177,N_3873,N_3919);
nor U4178 (N_4178,N_3112,N_3399);
nand U4179 (N_4179,N_3731,N_3895);
and U4180 (N_4180,N_3696,N_3766);
or U4181 (N_4181,N_3788,N_3440);
or U4182 (N_4182,N_3984,N_3002);
or U4183 (N_4183,N_3455,N_3116);
or U4184 (N_4184,N_3282,N_3787);
or U4185 (N_4185,N_3651,N_3029);
nor U4186 (N_4186,N_3125,N_3156);
and U4187 (N_4187,N_3579,N_3698);
or U4188 (N_4188,N_3416,N_3213);
nor U4189 (N_4189,N_3232,N_3202);
and U4190 (N_4190,N_3760,N_3019);
or U4191 (N_4191,N_3382,N_3689);
and U4192 (N_4192,N_3352,N_3060);
xor U4193 (N_4193,N_3404,N_3091);
and U4194 (N_4194,N_3769,N_3780);
nand U4195 (N_4195,N_3990,N_3242);
or U4196 (N_4196,N_3988,N_3368);
nand U4197 (N_4197,N_3395,N_3499);
nor U4198 (N_4198,N_3884,N_3292);
nor U4199 (N_4199,N_3070,N_3464);
nand U4200 (N_4200,N_3033,N_3188);
nor U4201 (N_4201,N_3333,N_3515);
nor U4202 (N_4202,N_3486,N_3705);
nand U4203 (N_4203,N_3833,N_3817);
or U4204 (N_4204,N_3736,N_3140);
and U4205 (N_4205,N_3385,N_3247);
or U4206 (N_4206,N_3796,N_3406);
or U4207 (N_4207,N_3995,N_3936);
and U4208 (N_4208,N_3795,N_3738);
nand U4209 (N_4209,N_3811,N_3252);
nor U4210 (N_4210,N_3634,N_3268);
and U4211 (N_4211,N_3185,N_3315);
or U4212 (N_4212,N_3943,N_3501);
nand U4213 (N_4213,N_3612,N_3073);
nor U4214 (N_4214,N_3208,N_3835);
or U4215 (N_4215,N_3905,N_3016);
nor U4216 (N_4216,N_3804,N_3401);
and U4217 (N_4217,N_3173,N_3831);
or U4218 (N_4218,N_3781,N_3853);
nand U4219 (N_4219,N_3136,N_3462);
nand U4220 (N_4220,N_3318,N_3563);
nor U4221 (N_4221,N_3653,N_3308);
nand U4222 (N_4222,N_3614,N_3514);
nor U4223 (N_4223,N_3728,N_3840);
or U4224 (N_4224,N_3391,N_3510);
nor U4225 (N_4225,N_3089,N_3149);
nand U4226 (N_4226,N_3686,N_3470);
nor U4227 (N_4227,N_3398,N_3164);
nand U4228 (N_4228,N_3751,N_3084);
and U4229 (N_4229,N_3042,N_3323);
and U4230 (N_4230,N_3604,N_3189);
nand U4231 (N_4231,N_3812,N_3433);
or U4232 (N_4232,N_3490,N_3552);
and U4233 (N_4233,N_3963,N_3043);
nor U4234 (N_4234,N_3683,N_3926);
or U4235 (N_4235,N_3600,N_3351);
xor U4236 (N_4236,N_3710,N_3859);
and U4237 (N_4237,N_3215,N_3130);
and U4238 (N_4238,N_3064,N_3733);
nand U4239 (N_4239,N_3198,N_3316);
nand U4240 (N_4240,N_3670,N_3658);
nor U4241 (N_4241,N_3374,N_3672);
nor U4242 (N_4242,N_3855,N_3941);
and U4243 (N_4243,N_3821,N_3371);
nand U4244 (N_4244,N_3656,N_3946);
nor U4245 (N_4245,N_3296,N_3850);
nand U4246 (N_4246,N_3244,N_3523);
or U4247 (N_4247,N_3757,N_3844);
and U4248 (N_4248,N_3050,N_3881);
and U4249 (N_4249,N_3447,N_3803);
nand U4250 (N_4250,N_3877,N_3624);
nand U4251 (N_4251,N_3967,N_3325);
nor U4252 (N_4252,N_3134,N_3266);
or U4253 (N_4253,N_3834,N_3643);
nand U4254 (N_4254,N_3893,N_3115);
or U4255 (N_4255,N_3965,N_3977);
or U4256 (N_4256,N_3993,N_3233);
xor U4257 (N_4257,N_3145,N_3580);
nor U4258 (N_4258,N_3593,N_3277);
nor U4259 (N_4259,N_3157,N_3273);
and U4260 (N_4260,N_3707,N_3028);
nand U4261 (N_4261,N_3026,N_3550);
nand U4262 (N_4262,N_3295,N_3297);
xnor U4263 (N_4263,N_3137,N_3601);
and U4264 (N_4264,N_3697,N_3545);
nor U4265 (N_4265,N_3594,N_3903);
nor U4266 (N_4266,N_3389,N_3311);
and U4267 (N_4267,N_3526,N_3585);
and U4268 (N_4268,N_3251,N_3179);
and U4269 (N_4269,N_3020,N_3306);
nand U4270 (N_4270,N_3017,N_3038);
and U4271 (N_4271,N_3516,N_3265);
and U4272 (N_4272,N_3059,N_3548);
and U4273 (N_4273,N_3236,N_3192);
and U4274 (N_4274,N_3771,N_3942);
nor U4275 (N_4275,N_3613,N_3761);
or U4276 (N_4276,N_3370,N_3715);
or U4277 (N_4277,N_3489,N_3369);
nor U4278 (N_4278,N_3283,N_3097);
nand U4279 (N_4279,N_3138,N_3122);
or U4280 (N_4280,N_3196,N_3053);
nor U4281 (N_4281,N_3979,N_3481);
nor U4282 (N_4282,N_3348,N_3448);
and U4283 (N_4283,N_3360,N_3354);
and U4284 (N_4284,N_3327,N_3756);
nand U4285 (N_4285,N_3169,N_3183);
and U4286 (N_4286,N_3258,N_3223);
or U4287 (N_4287,N_3420,N_3113);
or U4288 (N_4288,N_3246,N_3956);
and U4289 (N_4289,N_3141,N_3396);
nand U4290 (N_4290,N_3901,N_3347);
or U4291 (N_4291,N_3418,N_3546);
nor U4292 (N_4292,N_3438,N_3667);
and U4293 (N_4293,N_3882,N_3008);
and U4294 (N_4294,N_3003,N_3077);
and U4295 (N_4295,N_3493,N_3765);
and U4296 (N_4296,N_3040,N_3638);
nand U4297 (N_4297,N_3627,N_3224);
nor U4298 (N_4298,N_3495,N_3566);
nand U4299 (N_4299,N_3094,N_3639);
nand U4300 (N_4300,N_3007,N_3264);
nand U4301 (N_4301,N_3468,N_3344);
or U4302 (N_4302,N_3485,N_3923);
or U4303 (N_4303,N_3774,N_3547);
nand U4304 (N_4304,N_3676,N_3773);
nor U4305 (N_4305,N_3324,N_3810);
nor U4306 (N_4306,N_3309,N_3851);
or U4307 (N_4307,N_3891,N_3214);
nand U4308 (N_4308,N_3362,N_3088);
and U4309 (N_4309,N_3133,N_3472);
nand U4310 (N_4310,N_3358,N_3417);
xnor U4311 (N_4311,N_3649,N_3650);
nand U4312 (N_4312,N_3478,N_3818);
and U4313 (N_4313,N_3709,N_3573);
or U4314 (N_4314,N_3335,N_3887);
xor U4315 (N_4315,N_3848,N_3665);
nor U4316 (N_4316,N_3734,N_3456);
nand U4317 (N_4317,N_3127,N_3986);
and U4318 (N_4318,N_3458,N_3680);
nand U4319 (N_4319,N_3932,N_3997);
nand U4320 (N_4320,N_3270,N_3699);
and U4321 (N_4321,N_3533,N_3659);
or U4322 (N_4322,N_3254,N_3935);
and U4323 (N_4323,N_3457,N_3030);
or U4324 (N_4324,N_3915,N_3342);
nand U4325 (N_4325,N_3888,N_3980);
nor U4326 (N_4326,N_3465,N_3921);
or U4327 (N_4327,N_3074,N_3828);
nor U4328 (N_4328,N_3274,N_3503);
or U4329 (N_4329,N_3105,N_3163);
nor U4330 (N_4330,N_3471,N_3535);
nor U4331 (N_4331,N_3626,N_3725);
and U4332 (N_4332,N_3386,N_3167);
or U4333 (N_4333,N_3284,N_3720);
or U4334 (N_4334,N_3178,N_3816);
nor U4335 (N_4335,N_3908,N_3307);
nand U4336 (N_4336,N_3727,N_3827);
xnor U4337 (N_4337,N_3814,N_3857);
nand U4338 (N_4338,N_3763,N_3629);
or U4339 (N_4339,N_3496,N_3379);
or U4340 (N_4340,N_3502,N_3380);
and U4341 (N_4341,N_3556,N_3597);
or U4342 (N_4342,N_3906,N_3718);
nand U4343 (N_4343,N_3085,N_3578);
nand U4344 (N_4344,N_3621,N_3770);
or U4345 (N_4345,N_3513,N_3802);
and U4346 (N_4346,N_3206,N_3747);
nand U4347 (N_4347,N_3591,N_3959);
nor U4348 (N_4348,N_3971,N_3565);
or U4349 (N_4349,N_3193,N_3036);
and U4350 (N_4350,N_3712,N_3852);
and U4351 (N_4351,N_3469,N_3520);
nand U4352 (N_4352,N_3415,N_3782);
nor U4353 (N_4353,N_3717,N_3711);
nand U4354 (N_4354,N_3602,N_3245);
or U4355 (N_4355,N_3958,N_3588);
nor U4356 (N_4356,N_3910,N_3534);
nand U4357 (N_4357,N_3405,N_3180);
and U4358 (N_4358,N_3660,N_3161);
nand U4359 (N_4359,N_3532,N_3544);
and U4360 (N_4360,N_3900,N_3222);
or U4361 (N_4361,N_3092,N_3576);
and U4362 (N_4362,N_3182,N_3584);
nor U4363 (N_4363,N_3424,N_3726);
nand U4364 (N_4364,N_3739,N_3114);
nand U4365 (N_4365,N_3226,N_3078);
or U4366 (N_4366,N_3808,N_3809);
nand U4367 (N_4367,N_3436,N_3713);
or U4368 (N_4368,N_3973,N_3693);
or U4369 (N_4369,N_3381,N_3797);
nor U4370 (N_4370,N_3275,N_3011);
and U4371 (N_4371,N_3057,N_3066);
nor U4372 (N_4372,N_3652,N_3217);
or U4373 (N_4373,N_3508,N_3158);
and U4374 (N_4374,N_3729,N_3794);
and U4375 (N_4375,N_3722,N_3225);
and U4376 (N_4376,N_3126,N_3758);
nor U4377 (N_4377,N_3661,N_3319);
nand U4378 (N_4378,N_3845,N_3093);
nor U4379 (N_4379,N_3858,N_3021);
and U4380 (N_4380,N_3373,N_3562);
and U4381 (N_4381,N_3976,N_3086);
nor U4382 (N_4382,N_3201,N_3969);
nor U4383 (N_4383,N_3572,N_3950);
or U4384 (N_4384,N_3257,N_3972);
nor U4385 (N_4385,N_3955,N_3541);
nor U4386 (N_4386,N_3839,N_3234);
or U4387 (N_4387,N_3981,N_3949);
and U4388 (N_4388,N_3459,N_3590);
nand U4389 (N_4389,N_3779,N_3863);
nor U4390 (N_4390,N_3394,N_3421);
or U4391 (N_4391,N_3982,N_3087);
and U4392 (N_4392,N_3047,N_3837);
or U4393 (N_4393,N_3467,N_3740);
and U4394 (N_4394,N_3522,N_3790);
nand U4395 (N_4395,N_3049,N_3365);
nor U4396 (N_4396,N_3071,N_3843);
or U4397 (N_4397,N_3001,N_3025);
or U4398 (N_4398,N_3475,N_3452);
and U4399 (N_4399,N_3933,N_3885);
or U4400 (N_4400,N_3269,N_3150);
nand U4401 (N_4401,N_3759,N_3934);
nand U4402 (N_4402,N_3957,N_3124);
nand U4403 (N_4403,N_3239,N_3194);
and U4404 (N_4404,N_3506,N_3605);
or U4405 (N_4405,N_3312,N_3099);
nand U4406 (N_4406,N_3174,N_3356);
and U4407 (N_4407,N_3497,N_3824);
or U4408 (N_4408,N_3966,N_3451);
or U4409 (N_4409,N_3872,N_3635);
nor U4410 (N_4410,N_3152,N_3871);
or U4411 (N_4411,N_3477,N_3392);
and U4412 (N_4412,N_3677,N_3123);
or U4413 (N_4413,N_3328,N_3151);
and U4414 (N_4414,N_3911,N_3521);
and U4415 (N_4415,N_3237,N_3014);
and U4416 (N_4416,N_3700,N_3592);
nor U4417 (N_4417,N_3492,N_3536);
nand U4418 (N_4418,N_3611,N_3975);
xnor U4419 (N_4419,N_3186,N_3846);
xor U4420 (N_4420,N_3587,N_3960);
nand U4421 (N_4421,N_3861,N_3343);
or U4422 (N_4422,N_3166,N_3632);
or U4423 (N_4423,N_3387,N_3259);
nor U4424 (N_4424,N_3633,N_3184);
nand U4425 (N_4425,N_3642,N_3317);
nand U4426 (N_4426,N_3466,N_3894);
nor U4427 (N_4427,N_3701,N_3190);
or U4428 (N_4428,N_3195,N_3403);
or U4429 (N_4429,N_3162,N_3081);
or U4430 (N_4430,N_3664,N_3263);
or U4431 (N_4431,N_3938,N_3868);
nor U4432 (N_4432,N_3830,N_3181);
or U4433 (N_4433,N_3841,N_3527);
or U4434 (N_4434,N_3090,N_3742);
or U4435 (N_4435,N_3261,N_3069);
nor U4436 (N_4436,N_3961,N_3108);
and U4437 (N_4437,N_3784,N_3119);
and U4438 (N_4438,N_3388,N_3724);
and U4439 (N_4439,N_3359,N_3645);
and U4440 (N_4440,N_3483,N_3409);
nor U4441 (N_4441,N_3640,N_3569);
and U4442 (N_4442,N_3937,N_3445);
and U4443 (N_4443,N_3480,N_3860);
and U4444 (N_4444,N_3755,N_3832);
nand U4445 (N_4445,N_3743,N_3176);
nor U4446 (N_4446,N_3785,N_3798);
nand U4447 (N_4447,N_3849,N_3630);
or U4448 (N_4448,N_3939,N_3211);
nand U4449 (N_4449,N_3775,N_3663);
and U4450 (N_4450,N_3679,N_3061);
and U4451 (N_4451,N_3574,N_3512);
nand U4452 (N_4452,N_3688,N_3842);
and U4453 (N_4453,N_3551,N_3567);
nand U4454 (N_4454,N_3553,N_3005);
nand U4455 (N_4455,N_3160,N_3836);
or U4456 (N_4456,N_3999,N_3397);
and U4457 (N_4457,N_3430,N_3168);
nor U4458 (N_4458,N_3694,N_3620);
and U4459 (N_4459,N_3243,N_3778);
and U4460 (N_4460,N_3255,N_3807);
nand U4461 (N_4461,N_3175,N_3428);
or U4462 (N_4462,N_3147,N_3331);
nand U4463 (N_4463,N_3221,N_3383);
or U4464 (N_4464,N_3346,N_3494);
nand U4465 (N_4465,N_3617,N_3928);
nor U4466 (N_4466,N_3646,N_3666);
or U4467 (N_4467,N_3813,N_3479);
or U4468 (N_4468,N_3429,N_3056);
and U4469 (N_4469,N_3439,N_3083);
nor U4470 (N_4470,N_3453,N_3647);
nand U4471 (N_4471,N_3998,N_3376);
and U4472 (N_4472,N_3363,N_3098);
or U4473 (N_4473,N_3695,N_3210);
or U4474 (N_4474,N_3838,N_3992);
nor U4475 (N_4475,N_3648,N_3793);
or U4476 (N_4476,N_3628,N_3669);
nand U4477 (N_4477,N_3920,N_3596);
or U4478 (N_4478,N_3235,N_3799);
or U4479 (N_4479,N_3559,N_3554);
nor U4480 (N_4480,N_3500,N_3867);
and U4481 (N_4481,N_3367,N_3129);
or U4482 (N_4482,N_3706,N_3340);
nor U4483 (N_4483,N_3139,N_3586);
and U4484 (N_4484,N_3636,N_3024);
nand U4485 (N_4485,N_3207,N_3107);
and U4486 (N_4486,N_3745,N_3561);
or U4487 (N_4487,N_3364,N_3902);
nor U4488 (N_4488,N_3752,N_3407);
nor U4489 (N_4489,N_3260,N_3487);
and U4490 (N_4490,N_3062,N_3735);
nor U4491 (N_4491,N_3985,N_3219);
nor U4492 (N_4492,N_3598,N_3509);
nand U4493 (N_4493,N_3249,N_3410);
and U4494 (N_4494,N_3063,N_3044);
and U4495 (N_4495,N_3117,N_3216);
nand U4496 (N_4496,N_3599,N_3289);
nand U4497 (N_4497,N_3748,N_3987);
nor U4498 (N_4498,N_3408,N_3983);
nand U4499 (N_4499,N_3012,N_3944);
nor U4500 (N_4500,N_3771,N_3825);
or U4501 (N_4501,N_3949,N_3626);
and U4502 (N_4502,N_3974,N_3512);
nand U4503 (N_4503,N_3373,N_3165);
nor U4504 (N_4504,N_3129,N_3774);
and U4505 (N_4505,N_3124,N_3584);
and U4506 (N_4506,N_3982,N_3599);
and U4507 (N_4507,N_3234,N_3361);
and U4508 (N_4508,N_3203,N_3375);
and U4509 (N_4509,N_3299,N_3200);
nor U4510 (N_4510,N_3152,N_3043);
nand U4511 (N_4511,N_3129,N_3512);
xnor U4512 (N_4512,N_3633,N_3350);
xnor U4513 (N_4513,N_3952,N_3823);
nor U4514 (N_4514,N_3736,N_3512);
nor U4515 (N_4515,N_3728,N_3771);
nand U4516 (N_4516,N_3748,N_3306);
nand U4517 (N_4517,N_3587,N_3513);
nor U4518 (N_4518,N_3600,N_3576);
or U4519 (N_4519,N_3321,N_3128);
nor U4520 (N_4520,N_3756,N_3460);
nand U4521 (N_4521,N_3875,N_3465);
nor U4522 (N_4522,N_3074,N_3785);
and U4523 (N_4523,N_3108,N_3559);
nand U4524 (N_4524,N_3741,N_3495);
nand U4525 (N_4525,N_3273,N_3573);
nor U4526 (N_4526,N_3980,N_3048);
or U4527 (N_4527,N_3769,N_3851);
nand U4528 (N_4528,N_3655,N_3197);
or U4529 (N_4529,N_3491,N_3873);
nor U4530 (N_4530,N_3065,N_3657);
or U4531 (N_4531,N_3124,N_3063);
or U4532 (N_4532,N_3322,N_3422);
nor U4533 (N_4533,N_3175,N_3665);
and U4534 (N_4534,N_3471,N_3096);
nor U4535 (N_4535,N_3303,N_3305);
nand U4536 (N_4536,N_3484,N_3632);
nand U4537 (N_4537,N_3324,N_3056);
and U4538 (N_4538,N_3711,N_3099);
nand U4539 (N_4539,N_3293,N_3038);
nand U4540 (N_4540,N_3198,N_3099);
and U4541 (N_4541,N_3731,N_3190);
or U4542 (N_4542,N_3671,N_3591);
nor U4543 (N_4543,N_3807,N_3001);
and U4544 (N_4544,N_3072,N_3547);
and U4545 (N_4545,N_3920,N_3945);
nand U4546 (N_4546,N_3610,N_3830);
and U4547 (N_4547,N_3978,N_3316);
or U4548 (N_4548,N_3365,N_3505);
or U4549 (N_4549,N_3580,N_3963);
nand U4550 (N_4550,N_3396,N_3774);
nor U4551 (N_4551,N_3062,N_3976);
and U4552 (N_4552,N_3603,N_3652);
or U4553 (N_4553,N_3411,N_3884);
and U4554 (N_4554,N_3155,N_3635);
and U4555 (N_4555,N_3203,N_3229);
and U4556 (N_4556,N_3720,N_3671);
nor U4557 (N_4557,N_3541,N_3817);
xor U4558 (N_4558,N_3027,N_3369);
nand U4559 (N_4559,N_3321,N_3612);
or U4560 (N_4560,N_3908,N_3737);
or U4561 (N_4561,N_3857,N_3683);
nor U4562 (N_4562,N_3097,N_3262);
nor U4563 (N_4563,N_3845,N_3473);
nor U4564 (N_4564,N_3472,N_3356);
or U4565 (N_4565,N_3318,N_3425);
or U4566 (N_4566,N_3535,N_3974);
or U4567 (N_4567,N_3465,N_3359);
or U4568 (N_4568,N_3422,N_3780);
nor U4569 (N_4569,N_3596,N_3196);
nand U4570 (N_4570,N_3147,N_3350);
nand U4571 (N_4571,N_3850,N_3909);
nand U4572 (N_4572,N_3057,N_3573);
or U4573 (N_4573,N_3745,N_3139);
nand U4574 (N_4574,N_3379,N_3032);
or U4575 (N_4575,N_3039,N_3326);
nor U4576 (N_4576,N_3439,N_3550);
nand U4577 (N_4577,N_3526,N_3788);
nand U4578 (N_4578,N_3382,N_3338);
nand U4579 (N_4579,N_3992,N_3010);
or U4580 (N_4580,N_3617,N_3398);
and U4581 (N_4581,N_3968,N_3232);
nor U4582 (N_4582,N_3918,N_3075);
nor U4583 (N_4583,N_3290,N_3962);
nand U4584 (N_4584,N_3801,N_3992);
nor U4585 (N_4585,N_3793,N_3790);
or U4586 (N_4586,N_3735,N_3381);
or U4587 (N_4587,N_3860,N_3613);
and U4588 (N_4588,N_3898,N_3988);
or U4589 (N_4589,N_3886,N_3626);
nand U4590 (N_4590,N_3046,N_3933);
nor U4591 (N_4591,N_3458,N_3483);
or U4592 (N_4592,N_3817,N_3504);
nor U4593 (N_4593,N_3352,N_3478);
nand U4594 (N_4594,N_3023,N_3894);
and U4595 (N_4595,N_3938,N_3306);
and U4596 (N_4596,N_3790,N_3474);
nand U4597 (N_4597,N_3865,N_3708);
nor U4598 (N_4598,N_3341,N_3966);
and U4599 (N_4599,N_3229,N_3983);
or U4600 (N_4600,N_3965,N_3836);
nand U4601 (N_4601,N_3681,N_3149);
nand U4602 (N_4602,N_3358,N_3301);
nand U4603 (N_4603,N_3253,N_3649);
or U4604 (N_4604,N_3973,N_3578);
or U4605 (N_4605,N_3278,N_3279);
nand U4606 (N_4606,N_3542,N_3736);
and U4607 (N_4607,N_3157,N_3783);
nor U4608 (N_4608,N_3441,N_3387);
nand U4609 (N_4609,N_3525,N_3025);
and U4610 (N_4610,N_3403,N_3160);
nand U4611 (N_4611,N_3356,N_3850);
nor U4612 (N_4612,N_3761,N_3245);
nor U4613 (N_4613,N_3332,N_3350);
and U4614 (N_4614,N_3448,N_3171);
and U4615 (N_4615,N_3247,N_3782);
nor U4616 (N_4616,N_3611,N_3360);
nand U4617 (N_4617,N_3538,N_3226);
nand U4618 (N_4618,N_3677,N_3579);
and U4619 (N_4619,N_3151,N_3829);
xnor U4620 (N_4620,N_3077,N_3744);
and U4621 (N_4621,N_3522,N_3789);
nor U4622 (N_4622,N_3510,N_3780);
or U4623 (N_4623,N_3257,N_3441);
nor U4624 (N_4624,N_3002,N_3072);
nor U4625 (N_4625,N_3008,N_3795);
nand U4626 (N_4626,N_3707,N_3844);
and U4627 (N_4627,N_3091,N_3803);
and U4628 (N_4628,N_3109,N_3497);
nand U4629 (N_4629,N_3174,N_3058);
nor U4630 (N_4630,N_3990,N_3560);
and U4631 (N_4631,N_3011,N_3724);
or U4632 (N_4632,N_3043,N_3262);
and U4633 (N_4633,N_3962,N_3102);
nand U4634 (N_4634,N_3978,N_3682);
nor U4635 (N_4635,N_3676,N_3976);
and U4636 (N_4636,N_3948,N_3851);
or U4637 (N_4637,N_3431,N_3666);
or U4638 (N_4638,N_3573,N_3937);
or U4639 (N_4639,N_3535,N_3051);
xnor U4640 (N_4640,N_3121,N_3529);
or U4641 (N_4641,N_3277,N_3677);
nor U4642 (N_4642,N_3957,N_3495);
or U4643 (N_4643,N_3534,N_3784);
and U4644 (N_4644,N_3323,N_3523);
nor U4645 (N_4645,N_3713,N_3368);
nor U4646 (N_4646,N_3612,N_3237);
nor U4647 (N_4647,N_3120,N_3059);
nand U4648 (N_4648,N_3230,N_3821);
and U4649 (N_4649,N_3928,N_3959);
nor U4650 (N_4650,N_3859,N_3037);
or U4651 (N_4651,N_3168,N_3274);
and U4652 (N_4652,N_3872,N_3258);
or U4653 (N_4653,N_3005,N_3105);
or U4654 (N_4654,N_3538,N_3949);
nor U4655 (N_4655,N_3538,N_3630);
xor U4656 (N_4656,N_3187,N_3332);
or U4657 (N_4657,N_3049,N_3171);
nand U4658 (N_4658,N_3984,N_3135);
nand U4659 (N_4659,N_3119,N_3344);
and U4660 (N_4660,N_3489,N_3665);
or U4661 (N_4661,N_3297,N_3873);
nand U4662 (N_4662,N_3046,N_3831);
nand U4663 (N_4663,N_3451,N_3759);
or U4664 (N_4664,N_3657,N_3183);
and U4665 (N_4665,N_3440,N_3918);
nor U4666 (N_4666,N_3040,N_3149);
nor U4667 (N_4667,N_3415,N_3976);
or U4668 (N_4668,N_3464,N_3175);
and U4669 (N_4669,N_3516,N_3102);
nand U4670 (N_4670,N_3251,N_3741);
nand U4671 (N_4671,N_3320,N_3726);
and U4672 (N_4672,N_3988,N_3521);
nand U4673 (N_4673,N_3147,N_3178);
nand U4674 (N_4674,N_3362,N_3718);
or U4675 (N_4675,N_3256,N_3143);
or U4676 (N_4676,N_3100,N_3912);
and U4677 (N_4677,N_3661,N_3107);
nand U4678 (N_4678,N_3367,N_3995);
nand U4679 (N_4679,N_3558,N_3534);
nor U4680 (N_4680,N_3202,N_3990);
and U4681 (N_4681,N_3046,N_3123);
nor U4682 (N_4682,N_3804,N_3955);
nor U4683 (N_4683,N_3843,N_3322);
or U4684 (N_4684,N_3105,N_3247);
nand U4685 (N_4685,N_3970,N_3232);
nand U4686 (N_4686,N_3017,N_3773);
nor U4687 (N_4687,N_3598,N_3801);
or U4688 (N_4688,N_3218,N_3947);
nor U4689 (N_4689,N_3669,N_3350);
and U4690 (N_4690,N_3248,N_3502);
nand U4691 (N_4691,N_3204,N_3101);
nand U4692 (N_4692,N_3001,N_3290);
and U4693 (N_4693,N_3081,N_3509);
nand U4694 (N_4694,N_3227,N_3549);
xor U4695 (N_4695,N_3807,N_3327);
nand U4696 (N_4696,N_3209,N_3554);
and U4697 (N_4697,N_3345,N_3013);
nand U4698 (N_4698,N_3723,N_3803);
or U4699 (N_4699,N_3362,N_3010);
nor U4700 (N_4700,N_3151,N_3270);
nand U4701 (N_4701,N_3184,N_3536);
and U4702 (N_4702,N_3425,N_3328);
nand U4703 (N_4703,N_3865,N_3105);
or U4704 (N_4704,N_3742,N_3349);
nand U4705 (N_4705,N_3040,N_3396);
xor U4706 (N_4706,N_3809,N_3245);
nand U4707 (N_4707,N_3417,N_3993);
nand U4708 (N_4708,N_3026,N_3136);
nand U4709 (N_4709,N_3405,N_3009);
or U4710 (N_4710,N_3870,N_3754);
and U4711 (N_4711,N_3566,N_3899);
nor U4712 (N_4712,N_3929,N_3465);
or U4713 (N_4713,N_3219,N_3720);
nor U4714 (N_4714,N_3344,N_3267);
nand U4715 (N_4715,N_3539,N_3033);
and U4716 (N_4716,N_3151,N_3723);
nor U4717 (N_4717,N_3204,N_3107);
xnor U4718 (N_4718,N_3254,N_3559);
nand U4719 (N_4719,N_3552,N_3647);
nand U4720 (N_4720,N_3654,N_3487);
nor U4721 (N_4721,N_3979,N_3034);
nand U4722 (N_4722,N_3828,N_3241);
nor U4723 (N_4723,N_3228,N_3649);
and U4724 (N_4724,N_3950,N_3426);
and U4725 (N_4725,N_3424,N_3897);
and U4726 (N_4726,N_3788,N_3960);
nand U4727 (N_4727,N_3021,N_3915);
nand U4728 (N_4728,N_3202,N_3733);
or U4729 (N_4729,N_3876,N_3786);
or U4730 (N_4730,N_3492,N_3052);
nor U4731 (N_4731,N_3560,N_3394);
and U4732 (N_4732,N_3293,N_3345);
or U4733 (N_4733,N_3265,N_3497);
nand U4734 (N_4734,N_3877,N_3936);
nor U4735 (N_4735,N_3901,N_3284);
nor U4736 (N_4736,N_3358,N_3871);
and U4737 (N_4737,N_3405,N_3668);
nor U4738 (N_4738,N_3547,N_3896);
nor U4739 (N_4739,N_3629,N_3875);
or U4740 (N_4740,N_3061,N_3555);
nor U4741 (N_4741,N_3367,N_3030);
or U4742 (N_4742,N_3930,N_3713);
and U4743 (N_4743,N_3508,N_3099);
nor U4744 (N_4744,N_3867,N_3752);
and U4745 (N_4745,N_3289,N_3392);
nand U4746 (N_4746,N_3718,N_3266);
and U4747 (N_4747,N_3294,N_3830);
and U4748 (N_4748,N_3263,N_3897);
nor U4749 (N_4749,N_3011,N_3931);
nand U4750 (N_4750,N_3619,N_3585);
nand U4751 (N_4751,N_3313,N_3501);
nand U4752 (N_4752,N_3710,N_3286);
or U4753 (N_4753,N_3193,N_3867);
and U4754 (N_4754,N_3168,N_3566);
or U4755 (N_4755,N_3999,N_3998);
or U4756 (N_4756,N_3119,N_3008);
nor U4757 (N_4757,N_3960,N_3353);
or U4758 (N_4758,N_3385,N_3981);
and U4759 (N_4759,N_3578,N_3780);
xnor U4760 (N_4760,N_3270,N_3063);
nand U4761 (N_4761,N_3943,N_3036);
xnor U4762 (N_4762,N_3252,N_3531);
or U4763 (N_4763,N_3535,N_3302);
and U4764 (N_4764,N_3507,N_3211);
nor U4765 (N_4765,N_3878,N_3007);
nor U4766 (N_4766,N_3271,N_3844);
nor U4767 (N_4767,N_3740,N_3122);
nand U4768 (N_4768,N_3831,N_3929);
nor U4769 (N_4769,N_3823,N_3014);
and U4770 (N_4770,N_3524,N_3396);
or U4771 (N_4771,N_3227,N_3565);
and U4772 (N_4772,N_3482,N_3082);
or U4773 (N_4773,N_3096,N_3133);
nor U4774 (N_4774,N_3881,N_3222);
nor U4775 (N_4775,N_3670,N_3578);
and U4776 (N_4776,N_3998,N_3414);
or U4777 (N_4777,N_3958,N_3015);
or U4778 (N_4778,N_3495,N_3347);
nand U4779 (N_4779,N_3609,N_3451);
nand U4780 (N_4780,N_3252,N_3333);
nor U4781 (N_4781,N_3003,N_3517);
and U4782 (N_4782,N_3298,N_3508);
or U4783 (N_4783,N_3450,N_3820);
and U4784 (N_4784,N_3060,N_3514);
nand U4785 (N_4785,N_3201,N_3226);
and U4786 (N_4786,N_3030,N_3615);
or U4787 (N_4787,N_3695,N_3124);
or U4788 (N_4788,N_3398,N_3155);
nand U4789 (N_4789,N_3720,N_3122);
nor U4790 (N_4790,N_3877,N_3859);
nor U4791 (N_4791,N_3302,N_3195);
nor U4792 (N_4792,N_3347,N_3834);
or U4793 (N_4793,N_3437,N_3973);
nand U4794 (N_4794,N_3536,N_3326);
nand U4795 (N_4795,N_3124,N_3087);
nor U4796 (N_4796,N_3987,N_3117);
nand U4797 (N_4797,N_3385,N_3318);
nor U4798 (N_4798,N_3158,N_3413);
nand U4799 (N_4799,N_3974,N_3376);
nor U4800 (N_4800,N_3473,N_3470);
nand U4801 (N_4801,N_3155,N_3068);
or U4802 (N_4802,N_3506,N_3070);
and U4803 (N_4803,N_3324,N_3853);
or U4804 (N_4804,N_3913,N_3536);
and U4805 (N_4805,N_3227,N_3970);
nor U4806 (N_4806,N_3000,N_3940);
nor U4807 (N_4807,N_3861,N_3485);
or U4808 (N_4808,N_3283,N_3738);
or U4809 (N_4809,N_3777,N_3801);
and U4810 (N_4810,N_3959,N_3372);
nand U4811 (N_4811,N_3723,N_3473);
or U4812 (N_4812,N_3411,N_3319);
or U4813 (N_4813,N_3740,N_3301);
and U4814 (N_4814,N_3538,N_3322);
or U4815 (N_4815,N_3906,N_3946);
nand U4816 (N_4816,N_3948,N_3738);
nand U4817 (N_4817,N_3639,N_3224);
nor U4818 (N_4818,N_3839,N_3677);
nor U4819 (N_4819,N_3773,N_3640);
or U4820 (N_4820,N_3736,N_3920);
and U4821 (N_4821,N_3676,N_3811);
and U4822 (N_4822,N_3638,N_3204);
and U4823 (N_4823,N_3614,N_3345);
and U4824 (N_4824,N_3010,N_3780);
nand U4825 (N_4825,N_3886,N_3034);
nor U4826 (N_4826,N_3964,N_3623);
nand U4827 (N_4827,N_3440,N_3845);
or U4828 (N_4828,N_3749,N_3969);
nor U4829 (N_4829,N_3355,N_3913);
nand U4830 (N_4830,N_3025,N_3971);
nor U4831 (N_4831,N_3168,N_3333);
or U4832 (N_4832,N_3458,N_3498);
nor U4833 (N_4833,N_3200,N_3497);
or U4834 (N_4834,N_3956,N_3112);
or U4835 (N_4835,N_3956,N_3220);
nor U4836 (N_4836,N_3245,N_3452);
nand U4837 (N_4837,N_3132,N_3094);
and U4838 (N_4838,N_3348,N_3761);
nor U4839 (N_4839,N_3775,N_3169);
or U4840 (N_4840,N_3971,N_3120);
and U4841 (N_4841,N_3605,N_3412);
and U4842 (N_4842,N_3089,N_3349);
nand U4843 (N_4843,N_3169,N_3035);
and U4844 (N_4844,N_3987,N_3296);
and U4845 (N_4845,N_3764,N_3022);
or U4846 (N_4846,N_3756,N_3806);
nor U4847 (N_4847,N_3219,N_3344);
or U4848 (N_4848,N_3309,N_3296);
nand U4849 (N_4849,N_3234,N_3967);
and U4850 (N_4850,N_3947,N_3939);
nor U4851 (N_4851,N_3229,N_3007);
nor U4852 (N_4852,N_3723,N_3212);
or U4853 (N_4853,N_3049,N_3425);
and U4854 (N_4854,N_3933,N_3851);
or U4855 (N_4855,N_3820,N_3622);
nand U4856 (N_4856,N_3377,N_3437);
nand U4857 (N_4857,N_3236,N_3256);
or U4858 (N_4858,N_3447,N_3938);
and U4859 (N_4859,N_3079,N_3316);
and U4860 (N_4860,N_3766,N_3056);
nand U4861 (N_4861,N_3520,N_3144);
nor U4862 (N_4862,N_3662,N_3381);
and U4863 (N_4863,N_3564,N_3120);
or U4864 (N_4864,N_3505,N_3198);
nor U4865 (N_4865,N_3621,N_3522);
nor U4866 (N_4866,N_3279,N_3685);
or U4867 (N_4867,N_3844,N_3166);
and U4868 (N_4868,N_3995,N_3118);
or U4869 (N_4869,N_3065,N_3986);
nand U4870 (N_4870,N_3284,N_3231);
nor U4871 (N_4871,N_3382,N_3241);
nand U4872 (N_4872,N_3743,N_3419);
nor U4873 (N_4873,N_3325,N_3175);
nand U4874 (N_4874,N_3271,N_3267);
or U4875 (N_4875,N_3690,N_3962);
nor U4876 (N_4876,N_3006,N_3422);
and U4877 (N_4877,N_3636,N_3138);
nor U4878 (N_4878,N_3273,N_3979);
nand U4879 (N_4879,N_3408,N_3366);
and U4880 (N_4880,N_3117,N_3890);
nand U4881 (N_4881,N_3735,N_3184);
nand U4882 (N_4882,N_3333,N_3748);
nand U4883 (N_4883,N_3984,N_3896);
nor U4884 (N_4884,N_3017,N_3483);
nor U4885 (N_4885,N_3042,N_3720);
or U4886 (N_4886,N_3477,N_3151);
and U4887 (N_4887,N_3132,N_3536);
and U4888 (N_4888,N_3104,N_3959);
or U4889 (N_4889,N_3060,N_3804);
nor U4890 (N_4890,N_3703,N_3901);
nor U4891 (N_4891,N_3853,N_3033);
nor U4892 (N_4892,N_3244,N_3874);
nand U4893 (N_4893,N_3880,N_3494);
nor U4894 (N_4894,N_3973,N_3017);
or U4895 (N_4895,N_3800,N_3516);
nor U4896 (N_4896,N_3278,N_3863);
and U4897 (N_4897,N_3606,N_3103);
nor U4898 (N_4898,N_3066,N_3346);
nor U4899 (N_4899,N_3904,N_3280);
or U4900 (N_4900,N_3390,N_3129);
nor U4901 (N_4901,N_3519,N_3446);
nand U4902 (N_4902,N_3217,N_3676);
and U4903 (N_4903,N_3906,N_3306);
and U4904 (N_4904,N_3858,N_3470);
xnor U4905 (N_4905,N_3805,N_3667);
or U4906 (N_4906,N_3317,N_3366);
or U4907 (N_4907,N_3918,N_3346);
and U4908 (N_4908,N_3586,N_3269);
or U4909 (N_4909,N_3244,N_3887);
and U4910 (N_4910,N_3541,N_3314);
nor U4911 (N_4911,N_3607,N_3539);
or U4912 (N_4912,N_3386,N_3517);
or U4913 (N_4913,N_3291,N_3563);
and U4914 (N_4914,N_3107,N_3673);
nor U4915 (N_4915,N_3192,N_3781);
nand U4916 (N_4916,N_3214,N_3457);
nor U4917 (N_4917,N_3163,N_3615);
nand U4918 (N_4918,N_3119,N_3338);
or U4919 (N_4919,N_3105,N_3905);
nand U4920 (N_4920,N_3256,N_3295);
nand U4921 (N_4921,N_3518,N_3025);
nor U4922 (N_4922,N_3757,N_3247);
nand U4923 (N_4923,N_3252,N_3002);
or U4924 (N_4924,N_3703,N_3300);
nand U4925 (N_4925,N_3643,N_3856);
nand U4926 (N_4926,N_3844,N_3282);
nand U4927 (N_4927,N_3358,N_3433);
and U4928 (N_4928,N_3965,N_3673);
or U4929 (N_4929,N_3785,N_3209);
or U4930 (N_4930,N_3520,N_3230);
nand U4931 (N_4931,N_3091,N_3960);
nor U4932 (N_4932,N_3265,N_3196);
or U4933 (N_4933,N_3691,N_3037);
or U4934 (N_4934,N_3714,N_3427);
nand U4935 (N_4935,N_3893,N_3357);
nand U4936 (N_4936,N_3160,N_3856);
nand U4937 (N_4937,N_3911,N_3193);
nor U4938 (N_4938,N_3512,N_3236);
nor U4939 (N_4939,N_3705,N_3176);
nand U4940 (N_4940,N_3200,N_3675);
and U4941 (N_4941,N_3762,N_3984);
and U4942 (N_4942,N_3614,N_3775);
or U4943 (N_4943,N_3817,N_3732);
nor U4944 (N_4944,N_3990,N_3042);
nor U4945 (N_4945,N_3870,N_3152);
xnor U4946 (N_4946,N_3540,N_3764);
nand U4947 (N_4947,N_3044,N_3247);
nand U4948 (N_4948,N_3823,N_3780);
nand U4949 (N_4949,N_3521,N_3895);
nor U4950 (N_4950,N_3587,N_3883);
nor U4951 (N_4951,N_3985,N_3347);
or U4952 (N_4952,N_3278,N_3403);
or U4953 (N_4953,N_3755,N_3850);
or U4954 (N_4954,N_3974,N_3679);
nand U4955 (N_4955,N_3060,N_3206);
and U4956 (N_4956,N_3779,N_3044);
nor U4957 (N_4957,N_3176,N_3009);
nor U4958 (N_4958,N_3504,N_3609);
nand U4959 (N_4959,N_3572,N_3558);
or U4960 (N_4960,N_3942,N_3235);
and U4961 (N_4961,N_3475,N_3427);
or U4962 (N_4962,N_3125,N_3924);
nand U4963 (N_4963,N_3509,N_3998);
nor U4964 (N_4964,N_3862,N_3658);
or U4965 (N_4965,N_3591,N_3783);
and U4966 (N_4966,N_3647,N_3307);
nand U4967 (N_4967,N_3383,N_3718);
nand U4968 (N_4968,N_3427,N_3652);
or U4969 (N_4969,N_3961,N_3030);
nor U4970 (N_4970,N_3258,N_3501);
nand U4971 (N_4971,N_3443,N_3458);
or U4972 (N_4972,N_3861,N_3298);
nor U4973 (N_4973,N_3940,N_3004);
nor U4974 (N_4974,N_3699,N_3663);
or U4975 (N_4975,N_3957,N_3304);
and U4976 (N_4976,N_3678,N_3486);
nor U4977 (N_4977,N_3941,N_3406);
or U4978 (N_4978,N_3162,N_3503);
nand U4979 (N_4979,N_3237,N_3171);
and U4980 (N_4980,N_3021,N_3991);
nand U4981 (N_4981,N_3223,N_3611);
and U4982 (N_4982,N_3367,N_3027);
and U4983 (N_4983,N_3206,N_3485);
nand U4984 (N_4984,N_3961,N_3596);
nand U4985 (N_4985,N_3661,N_3498);
nand U4986 (N_4986,N_3382,N_3879);
or U4987 (N_4987,N_3198,N_3489);
nor U4988 (N_4988,N_3794,N_3903);
nor U4989 (N_4989,N_3593,N_3333);
and U4990 (N_4990,N_3274,N_3913);
or U4991 (N_4991,N_3875,N_3329);
and U4992 (N_4992,N_3430,N_3744);
nor U4993 (N_4993,N_3944,N_3564);
nor U4994 (N_4994,N_3897,N_3341);
nor U4995 (N_4995,N_3017,N_3119);
nor U4996 (N_4996,N_3379,N_3601);
or U4997 (N_4997,N_3749,N_3699);
or U4998 (N_4998,N_3293,N_3674);
nand U4999 (N_4999,N_3669,N_3231);
and UO_0 (O_0,N_4501,N_4612);
nor UO_1 (O_1,N_4001,N_4344);
and UO_2 (O_2,N_4912,N_4594);
or UO_3 (O_3,N_4458,N_4216);
and UO_4 (O_4,N_4184,N_4848);
or UO_5 (O_5,N_4143,N_4101);
and UO_6 (O_6,N_4632,N_4250);
and UO_7 (O_7,N_4338,N_4491);
and UO_8 (O_8,N_4092,N_4439);
and UO_9 (O_9,N_4111,N_4931);
xnor UO_10 (O_10,N_4069,N_4644);
nor UO_11 (O_11,N_4790,N_4263);
or UO_12 (O_12,N_4026,N_4811);
or UO_13 (O_13,N_4191,N_4681);
or UO_14 (O_14,N_4788,N_4964);
nor UO_15 (O_15,N_4292,N_4479);
and UO_16 (O_16,N_4300,N_4232);
nand UO_17 (O_17,N_4158,N_4499);
or UO_18 (O_18,N_4924,N_4684);
or UO_19 (O_19,N_4537,N_4055);
and UO_20 (O_20,N_4324,N_4102);
nand UO_21 (O_21,N_4891,N_4041);
and UO_22 (O_22,N_4999,N_4951);
nor UO_23 (O_23,N_4226,N_4602);
nand UO_24 (O_24,N_4792,N_4469);
nor UO_25 (O_25,N_4084,N_4463);
or UO_26 (O_26,N_4677,N_4820);
nor UO_27 (O_27,N_4554,N_4450);
or UO_28 (O_28,N_4078,N_4757);
nor UO_29 (O_29,N_4878,N_4492);
nand UO_30 (O_30,N_4853,N_4736);
nor UO_31 (O_31,N_4911,N_4424);
and UO_32 (O_32,N_4569,N_4406);
nand UO_33 (O_33,N_4875,N_4618);
or UO_34 (O_34,N_4900,N_4401);
and UO_35 (O_35,N_4634,N_4855);
nor UO_36 (O_36,N_4861,N_4393);
or UO_37 (O_37,N_4504,N_4438);
or UO_38 (O_38,N_4833,N_4986);
and UO_39 (O_39,N_4805,N_4573);
nor UO_40 (O_40,N_4712,N_4770);
and UO_41 (O_41,N_4284,N_4920);
nor UO_42 (O_42,N_4199,N_4630);
nand UO_43 (O_43,N_4601,N_4654);
nand UO_44 (O_44,N_4732,N_4985);
nor UO_45 (O_45,N_4091,N_4222);
nand UO_46 (O_46,N_4633,N_4272);
nor UO_47 (O_47,N_4256,N_4694);
nor UO_48 (O_48,N_4082,N_4160);
or UO_49 (O_49,N_4154,N_4345);
and UO_50 (O_50,N_4433,N_4476);
or UO_51 (O_51,N_4416,N_4703);
or UO_52 (O_52,N_4490,N_4827);
nand UO_53 (O_53,N_4052,N_4752);
or UO_54 (O_54,N_4954,N_4390);
and UO_55 (O_55,N_4747,N_4536);
or UO_56 (O_56,N_4238,N_4690);
or UO_57 (O_57,N_4067,N_4007);
and UO_58 (O_58,N_4127,N_4157);
nand UO_59 (O_59,N_4593,N_4898);
and UO_60 (O_60,N_4497,N_4806);
and UO_61 (O_61,N_4723,N_4085);
or UO_62 (O_62,N_4921,N_4362);
nand UO_63 (O_63,N_4043,N_4707);
or UO_64 (O_64,N_4139,N_4136);
nand UO_65 (O_65,N_4236,N_4702);
or UO_66 (O_66,N_4452,N_4231);
nor UO_67 (O_67,N_4493,N_4872);
or UO_68 (O_68,N_4600,N_4759);
or UO_69 (O_69,N_4813,N_4847);
and UO_70 (O_70,N_4241,N_4242);
or UO_71 (O_71,N_4065,N_4926);
or UO_72 (O_72,N_4934,N_4112);
or UO_73 (O_73,N_4328,N_4560);
and UO_74 (O_74,N_4066,N_4196);
nor UO_75 (O_75,N_4090,N_4419);
and UO_76 (O_76,N_4795,N_4611);
nand UO_77 (O_77,N_4777,N_4555);
nand UO_78 (O_78,N_4378,N_4763);
nand UO_79 (O_79,N_4755,N_4247);
nand UO_80 (O_80,N_4275,N_4444);
nand UO_81 (O_81,N_4040,N_4693);
nand UO_82 (O_82,N_4809,N_4761);
nand UO_83 (O_83,N_4371,N_4787);
nand UO_84 (O_84,N_4538,N_4525);
nand UO_85 (O_85,N_4008,N_4756);
or UO_86 (O_86,N_4956,N_4183);
nand UO_87 (O_87,N_4530,N_4412);
and UO_88 (O_88,N_4322,N_4507);
nor UO_89 (O_89,N_4024,N_4987);
or UO_90 (O_90,N_4505,N_4015);
and UO_91 (O_91,N_4034,N_4613);
nor UO_92 (O_92,N_4266,N_4198);
nand UO_93 (O_93,N_4983,N_4754);
nand UO_94 (O_94,N_4385,N_4974);
nor UO_95 (O_95,N_4482,N_4785);
nor UO_96 (O_96,N_4355,N_4186);
or UO_97 (O_97,N_4121,N_4223);
or UO_98 (O_98,N_4816,N_4887);
xor UO_99 (O_99,N_4529,N_4725);
nor UO_100 (O_100,N_4152,N_4904);
and UO_101 (O_101,N_4359,N_4445);
and UO_102 (O_102,N_4721,N_4583);
nor UO_103 (O_103,N_4151,N_4510);
or UO_104 (O_104,N_4994,N_4076);
and UO_105 (O_105,N_4133,N_4739);
or UO_106 (O_106,N_4435,N_4044);
and UO_107 (O_107,N_4443,N_4549);
or UO_108 (O_108,N_4030,N_4860);
nor UO_109 (O_109,N_4336,N_4882);
and UO_110 (O_110,N_4080,N_4387);
nor UO_111 (O_111,N_4290,N_4749);
nor UO_112 (O_112,N_4957,N_4126);
and UO_113 (O_113,N_4998,N_4360);
and UO_114 (O_114,N_4706,N_4886);
nor UO_115 (O_115,N_4147,N_4893);
nor UO_116 (O_116,N_4683,N_4701);
or UO_117 (O_117,N_4794,N_4532);
nand UO_118 (O_118,N_4356,N_4029);
nand UO_119 (O_119,N_4096,N_4866);
nand UO_120 (O_120,N_4695,N_4699);
nor UO_121 (O_121,N_4167,N_4871);
or UO_122 (O_122,N_4810,N_4148);
and UO_123 (O_123,N_4016,N_4724);
or UO_124 (O_124,N_4221,N_4545);
nor UO_125 (O_125,N_4441,N_4648);
or UO_126 (O_126,N_4726,N_4837);
and UO_127 (O_127,N_4405,N_4698);
or UO_128 (O_128,N_4006,N_4367);
or UO_129 (O_129,N_4233,N_4310);
nand UO_130 (O_130,N_4487,N_4864);
nand UO_131 (O_131,N_4850,N_4046);
and UO_132 (O_132,N_4192,N_4516);
nor UO_133 (O_133,N_4717,N_4835);
or UO_134 (O_134,N_4308,N_4959);
or UO_135 (O_135,N_4885,N_4470);
nor UO_136 (O_136,N_4819,N_4834);
and UO_137 (O_137,N_4234,N_4365);
nor UO_138 (O_138,N_4585,N_4451);
nor UO_139 (O_139,N_4420,N_4169);
nand UO_140 (O_140,N_4341,N_4282);
nor UO_141 (O_141,N_4289,N_4313);
and UO_142 (O_142,N_4047,N_4201);
nand UO_143 (O_143,N_4989,N_4631);
and UO_144 (O_144,N_4992,N_4166);
nor UO_145 (O_145,N_4141,N_4366);
nor UO_146 (O_146,N_4624,N_4392);
nor UO_147 (O_147,N_4446,N_4075);
nor UO_148 (O_148,N_4863,N_4262);
or UO_149 (O_149,N_4170,N_4804);
nor UO_150 (O_150,N_4590,N_4347);
nor UO_151 (O_151,N_4927,N_4682);
or UO_152 (O_152,N_4273,N_4175);
nor UO_153 (O_153,N_4018,N_4454);
and UO_154 (O_154,N_4259,N_4883);
nor UO_155 (O_155,N_4291,N_4975);
nand UO_156 (O_156,N_4851,N_4010);
nor UO_157 (O_157,N_4017,N_4421);
nand UO_158 (O_158,N_4945,N_4908);
nand UO_159 (O_159,N_4815,N_4379);
or UO_160 (O_160,N_4824,N_4870);
or UO_161 (O_161,N_4063,N_4636);
or UO_162 (O_162,N_4240,N_4219);
or UO_163 (O_163,N_4722,N_4000);
xor UO_164 (O_164,N_4981,N_4255);
and UO_165 (O_165,N_4249,N_4727);
nand UO_166 (O_166,N_4025,N_4838);
nand UO_167 (O_167,N_4966,N_4786);
or UO_168 (O_168,N_4937,N_4942);
nor UO_169 (O_169,N_4674,N_4205);
nor UO_170 (O_170,N_4836,N_4320);
nor UO_171 (O_171,N_4528,N_4544);
and UO_172 (O_172,N_4980,N_4696);
nand UO_173 (O_173,N_4400,N_4830);
or UO_174 (O_174,N_4666,N_4109);
nor UO_175 (O_175,N_4281,N_4514);
nand UO_176 (O_176,N_4543,N_4649);
nor UO_177 (O_177,N_4991,N_4656);
and UO_178 (O_178,N_4062,N_4116);
or UO_179 (O_179,N_4880,N_4558);
and UO_180 (O_180,N_4404,N_4628);
or UO_181 (O_181,N_4352,N_4688);
nand UO_182 (O_182,N_4892,N_4896);
nor UO_183 (O_183,N_4839,N_4115);
and UO_184 (O_184,N_4224,N_4910);
nor UO_185 (O_185,N_4088,N_4070);
or UO_186 (O_186,N_4697,N_4417);
or UO_187 (O_187,N_4485,N_4735);
nor UO_188 (O_188,N_4572,N_4764);
and UO_189 (O_189,N_4331,N_4728);
nand UO_190 (O_190,N_4407,N_4237);
nand UO_191 (O_191,N_4267,N_4260);
nor UO_192 (O_192,N_4350,N_4386);
nor UO_193 (O_193,N_4276,N_4997);
nand UO_194 (O_194,N_4168,N_4494);
and UO_195 (O_195,N_4335,N_4426);
and UO_196 (O_196,N_4559,N_4225);
nor UO_197 (O_197,N_4459,N_4261);
and UO_198 (O_198,N_4581,N_4700);
or UO_199 (O_199,N_4103,N_4229);
nand UO_200 (O_200,N_4467,N_4879);
nand UO_201 (O_201,N_4120,N_4823);
nand UO_202 (O_202,N_4597,N_4039);
nand UO_203 (O_203,N_4354,N_4840);
nor UO_204 (O_204,N_4771,N_4180);
nand UO_205 (O_205,N_4129,N_4596);
and UO_206 (O_206,N_4709,N_4132);
nand UO_207 (O_207,N_4265,N_4181);
nand UO_208 (O_208,N_4174,N_4375);
or UO_209 (O_209,N_4551,N_4570);
nand UO_210 (O_210,N_4852,N_4639);
nand UO_211 (O_211,N_4455,N_4162);
nand UO_212 (O_212,N_4766,N_4302);
nand UO_213 (O_213,N_4298,N_4037);
or UO_214 (O_214,N_4213,N_4965);
and UO_215 (O_215,N_4311,N_4780);
and UO_216 (O_216,N_4486,N_4427);
nor UO_217 (O_217,N_4577,N_4217);
nor UO_218 (O_218,N_4916,N_4933);
and UO_219 (O_219,N_4932,N_4337);
and UO_220 (O_220,N_4408,N_4033);
nor UO_221 (O_221,N_4899,N_4969);
and UO_222 (O_222,N_4049,N_4915);
nand UO_223 (O_223,N_4753,N_4145);
nand UO_224 (O_224,N_4961,N_4220);
nand UO_225 (O_225,N_4193,N_4901);
nand UO_226 (O_226,N_4442,N_4607);
nand UO_227 (O_227,N_4483,N_4472);
or UO_228 (O_228,N_4527,N_4422);
nor UO_229 (O_229,N_4663,N_4984);
or UO_230 (O_230,N_4032,N_4844);
nor UO_231 (O_231,N_4051,N_4552);
nor UO_232 (O_232,N_4429,N_4448);
or UO_233 (O_233,N_4758,N_4332);
or UO_234 (O_234,N_4218,N_4351);
or UO_235 (O_235,N_4620,N_4048);
or UO_236 (O_236,N_4673,N_4176);
nor UO_237 (O_237,N_4968,N_4941);
nor UO_238 (O_238,N_4161,N_4626);
nand UO_239 (O_239,N_4520,N_4077);
or UO_240 (O_240,N_4973,N_4647);
nand UO_241 (O_241,N_4056,N_4097);
nor UO_242 (O_242,N_4153,N_4720);
nand UO_243 (O_243,N_4678,N_4163);
and UO_244 (O_244,N_4079,N_4917);
nor UO_245 (O_245,N_4312,N_4149);
or UO_246 (O_246,N_4477,N_4667);
nand UO_247 (O_247,N_4606,N_4603);
nand UO_248 (O_248,N_4093,N_4958);
nand UO_249 (O_249,N_4928,N_4150);
and UO_250 (O_250,N_4509,N_4449);
and UO_251 (O_251,N_4142,N_4475);
nor UO_252 (O_252,N_4370,N_4664);
nor UO_253 (O_253,N_4645,N_4988);
and UO_254 (O_254,N_4784,N_4277);
nor UO_255 (O_255,N_4358,N_4203);
or UO_256 (O_256,N_4854,N_4123);
nor UO_257 (O_257,N_4481,N_4506);
or UO_258 (O_258,N_4003,N_4939);
and UO_259 (O_259,N_4253,N_4227);
and UO_260 (O_260,N_4104,N_4173);
nand UO_261 (O_261,N_4087,N_4436);
nor UO_262 (O_262,N_4579,N_4005);
or UO_263 (O_263,N_4762,N_4995);
or UO_264 (O_264,N_4881,N_4778);
or UO_265 (O_265,N_4553,N_4296);
nor UO_266 (O_266,N_4189,N_4464);
and UO_267 (O_267,N_4542,N_4923);
and UO_268 (O_268,N_4742,N_4270);
or UO_269 (O_269,N_4897,N_4394);
and UO_270 (O_270,N_4676,N_4867);
nand UO_271 (O_271,N_4307,N_4212);
and UO_272 (O_272,N_4710,N_4769);
or UO_273 (O_273,N_4172,N_4598);
nand UO_274 (O_274,N_4114,N_4019);
or UO_275 (O_275,N_4230,N_4658);
and UO_276 (O_276,N_4615,N_4204);
or UO_277 (O_277,N_4306,N_4182);
nand UO_278 (O_278,N_4021,N_4369);
or UO_279 (O_279,N_4295,N_4629);
nor UO_280 (O_280,N_4976,N_4605);
nand UO_281 (O_281,N_4713,N_4465);
nand UO_282 (O_282,N_4135,N_4869);
nor UO_283 (O_283,N_4190,N_4905);
nand UO_284 (O_284,N_4868,N_4380);
nor UO_285 (O_285,N_4488,N_4215);
nand UO_286 (O_286,N_4094,N_4943);
nor UO_287 (O_287,N_4100,N_4319);
nand UO_288 (O_288,N_4550,N_4675);
and UO_289 (O_289,N_4361,N_4944);
xor UO_290 (O_290,N_4567,N_4540);
and UO_291 (O_291,N_4089,N_4478);
nor UO_292 (O_292,N_4705,N_4202);
or UO_293 (O_293,N_4519,N_4963);
nand UO_294 (O_294,N_4274,N_4125);
or UO_295 (O_295,N_4171,N_4803);
and UO_296 (O_296,N_4789,N_4244);
xor UO_297 (O_297,N_4164,N_4760);
and UO_298 (O_298,N_4188,N_4971);
nor UO_299 (O_299,N_4680,N_4745);
or UO_300 (O_300,N_4619,N_4297);
nand UO_301 (O_301,N_4278,N_4748);
or UO_302 (O_302,N_4144,N_4327);
nand UO_303 (O_303,N_4178,N_4978);
nor UO_304 (O_304,N_4918,N_4418);
nand UO_305 (O_305,N_4309,N_4413);
nor UO_306 (O_306,N_4305,N_4246);
and UO_307 (O_307,N_4779,N_4522);
nand UO_308 (O_308,N_4773,N_4425);
and UO_309 (O_309,N_4595,N_4128);
nand UO_310 (O_310,N_4134,N_4431);
or UO_311 (O_311,N_4800,N_4642);
nand UO_312 (O_312,N_4765,N_4556);
nor UO_313 (O_313,N_4108,N_4257);
nand UO_314 (O_314,N_4716,N_4635);
or UO_315 (O_315,N_4523,N_4329);
and UO_316 (O_316,N_4890,N_4317);
and UO_317 (O_317,N_4589,N_4858);
nand UO_318 (O_318,N_4099,N_4107);
or UO_319 (O_319,N_4617,N_4643);
nor UO_320 (O_320,N_4660,N_4251);
nand UO_321 (O_321,N_4825,N_4208);
nor UO_322 (O_322,N_4410,N_4614);
or UO_323 (O_323,N_4856,N_4691);
nor UO_324 (O_324,N_4797,N_4894);
nor UO_325 (O_325,N_4130,N_4744);
and UO_326 (O_326,N_4110,N_4381);
nor UO_327 (O_327,N_4832,N_4767);
nand UO_328 (O_328,N_4403,N_4563);
or UO_329 (O_329,N_4623,N_4258);
nand UO_330 (O_330,N_4211,N_4609);
nand UO_331 (O_331,N_4402,N_4960);
nor UO_332 (O_332,N_4072,N_4105);
nand UO_333 (O_333,N_4907,N_4318);
and UO_334 (O_334,N_4384,N_4561);
nor UO_335 (O_335,N_4807,N_4746);
nor UO_336 (O_336,N_4750,N_4179);
or UO_337 (O_337,N_4131,N_4373);
and UO_338 (O_338,N_4498,N_4177);
nand UO_339 (O_339,N_4357,N_4415);
nand UO_340 (O_340,N_4254,N_4798);
and UO_341 (O_341,N_4002,N_4061);
nor UO_342 (O_342,N_4252,N_4972);
nand UO_343 (O_343,N_4457,N_4977);
or UO_344 (O_344,N_4325,N_4802);
and UO_345 (O_345,N_4214,N_4004);
or UO_346 (O_346,N_4098,N_4165);
nand UO_347 (O_347,N_4489,N_4437);
nand UO_348 (O_348,N_4339,N_4083);
and UO_349 (O_349,N_4929,N_4304);
or UO_350 (O_350,N_4627,N_4474);
nand UO_351 (O_351,N_4315,N_4245);
and UO_352 (O_352,N_4708,N_4940);
and UO_353 (O_353,N_4653,N_4187);
or UO_354 (O_354,N_4197,N_4849);
and UO_355 (O_355,N_4146,N_4970);
nor UO_356 (O_356,N_4389,N_4718);
and UO_357 (O_357,N_4565,N_4430);
nand UO_358 (O_358,N_4608,N_4036);
nand UO_359 (O_359,N_4862,N_4195);
or UO_360 (O_360,N_4533,N_4671);
and UO_361 (O_361,N_4409,N_4138);
nor UO_362 (O_362,N_4826,N_4580);
xor UO_363 (O_363,N_4468,N_4466);
nor UO_364 (O_364,N_4925,N_4859);
or UO_365 (O_365,N_4122,N_4496);
and UO_366 (O_366,N_4460,N_4294);
nor UO_367 (O_367,N_4814,N_4353);
and UO_368 (O_368,N_4023,N_4081);
and UO_369 (O_369,N_4471,N_4651);
nor UO_370 (O_370,N_4391,N_4228);
and UO_371 (O_371,N_4521,N_4316);
nand UO_372 (O_372,N_4776,N_4562);
nor UO_373 (O_373,N_4397,N_4377);
and UO_374 (O_374,N_4948,N_4616);
nand UO_375 (O_375,N_4064,N_4264);
or UO_376 (O_376,N_4495,N_4326);
nand UO_377 (O_377,N_4622,N_4652);
nor UO_378 (O_378,N_4734,N_4428);
nand UO_379 (O_379,N_4159,N_4035);
or UO_380 (O_380,N_4374,N_4591);
and UO_381 (O_381,N_4364,N_4637);
and UO_382 (O_382,N_4679,N_4564);
nand UO_383 (O_383,N_4743,N_4348);
nor UO_384 (O_384,N_4207,N_4657);
nor UO_385 (O_385,N_4395,N_4053);
and UO_386 (O_386,N_4117,N_4022);
nor UO_387 (O_387,N_4730,N_4368);
and UO_388 (O_388,N_4740,N_4845);
and UO_389 (O_389,N_4140,N_4655);
nor UO_390 (O_390,N_4547,N_4668);
or UO_391 (O_391,N_4922,N_4936);
or UO_392 (O_392,N_4330,N_4799);
or UO_393 (O_393,N_4383,N_4531);
or UO_394 (O_394,N_4054,N_4587);
nand UO_395 (O_395,N_4071,N_4349);
nand UO_396 (O_396,N_4511,N_4733);
and UO_397 (O_397,N_4793,N_4020);
and UO_398 (O_398,N_4578,N_4124);
nor UO_399 (O_399,N_4566,N_4650);
and UO_400 (O_400,N_4685,N_4812);
and UO_401 (O_401,N_4775,N_4950);
and UO_402 (O_402,N_4946,N_4582);
and UO_403 (O_403,N_4588,N_4038);
nand UO_404 (O_404,N_4641,N_4888);
xnor UO_405 (O_405,N_4791,N_4661);
nand UO_406 (O_406,N_4571,N_4073);
nor UO_407 (O_407,N_4646,N_4239);
or UO_408 (O_408,N_4423,N_4301);
and UO_409 (O_409,N_4271,N_4669);
and UO_410 (O_410,N_4738,N_4512);
nand UO_411 (O_411,N_4399,N_4119);
and UO_412 (O_412,N_4209,N_4517);
nor UO_413 (O_413,N_4280,N_4287);
and UO_414 (O_414,N_4503,N_4382);
or UO_415 (O_415,N_4515,N_4293);
and UO_416 (O_416,N_4938,N_4783);
nand UO_417 (O_417,N_4576,N_4568);
and UO_418 (O_418,N_4884,N_4828);
nor UO_419 (O_419,N_4027,N_4074);
and UO_420 (O_420,N_4914,N_4243);
nor UO_421 (O_421,N_4947,N_4058);
nand UO_422 (O_422,N_4843,N_4952);
or UO_423 (O_423,N_4333,N_4095);
nand UO_424 (O_424,N_4411,N_4772);
nor UO_425 (O_425,N_4206,N_4106);
nor UO_426 (O_426,N_4913,N_4518);
or UO_427 (O_427,N_4500,N_4996);
nor UO_428 (O_428,N_4299,N_4751);
nor UO_429 (O_429,N_4876,N_4796);
nor UO_430 (O_430,N_4113,N_4672);
nand UO_431 (O_431,N_4935,N_4137);
or UO_432 (O_432,N_4895,N_4781);
or UO_433 (O_433,N_4604,N_4774);
nor UO_434 (O_434,N_4156,N_4068);
nand UO_435 (O_435,N_4801,N_4513);
nand UO_436 (O_436,N_4737,N_4342);
and UO_437 (O_437,N_4414,N_4692);
and UO_438 (O_438,N_4930,N_4993);
or UO_439 (O_439,N_4906,N_4817);
or UO_440 (O_440,N_4621,N_4714);
or UO_441 (O_441,N_4268,N_4323);
or UO_442 (O_442,N_4548,N_4059);
nand UO_443 (O_443,N_4715,N_4434);
or UO_444 (O_444,N_4821,N_4768);
nor UO_445 (O_445,N_4955,N_4846);
and UO_446 (O_446,N_4874,N_4502);
nor UO_447 (O_447,N_4283,N_4508);
nor UO_448 (O_448,N_4979,N_4575);
nand UO_449 (O_449,N_4346,N_4456);
nor UO_450 (O_450,N_4711,N_4831);
nor UO_451 (O_451,N_4013,N_4541);
or UO_452 (O_452,N_4808,N_4060);
nand UO_453 (O_453,N_4461,N_4829);
nor UO_454 (O_454,N_4248,N_4288);
and UO_455 (O_455,N_4269,N_4841);
nor UO_456 (O_456,N_4953,N_4398);
and UO_457 (O_457,N_4210,N_4729);
nor UO_458 (O_458,N_4155,N_4586);
and UO_459 (O_459,N_4086,N_4534);
nand UO_460 (O_460,N_4057,N_4012);
or UO_461 (O_461,N_4118,N_4902);
nor UO_462 (O_462,N_4574,N_4185);
and UO_463 (O_463,N_4967,N_4050);
or UO_464 (O_464,N_4285,N_4686);
or UO_465 (O_465,N_4731,N_4376);
or UO_466 (O_466,N_4235,N_4625);
nor UO_467 (O_467,N_4982,N_4539);
nor UO_468 (O_468,N_4432,N_4962);
nor UO_469 (O_469,N_4194,N_4687);
nand UO_470 (O_470,N_4865,N_4321);
or UO_471 (O_471,N_4009,N_4042);
or UO_472 (O_472,N_4610,N_4546);
nor UO_473 (O_473,N_4334,N_4903);
and UO_474 (O_474,N_4877,N_4372);
nor UO_475 (O_475,N_4665,N_4447);
nand UO_476 (O_476,N_4363,N_4857);
and UO_477 (O_477,N_4480,N_4200);
nand UO_478 (O_478,N_4028,N_4662);
or UO_479 (O_479,N_4704,N_4484);
xnor UO_480 (O_480,N_4524,N_4842);
or UO_481 (O_481,N_4031,N_4473);
and UO_482 (O_482,N_4719,N_4741);
or UO_483 (O_483,N_4990,N_4822);
nand UO_484 (O_484,N_4640,N_4314);
nor UO_485 (O_485,N_4818,N_4388);
nand UO_486 (O_486,N_4659,N_4889);
or UO_487 (O_487,N_4909,N_4303);
and UO_488 (O_488,N_4949,N_4592);
or UO_489 (O_489,N_4584,N_4873);
nor UO_490 (O_490,N_4599,N_4014);
or UO_491 (O_491,N_4045,N_4462);
nand UO_492 (O_492,N_4440,N_4286);
or UO_493 (O_493,N_4782,N_4670);
or UO_494 (O_494,N_4638,N_4535);
or UO_495 (O_495,N_4526,N_4279);
nor UO_496 (O_496,N_4343,N_4919);
nand UO_497 (O_497,N_4340,N_4689);
and UO_498 (O_498,N_4557,N_4011);
nor UO_499 (O_499,N_4396,N_4453);
nor UO_500 (O_500,N_4197,N_4950);
nand UO_501 (O_501,N_4548,N_4656);
and UO_502 (O_502,N_4002,N_4573);
and UO_503 (O_503,N_4096,N_4270);
nand UO_504 (O_504,N_4326,N_4600);
nor UO_505 (O_505,N_4812,N_4616);
nor UO_506 (O_506,N_4569,N_4166);
and UO_507 (O_507,N_4217,N_4618);
xnor UO_508 (O_508,N_4743,N_4356);
nand UO_509 (O_509,N_4142,N_4585);
or UO_510 (O_510,N_4326,N_4349);
nand UO_511 (O_511,N_4522,N_4850);
nor UO_512 (O_512,N_4752,N_4719);
or UO_513 (O_513,N_4563,N_4713);
nor UO_514 (O_514,N_4983,N_4808);
nor UO_515 (O_515,N_4467,N_4889);
nor UO_516 (O_516,N_4799,N_4090);
and UO_517 (O_517,N_4301,N_4357);
nand UO_518 (O_518,N_4250,N_4099);
nor UO_519 (O_519,N_4833,N_4616);
or UO_520 (O_520,N_4448,N_4895);
nand UO_521 (O_521,N_4182,N_4719);
or UO_522 (O_522,N_4179,N_4576);
nand UO_523 (O_523,N_4283,N_4168);
or UO_524 (O_524,N_4422,N_4065);
xor UO_525 (O_525,N_4991,N_4867);
nor UO_526 (O_526,N_4034,N_4826);
or UO_527 (O_527,N_4413,N_4111);
nand UO_528 (O_528,N_4062,N_4871);
or UO_529 (O_529,N_4076,N_4818);
nand UO_530 (O_530,N_4365,N_4196);
nor UO_531 (O_531,N_4510,N_4970);
nand UO_532 (O_532,N_4050,N_4951);
nand UO_533 (O_533,N_4857,N_4937);
nor UO_534 (O_534,N_4635,N_4210);
and UO_535 (O_535,N_4413,N_4923);
nor UO_536 (O_536,N_4638,N_4332);
or UO_537 (O_537,N_4164,N_4877);
and UO_538 (O_538,N_4729,N_4092);
or UO_539 (O_539,N_4018,N_4991);
nor UO_540 (O_540,N_4287,N_4895);
and UO_541 (O_541,N_4122,N_4263);
nor UO_542 (O_542,N_4060,N_4378);
and UO_543 (O_543,N_4374,N_4760);
nand UO_544 (O_544,N_4652,N_4628);
and UO_545 (O_545,N_4295,N_4769);
nand UO_546 (O_546,N_4590,N_4409);
and UO_547 (O_547,N_4741,N_4493);
nand UO_548 (O_548,N_4712,N_4983);
nor UO_549 (O_549,N_4026,N_4540);
and UO_550 (O_550,N_4770,N_4132);
nand UO_551 (O_551,N_4349,N_4619);
and UO_552 (O_552,N_4737,N_4909);
nor UO_553 (O_553,N_4583,N_4980);
nor UO_554 (O_554,N_4991,N_4691);
nor UO_555 (O_555,N_4744,N_4596);
or UO_556 (O_556,N_4151,N_4245);
or UO_557 (O_557,N_4001,N_4378);
and UO_558 (O_558,N_4382,N_4641);
and UO_559 (O_559,N_4193,N_4089);
or UO_560 (O_560,N_4908,N_4517);
nand UO_561 (O_561,N_4269,N_4848);
nor UO_562 (O_562,N_4330,N_4827);
or UO_563 (O_563,N_4243,N_4872);
or UO_564 (O_564,N_4172,N_4250);
and UO_565 (O_565,N_4596,N_4639);
nand UO_566 (O_566,N_4536,N_4686);
nand UO_567 (O_567,N_4432,N_4544);
nor UO_568 (O_568,N_4928,N_4234);
and UO_569 (O_569,N_4287,N_4830);
or UO_570 (O_570,N_4095,N_4998);
nand UO_571 (O_571,N_4361,N_4379);
or UO_572 (O_572,N_4812,N_4769);
nor UO_573 (O_573,N_4676,N_4301);
and UO_574 (O_574,N_4428,N_4368);
and UO_575 (O_575,N_4041,N_4313);
or UO_576 (O_576,N_4156,N_4874);
nand UO_577 (O_577,N_4238,N_4176);
and UO_578 (O_578,N_4985,N_4844);
nor UO_579 (O_579,N_4888,N_4378);
or UO_580 (O_580,N_4866,N_4343);
nor UO_581 (O_581,N_4708,N_4748);
or UO_582 (O_582,N_4356,N_4723);
and UO_583 (O_583,N_4429,N_4410);
xor UO_584 (O_584,N_4160,N_4194);
nand UO_585 (O_585,N_4723,N_4495);
xnor UO_586 (O_586,N_4854,N_4544);
or UO_587 (O_587,N_4877,N_4481);
or UO_588 (O_588,N_4497,N_4975);
nand UO_589 (O_589,N_4615,N_4851);
nand UO_590 (O_590,N_4752,N_4106);
nand UO_591 (O_591,N_4460,N_4803);
nand UO_592 (O_592,N_4797,N_4839);
and UO_593 (O_593,N_4141,N_4011);
nor UO_594 (O_594,N_4979,N_4492);
nand UO_595 (O_595,N_4979,N_4268);
nand UO_596 (O_596,N_4966,N_4976);
nor UO_597 (O_597,N_4790,N_4715);
and UO_598 (O_598,N_4093,N_4694);
nor UO_599 (O_599,N_4475,N_4557);
or UO_600 (O_600,N_4603,N_4510);
nor UO_601 (O_601,N_4666,N_4712);
or UO_602 (O_602,N_4560,N_4775);
nor UO_603 (O_603,N_4460,N_4206);
nand UO_604 (O_604,N_4194,N_4366);
nor UO_605 (O_605,N_4294,N_4451);
and UO_606 (O_606,N_4872,N_4098);
nor UO_607 (O_607,N_4227,N_4097);
or UO_608 (O_608,N_4078,N_4769);
and UO_609 (O_609,N_4432,N_4522);
or UO_610 (O_610,N_4645,N_4159);
nor UO_611 (O_611,N_4969,N_4153);
or UO_612 (O_612,N_4238,N_4192);
or UO_613 (O_613,N_4685,N_4320);
nor UO_614 (O_614,N_4501,N_4838);
nand UO_615 (O_615,N_4373,N_4842);
xnor UO_616 (O_616,N_4046,N_4167);
or UO_617 (O_617,N_4630,N_4588);
or UO_618 (O_618,N_4476,N_4535);
nor UO_619 (O_619,N_4811,N_4493);
and UO_620 (O_620,N_4521,N_4115);
or UO_621 (O_621,N_4162,N_4629);
nand UO_622 (O_622,N_4276,N_4378);
nand UO_623 (O_623,N_4259,N_4812);
nand UO_624 (O_624,N_4015,N_4771);
or UO_625 (O_625,N_4425,N_4352);
nor UO_626 (O_626,N_4711,N_4016);
nand UO_627 (O_627,N_4278,N_4849);
nor UO_628 (O_628,N_4352,N_4067);
or UO_629 (O_629,N_4392,N_4015);
and UO_630 (O_630,N_4743,N_4579);
nor UO_631 (O_631,N_4606,N_4395);
or UO_632 (O_632,N_4945,N_4469);
nand UO_633 (O_633,N_4887,N_4075);
and UO_634 (O_634,N_4371,N_4447);
nor UO_635 (O_635,N_4788,N_4650);
nor UO_636 (O_636,N_4354,N_4640);
or UO_637 (O_637,N_4808,N_4110);
nor UO_638 (O_638,N_4022,N_4819);
nand UO_639 (O_639,N_4187,N_4424);
nor UO_640 (O_640,N_4555,N_4370);
nand UO_641 (O_641,N_4818,N_4886);
or UO_642 (O_642,N_4251,N_4758);
nor UO_643 (O_643,N_4834,N_4766);
and UO_644 (O_644,N_4879,N_4138);
or UO_645 (O_645,N_4378,N_4776);
and UO_646 (O_646,N_4455,N_4368);
nor UO_647 (O_647,N_4981,N_4608);
nand UO_648 (O_648,N_4899,N_4700);
or UO_649 (O_649,N_4242,N_4611);
or UO_650 (O_650,N_4068,N_4969);
or UO_651 (O_651,N_4754,N_4203);
nor UO_652 (O_652,N_4890,N_4789);
nor UO_653 (O_653,N_4346,N_4470);
or UO_654 (O_654,N_4990,N_4246);
and UO_655 (O_655,N_4526,N_4656);
or UO_656 (O_656,N_4417,N_4634);
and UO_657 (O_657,N_4812,N_4153);
nand UO_658 (O_658,N_4135,N_4251);
nor UO_659 (O_659,N_4426,N_4676);
or UO_660 (O_660,N_4017,N_4198);
nand UO_661 (O_661,N_4420,N_4706);
or UO_662 (O_662,N_4812,N_4408);
nor UO_663 (O_663,N_4729,N_4268);
and UO_664 (O_664,N_4091,N_4971);
or UO_665 (O_665,N_4021,N_4219);
nor UO_666 (O_666,N_4459,N_4658);
nor UO_667 (O_667,N_4224,N_4903);
or UO_668 (O_668,N_4976,N_4705);
or UO_669 (O_669,N_4755,N_4989);
and UO_670 (O_670,N_4374,N_4502);
or UO_671 (O_671,N_4556,N_4376);
or UO_672 (O_672,N_4177,N_4205);
nor UO_673 (O_673,N_4679,N_4105);
xnor UO_674 (O_674,N_4531,N_4426);
or UO_675 (O_675,N_4142,N_4965);
nor UO_676 (O_676,N_4966,N_4059);
or UO_677 (O_677,N_4990,N_4719);
nor UO_678 (O_678,N_4114,N_4294);
nor UO_679 (O_679,N_4187,N_4559);
and UO_680 (O_680,N_4514,N_4531);
or UO_681 (O_681,N_4689,N_4850);
xnor UO_682 (O_682,N_4675,N_4008);
or UO_683 (O_683,N_4710,N_4241);
and UO_684 (O_684,N_4124,N_4017);
or UO_685 (O_685,N_4193,N_4698);
and UO_686 (O_686,N_4945,N_4063);
nand UO_687 (O_687,N_4771,N_4858);
and UO_688 (O_688,N_4228,N_4262);
and UO_689 (O_689,N_4376,N_4946);
nor UO_690 (O_690,N_4435,N_4077);
and UO_691 (O_691,N_4249,N_4540);
or UO_692 (O_692,N_4237,N_4918);
nor UO_693 (O_693,N_4368,N_4905);
nand UO_694 (O_694,N_4268,N_4087);
and UO_695 (O_695,N_4792,N_4686);
or UO_696 (O_696,N_4116,N_4859);
nand UO_697 (O_697,N_4388,N_4008);
or UO_698 (O_698,N_4453,N_4405);
or UO_699 (O_699,N_4380,N_4848);
nor UO_700 (O_700,N_4113,N_4525);
nand UO_701 (O_701,N_4733,N_4086);
or UO_702 (O_702,N_4074,N_4461);
or UO_703 (O_703,N_4408,N_4693);
and UO_704 (O_704,N_4845,N_4134);
and UO_705 (O_705,N_4395,N_4244);
nand UO_706 (O_706,N_4703,N_4017);
nor UO_707 (O_707,N_4014,N_4956);
or UO_708 (O_708,N_4732,N_4457);
and UO_709 (O_709,N_4355,N_4356);
nand UO_710 (O_710,N_4641,N_4403);
nor UO_711 (O_711,N_4349,N_4556);
nand UO_712 (O_712,N_4189,N_4016);
nand UO_713 (O_713,N_4031,N_4406);
nand UO_714 (O_714,N_4657,N_4708);
xor UO_715 (O_715,N_4592,N_4895);
and UO_716 (O_716,N_4816,N_4099);
or UO_717 (O_717,N_4716,N_4649);
nor UO_718 (O_718,N_4980,N_4015);
and UO_719 (O_719,N_4598,N_4405);
nand UO_720 (O_720,N_4413,N_4876);
and UO_721 (O_721,N_4969,N_4559);
or UO_722 (O_722,N_4496,N_4392);
nor UO_723 (O_723,N_4310,N_4231);
or UO_724 (O_724,N_4047,N_4353);
or UO_725 (O_725,N_4342,N_4142);
or UO_726 (O_726,N_4033,N_4988);
and UO_727 (O_727,N_4062,N_4681);
or UO_728 (O_728,N_4785,N_4756);
nand UO_729 (O_729,N_4862,N_4545);
nor UO_730 (O_730,N_4035,N_4576);
and UO_731 (O_731,N_4172,N_4672);
nand UO_732 (O_732,N_4516,N_4080);
nor UO_733 (O_733,N_4044,N_4815);
and UO_734 (O_734,N_4008,N_4265);
or UO_735 (O_735,N_4346,N_4202);
or UO_736 (O_736,N_4232,N_4508);
and UO_737 (O_737,N_4368,N_4301);
nor UO_738 (O_738,N_4924,N_4242);
and UO_739 (O_739,N_4225,N_4465);
nand UO_740 (O_740,N_4406,N_4242);
nor UO_741 (O_741,N_4547,N_4787);
or UO_742 (O_742,N_4593,N_4087);
nand UO_743 (O_743,N_4739,N_4983);
nand UO_744 (O_744,N_4823,N_4852);
and UO_745 (O_745,N_4434,N_4890);
or UO_746 (O_746,N_4797,N_4046);
and UO_747 (O_747,N_4594,N_4609);
or UO_748 (O_748,N_4605,N_4360);
nand UO_749 (O_749,N_4685,N_4456);
or UO_750 (O_750,N_4489,N_4338);
or UO_751 (O_751,N_4567,N_4002);
or UO_752 (O_752,N_4051,N_4333);
nor UO_753 (O_753,N_4176,N_4977);
or UO_754 (O_754,N_4506,N_4111);
or UO_755 (O_755,N_4457,N_4059);
nand UO_756 (O_756,N_4691,N_4811);
and UO_757 (O_757,N_4323,N_4333);
and UO_758 (O_758,N_4569,N_4768);
nor UO_759 (O_759,N_4113,N_4088);
or UO_760 (O_760,N_4085,N_4548);
nor UO_761 (O_761,N_4048,N_4930);
or UO_762 (O_762,N_4754,N_4871);
or UO_763 (O_763,N_4909,N_4289);
nor UO_764 (O_764,N_4701,N_4852);
nor UO_765 (O_765,N_4118,N_4165);
nand UO_766 (O_766,N_4330,N_4471);
or UO_767 (O_767,N_4283,N_4186);
nand UO_768 (O_768,N_4772,N_4019);
or UO_769 (O_769,N_4284,N_4801);
nor UO_770 (O_770,N_4009,N_4487);
nand UO_771 (O_771,N_4403,N_4670);
nor UO_772 (O_772,N_4299,N_4356);
and UO_773 (O_773,N_4592,N_4656);
nand UO_774 (O_774,N_4215,N_4108);
or UO_775 (O_775,N_4754,N_4652);
nor UO_776 (O_776,N_4608,N_4547);
and UO_777 (O_777,N_4743,N_4036);
or UO_778 (O_778,N_4223,N_4171);
nor UO_779 (O_779,N_4598,N_4840);
or UO_780 (O_780,N_4580,N_4213);
or UO_781 (O_781,N_4113,N_4641);
nand UO_782 (O_782,N_4227,N_4674);
nand UO_783 (O_783,N_4975,N_4946);
and UO_784 (O_784,N_4197,N_4459);
or UO_785 (O_785,N_4786,N_4900);
nor UO_786 (O_786,N_4001,N_4214);
nor UO_787 (O_787,N_4447,N_4033);
or UO_788 (O_788,N_4395,N_4345);
or UO_789 (O_789,N_4355,N_4517);
nand UO_790 (O_790,N_4258,N_4137);
and UO_791 (O_791,N_4059,N_4576);
nor UO_792 (O_792,N_4073,N_4328);
and UO_793 (O_793,N_4114,N_4266);
and UO_794 (O_794,N_4012,N_4120);
nand UO_795 (O_795,N_4491,N_4513);
nand UO_796 (O_796,N_4538,N_4775);
nor UO_797 (O_797,N_4955,N_4384);
nor UO_798 (O_798,N_4352,N_4659);
nor UO_799 (O_799,N_4631,N_4135);
nand UO_800 (O_800,N_4566,N_4882);
and UO_801 (O_801,N_4264,N_4554);
or UO_802 (O_802,N_4901,N_4203);
nand UO_803 (O_803,N_4990,N_4041);
or UO_804 (O_804,N_4167,N_4961);
nor UO_805 (O_805,N_4850,N_4495);
or UO_806 (O_806,N_4624,N_4861);
nor UO_807 (O_807,N_4326,N_4873);
nor UO_808 (O_808,N_4819,N_4838);
nand UO_809 (O_809,N_4019,N_4745);
or UO_810 (O_810,N_4657,N_4614);
nand UO_811 (O_811,N_4629,N_4568);
or UO_812 (O_812,N_4084,N_4965);
and UO_813 (O_813,N_4880,N_4961);
and UO_814 (O_814,N_4850,N_4705);
or UO_815 (O_815,N_4262,N_4276);
nand UO_816 (O_816,N_4064,N_4095);
or UO_817 (O_817,N_4941,N_4759);
and UO_818 (O_818,N_4466,N_4676);
nor UO_819 (O_819,N_4161,N_4018);
nand UO_820 (O_820,N_4909,N_4845);
nor UO_821 (O_821,N_4659,N_4423);
or UO_822 (O_822,N_4886,N_4872);
nor UO_823 (O_823,N_4933,N_4547);
nand UO_824 (O_824,N_4856,N_4178);
nand UO_825 (O_825,N_4685,N_4484);
nor UO_826 (O_826,N_4315,N_4446);
and UO_827 (O_827,N_4902,N_4607);
nor UO_828 (O_828,N_4990,N_4165);
nor UO_829 (O_829,N_4521,N_4574);
nand UO_830 (O_830,N_4270,N_4243);
xor UO_831 (O_831,N_4272,N_4408);
or UO_832 (O_832,N_4580,N_4546);
or UO_833 (O_833,N_4023,N_4911);
or UO_834 (O_834,N_4770,N_4767);
or UO_835 (O_835,N_4375,N_4179);
nand UO_836 (O_836,N_4188,N_4828);
nand UO_837 (O_837,N_4694,N_4568);
nor UO_838 (O_838,N_4397,N_4272);
nor UO_839 (O_839,N_4933,N_4958);
or UO_840 (O_840,N_4997,N_4530);
or UO_841 (O_841,N_4001,N_4482);
nand UO_842 (O_842,N_4362,N_4784);
and UO_843 (O_843,N_4273,N_4850);
or UO_844 (O_844,N_4061,N_4973);
and UO_845 (O_845,N_4585,N_4106);
or UO_846 (O_846,N_4371,N_4860);
nor UO_847 (O_847,N_4952,N_4188);
nor UO_848 (O_848,N_4952,N_4040);
and UO_849 (O_849,N_4199,N_4707);
nor UO_850 (O_850,N_4633,N_4120);
nand UO_851 (O_851,N_4481,N_4519);
and UO_852 (O_852,N_4618,N_4836);
nor UO_853 (O_853,N_4436,N_4361);
xor UO_854 (O_854,N_4182,N_4421);
nor UO_855 (O_855,N_4031,N_4614);
or UO_856 (O_856,N_4507,N_4434);
or UO_857 (O_857,N_4139,N_4993);
or UO_858 (O_858,N_4479,N_4683);
or UO_859 (O_859,N_4835,N_4257);
or UO_860 (O_860,N_4147,N_4617);
or UO_861 (O_861,N_4289,N_4959);
nand UO_862 (O_862,N_4454,N_4627);
and UO_863 (O_863,N_4269,N_4198);
or UO_864 (O_864,N_4012,N_4724);
or UO_865 (O_865,N_4649,N_4841);
xor UO_866 (O_866,N_4021,N_4431);
and UO_867 (O_867,N_4014,N_4251);
and UO_868 (O_868,N_4984,N_4488);
and UO_869 (O_869,N_4938,N_4879);
and UO_870 (O_870,N_4340,N_4430);
or UO_871 (O_871,N_4836,N_4191);
and UO_872 (O_872,N_4910,N_4465);
nor UO_873 (O_873,N_4304,N_4001);
nor UO_874 (O_874,N_4649,N_4515);
or UO_875 (O_875,N_4093,N_4431);
nand UO_876 (O_876,N_4194,N_4900);
and UO_877 (O_877,N_4337,N_4252);
or UO_878 (O_878,N_4682,N_4694);
nor UO_879 (O_879,N_4418,N_4137);
and UO_880 (O_880,N_4042,N_4624);
and UO_881 (O_881,N_4746,N_4608);
and UO_882 (O_882,N_4037,N_4993);
nor UO_883 (O_883,N_4863,N_4121);
or UO_884 (O_884,N_4140,N_4696);
or UO_885 (O_885,N_4601,N_4551);
or UO_886 (O_886,N_4224,N_4743);
xnor UO_887 (O_887,N_4540,N_4275);
nand UO_888 (O_888,N_4178,N_4407);
or UO_889 (O_889,N_4973,N_4919);
or UO_890 (O_890,N_4006,N_4201);
nand UO_891 (O_891,N_4344,N_4299);
and UO_892 (O_892,N_4677,N_4745);
nand UO_893 (O_893,N_4121,N_4164);
nand UO_894 (O_894,N_4944,N_4279);
nor UO_895 (O_895,N_4941,N_4766);
nand UO_896 (O_896,N_4331,N_4425);
and UO_897 (O_897,N_4889,N_4898);
nand UO_898 (O_898,N_4737,N_4271);
nor UO_899 (O_899,N_4965,N_4418);
nor UO_900 (O_900,N_4173,N_4417);
nor UO_901 (O_901,N_4644,N_4364);
nand UO_902 (O_902,N_4699,N_4079);
nor UO_903 (O_903,N_4738,N_4927);
nand UO_904 (O_904,N_4303,N_4049);
nand UO_905 (O_905,N_4069,N_4723);
nand UO_906 (O_906,N_4043,N_4941);
xnor UO_907 (O_907,N_4400,N_4480);
or UO_908 (O_908,N_4971,N_4514);
nor UO_909 (O_909,N_4796,N_4360);
nand UO_910 (O_910,N_4386,N_4899);
nor UO_911 (O_911,N_4814,N_4467);
or UO_912 (O_912,N_4298,N_4144);
nand UO_913 (O_913,N_4320,N_4777);
and UO_914 (O_914,N_4630,N_4621);
nand UO_915 (O_915,N_4960,N_4728);
nand UO_916 (O_916,N_4907,N_4929);
nand UO_917 (O_917,N_4068,N_4225);
nand UO_918 (O_918,N_4966,N_4427);
nand UO_919 (O_919,N_4340,N_4549);
or UO_920 (O_920,N_4748,N_4966);
nor UO_921 (O_921,N_4638,N_4959);
and UO_922 (O_922,N_4650,N_4667);
and UO_923 (O_923,N_4416,N_4088);
and UO_924 (O_924,N_4979,N_4819);
nand UO_925 (O_925,N_4039,N_4685);
and UO_926 (O_926,N_4207,N_4978);
and UO_927 (O_927,N_4249,N_4159);
or UO_928 (O_928,N_4403,N_4430);
or UO_929 (O_929,N_4658,N_4582);
and UO_930 (O_930,N_4853,N_4406);
nor UO_931 (O_931,N_4203,N_4834);
nor UO_932 (O_932,N_4433,N_4348);
nand UO_933 (O_933,N_4597,N_4396);
or UO_934 (O_934,N_4585,N_4773);
nand UO_935 (O_935,N_4613,N_4698);
and UO_936 (O_936,N_4176,N_4907);
or UO_937 (O_937,N_4387,N_4828);
xnor UO_938 (O_938,N_4394,N_4295);
nand UO_939 (O_939,N_4379,N_4258);
and UO_940 (O_940,N_4196,N_4158);
or UO_941 (O_941,N_4112,N_4311);
and UO_942 (O_942,N_4798,N_4106);
nand UO_943 (O_943,N_4244,N_4797);
and UO_944 (O_944,N_4077,N_4936);
and UO_945 (O_945,N_4534,N_4564);
or UO_946 (O_946,N_4613,N_4357);
and UO_947 (O_947,N_4300,N_4758);
nor UO_948 (O_948,N_4837,N_4408);
nor UO_949 (O_949,N_4208,N_4206);
nand UO_950 (O_950,N_4729,N_4371);
nand UO_951 (O_951,N_4995,N_4608);
nand UO_952 (O_952,N_4020,N_4872);
nor UO_953 (O_953,N_4972,N_4642);
and UO_954 (O_954,N_4153,N_4025);
nand UO_955 (O_955,N_4950,N_4603);
nor UO_956 (O_956,N_4944,N_4846);
and UO_957 (O_957,N_4025,N_4624);
nand UO_958 (O_958,N_4699,N_4212);
nor UO_959 (O_959,N_4815,N_4221);
nor UO_960 (O_960,N_4386,N_4591);
and UO_961 (O_961,N_4557,N_4574);
nor UO_962 (O_962,N_4781,N_4613);
nor UO_963 (O_963,N_4467,N_4954);
or UO_964 (O_964,N_4789,N_4623);
or UO_965 (O_965,N_4432,N_4924);
and UO_966 (O_966,N_4353,N_4794);
nand UO_967 (O_967,N_4712,N_4067);
nor UO_968 (O_968,N_4841,N_4615);
or UO_969 (O_969,N_4015,N_4769);
and UO_970 (O_970,N_4404,N_4000);
and UO_971 (O_971,N_4406,N_4260);
and UO_972 (O_972,N_4404,N_4741);
nor UO_973 (O_973,N_4979,N_4328);
or UO_974 (O_974,N_4663,N_4390);
nand UO_975 (O_975,N_4802,N_4439);
nor UO_976 (O_976,N_4802,N_4097);
or UO_977 (O_977,N_4223,N_4222);
nand UO_978 (O_978,N_4045,N_4071);
and UO_979 (O_979,N_4670,N_4543);
and UO_980 (O_980,N_4932,N_4978);
nor UO_981 (O_981,N_4185,N_4205);
or UO_982 (O_982,N_4460,N_4379);
or UO_983 (O_983,N_4426,N_4517);
and UO_984 (O_984,N_4026,N_4898);
and UO_985 (O_985,N_4417,N_4653);
nand UO_986 (O_986,N_4048,N_4450);
or UO_987 (O_987,N_4508,N_4850);
nor UO_988 (O_988,N_4909,N_4731);
or UO_989 (O_989,N_4956,N_4946);
nor UO_990 (O_990,N_4303,N_4985);
and UO_991 (O_991,N_4388,N_4718);
nor UO_992 (O_992,N_4466,N_4819);
and UO_993 (O_993,N_4817,N_4394);
nor UO_994 (O_994,N_4556,N_4236);
nand UO_995 (O_995,N_4611,N_4660);
and UO_996 (O_996,N_4904,N_4203);
and UO_997 (O_997,N_4603,N_4694);
nand UO_998 (O_998,N_4515,N_4303);
and UO_999 (O_999,N_4465,N_4574);
endmodule