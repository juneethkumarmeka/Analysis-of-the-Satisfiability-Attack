module basic_5000_50000_5000_10_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nand U0 (N_0,In_635,In_719);
xor U1 (N_1,In_683,In_887);
xnor U2 (N_2,In_2135,In_2220);
nand U3 (N_3,In_2642,In_3767);
or U4 (N_4,In_99,In_4692);
nand U5 (N_5,In_2384,In_4785);
nor U6 (N_6,In_707,In_3322);
xor U7 (N_7,In_3392,In_374);
nor U8 (N_8,In_850,In_975);
nor U9 (N_9,In_3250,In_250);
or U10 (N_10,In_3997,In_1437);
nand U11 (N_11,In_3843,In_1261);
nor U12 (N_12,In_4039,In_3396);
xnor U13 (N_13,In_417,In_4061);
and U14 (N_14,In_2914,In_2728);
nand U15 (N_15,In_1045,In_821);
and U16 (N_16,In_2857,In_3492);
xor U17 (N_17,In_3548,In_1600);
xnor U18 (N_18,In_4859,In_1737);
or U19 (N_19,In_3083,In_4670);
and U20 (N_20,In_4870,In_3160);
and U21 (N_21,In_4251,In_2791);
nand U22 (N_22,In_2569,In_4338);
nor U23 (N_23,In_2363,In_3431);
and U24 (N_24,In_336,In_997);
xnor U25 (N_25,In_1881,In_630);
and U26 (N_26,In_4815,In_1703);
and U27 (N_27,In_1263,In_1072);
nand U28 (N_28,In_4408,In_4745);
nor U29 (N_29,In_2688,In_1351);
nor U30 (N_30,In_1053,In_599);
and U31 (N_31,In_4685,In_1021);
and U32 (N_32,In_908,In_1741);
or U33 (N_33,In_991,In_1557);
and U34 (N_34,In_1893,In_3463);
and U35 (N_35,In_202,In_3712);
and U36 (N_36,In_2831,In_3954);
nand U37 (N_37,In_1055,In_1944);
and U38 (N_38,In_2338,In_382);
or U39 (N_39,In_4106,In_3015);
xnor U40 (N_40,In_3986,In_807);
nor U41 (N_41,In_4849,In_4111);
nor U42 (N_42,In_1791,In_824);
nor U43 (N_43,In_1672,In_1398);
nor U44 (N_44,In_1237,In_4081);
or U45 (N_45,In_3452,In_1473);
nand U46 (N_46,In_3402,In_3389);
and U47 (N_47,In_4919,In_461);
nor U48 (N_48,In_1930,In_189);
nand U49 (N_49,In_1457,In_1613);
nor U50 (N_50,In_3519,In_4454);
xnor U51 (N_51,In_2621,In_3706);
or U52 (N_52,In_3564,In_1408);
nand U53 (N_53,In_75,In_4392);
and U54 (N_54,In_403,In_3221);
xnor U55 (N_55,In_1866,In_4292);
nand U56 (N_56,In_4598,In_199);
xnor U57 (N_57,In_4606,In_4154);
nor U58 (N_58,In_3258,In_2798);
nor U59 (N_59,In_642,In_2833);
nand U60 (N_60,In_2182,In_2361);
nor U61 (N_61,In_866,In_2223);
and U62 (N_62,In_4256,In_1979);
nor U63 (N_63,In_1358,In_1477);
xor U64 (N_64,In_3691,In_4427);
xnor U65 (N_65,In_3632,In_1594);
xor U66 (N_66,In_2360,In_2002);
or U67 (N_67,In_2753,In_3302);
xor U68 (N_68,In_1680,In_1647);
nand U69 (N_69,In_3298,In_4534);
nand U70 (N_70,In_3465,In_43);
or U71 (N_71,In_4040,In_3569);
nor U72 (N_72,In_3567,In_3067);
or U73 (N_73,In_2518,In_4314);
and U74 (N_74,In_302,In_2139);
nor U75 (N_75,In_3466,In_1331);
nor U76 (N_76,In_4986,In_28);
and U77 (N_77,In_3011,In_1921);
nor U78 (N_78,In_1714,In_3399);
or U79 (N_79,In_4973,In_1056);
nand U80 (N_80,In_1880,In_2354);
xor U81 (N_81,In_1831,In_1100);
xnor U82 (N_82,In_2564,In_973);
and U83 (N_83,In_4827,In_1926);
and U84 (N_84,In_4577,In_1622);
nand U85 (N_85,In_393,In_2699);
and U86 (N_86,In_4136,In_1621);
nand U87 (N_87,In_3869,In_3175);
or U88 (N_88,In_2409,In_1505);
nand U89 (N_89,In_1538,In_1214);
xnor U90 (N_90,In_24,In_3588);
or U91 (N_91,In_3897,In_938);
nor U92 (N_92,In_2199,In_1368);
or U93 (N_93,In_4344,In_4053);
and U94 (N_94,In_1834,In_3561);
nor U95 (N_95,In_2365,In_774);
nand U96 (N_96,In_1489,In_3848);
nor U97 (N_97,In_1363,In_3647);
nor U98 (N_98,In_4376,In_4492);
or U99 (N_99,In_3711,In_4934);
or U100 (N_100,In_373,In_3599);
nor U101 (N_101,In_387,In_112);
nor U102 (N_102,In_34,In_465);
nand U103 (N_103,In_1932,In_2230);
nor U104 (N_104,In_547,In_3806);
xnor U105 (N_105,In_1707,In_2531);
nand U106 (N_106,In_2161,In_1438);
nand U107 (N_107,In_4303,In_4916);
and U108 (N_108,In_4962,In_2284);
xnor U109 (N_109,In_962,In_4991);
and U110 (N_110,In_2962,In_4412);
nor U111 (N_111,In_2647,In_3433);
and U112 (N_112,In_262,In_355);
and U113 (N_113,In_756,In_2969);
or U114 (N_114,In_3746,In_1789);
and U115 (N_115,In_1440,In_2555);
and U116 (N_116,In_2836,In_2341);
xnor U117 (N_117,In_2378,In_2867);
nand U118 (N_118,In_3984,In_226);
or U119 (N_119,In_1292,In_1362);
nor U120 (N_120,In_659,In_605);
nor U121 (N_121,In_3728,In_3337);
and U122 (N_122,In_15,In_1427);
and U123 (N_123,In_3601,In_1794);
xnor U124 (N_124,In_3040,In_3085);
or U125 (N_125,In_67,In_1446);
or U126 (N_126,In_3248,In_1959);
nor U127 (N_127,In_2662,In_231);
nand U128 (N_128,In_4539,In_3764);
nand U129 (N_129,In_1805,In_1819);
nand U130 (N_130,In_4620,In_4956);
and U131 (N_131,In_4621,In_2150);
nand U132 (N_132,In_2896,In_1273);
nor U133 (N_133,In_3730,In_1463);
nor U134 (N_134,In_4034,In_2918);
xor U135 (N_135,In_4947,In_2895);
xor U136 (N_136,In_1009,In_2392);
nand U137 (N_137,In_4803,In_4082);
xor U138 (N_138,In_639,In_2674);
nor U139 (N_139,In_2576,In_4832);
nand U140 (N_140,In_4470,In_3971);
nand U141 (N_141,In_3211,In_3798);
nand U142 (N_142,In_4382,In_3208);
and U143 (N_143,In_1821,In_1164);
nor U144 (N_144,In_2934,In_1658);
nor U145 (N_145,In_4861,In_2399);
nor U146 (N_146,In_1887,In_3851);
nor U147 (N_147,In_45,In_197);
xnor U148 (N_148,In_1493,In_1920);
and U149 (N_149,In_353,In_1911);
xnor U150 (N_150,In_3371,In_532);
xnor U151 (N_151,In_4591,In_2508);
and U152 (N_152,In_2710,In_1601);
xor U153 (N_153,In_107,In_4613);
nor U154 (N_154,In_2056,In_346);
and U155 (N_155,In_677,In_668);
xnor U156 (N_156,In_647,In_3308);
nor U157 (N_157,In_3150,In_4269);
xor U158 (N_158,In_1704,In_2007);
or U159 (N_159,In_3339,In_606);
nand U160 (N_160,In_4547,In_3753);
nor U161 (N_161,In_4864,In_185);
xnor U162 (N_162,In_1767,In_1595);
nand U163 (N_163,In_1572,In_4065);
nor U164 (N_164,In_2034,In_44);
or U165 (N_165,In_2677,In_2610);
nand U166 (N_166,In_2093,In_3629);
and U167 (N_167,In_1384,In_2407);
xor U168 (N_168,In_170,In_3607);
or U169 (N_169,In_3428,In_289);
and U170 (N_170,In_701,In_4019);
nand U171 (N_171,In_1695,In_1059);
nor U172 (N_172,In_2130,In_3158);
xor U173 (N_173,In_1002,In_4459);
nand U174 (N_174,In_1439,In_20);
xor U175 (N_175,In_4033,In_4263);
or U176 (N_176,In_4545,In_3750);
or U177 (N_177,In_3779,In_1983);
or U178 (N_178,In_4489,In_1651);
and U179 (N_179,In_1078,In_2281);
xor U180 (N_180,In_2917,In_2371);
or U181 (N_181,In_3482,In_2208);
xnor U182 (N_182,In_1186,In_58);
and U183 (N_183,In_3889,In_1373);
nor U184 (N_184,In_4367,In_1949);
nand U185 (N_185,In_3039,In_921);
or U186 (N_186,In_3542,In_445);
nand U187 (N_187,In_438,In_1156);
nand U188 (N_188,In_504,In_4103);
and U189 (N_189,In_492,In_4520);
xor U190 (N_190,In_1765,In_1141);
nor U191 (N_191,In_4596,In_2043);
nor U192 (N_192,In_2079,In_2071);
xnor U193 (N_193,In_180,In_4942);
xnor U194 (N_194,In_1654,In_514);
nand U195 (N_195,In_1648,In_1635);
nand U196 (N_196,In_4233,In_2140);
and U197 (N_197,In_4067,In_3789);
and U198 (N_198,In_545,In_4578);
and U199 (N_199,In_4333,In_260);
and U200 (N_200,In_1213,In_69);
nand U201 (N_201,In_3066,In_95);
nand U202 (N_202,In_4299,In_2709);
nor U203 (N_203,In_832,In_3416);
xnor U204 (N_204,In_2579,In_4373);
or U205 (N_205,In_1945,In_3376);
xnor U206 (N_206,In_1646,In_4298);
nor U207 (N_207,In_793,In_2800);
xnor U208 (N_208,In_1504,In_415);
xnor U209 (N_209,In_4654,In_503);
nor U210 (N_210,In_4610,In_2608);
xnor U211 (N_211,In_3604,In_1468);
nor U212 (N_212,In_2990,In_1191);
or U213 (N_213,In_2910,In_3552);
and U214 (N_214,In_436,In_2243);
nor U215 (N_215,In_3448,In_4920);
nor U216 (N_216,In_4209,In_4754);
and U217 (N_217,In_1091,In_478);
nor U218 (N_218,In_2872,In_3804);
xnor U219 (N_219,In_3235,In_378);
nand U220 (N_220,In_4167,In_3594);
or U221 (N_221,In_3923,In_1041);
nand U222 (N_222,In_2435,In_2953);
and U223 (N_223,In_142,In_2368);
or U224 (N_224,In_2442,In_1062);
xor U225 (N_225,In_2205,In_3);
xnor U226 (N_226,In_2922,In_2692);
and U227 (N_227,In_4502,In_66);
xnor U228 (N_228,In_3027,In_2242);
and U229 (N_229,In_4930,In_3756);
and U230 (N_230,In_4965,In_1749);
nand U231 (N_231,In_3687,In_2095);
or U232 (N_232,In_2351,In_527);
nor U233 (N_233,In_2604,In_3377);
or U234 (N_234,In_4132,In_2129);
nand U235 (N_235,In_3685,In_2852);
nand U236 (N_236,In_1770,In_3579);
nor U237 (N_237,In_812,In_2479);
xor U238 (N_238,In_3709,In_3538);
xnor U239 (N_239,In_3197,In_704);
nor U240 (N_240,In_3627,In_2817);
nor U241 (N_241,In_1873,In_2186);
nand U242 (N_242,In_3895,In_2722);
xor U243 (N_243,In_645,In_156);
nor U244 (N_244,In_777,In_3704);
xnor U245 (N_245,In_2102,In_316);
nand U246 (N_246,In_3582,In_828);
and U247 (N_247,In_4366,In_2276);
nor U248 (N_248,In_4980,In_716);
and U249 (N_249,In_240,In_2425);
nor U250 (N_250,In_3340,In_752);
or U251 (N_251,In_3935,In_1968);
or U252 (N_252,In_2445,In_4301);
nand U253 (N_253,In_4755,In_4463);
nor U254 (N_254,In_1725,In_1294);
nand U255 (N_255,In_1220,In_1938);
or U256 (N_256,In_3560,In_2000);
xnor U257 (N_257,In_3877,In_1951);
xor U258 (N_258,In_2645,In_826);
xor U259 (N_259,In_1700,In_386);
nand U260 (N_260,In_4883,In_4164);
xor U261 (N_261,In_4813,In_2596);
xor U262 (N_262,In_3132,In_4425);
nor U263 (N_263,In_1242,In_219);
nand U264 (N_264,In_1040,In_1476);
or U265 (N_265,In_1432,In_4026);
and U266 (N_266,In_2156,In_3682);
nand U267 (N_267,In_778,In_2785);
and U268 (N_268,In_1839,In_4566);
nand U269 (N_269,In_688,In_1169);
or U270 (N_270,In_4787,In_4588);
and U271 (N_271,In_2454,In_4519);
or U272 (N_272,In_2027,In_2359);
nand U273 (N_273,In_1752,In_3219);
nor U274 (N_274,In_1809,In_1174);
nor U275 (N_275,In_1318,In_1499);
xnor U276 (N_276,In_3405,In_914);
xor U277 (N_277,In_990,In_3525);
and U278 (N_278,In_4702,In_398);
nand U279 (N_279,In_1643,In_912);
nand U280 (N_280,In_3269,In_3342);
nand U281 (N_281,In_1708,In_1037);
and U282 (N_282,In_855,In_182);
xnor U283 (N_283,In_4445,In_3577);
nor U284 (N_284,In_811,In_817);
or U285 (N_285,In_1515,In_1496);
or U286 (N_286,In_3044,In_4735);
xor U287 (N_287,In_2319,In_770);
nand U288 (N_288,In_1296,In_2385);
nor U289 (N_289,In_4464,In_3016);
nand U290 (N_290,In_1867,In_2117);
nand U291 (N_291,In_3179,In_3671);
nor U292 (N_292,In_4417,In_3257);
or U293 (N_293,In_4901,In_2424);
nand U294 (N_294,In_2013,In_1792);
or U295 (N_295,In_651,In_711);
nand U296 (N_296,In_4310,In_731);
nand U297 (N_297,In_3109,In_693);
and U298 (N_298,In_781,In_169);
nor U299 (N_299,In_2024,In_1067);
nor U300 (N_300,In_2394,In_2201);
nor U301 (N_301,In_372,In_4092);
xor U302 (N_302,In_4955,In_2077);
or U303 (N_303,In_3666,In_2553);
or U304 (N_304,In_528,In_4237);
or U305 (N_305,In_4678,In_2684);
xor U306 (N_306,In_3763,In_3360);
and U307 (N_307,In_224,In_2404);
nand U308 (N_308,In_276,In_4892);
and U309 (N_309,In_3595,In_4918);
nand U310 (N_310,In_4498,In_2822);
or U311 (N_311,In_3633,In_3035);
or U312 (N_312,In_4634,In_2966);
or U313 (N_313,In_758,In_845);
xor U314 (N_314,In_837,In_1085);
nand U315 (N_315,In_4949,In_531);
nor U316 (N_316,In_1478,In_4083);
nand U317 (N_317,In_1954,In_4887);
xnor U318 (N_318,In_2731,In_2290);
or U319 (N_319,In_2561,In_3196);
nand U320 (N_320,In_2902,In_541);
xor U321 (N_321,In_697,In_2939);
xnor U322 (N_322,In_4329,In_1309);
xor U323 (N_323,In_2040,In_3566);
nor U324 (N_324,In_4889,In_520);
and U325 (N_325,In_2159,In_2776);
nand U326 (N_326,In_419,In_1071);
or U327 (N_327,In_1211,In_1375);
xor U328 (N_328,In_2317,In_2214);
nand U329 (N_329,In_4352,In_3977);
and U330 (N_330,In_2315,In_949);
and U331 (N_331,In_2883,In_1715);
nor U332 (N_332,In_2861,In_315);
xnor U333 (N_333,In_1806,In_4840);
nor U334 (N_334,In_4770,In_994);
nor U335 (N_335,In_4385,In_1003);
nand U336 (N_336,In_3498,In_2189);
nor U337 (N_337,In_1563,In_2998);
xnor U338 (N_338,In_958,In_3426);
nand U339 (N_339,In_116,In_4176);
xor U340 (N_340,In_1987,In_1026);
and U341 (N_341,In_2860,In_2698);
nand U342 (N_342,In_248,In_2331);
xor U343 (N_343,In_2682,In_1555);
xor U344 (N_344,In_4434,In_4663);
xor U345 (N_345,In_2413,In_815);
nor U346 (N_346,In_810,In_1245);
or U347 (N_347,In_2778,In_1144);
xor U348 (N_348,In_2629,In_4726);
nand U349 (N_349,In_3981,In_4527);
nor U350 (N_350,In_2680,In_3727);
nor U351 (N_351,In_2643,In_563);
nand U352 (N_352,In_872,In_4643);
and U353 (N_353,In_1204,In_2761);
and U354 (N_354,In_3424,In_4676);
and U355 (N_355,In_1787,In_4667);
and U356 (N_356,In_3778,In_4325);
xnor U357 (N_357,In_4121,In_2572);
nand U358 (N_358,In_3831,In_1352);
and U359 (N_359,In_4543,In_65);
xnor U360 (N_360,In_2874,In_2949);
nand U361 (N_361,In_834,In_4494);
or U362 (N_362,In_388,In_1198);
xnor U363 (N_363,In_576,In_2188);
nor U364 (N_364,In_995,In_1000);
nor U365 (N_365,In_2879,In_76);
nor U366 (N_366,In_4641,In_4473);
nand U367 (N_367,In_3052,In_1533);
nor U368 (N_368,In_2307,In_820);
or U369 (N_369,In_4438,In_2306);
xnor U370 (N_370,In_943,In_2641);
xor U371 (N_371,In_1514,In_1995);
xnor U372 (N_372,In_1286,In_3019);
xnor U373 (N_373,In_1339,In_3184);
nand U374 (N_374,In_1024,In_3456);
xor U375 (N_375,In_853,In_2975);
nand U376 (N_376,In_2630,In_1014);
or U377 (N_377,In_927,In_3624);
nand U378 (N_378,In_579,In_1537);
nand U379 (N_379,In_4761,In_1520);
xor U380 (N_380,In_3411,In_4509);
xnor U381 (N_381,In_4038,In_1685);
and U382 (N_382,In_350,In_228);
xnor U383 (N_383,In_190,In_4261);
nor U384 (N_384,In_2176,In_787);
nor U385 (N_385,In_4000,In_2370);
and U386 (N_386,In_2376,In_1369);
xnor U387 (N_387,In_2971,In_3590);
nand U388 (N_388,In_3803,In_3978);
nand U389 (N_389,In_733,In_1625);
xnor U390 (N_390,In_968,In_4495);
nor U391 (N_391,In_4122,In_4377);
nand U392 (N_392,In_4798,In_236);
nand U393 (N_393,In_2035,In_4626);
and U394 (N_394,In_2416,In_3353);
or U395 (N_395,In_2033,In_1025);
xor U396 (N_396,In_3755,In_3982);
and U397 (N_397,In_3589,In_964);
nor U398 (N_398,In_420,In_749);
or U399 (N_399,In_1645,In_1051);
xor U400 (N_400,In_662,In_925);
xor U401 (N_401,In_2515,In_4064);
nor U402 (N_402,In_2146,In_1280);
nor U403 (N_403,In_1034,In_3245);
nor U404 (N_404,In_1094,In_4854);
nand U405 (N_405,In_1152,In_2167);
and U406 (N_406,In_4897,In_3325);
nand U407 (N_407,In_2237,In_1084);
nor U408 (N_408,In_3773,In_3268);
or U409 (N_409,In_2429,In_739);
or U410 (N_410,In_2485,In_3926);
nor U411 (N_411,In_2719,In_1740);
xor U412 (N_412,In_4902,In_3677);
or U413 (N_413,In_4953,In_2658);
nor U414 (N_414,In_4576,In_2327);
and U415 (N_415,In_4137,In_3850);
or U416 (N_416,In_3591,In_1166);
or U417 (N_417,In_4911,In_1394);
nor U418 (N_418,In_513,In_4278);
nor U419 (N_419,In_4128,In_3177);
nor U420 (N_420,In_3295,In_4822);
and U421 (N_421,In_2585,In_3506);
nand U422 (N_422,In_4469,In_4364);
nand U423 (N_423,In_608,In_2732);
and U424 (N_424,In_4531,In_3661);
nand U425 (N_425,In_1020,In_171);
and U426 (N_426,In_3146,In_3081);
and U427 (N_427,In_3274,In_4675);
xnor U428 (N_428,In_4096,In_4486);
nor U429 (N_429,In_4885,In_3111);
nand U430 (N_430,In_2248,In_1813);
and U431 (N_431,In_4485,In_2651);
nand U432 (N_432,In_2443,In_4259);
or U433 (N_433,In_2105,In_4305);
or U434 (N_434,In_4191,In_3190);
xor U435 (N_435,In_473,In_102);
xnor U436 (N_436,In_629,In_4243);
nor U437 (N_437,In_4172,In_214);
nor U438 (N_438,In_3675,In_3287);
xnor U439 (N_439,In_4085,In_1933);
nand U440 (N_440,In_1902,In_4479);
or U441 (N_441,In_4639,In_3883);
nand U442 (N_442,In_4126,In_1603);
and U443 (N_443,In_3075,In_2134);
or U444 (N_444,In_3681,In_729);
or U445 (N_445,In_1350,In_1561);
nor U446 (N_446,In_1,In_2968);
or U447 (N_447,In_4347,In_1293);
nand U448 (N_448,In_3306,In_3719);
nor U449 (N_449,In_397,In_2391);
nor U450 (N_450,In_4597,In_3210);
or U451 (N_451,In_1682,In_4656);
xor U452 (N_452,In_673,In_2401);
xnor U453 (N_453,In_1733,In_4593);
xnor U454 (N_454,In_1535,In_4169);
nand U455 (N_455,In_2241,In_1846);
xnor U456 (N_456,In_4720,In_4435);
xnor U457 (N_457,In_4027,In_2157);
or U458 (N_458,In_2301,In_2125);
and U459 (N_459,In_3815,In_734);
nor U460 (N_460,In_664,In_4341);
nand U461 (N_461,In_2137,In_4286);
nor U462 (N_462,In_2963,In_3860);
nor U463 (N_463,In_4821,In_81);
xor U464 (N_464,In_383,In_2067);
and U465 (N_465,In_1173,In_1592);
and U466 (N_466,In_3319,In_4940);
and U467 (N_467,In_2568,In_1189);
nand U468 (N_468,In_4936,In_2469);
or U469 (N_469,In_1104,In_3267);
nor U470 (N_470,In_4561,In_4878);
nand U471 (N_471,In_4046,In_3404);
nand U472 (N_472,In_3775,In_104);
and U473 (N_473,In_1524,In_4188);
and U474 (N_474,In_4196,In_4623);
nand U475 (N_475,In_998,In_621);
nand U476 (N_476,In_633,In_1689);
and U477 (N_477,In_2877,In_1497);
or U478 (N_478,In_2127,In_3422);
nor U479 (N_479,In_3749,In_4680);
xnor U480 (N_480,In_2495,In_4684);
nor U481 (N_481,In_412,In_4059);
nor U482 (N_482,In_2239,In_4133);
xor U483 (N_483,In_286,In_1076);
and U484 (N_484,In_357,In_3133);
and U485 (N_485,In_1730,In_2374);
nand U486 (N_486,In_4941,In_4015);
nand U487 (N_487,In_1482,In_2350);
xnor U488 (N_488,In_1364,In_4193);
xor U489 (N_489,In_1259,In_2899);
nand U490 (N_490,In_4742,In_358);
or U491 (N_491,In_4699,In_4114);
and U492 (N_492,In_148,In_940);
or U493 (N_493,In_1033,In_3143);
nand U494 (N_494,In_235,In_3408);
and U495 (N_495,In_2560,In_4521);
xor U496 (N_496,In_1249,In_1306);
or U497 (N_497,In_2916,In_3908);
nor U498 (N_498,In_3122,In_2841);
and U499 (N_499,In_3374,In_3264);
or U500 (N_500,In_2053,In_4267);
and U501 (N_501,In_1413,In_2291);
xnor U502 (N_502,In_487,In_1623);
and U503 (N_503,In_239,In_3009);
xor U504 (N_504,In_1953,In_3136);
and U505 (N_505,In_1738,In_3406);
or U506 (N_506,In_3752,In_2633);
or U507 (N_507,In_3754,In_1079);
or U508 (N_508,In_3317,In_4728);
and U509 (N_509,In_3639,In_354);
xor U510 (N_510,In_1417,In_343);
nor U511 (N_511,In_637,In_4627);
nor U512 (N_512,In_338,In_4369);
or U513 (N_513,In_4748,In_3380);
nor U514 (N_514,In_1074,In_1855);
nor U515 (N_515,In_1030,In_4115);
xor U516 (N_516,In_3403,In_3247);
and U517 (N_517,In_4612,In_2249);
nand U518 (N_518,In_1650,In_3533);
and U519 (N_519,In_2908,In_3414);
nand U520 (N_520,In_3151,In_3313);
or U521 (N_521,In_188,In_4913);
xnor U522 (N_522,In_3028,In_139);
and U523 (N_523,In_3885,In_4244);
nand U524 (N_524,In_4482,In_740);
xor U525 (N_525,In_3417,In_4758);
and U526 (N_526,In_1901,In_2449);
or U527 (N_527,In_2639,In_2533);
or U528 (N_528,In_2891,In_2727);
nand U529 (N_529,In_3300,In_4683);
nor U530 (N_530,In_4618,In_474);
and U531 (N_531,In_2563,In_464);
nand U532 (N_532,In_748,In_2078);
and U533 (N_533,In_4322,In_4817);
nor U534 (N_534,In_808,In_1274);
or U535 (N_535,In_4603,In_4769);
nor U536 (N_536,In_2799,In_173);
xnor U537 (N_537,In_2780,In_1955);
or U538 (N_538,In_2254,In_755);
nand U539 (N_539,In_3943,In_488);
or U540 (N_540,In_4231,In_1196);
or U541 (N_541,In_2037,In_1167);
and U542 (N_542,In_1070,In_4850);
and U543 (N_543,In_3635,In_2687);
xnor U544 (N_544,In_3858,In_3323);
or U545 (N_545,In_2951,In_1228);
or U546 (N_546,In_4960,In_879);
nand U547 (N_547,In_2106,In_2521);
nor U548 (N_548,In_2268,In_10);
xor U549 (N_549,In_3959,In_4087);
nor U550 (N_550,In_1137,In_2679);
xor U551 (N_551,In_1582,In_1447);
or U552 (N_552,In_1876,In_3014);
nor U553 (N_553,In_4468,In_1862);
xnor U554 (N_554,In_4957,In_481);
or U555 (N_555,In_1606,In_3173);
and U556 (N_556,In_1567,In_1066);
nand U557 (N_557,In_368,In_911);
or U558 (N_558,In_4995,In_4008);
or U559 (N_559,In_3558,In_3799);
and U560 (N_560,In_2826,In_512);
or U561 (N_561,In_2014,In_3619);
and U562 (N_562,In_2048,In_4910);
nand U563 (N_563,In_351,In_2562);
nor U564 (N_564,In_4514,In_3462);
xor U565 (N_565,In_3611,In_2029);
or U566 (N_566,In_3030,In_1370);
nand U567 (N_567,In_1233,In_3383);
xor U568 (N_568,In_1462,In_2516);
xor U569 (N_569,In_784,In_1207);
nor U570 (N_570,In_3225,In_1577);
or U571 (N_571,In_1126,In_4528);
xor U572 (N_572,In_1547,In_2648);
and U573 (N_573,In_4441,In_4694);
nor U574 (N_574,In_1005,In_3008);
xor U575 (N_575,In_4510,In_5);
nand U576 (N_576,In_3929,In_2313);
and U577 (N_577,In_2072,In_4563);
and U578 (N_578,In_1264,In_1361);
xor U579 (N_579,In_2348,In_959);
or U580 (N_580,In_1684,In_4493);
and U581 (N_581,In_2163,In_4776);
or U582 (N_582,In_3097,In_4952);
and U583 (N_583,In_4195,In_3435);
and U584 (N_584,In_1895,In_1268);
xnor U585 (N_585,In_3129,In_610);
and U586 (N_586,In_283,In_3203);
nor U587 (N_587,In_4224,In_2557);
xor U588 (N_588,In_905,In_4744);
nand U589 (N_589,In_1970,In_3597);
nor U590 (N_590,In_3650,In_1702);
nand U591 (N_591,In_4160,In_4311);
xor U592 (N_592,In_103,In_2797);
nand U593 (N_593,In_3827,In_3013);
or U594 (N_594,In_4607,In_4055);
nor U595 (N_595,In_3970,In_4963);
nand U596 (N_596,In_3022,In_4651);
or U597 (N_597,In_891,In_2567);
or U598 (N_598,In_1206,In_3148);
and U599 (N_599,In_3444,In_4734);
and U600 (N_600,In_4704,In_2369);
nor U601 (N_601,In_1967,In_2064);
nand U602 (N_602,In_3847,In_4396);
and U603 (N_603,In_1082,In_3707);
and U604 (N_604,In_2549,In_124);
nor U605 (N_605,In_3007,In_3320);
nand U606 (N_606,In_1086,In_455);
and U607 (N_607,In_842,In_4429);
xor U608 (N_608,In_1627,In_1039);
nor U609 (N_609,In_2155,In_2673);
or U610 (N_610,In_1460,In_4512);
or U611 (N_611,In_2810,In_2906);
nor U612 (N_612,In_4615,In_881);
xnor U613 (N_613,In_1410,In_1912);
and U614 (N_614,In_2609,In_4567);
and U615 (N_615,In_4739,In_1265);
nand U616 (N_616,In_1122,In_4775);
nand U617 (N_617,In_1888,In_3114);
nor U618 (N_618,In_3575,In_4042);
or U619 (N_619,In_1190,In_3505);
xor U620 (N_620,In_4779,In_1964);
and U621 (N_621,In_1355,In_4125);
or U622 (N_622,In_132,In_4809);
or U623 (N_623,In_1583,In_1184);
nand U624 (N_624,In_1433,In_3189);
and U625 (N_625,In_3504,In_591);
nand U626 (N_626,In_2339,In_94);
or U627 (N_627,In_2991,In_1756);
nor U628 (N_628,In_3862,In_2801);
nor U629 (N_629,In_3441,In_480);
or U630 (N_630,In_2723,In_2439);
or U631 (N_631,In_4323,In_3968);
xor U632 (N_632,In_3725,In_2280);
or U633 (N_633,In_3213,In_2388);
or U634 (N_634,In_3948,In_4181);
and U635 (N_635,In_1275,In_3509);
nand U636 (N_636,In_2956,In_3690);
or U637 (N_637,In_4319,In_2943);
nand U638 (N_638,In_2502,In_2195);
xor U639 (N_639,In_4524,In_1729);
xor U640 (N_640,In_1996,In_3123);
nand U641 (N_641,In_1785,In_4592);
nand U642 (N_642,In_607,In_2049);
nand U643 (N_643,In_2905,In_462);
xor U644 (N_644,In_4933,In_4357);
xor U645 (N_645,In_1498,In_376);
xor U646 (N_646,In_1448,In_2087);
nand U647 (N_647,In_823,In_2065);
or U648 (N_648,In_3584,In_249);
or U649 (N_649,In_916,In_4437);
and U650 (N_650,In_773,In_4846);
or U651 (N_651,In_1965,In_3464);
nor U652 (N_652,In_1154,In_1958);
nor U653 (N_653,In_1090,In_865);
or U654 (N_654,In_1940,In_2467);
or U655 (N_655,In_1948,In_2403);
or U656 (N_656,In_4477,In_4077);
or U657 (N_657,In_4569,In_2884);
and U658 (N_658,In_341,In_2944);
xor U659 (N_659,In_3880,In_196);
or U660 (N_660,In_4671,In_1305);
and U661 (N_661,In_3521,In_4990);
and U662 (N_662,In_1963,In_2184);
or U663 (N_663,In_3098,In_4937);
nand U664 (N_664,In_3029,In_833);
xor U665 (N_665,In_1517,In_1128);
nand U666 (N_666,In_126,In_4797);
nand U667 (N_667,In_3737,In_360);
nor U668 (N_668,In_3940,In_1120);
nor U669 (N_669,In_1896,In_1936);
nand U670 (N_670,In_2929,In_741);
nor U671 (N_671,In_4226,In_3537);
xor U672 (N_672,In_1576,In_35);
or U673 (N_673,In_470,In_918);
and U674 (N_674,In_3063,In_671);
nand U675 (N_675,In_1253,In_381);
or U676 (N_676,In_3366,In_2433);
or U677 (N_677,In_345,In_4824);
nand U678 (N_678,In_1565,In_1775);
or U679 (N_679,In_1208,In_2747);
nand U680 (N_680,In_391,In_1990);
xnor U681 (N_681,In_4935,In_210);
and U682 (N_682,In_1641,In_663);
xor U683 (N_683,In_2685,In_3873);
or U684 (N_684,In_297,In_4407);
xnor U685 (N_685,In_3899,In_409);
nand U686 (N_686,In_4374,In_500);
nand U687 (N_687,In_3503,In_1927);
nand U688 (N_688,In_1797,In_2364);
xnor U689 (N_689,In_4294,In_3303);
or U690 (N_690,In_2355,In_3892);
and U691 (N_691,In_1856,In_4254);
nand U692 (N_692,In_2221,In_413);
xor U693 (N_693,In_437,In_1288);
xor U694 (N_694,In_3092,In_710);
xnor U695 (N_695,In_4915,In_3648);
nor U696 (N_696,In_317,In_1751);
nand U697 (N_697,In_136,In_1112);
nand U698 (N_698,In_4143,In_3623);
and U699 (N_699,In_4833,In_2311);
xor U700 (N_700,In_582,In_3696);
xor U701 (N_701,In_878,In_3640);
and U702 (N_702,In_738,In_2725);
nor U703 (N_703,In_2224,In_4862);
xnor U704 (N_704,In_1508,In_899);
or U705 (N_705,In_2038,In_4647);
nor U706 (N_706,In_1728,In_1711);
nand U707 (N_707,In_790,In_3476);
nor U708 (N_708,In_3137,In_1469);
and U709 (N_709,In_1042,In_3472);
or U710 (N_710,In_1093,In_100);
nor U711 (N_711,In_4093,In_676);
or U712 (N_712,In_507,In_2162);
and U713 (N_713,In_1999,In_2661);
or U714 (N_714,In_971,In_2103);
nor U715 (N_715,In_4984,In_2179);
and U716 (N_716,In_2507,In_2410);
xnor U717 (N_717,In_3985,In_2566);
and U718 (N_718,In_1673,In_2885);
or U719 (N_719,In_2377,In_3936);
nor U720 (N_720,In_2231,In_4239);
and U721 (N_721,In_2329,In_4896);
xnor U722 (N_722,In_1278,In_322);
or U723 (N_723,In_3367,In_2794);
or U724 (N_724,In_3865,In_3185);
or U725 (N_725,In_1519,In_1349);
and U726 (N_726,In_4379,In_258);
xor U727 (N_727,In_3144,In_166);
nor U728 (N_728,In_4823,In_4003);
and U729 (N_729,In_129,In_1800);
xnor U730 (N_730,In_4031,In_4970);
nand U731 (N_731,In_11,In_241);
nand U732 (N_732,In_4608,In_3261);
nor U733 (N_733,In_675,In_3357);
and U734 (N_734,In_952,In_266);
and U735 (N_735,In_3995,In_2584);
xnor U736 (N_736,In_3385,In_3156);
xor U737 (N_737,In_3625,In_4194);
or U738 (N_738,In_1574,In_212);
and U739 (N_739,In_2539,In_895);
xnor U740 (N_740,In_1942,In_4834);
xor U741 (N_741,In_3262,In_1379);
or U742 (N_742,In_2349,In_4882);
and U743 (N_743,In_3234,In_88);
nor U744 (N_744,In_852,In_1329);
nor U745 (N_745,In_4535,In_4242);
and U746 (N_746,In_2259,In_3421);
and U747 (N_747,In_4490,In_1324);
nand U748 (N_748,In_546,In_4342);
xor U749 (N_749,In_941,In_2450);
or U750 (N_750,In_476,In_22);
and U751 (N_751,In_655,In_4018);
nor U752 (N_752,In_3568,In_3355);
or U753 (N_753,In_4308,In_1134);
and U754 (N_754,In_2004,In_1947);
nor U755 (N_755,In_4011,In_1153);
xor U756 (N_756,In_2702,In_2748);
xnor U757 (N_757,In_4552,In_3649);
xnor U758 (N_758,In_4462,In_439);
or U759 (N_759,In_3988,In_841);
xnor U760 (N_760,In_4966,In_1795);
and U761 (N_761,In_349,In_2444);
nand U762 (N_762,In_4197,In_1248);
nor U763 (N_763,In_2383,In_2784);
or U764 (N_764,In_4879,In_3951);
and U765 (N_765,In_2256,In_2304);
and U766 (N_766,In_457,In_4570);
nand U767 (N_767,In_402,In_4375);
nand U768 (N_768,In_2954,In_2570);
and U769 (N_769,In_2795,In_3794);
nor U770 (N_770,In_38,In_4944);
nand U771 (N_771,In_3291,In_163);
and U772 (N_772,In_1546,In_2379);
nand U773 (N_773,In_3471,In_4022);
or U774 (N_774,In_4698,In_4795);
or U775 (N_775,In_1709,In_1019);
and U776 (N_776,In_339,In_328);
nand U777 (N_777,In_4413,In_1317);
or U778 (N_778,In_3578,In_2530);
or U779 (N_779,In_1031,In_3478);
nor U780 (N_780,In_2589,In_2393);
xor U781 (N_781,In_1534,In_1057);
xor U782 (N_782,In_1371,In_3000);
or U783 (N_783,In_1726,In_3510);
or U784 (N_784,In_1599,In_3820);
or U785 (N_785,In_1089,In_3857);
xnor U786 (N_786,In_4789,In_2468);
xnor U787 (N_787,In_2599,In_2362);
nor U788 (N_788,In_3670,In_3508);
or U789 (N_789,In_4148,In_2158);
nand U790 (N_790,In_835,In_4782);
nor U791 (N_791,In_2207,In_3186);
xnor U792 (N_792,In_2375,In_4240);
and U793 (N_793,In_1596,In_4914);
or U794 (N_794,In_4974,In_367);
nand U795 (N_795,In_4217,In_2779);
or U796 (N_796,In_979,In_764);
and U797 (N_797,In_290,In_486);
or U798 (N_798,In_3110,In_1357);
nand U799 (N_799,In_4442,In_2164);
and U800 (N_800,In_2405,In_3733);
nand U801 (N_801,In_1973,In_2538);
or U802 (N_802,In_2668,In_4853);
nand U803 (N_803,In_2213,In_1127);
and U804 (N_804,In_2253,In_3545);
xnor U805 (N_805,In_1928,In_1474);
xnor U806 (N_806,In_265,In_2458);
or U807 (N_807,In_211,In_3350);
and U808 (N_808,In_611,In_1528);
xor U809 (N_809,In_4088,In_699);
nor U810 (N_810,In_1889,In_2165);
nand U811 (N_811,In_730,In_623);
and U812 (N_812,In_3370,In_3076);
xnor U813 (N_813,In_2613,In_555);
or U814 (N_814,In_3334,In_1063);
nor U815 (N_815,In_3960,In_2019);
nand U816 (N_816,In_3761,In_1231);
xor U817 (N_817,In_4646,In_1124);
xor U818 (N_818,In_2187,In_4135);
and U819 (N_819,In_3828,In_3501);
or U820 (N_820,In_3115,In_883);
or U821 (N_821,In_3634,In_279);
nand U822 (N_822,In_2691,In_867);
and U823 (N_823,In_4036,In_1773);
nand U824 (N_824,In_1282,In_2022);
and U825 (N_825,In_0,In_715);
nor U826 (N_826,In_4219,In_2238);
or U827 (N_827,In_3064,In_1312);
xnor U828 (N_828,In_4110,In_4497);
or U829 (N_829,In_2558,In_2957);
xor U830 (N_830,In_1639,In_3663);
and U831 (N_831,In_2924,In_2172);
or U832 (N_832,In_2250,In_509);
nor U833 (N_833,In_4474,In_1743);
or U834 (N_834,In_3330,In_3181);
xor U835 (N_835,In_119,In_3751);
or U836 (N_836,In_37,In_2919);
xnor U837 (N_837,In_2933,In_3058);
or U838 (N_838,In_1337,In_3381);
xnor U839 (N_839,In_780,In_1644);
xnor U840 (N_840,In_2614,In_646);
nor U841 (N_841,In_3401,In_3906);
xor U842 (N_842,In_4288,In_1359);
nor U843 (N_843,In_4354,In_1027);
and U844 (N_844,In_3792,In_981);
and U845 (N_845,In_3217,In_1863);
nor U846 (N_846,In_3487,In_3614);
nor U847 (N_847,In_3093,In_1008);
xor U848 (N_848,In_2066,In_1121);
xnor U849 (N_849,In_4372,In_2494);
nand U850 (N_850,In_4582,In_4976);
or U851 (N_851,In_3976,In_1386);
nor U852 (N_852,In_3361,In_3630);
nand U853 (N_853,In_1320,In_4816);
xnor U854 (N_854,In_1392,In_4587);
nor U855 (N_855,In_344,In_3051);
nor U856 (N_856,In_2965,In_2517);
nor U857 (N_857,In_4467,In_1982);
nand U858 (N_858,In_4810,In_2367);
nand U859 (N_859,In_4526,In_4788);
nand U860 (N_860,In_2788,In_2950);
and U861 (N_861,In_4579,In_1854);
or U862 (N_862,In_2147,In_1946);
or U863 (N_863,In_3683,In_3972);
nand U864 (N_864,In_3724,In_3279);
and U865 (N_865,In_1762,In_901);
and U866 (N_866,In_3859,In_3788);
or U867 (N_867,In_57,In_3227);
or U868 (N_868,In_3288,In_3620);
xnor U869 (N_869,In_759,In_2670);
nand U870 (N_870,In_3231,In_1103);
or U871 (N_871,In_4805,In_4245);
xnor U872 (N_872,In_4179,In_2173);
nand U873 (N_873,In_1441,In_2247);
or U874 (N_874,In_1402,In_4365);
and U875 (N_875,In_2824,In_234);
nor U876 (N_876,In_4875,In_533);
nor U877 (N_877,In_3212,In_2540);
nand U878 (N_878,In_1354,In_526);
and U879 (N_879,In_4401,In_1619);
or U880 (N_880,In_4161,In_229);
nand U881 (N_881,In_2265,In_1992);
or U882 (N_882,In_1835,In_4706);
or U883 (N_883,In_4622,In_2493);
and U884 (N_884,In_2200,In_1050);
xor U885 (N_885,In_1742,In_3786);
and U886 (N_886,In_1283,In_2847);
or U887 (N_887,In_4381,In_4021);
or U888 (N_888,In_3965,In_3718);
or U889 (N_889,In_4391,In_4162);
and U890 (N_890,In_108,In_1406);
and U891 (N_891,In_3373,In_79);
nor U892 (N_892,In_3921,In_2289);
nand U893 (N_893,In_3147,In_2839);
or U894 (N_894,In_1553,In_4400);
nor U895 (N_895,In_3010,In_2980);
xnor U896 (N_896,In_1986,In_2793);
and U897 (N_897,In_2875,In_4929);
nor U898 (N_898,In_4016,In_2194);
nor U899 (N_899,In_1937,In_1562);
and U900 (N_900,In_1348,In_3050);
xnor U901 (N_901,In_2168,In_2236);
nand U902 (N_902,In_4573,In_1223);
or U903 (N_903,In_2669,In_4600);
xnor U904 (N_904,In_1810,In_4530);
nand U905 (N_905,In_1132,In_4145);
and U906 (N_906,In_4905,In_2911);
nand U907 (N_907,In_1080,In_3636);
xor U908 (N_908,In_1894,In_3530);
nor U909 (N_909,In_174,In_2701);
nor U910 (N_910,In_3281,In_1816);
or U911 (N_911,In_1250,In_586);
nor U912 (N_912,In_4954,In_1811);
xor U913 (N_913,In_2332,In_2894);
or U914 (N_914,In_1172,In_146);
nand U915 (N_915,In_4866,In_4837);
and U916 (N_916,In_2466,In_2461);
nor U917 (N_917,In_3631,In_766);
and U918 (N_918,In_1313,In_4118);
nor U919 (N_919,In_151,In_1843);
nand U920 (N_920,In_3468,In_1422);
nor U921 (N_921,In_4300,In_4496);
and U922 (N_922,In_4326,In_1628);
nand U923 (N_923,In_1763,In_2325);
nor U924 (N_924,In_4102,In_1612);
nand U925 (N_925,In_3695,In_144);
nor U926 (N_926,In_1683,In_4199);
nand U927 (N_927,In_4073,In_3893);
xor U928 (N_928,In_1131,In_1252);
nand U929 (N_929,In_1906,In_3780);
nand U930 (N_930,In_3450,In_2119);
or U931 (N_931,In_3581,In_3991);
and U932 (N_932,In_960,In_1227);
or U933 (N_933,In_3659,In_584);
nor U934 (N_934,In_3844,In_3652);
xor U935 (N_935,In_1769,In_4484);
and U936 (N_936,In_3199,In_4987);
or U937 (N_937,In_2437,In_3393);
xor U938 (N_938,In_4773,In_3502);
xnor U939 (N_939,In_2411,In_2009);
or U940 (N_940,In_2366,In_4466);
xor U941 (N_941,In_3356,In_3240);
nor U942 (N_942,In_1399,In_3710);
and U943 (N_943,In_577,In_750);
nand U944 (N_944,In_1110,In_4156);
xnor U945 (N_945,In_3419,In_340);
nand U946 (N_946,In_3216,In_2142);
nand U947 (N_947,In_3835,In_1116);
nor U948 (N_948,In_2806,In_3047);
xor U949 (N_949,In_4863,In_3824);
nor U950 (N_950,In_2663,In_1712);
xnor U951 (N_951,In_2036,In_2011);
or U952 (N_952,In_721,In_3522);
or U953 (N_953,In_772,In_3866);
xnor U954 (N_954,In_1230,In_2590);
nor U955 (N_955,In_3928,In_2892);
xor U956 (N_956,In_4349,In_2174);
nand U957 (N_957,In_1185,In_1922);
or U958 (N_958,In_4075,In_2426);
or U959 (N_959,In_3800,In_657);
nor U960 (N_960,In_1516,In_3469);
and U961 (N_961,In_2086,In_1777);
or U962 (N_962,In_4912,In_4138);
xor U963 (N_963,In_312,In_1585);
nor U964 (N_964,In_1133,In_928);
or U965 (N_965,In_4948,In_2257);
xor U966 (N_966,In_572,In_2353);
nand U967 (N_967,In_1923,In_1607);
nor U968 (N_968,In_574,In_4924);
and U969 (N_969,In_1284,In_347);
nor U970 (N_970,In_2309,In_2573);
nand U971 (N_971,In_1099,In_2003);
or U972 (N_972,In_2724,In_2081);
xnor U973 (N_973,In_2432,In_517);
nor U974 (N_974,In_333,In_4348);
or U975 (N_975,In_963,In_1731);
or U976 (N_976,In_2012,In_3949);
and U977 (N_977,In_2151,In_1506);
or U978 (N_978,In_314,In_1564);
nand U979 (N_979,In_1038,In_1931);
xnor U980 (N_980,In_4943,In_4652);
nor U981 (N_981,In_3919,In_1541);
nand U982 (N_982,In_3205,In_2270);
and U983 (N_983,In_3598,In_2703);
or U984 (N_984,In_329,In_3628);
xor U985 (N_985,In_1429,In_2925);
and U986 (N_986,In_636,In_1118);
nand U987 (N_987,In_62,In_3107);
and U988 (N_988,In_1823,In_2357);
or U989 (N_989,In_1586,In_2635);
or U990 (N_990,In_42,In_1698);
nand U991 (N_991,In_2121,In_1325);
nand U992 (N_992,In_3962,In_2932);
nor U993 (N_993,In_3797,In_3743);
and U994 (N_994,In_4071,In_2941);
or U995 (N_995,In_186,In_2132);
xnor U996 (N_996,In_274,In_3265);
xnor U997 (N_997,In_2042,In_84);
and U998 (N_998,In_1884,In_1251);
xnor U999 (N_999,In_3532,In_818);
nand U1000 (N_1000,In_4522,In_2926);
or U1001 (N_1001,In_3176,In_874);
xor U1002 (N_1002,In_1851,In_4264);
xor U1003 (N_1003,In_2500,In_844);
nand U1004 (N_1004,In_893,In_2123);
xor U1005 (N_1005,In_3395,In_21);
nor U1006 (N_1006,In_218,In_1604);
nor U1007 (N_1007,In_728,In_4272);
xnor U1008 (N_1008,In_4888,In_3879);
xor U1009 (N_1009,In_604,In_3460);
xnor U1010 (N_1010,In_2219,In_3358);
nand U1011 (N_1011,In_1614,In_1247);
or U1012 (N_1012,In_687,In_609);
or U1013 (N_1013,In_1376,In_4835);
and U1014 (N_1014,In_1657,In_4807);
nand U1015 (N_1015,In_3163,In_4981);
xnor U1016 (N_1016,In_1016,In_1488);
nand U1017 (N_1017,In_722,In_3841);
xnor U1018 (N_1018,In_1828,In_4320);
nand U1019 (N_1019,In_2804,In_3747);
xnor U1020 (N_1020,In_1890,In_1713);
and U1021 (N_1021,In_2813,In_1917);
nor U1022 (N_1022,In_2320,In_594);
or U1023 (N_1023,In_4765,In_4792);
nand U1024 (N_1024,In_890,In_3096);
or U1025 (N_1025,In_3138,In_1006);
or U1026 (N_1026,In_4979,In_2447);
nor U1027 (N_1027,In_4218,In_1415);
xor U1028 (N_1028,In_2490,In_2226);
and U1029 (N_1029,In_1660,In_4869);
xnor U1030 (N_1030,In_40,In_4542);
xnor U1031 (N_1031,In_2481,In_3457);
or U1032 (N_1032,In_4229,In_4668);
nor U1033 (N_1033,In_3587,In_1758);
nor U1034 (N_1034,In_3384,In_694);
and U1035 (N_1035,In_53,In_2617);
nor U1036 (N_1036,In_1620,In_4565);
and U1037 (N_1037,In_2715,In_634);
or U1038 (N_1038,In_1509,In_900);
and U1039 (N_1039,In_3766,In_4183);
nand U1040 (N_1040,In_618,In_1649);
nand U1041 (N_1041,In_4423,In_3391);
and U1042 (N_1042,In_2977,In_3702);
nand U1043 (N_1043,In_1836,In_843);
nand U1044 (N_1044,In_380,In_3104);
xnor U1045 (N_1045,In_2109,In_1240);
and U1046 (N_1046,In_3207,In_4529);
nor U1047 (N_1047,In_4891,In_4968);
nand U1048 (N_1048,In_2116,In_318);
nand U1049 (N_1049,In_3459,In_128);
or U1050 (N_1050,In_2808,In_1858);
xor U1051 (N_1051,In_3071,In_242);
and U1052 (N_1052,In_522,In_2729);
or U1053 (N_1053,In_4414,In_1760);
nor U1054 (N_1054,In_1977,In_3347);
and U1055 (N_1055,In_665,In_9);
or U1056 (N_1056,In_3646,In_2459);
and U1057 (N_1057,In_2897,In_1908);
nand U1058 (N_1058,In_3241,In_3121);
and U1059 (N_1059,In_3284,In_4724);
nor U1060 (N_1060,In_3400,In_744);
nor U1061 (N_1061,In_4746,In_4455);
nor U1062 (N_1062,In_3987,In_2601);
or U1063 (N_1063,In_2853,In_1342);
or U1064 (N_1064,In_1087,In_1720);
xnor U1065 (N_1065,In_1149,In_3020);
xor U1066 (N_1066,In_110,In_4291);
nor U1067 (N_1067,In_570,In_1419);
and U1068 (N_1068,In_1848,In_2111);
or U1069 (N_1069,In_3124,In_3451);
xor U1070 (N_1070,In_3574,In_3479);
nand U1071 (N_1071,In_4134,In_4616);
and U1072 (N_1072,In_3301,In_3868);
or U1073 (N_1073,In_2821,In_2654);
nand U1074 (N_1074,In_2133,In_4750);
xnor U1075 (N_1075,In_3335,In_4630);
and U1076 (N_1076,In_4295,In_3024);
or U1077 (N_1077,In_1744,In_14);
and U1078 (N_1078,In_3170,In_2607);
and U1079 (N_1079,In_4180,In_1310);
nor U1080 (N_1080,In_432,In_31);
nor U1081 (N_1081,In_603,In_2690);
nand U1082 (N_1082,In_3495,In_17);
nand U1083 (N_1083,In_193,In_3442);
xnor U1084 (N_1084,In_4208,In_2486);
or U1085 (N_1085,In_4674,In_1199);
nor U1086 (N_1086,In_4187,In_3606);
and U1087 (N_1087,In_2597,In_3523);
nand U1088 (N_1088,In_2866,In_2697);
and U1089 (N_1089,In_1734,In_3520);
and U1090 (N_1090,In_2496,In_2512);
nor U1091 (N_1091,In_3455,In_3613);
xor U1092 (N_1092,In_953,In_1551);
xor U1093 (N_1093,In_3760,In_2519);
or U1094 (N_1094,In_654,In_3309);
and U1095 (N_1095,In_869,In_1830);
and U1096 (N_1096,In_452,In_4690);
xnor U1097 (N_1097,In_4540,In_4265);
and U1098 (N_1098,In_2324,In_1109);
xnor U1099 (N_1099,In_36,In_3486);
nor U1100 (N_1100,In_1782,In_4617);
nor U1101 (N_1101,In_3876,In_2052);
and U1102 (N_1102,In_1068,In_2460);
xor U1103 (N_1103,In_1140,In_4094);
xor U1104 (N_1104,In_2212,In_1918);
and U1105 (N_1105,In_2942,In_2335);
nor U1106 (N_1106,In_3518,In_4388);
and U1107 (N_1107,In_3990,In_3178);
nand U1108 (N_1108,In_3667,In_854);
nor U1109 (N_1109,In_1270,In_4105);
or U1110 (N_1110,In_3903,In_395);
nor U1111 (N_1111,In_2415,In_1724);
nand U1112 (N_1112,In_1495,In_2487);
and U1113 (N_1113,In_2476,In_3443);
nor U1114 (N_1114,In_4049,In_7);
nor U1115 (N_1115,In_1929,In_3947);
xor U1116 (N_1116,In_440,In_2946);
xor U1117 (N_1117,In_1272,In_1036);
nand U1118 (N_1118,In_2482,In_4358);
xnor U1119 (N_1119,In_1786,In_4221);
nand U1120 (N_1120,In_983,In_4166);
nor U1121 (N_1121,In_268,In_880);
or U1122 (N_1122,In_1686,In_4828);
nor U1123 (N_1123,In_301,In_4583);
nand U1124 (N_1124,In_4343,In_18);
nor U1125 (N_1125,In_3676,In_1256);
xor U1126 (N_1126,In_2303,In_2030);
nand U1127 (N_1127,In_4079,In_1807);
nand U1128 (N_1128,In_1960,In_3224);
nor U1129 (N_1129,In_3744,In_4640);
xor U1130 (N_1130,In_1287,In_3722);
or U1131 (N_1131,In_3070,In_4867);
or U1132 (N_1132,In_1106,In_2235);
or U1133 (N_1133,In_1674,In_1236);
xor U1134 (N_1134,In_4518,In_4395);
and U1135 (N_1135,In_2718,In_4664);
nand U1136 (N_1136,In_1747,In_3853);
or U1137 (N_1137,In_1723,In_1061);
or U1138 (N_1138,In_3791,In_3699);
nand U1139 (N_1139,In_2233,In_552);
or U1140 (N_1140,In_3529,In_4696);
or U1141 (N_1141,In_2744,In_4722);
nor U1142 (N_1142,In_167,In_256);
or U1143 (N_1143,In_3891,In_904);
or U1144 (N_1144,In_628,In_2823);
nor U1145 (N_1145,In_342,In_4589);
and U1146 (N_1146,In_1395,In_680);
xor U1147 (N_1147,In_2488,In_1716);
nand U1148 (N_1148,In_1818,In_4378);
xor U1149 (N_1149,In_622,In_1420);
nand U1150 (N_1150,In_406,In_3580);
xor U1151 (N_1151,In_4268,In_1913);
xnor U1152 (N_1152,In_4001,In_2624);
and U1153 (N_1153,In_4819,In_3420);
xor U1154 (N_1154,In_3025,In_3484);
or U1155 (N_1155,In_4481,In_1569);
and U1156 (N_1156,In_4682,In_2796);
and U1157 (N_1157,In_203,In_3105);
nor U1158 (N_1158,In_1845,In_1271);
xnor U1159 (N_1159,In_4904,In_4283);
xor U1160 (N_1160,In_511,In_1205);
or U1161 (N_1161,In_1114,In_2211);
nand U1162 (N_1162,In_1334,In_3113);
nor U1163 (N_1163,In_4155,In_2175);
nand U1164 (N_1164,In_3139,In_4855);
and U1165 (N_1165,In_4669,In_435);
nor U1166 (N_1166,In_3953,In_230);
or U1167 (N_1167,In_1260,In_3946);
nand U1168 (N_1168,In_4723,In_2586);
xnor U1169 (N_1169,In_335,In_1750);
nor U1170 (N_1170,In_2602,In_3952);
or U1171 (N_1171,In_164,In_656);
xnor U1172 (N_1172,In_4555,In_2714);
nand U1173 (N_1173,In_4147,In_1827);
nand U1174 (N_1174,In_1178,In_3161);
and U1175 (N_1175,In_4480,In_551);
and U1176 (N_1176,In_2059,In_3811);
or U1177 (N_1177,In_2473,In_987);
nand U1178 (N_1178,In_2632,In_3655);
and U1179 (N_1179,In_4389,In_113);
and U1180 (N_1180,In_4753,In_232);
and U1181 (N_1181,In_1693,In_3142);
nor U1182 (N_1182,In_705,In_3787);
and U1183 (N_1183,In_1860,In_2745);
nand U1184 (N_1184,In_3846,In_2982);
or U1185 (N_1185,In_678,In_3642);
xor U1186 (N_1186,In_2912,In_2848);
and U1187 (N_1187,In_3461,In_3017);
nand U1188 (N_1188,In_2815,In_2534);
nor U1189 (N_1189,In_3192,In_4158);
nor U1190 (N_1190,In_1203,In_1526);
or U1191 (N_1191,In_4642,In_3609);
and U1192 (N_1192,In_4931,In_1304);
nor U1193 (N_1193,In_779,In_1642);
nor U1194 (N_1194,In_217,In_4274);
xor U1195 (N_1195,In_3157,In_331);
and U1196 (N_1196,In_3825,In_4273);
and U1197 (N_1197,In_3413,In_3616);
or U1198 (N_1198,In_1598,In_2143);
or U1199 (N_1199,In_4409,In_1925);
and U1200 (N_1200,In_1512,In_1165);
and U1201 (N_1201,In_775,In_64);
and U1202 (N_1202,In_650,In_505);
and U1203 (N_1203,In_4781,In_200);
nand U1204 (N_1204,In_3126,In_4655);
or U1205 (N_1205,In_1882,In_4253);
nand U1206 (N_1206,In_3802,In_4614);
nand U1207 (N_1207,In_3454,In_1175);
nor U1208 (N_1208,In_573,In_578);
nand U1209 (N_1209,In_23,In_2730);
nor U1210 (N_1210,In_3872,In_361);
nand U1211 (N_1211,In_2005,In_2581);
nor U1212 (N_1212,In_3191,In_2605);
and U1213 (N_1213,In_993,In_3942);
nand U1214 (N_1214,In_479,In_1681);
xor U1215 (N_1215,In_3849,In_3665);
or U1216 (N_1216,In_1589,In_4080);
nor U1217 (N_1217,In_3072,In_2193);
and U1218 (N_1218,In_2148,In_4895);
and U1219 (N_1219,In_4207,In_760);
xnor U1220 (N_1220,In_1336,In_1915);
nand U1221 (N_1221,In_1874,In_4387);
nand U1222 (N_1222,In_1994,In_4362);
xor U1223 (N_1223,In_992,In_4633);
xnor U1224 (N_1224,In_3407,In_753);
xnor U1225 (N_1225,In_1257,In_2278);
or U1226 (N_1226,In_4657,In_3032);
and U1227 (N_1227,In_4168,In_4766);
or U1228 (N_1228,In_183,In_4116);
nor U1229 (N_1229,In_3223,In_1217);
nand U1230 (N_1230,In_1609,In_2283);
nand U1231 (N_1231,In_3714,In_583);
nand U1232 (N_1232,In_1671,In_2759);
or U1233 (N_1233,In_3932,In_2330);
nor U1234 (N_1234,In_2108,In_4605);
nand U1235 (N_1235,In_1939,In_4097);
xnor U1236 (N_1236,In_2001,In_137);
and U1237 (N_1237,In_3511,In_1367);
nand U1238 (N_1238,In_652,In_3894);
and U1239 (N_1239,In_1246,In_670);
nand U1240 (N_1240,In_2234,In_134);
or U1241 (N_1241,In_2528,In_2154);
or U1242 (N_1242,In_1158,In_4660);
or U1243 (N_1243,In_4845,In_4868);
and U1244 (N_1244,In_1157,In_4017);
nor U1245 (N_1245,In_3834,In_2340);
and U1246 (N_1246,In_4327,In_1991);
xnor U1247 (N_1247,In_1195,In_568);
nor U1248 (N_1248,In_2085,In_3660);
xnor U1249 (N_1249,In_4731,In_327);
nor U1250 (N_1250,In_433,In_4783);
nor U1251 (N_1251,In_2216,In_4432);
or U1252 (N_1252,In_2293,In_1677);
nand U1253 (N_1253,In_1822,In_2483);
nor U1254 (N_1254,In_2952,In_3209);
or U1255 (N_1255,In_2931,In_33);
nand U1256 (N_1256,In_198,In_424);
xor U1257 (N_1257,In_3565,In_4225);
or U1258 (N_1258,In_3759,In_4010);
nor U1259 (N_1259,In_1194,In_727);
and U1260 (N_1260,In_4297,In_4880);
or U1261 (N_1261,In_1151,In_4465);
and U1262 (N_1262,In_682,In_4206);
or U1263 (N_1263,In_1852,In_926);
and U1264 (N_1264,In_3187,In_2314);
xnor U1265 (N_1265,In_3732,In_4063);
and U1266 (N_1266,In_1510,In_4843);
or U1267 (N_1267,In_2260,In_2575);
and U1268 (N_1268,In_1559,In_2395);
nand U1269 (N_1269,In_1844,In_935);
or U1270 (N_1270,In_4089,In_2660);
nand U1271 (N_1271,In_3808,In_50);
xor U1272 (N_1272,In_4041,In_3128);
nand U1273 (N_1273,In_3214,In_155);
or U1274 (N_1274,In_4198,In_2775);
xor U1275 (N_1275,In_3605,In_4443);
xor U1276 (N_1276,In_363,In_1675);
nand U1277 (N_1277,In_689,In_1254);
nand U1278 (N_1278,In_876,In_3314);
nor U1279 (N_1279,In_858,In_3867);
nand U1280 (N_1280,In_698,In_988);
and U1281 (N_1281,In_4686,In_194);
xor U1282 (N_1282,In_3049,In_1123);
nor U1283 (N_1283,In_2057,In_3583);
or U1284 (N_1284,In_2631,In_1044);
or U1285 (N_1285,In_1046,In_2829);
nor U1286 (N_1286,In_4900,In_1525);
nor U1287 (N_1287,In_3641,In_1801);
nand U1288 (N_1288,In_4923,In_3626);
nor U1289 (N_1289,In_3668,In_873);
or U1290 (N_1290,In_955,In_3275);
nor U1291 (N_1291,In_684,In_2455);
and U1292 (N_1292,In_2756,In_293);
nor U1293 (N_1293,In_411,In_4687);
nand U1294 (N_1294,In_2983,In_325);
nand U1295 (N_1295,In_4227,In_1012);
xor U1296 (N_1296,In_2527,In_1241);
nor U1297 (N_1297,In_2959,In_4500);
nand U1298 (N_1298,In_4024,In_4881);
and U1299 (N_1299,In_859,In_1779);
nand U1300 (N_1300,In_767,In_4234);
nor U1301 (N_1301,In_1218,In_496);
nor U1302 (N_1302,In_4771,In_1049);
xnor U1303 (N_1303,In_3818,In_2492);
and U1304 (N_1304,In_272,In_703);
nor U1305 (N_1305,In_2373,In_3563);
nor U1306 (N_1306,In_207,In_3909);
xnor U1307 (N_1307,In_2272,In_4163);
nor U1308 (N_1308,In_3961,In_1838);
or U1309 (N_1309,In_498,In_1865);
and U1310 (N_1310,In_709,In_4725);
or U1311 (N_1311,In_4718,In_2141);
and U1312 (N_1312,In_3282,In_3324);
nand U1313 (N_1313,In_2882,In_1043);
xnor U1314 (N_1314,In_3333,In_4013);
nor U1315 (N_1315,In_1966,In_2840);
nand U1316 (N_1316,In_3924,In_2074);
xnor U1317 (N_1317,In_3467,In_862);
nand U1318 (N_1318,In_2489,In_3046);
or U1319 (N_1319,In_1381,In_71);
nor U1320 (N_1320,In_281,In_2726);
xnor U1321 (N_1321,In_2717,In_2984);
xnor U1322 (N_1322,In_1302,In_4768);
nand U1323 (N_1323,In_4985,In_2625);
nand U1324 (N_1324,In_61,In_1549);
or U1325 (N_1325,In_2092,In_4420);
or U1326 (N_1326,In_690,In_1382);
and U1327 (N_1327,In_700,In_954);
or U1328 (N_1328,In_2556,In_285);
nand U1329 (N_1329,In_2750,In_4318);
nor U1330 (N_1330,In_3130,In_3980);
nand U1331 (N_1331,In_530,In_1279);
or U1332 (N_1332,In_1803,In_1022);
and U1333 (N_1333,In_2878,In_223);
and U1334 (N_1334,In_407,In_2720);
nor U1335 (N_1335,In_2864,In_3678);
nor U1336 (N_1336,In_3551,In_3289);
nor U1337 (N_1337,In_4536,In_2097);
nand U1338 (N_1338,In_2986,In_2930);
xnor U1339 (N_1339,In_2903,In_3409);
and U1340 (N_1340,In_757,In_1423);
nor U1341 (N_1341,In_540,In_1341);
or U1342 (N_1342,In_4215,In_4631);
or U1343 (N_1343,In_4235,In_2101);
and U1344 (N_1344,In_2849,In_4740);
nor U1345 (N_1345,In_4511,In_3285);
nand U1346 (N_1346,In_1450,In_3686);
or U1347 (N_1347,In_1688,In_907);
and U1348 (N_1348,In_3003,In_1451);
and U1349 (N_1349,In_1664,In_3368);
nand U1350 (N_1350,In_2636,In_892);
nand U1351 (N_1351,In_1721,In_1618);
or U1352 (N_1352,In_1285,In_1841);
or U1353 (N_1353,In_863,In_41);
and U1354 (N_1354,In_1171,In_3527);
xor U1355 (N_1355,In_3572,In_4213);
or U1356 (N_1356,In_2678,In_2546);
xor U1357 (N_1357,In_3318,In_1799);
nor U1358 (N_1358,In_1975,In_1802);
or U1359 (N_1359,In_1500,In_3440);
xor U1360 (N_1360,In_2465,In_3332);
nor U1361 (N_1361,In_553,In_332);
nor U1362 (N_1362,In_4222,In_4727);
nand U1363 (N_1363,In_2774,In_1142);
and U1364 (N_1364,In_401,In_2644);
xnor U1365 (N_1365,In_1850,In_1483);
and U1366 (N_1366,In_3555,In_2297);
or U1367 (N_1367,In_52,In_1655);
or U1368 (N_1368,In_1941,In_4317);
or U1369 (N_1369,In_441,In_1035);
nor U1370 (N_1370,In_2522,In_2171);
nand U1371 (N_1371,In_4029,In_3470);
or U1372 (N_1372,In_2,In_3957);
nor U1373 (N_1373,In_933,In_2382);
xor U1374 (N_1374,In_4688,In_1077);
or U1375 (N_1375,In_3573,In_1192);
xor U1376 (N_1376,In_3771,In_2408);
xnor U1377 (N_1377,In_2113,In_672);
or U1378 (N_1378,In_1971,In_1748);
nand U1379 (N_1379,In_2620,In_4865);
or U1380 (N_1380,In_2655,In_3544);
nand U1381 (N_1381,In_2961,In_2017);
nor U1382 (N_1382,In_1481,In_4426);
nor U1383 (N_1383,In_1326,In_1428);
or U1384 (N_1384,In_123,In_1209);
and U1385 (N_1385,In_4284,In_3554);
and U1386 (N_1386,In_3705,In_3386);
and U1387 (N_1387,In_2251,In_4697);
or U1388 (N_1388,In_2880,In_2296);
nand U1389 (N_1389,In_1238,In_3726);
and U1390 (N_1390,In_444,In_1909);
or U1391 (N_1391,In_4786,In_3149);
xor U1392 (N_1392,In_288,In_2084);
nand U1393 (N_1393,In_934,In_1745);
and U1394 (N_1394,In_364,In_4149);
xnor U1395 (N_1395,In_805,In_2088);
or U1396 (N_1396,In_2160,In_4202);
and U1397 (N_1397,In_4223,In_2028);
and U1398 (N_1398,In_3293,In_308);
and U1399 (N_1399,In_1790,In_4997);
or U1400 (N_1400,In_4475,In_2288);
xnor U1401 (N_1401,In_4051,In_1511);
nand U1402 (N_1402,In_4247,In_1338);
nand U1403 (N_1403,In_3183,In_1484);
nor U1404 (N_1404,In_447,In_1388);
nand U1405 (N_1405,In_1536,In_1028);
nand U1406 (N_1406,In_1571,In_796);
or U1407 (N_1407,In_1853,In_1289);
nand U1408 (N_1408,In_3603,In_735);
and U1409 (N_1409,In_882,In_4281);
or U1410 (N_1410,In_3694,In_3911);
nand U1411 (N_1411,In_3119,In_4174);
and U1412 (N_1412,In_1372,In_2598);
or U1413 (N_1413,In_4361,In_523);
or U1414 (N_1414,In_674,In_4005);
and U1415 (N_1415,In_485,In_3941);
xnor U1416 (N_1416,In_1602,In_3541);
nor U1417 (N_1417,In_4876,In_587);
xor U1418 (N_1418,In_931,In_2279);
nor U1419 (N_1419,In_1840,In_4399);
xor U1420 (N_1420,In_3494,In_2114);
and U1421 (N_1421,In_1558,In_2854);
xnor U1422 (N_1422,In_2457,In_4715);
or U1423 (N_1423,In_4928,In_2402);
and U1424 (N_1424,In_3989,In_2855);
or U1425 (N_1425,In_122,In_3489);
or U1426 (N_1426,In_4763,In_4390);
or U1427 (N_1427,In_3934,In_4421);
xor U1428 (N_1428,In_884,In_2792);
nand U1429 (N_1429,In_2921,In_2264);
nor U1430 (N_1430,In_754,In_3260);
and U1431 (N_1431,In_518,In_2390);
nand U1432 (N_1432,In_115,In_3586);
or U1433 (N_1433,In_4101,In_4751);
xor U1434 (N_1434,In_732,In_691);
nand U1435 (N_1435,In_4120,In_153);
nor U1436 (N_1436,In_913,In_2274);
or U1437 (N_1437,In_2144,In_4277);
nor U1438 (N_1438,In_1857,In_3481);
xnor U1439 (N_1439,In_4257,In_2318);
and U1440 (N_1440,In_4488,In_1820);
or U1441 (N_1441,In_3526,In_4057);
xnor U1442 (N_1442,In_2255,In_3917);
xor U1443 (N_1443,In_2816,In_2606);
or U1444 (N_1444,In_4499,In_1566);
or U1445 (N_1445,In_3875,In_3973);
xor U1446 (N_1446,In_4791,In_4558);
nand U1447 (N_1447,In_3202,In_3094);
or U1448 (N_1448,In_4922,In_161);
or U1449 (N_1449,In_1013,In_1366);
and U1450 (N_1450,In_68,In_2245);
or U1451 (N_1451,In_3060,In_769);
and U1452 (N_1452,In_2131,In_1225);
and U1453 (N_1453,In_1833,In_4700);
or U1454 (N_1454,In_2252,In_3956);
nand U1455 (N_1455,In_32,In_3048);
nand U1456 (N_1456,In_4677,In_267);
xor U1457 (N_1457,In_4249,In_2090);
or U1458 (N_1458,In_2611,In_2987);
nand U1459 (N_1459,In_937,In_543);
nand U1460 (N_1460,In_4020,In_3006);
xor U1461 (N_1461,In_159,In_4404);
xnor U1462 (N_1462,In_215,In_4890);
nand U1463 (N_1463,In_1234,In_3819);
nand U1464 (N_1464,In_4332,In_4716);
xnor U1465 (N_1465,In_2421,In_1766);
xnor U1466 (N_1466,In_2010,In_4066);
nor U1467 (N_1467,In_2041,In_4559);
nor U1468 (N_1468,In_2993,In_1064);
nand U1469 (N_1469,In_2869,In_472);
nor U1470 (N_1470,In_3140,In_3769);
nor U1471 (N_1471,In_1295,In_2554);
nor U1472 (N_1472,In_2901,In_708);
or U1473 (N_1473,In_3864,In_80);
or U1474 (N_1474,In_3920,In_717);
xnor U1475 (N_1475,In_945,In_3602);
nand U1476 (N_1476,In_2021,In_567);
nand U1477 (N_1477,In_626,In_4359);
xnor U1478 (N_1478,In_4917,In_261);
nand U1479 (N_1479,In_1605,In_2696);
nor U1480 (N_1480,In_453,In_86);
nor U1481 (N_1481,In_4925,In_2913);
and U1482 (N_1482,In_1486,In_565);
or U1483 (N_1483,In_4324,In_2577);
nand U1484 (N_1484,In_4802,In_564);
xor U1485 (N_1485,In_1550,In_3723);
xor U1486 (N_1486,In_294,In_2595);
or U1487 (N_1487,In_3436,In_3781);
and U1488 (N_1488,In_596,In_269);
xnor U1489 (N_1489,In_2118,In_4360);
nand U1490 (N_1490,In_4852,In_2582);
nor U1491 (N_1491,In_1346,In_643);
and U1492 (N_1492,In_1244,In_2979);
or U1493 (N_1493,In_1753,In_4778);
nand U1494 (N_1494,In_589,In_3701);
xor U1495 (N_1495,In_1885,In_3812);
and U1496 (N_1496,In_4525,In_1771);
nand U1497 (N_1497,In_1632,In_2337);
and U1498 (N_1498,In_4774,In_4993);
or U1499 (N_1499,In_2686,In_3087);
xor U1500 (N_1500,In_2667,In_3074);
nand U1501 (N_1501,In_1663,In_1107);
and U1502 (N_1502,In_1530,In_2976);
and U1503 (N_1503,In_1540,In_1696);
nand U1504 (N_1504,In_4998,In_538);
or U1505 (N_1505,In_1849,In_3412);
nand U1506 (N_1506,In_400,In_792);
and U1507 (N_1507,In_4908,In_2634);
or U1508 (N_1508,In_3821,In_1900);
nand U1509 (N_1509,In_3276,In_1610);
and U1510 (N_1510,In_798,In_4009);
nor U1511 (N_1511,In_4236,In_4458);
xnor U1512 (N_1512,In_495,In_1162);
xnor U1513 (N_1513,In_1139,In_4959);
or U1514 (N_1514,In_4182,In_2400);
nand U1515 (N_1515,In_2381,In_3535);
and U1516 (N_1516,In_1668,In_4975);
nand U1517 (N_1517,In_3354,In_4450);
nor U1518 (N_1518,In_4950,In_3550);
or U1519 (N_1519,In_4513,In_1543);
or U1520 (N_1520,In_2076,In_2025);
nor U1521 (N_1521,In_4330,In_1315);
nor U1522 (N_1522,In_889,In_4594);
nand U1523 (N_1523,In_2592,In_3736);
xnor U1524 (N_1524,In_4780,In_2876);
or U1525 (N_1525,In_3829,In_1333);
and U1526 (N_1526,In_1578,In_803);
nand U1527 (N_1527,In_4794,In_3793);
xor U1528 (N_1528,In_216,In_2323);
xnor U1529 (N_1529,In_525,In_2506);
xor U1530 (N_1530,In_247,In_1290);
nor U1531 (N_1531,In_3091,In_4662);
nand U1532 (N_1532,In_4402,In_620);
xor U1533 (N_1533,In_410,In_12);
nand U1534 (N_1534,In_2945,In_1962);
or U1535 (N_1535,In_2616,In_2177);
xnor U1536 (N_1536,In_3901,In_60);
nor U1537 (N_1537,In_3777,In_191);
xor U1538 (N_1538,In_392,In_3226);
or U1539 (N_1539,In_4287,In_1096);
or U1540 (N_1540,In_4958,In_133);
xor U1541 (N_1541,In_966,In_2183);
or U1542 (N_1542,In_1796,In_4131);
nor U1543 (N_1543,In_2704,In_3662);
or U1544 (N_1544,In_3086,In_1631);
or U1545 (N_1545,In_2865,In_588);
nand U1546 (N_1546,In_2504,In_1444);
and U1547 (N_1547,In_2771,In_947);
and U1548 (N_1548,In_939,In_4368);
and U1549 (N_1549,In_2228,In_284);
nand U1550 (N_1550,In_1409,In_4052);
xor U1551 (N_1551,In_56,In_1697);
and U1552 (N_1552,In_3034,In_1652);
xor U1553 (N_1553,In_3708,In_326);
or U1554 (N_1554,In_4703,In_2600);
xnor U1555 (N_1555,In_3768,In_4069);
or U1556 (N_1556,In_932,In_1083);
or U1557 (N_1557,In_2947,In_257);
or U1558 (N_1558,In_2328,In_3165);
and U1559 (N_1559,In_2828,In_3485);
and U1560 (N_1560,In_2292,In_4549);
and U1561 (N_1561,In_138,In_3693);
nand U1562 (N_1562,In_246,In_894);
xnor U1563 (N_1563,In_4262,In_2499);
and U1564 (N_1564,In_3717,In_822);
nand U1565 (N_1565,In_562,In_423);
nand U1566 (N_1566,In_4448,In_4422);
xor U1567 (N_1567,In_1667,In_3713);
nor U1568 (N_1568,In_125,In_644);
nor U1569 (N_1569,In_4315,In_3326);
nor U1570 (N_1570,In_2020,In_2396);
and U1571 (N_1571,In_3638,In_942);
and U1572 (N_1572,In_3372,In_4557);
nor U1573 (N_1573,In_4601,In_661);
or U1574 (N_1574,In_4921,In_847);
nand U1575 (N_1575,In_930,In_2427);
xor U1576 (N_1576,In_2825,In_1666);
and U1577 (N_1577,In_800,In_4857);
and U1578 (N_1578,In_4635,In_2571);
xnor U1579 (N_1579,In_3369,In_3108);
nand U1580 (N_1580,In_3206,In_2229);
xor U1581 (N_1581,In_4436,In_176);
nor U1582 (N_1582,In_371,In_2352);
or U1583 (N_1583,In_1168,In_936);
or U1584 (N_1584,In_4025,In_29);
xor U1585 (N_1585,In_2652,In_1542);
and U1586 (N_1586,In_1130,In_3955);
nor U1587 (N_1587,In_2862,In_2881);
nor U1588 (N_1588,In_259,In_2510);
nand U1589 (N_1589,In_4757,In_1570);
nor U1590 (N_1590,In_2681,In_3043);
xnor U1591 (N_1591,In_2523,In_4648);
xnor U1592 (N_1592,In_3195,In_3540);
nor U1593 (N_1593,In_4293,In_2683);
xor U1594 (N_1594,In_4560,In_600);
or U1595 (N_1595,In_3979,In_3259);
and U1596 (N_1596,In_4478,In_47);
nor U1597 (N_1597,In_593,In_4);
nor U1598 (N_1598,In_797,In_2436);
xor U1599 (N_1599,In_3447,In_4047);
xor U1600 (N_1600,In_4449,In_4586);
nor U1601 (N_1601,In_590,In_2322);
or U1602 (N_1602,In_4012,In_2994);
or U1603 (N_1603,In_2777,In_857);
nand U1604 (N_1604,In_2626,In_287);
nor U1605 (N_1605,In_3344,In_3994);
or U1606 (N_1606,In_365,In_418);
and U1607 (N_1607,In_2333,In_4961);
and U1608 (N_1608,In_2734,In_1545);
nor U1609 (N_1609,In_4806,In_13);
nor U1610 (N_1610,In_1998,In_746);
or U1611 (N_1611,In_3059,In_1626);
nand U1612 (N_1612,In_3193,In_497);
nor U1613 (N_1613,In_2992,In_2032);
nor U1614 (N_1614,In_2541,In_3657);
xor U1615 (N_1615,In_1435,In_2203);
nand U1616 (N_1616,In_4127,In_1892);
xnor U1617 (N_1617,In_2082,In_4037);
or U1618 (N_1618,In_2695,In_1007);
and U1619 (N_1619,In_2326,In_2850);
or U1620 (N_1620,In_2452,In_3507);
nor U1621 (N_1621,In_2286,In_4762);
and U1622 (N_1622,In_2803,In_2063);
and U1623 (N_1623,In_1092,In_3975);
nand U1624 (N_1624,In_4072,In_3644);
nor U1625 (N_1625,In_3307,In_3363);
and U1626 (N_1626,In_2712,In_1179);
or U1627 (N_1627,In_3397,In_2055);
or U1628 (N_1628,In_801,In_2574);
or U1629 (N_1629,In_1636,In_3782);
nand U1630 (N_1630,In_3033,In_875);
nand U1631 (N_1631,In_4192,In_2856);
xor U1632 (N_1632,In_3612,In_233);
or U1633 (N_1633,In_4992,In_1426);
and U1634 (N_1634,In_54,In_3783);
nand U1635 (N_1635,In_1161,In_221);
and U1636 (N_1636,In_3913,In_1299);
and U1637 (N_1637,In_3922,In_910);
nor U1638 (N_1638,In_3263,In_3100);
nor U1639 (N_1639,In_1378,In_1826);
or U1640 (N_1640,In_702,In_1018);
nand U1641 (N_1641,In_1518,In_1216);
nor U1642 (N_1642,In_3430,In_1430);
and U1643 (N_1643,In_946,In_2752);
xor U1644 (N_1644,In_3762,In_3327);
xor U1645 (N_1645,In_3429,In_1842);
or U1646 (N_1646,In_4350,In_4814);
nor U1647 (N_1647,In_4141,In_4826);
and U1648 (N_1648,In_1136,In_2843);
and U1649 (N_1649,In_1859,In_2741);
or U1650 (N_1650,In_2185,In_4672);
xnor U1651 (N_1651,In_4220,In_244);
xor U1652 (N_1652,In_1615,In_489);
or U1653 (N_1653,In_561,In_1277);
xor U1654 (N_1654,In_4056,In_2650);
or U1655 (N_1655,In_477,In_3041);
or U1656 (N_1656,In_2058,In_1391);
or U1657 (N_1657,In_2638,In_679);
or U1658 (N_1658,In_4152,In_4084);
nand U1659 (N_1659,In_1239,In_2462);
xor U1660 (N_1660,In_3562,In_906);
or U1661 (N_1661,In_4838,In_2765);
and U1662 (N_1662,In_4665,In_404);
or U1663 (N_1663,In_2099,In_1717);
nand U1664 (N_1664,In_980,In_3038);
and U1665 (N_1665,In_3125,In_814);
or U1666 (N_1666,In_3031,In_3004);
and U1667 (N_1667,In_2098,In_3180);
nor U1668 (N_1668,In_785,In_4977);
nand U1669 (N_1669,In_3731,In_3228);
and U1670 (N_1670,In_816,In_3742);
or U1671 (N_1671,In_2845,In_483);
or U1672 (N_1672,In_614,In_1678);
or U1673 (N_1673,In_3882,In_3854);
or U1674 (N_1674,In_624,In_4632);
nor U1675 (N_1675,In_4903,In_3018);
and U1676 (N_1676,In_131,In_3674);
and U1677 (N_1677,In_4419,In_619);
and U1678 (N_1678,In_3394,In_1691);
or U1679 (N_1679,In_3079,In_4551);
or U1680 (N_1680,In_2471,In_534);
xor U1681 (N_1681,In_109,In_1988);
xor U1682 (N_1682,In_1197,In_1119);
nor U1683 (N_1683,In_369,In_601);
xnor U1684 (N_1684,In_4945,In_3735);
xnor U1685 (N_1685,In_3434,In_3237);
nor U1686 (N_1686,In_2886,In_549);
or U1687 (N_1687,In_2026,In_3037);
nand U1688 (N_1688,In_4501,In_2448);
nand U1689 (N_1689,In_1436,In_4140);
nor U1690 (N_1690,In_4839,In_3878);
xor U1691 (N_1691,In_4112,In_4201);
nor U1692 (N_1692,In_1579,In_3162);
or U1693 (N_1693,In_1424,In_106);
nor U1694 (N_1694,In_1507,In_1380);
or U1695 (N_1695,In_466,In_4260);
xor U1696 (N_1696,In_3905,In_201);
and U1697 (N_1697,In_2018,In_187);
nand U1698 (N_1698,In_416,In_83);
or U1699 (N_1699,In_389,In_70);
and U1700 (N_1700,In_4340,In_1115);
nand U1701 (N_1701,In_4711,In_838);
nor U1702 (N_1702,In_4398,In_2047);
or U1703 (N_1703,In_3021,In_3338);
nand U1704 (N_1704,In_2210,In_4714);
xor U1705 (N_1705,In_1532,In_1847);
xor U1706 (N_1706,In_1467,In_2672);
and U1707 (N_1707,In_3600,In_1872);
xor U1708 (N_1708,In_4927,In_1397);
nor U1709 (N_1709,In_2334,In_2080);
nor U1710 (N_1710,In_4457,In_3423);
nor U1711 (N_1711,In_3688,In_2623);
or U1712 (N_1712,In_3593,In_4829);
xnor U1713 (N_1713,In_2342,In_1861);
nor U1714 (N_1714,In_3135,In_2964);
nor U1715 (N_1715,In_2136,In_3758);
or U1716 (N_1716,In_4772,In_4159);
nor U1717 (N_1717,In_4252,In_3103);
nor U1718 (N_1718,In_2209,In_2356);
or U1719 (N_1719,In_1788,In_3716);
or U1720 (N_1720,In_3944,In_321);
nor U1721 (N_1721,In_1957,In_658);
xnor U1722 (N_1722,In_3515,In_3963);
xnor U1723 (N_1723,In_2277,In_3615);
nor U1724 (N_1724,In_782,In_4532);
and U1725 (N_1725,In_585,In_1443);
nand U1726 (N_1726,In_3534,In_2811);
xor U1727 (N_1727,In_3244,In_2768);
and U1728 (N_1728,In_1501,In_4666);
nor U1729 (N_1729,In_1554,In_1961);
nand U1730 (N_1730,In_89,In_1699);
xor U1731 (N_1731,In_1401,In_4290);
or U1732 (N_1732,In_27,In_1060);
xnor U1733 (N_1733,In_1345,In_2757);
nor U1734 (N_1734,In_3204,In_3805);
xnor U1735 (N_1735,In_3328,In_1670);
nand U1736 (N_1736,In_3871,In_3218);
or U1737 (N_1737,In_4729,In_868);
nor U1738 (N_1738,In_4747,In_2830);
xor U1739 (N_1739,In_4383,In_1385);
xnor U1740 (N_1740,In_771,In_1470);
or U1741 (N_1741,In_1513,In_2738);
nand U1742 (N_1742,In_3233,In_442);
and U1743 (N_1743,In_2665,In_3837);
nor U1744 (N_1744,In_2772,In_59);
nor U1745 (N_1745,In_1878,In_4334);
or U1746 (N_1746,In_1180,In_3888);
and U1747 (N_1747,In_4393,In_2312);
nor U1748 (N_1748,In_1943,In_763);
nand U1749 (N_1749,In_1661,In_4232);
xnor U1750 (N_1750,In_1389,In_96);
and U1751 (N_1751,In_1215,In_542);
or U1752 (N_1752,In_3907,In_3816);
nor U1753 (N_1753,In_3539,In_19);
nand U1754 (N_1754,In_4659,In_243);
and U1755 (N_1755,In_4394,In_4054);
nor U1756 (N_1756,In_2501,In_3375);
nor U1757 (N_1757,In_4893,In_1269);
or U1758 (N_1758,In_3912,In_4658);
and U1759 (N_1759,In_1343,In_2675);
nand U1760 (N_1760,In_2763,In_4030);
nand U1761 (N_1761,In_4799,In_3915);
nand U1762 (N_1762,In_1552,In_3292);
nor U1763 (N_1763,In_3814,In_836);
nor U1764 (N_1764,In_4541,In_631);
xor U1765 (N_1765,In_320,In_1307);
nand U1766 (N_1766,In_544,In_3222);
or U1767 (N_1767,In_747,In_4650);
xnor U1768 (N_1768,In_4405,In_2006);
xor U1769 (N_1769,In_484,In_1950);
or U1770 (N_1770,In_3445,In_1556);
nor U1771 (N_1771,In_482,In_1456);
nor U1772 (N_1772,In_944,In_4760);
or U1773 (N_1773,In_1222,In_2414);
xor U1774 (N_1774,In_4171,In_4113);
nand U1775 (N_1775,In_2464,In_888);
or U1776 (N_1776,In_73,In_3823);
and U1777 (N_1777,In_2529,In_4884);
nand U1778 (N_1778,In_2100,In_2428);
nand U1779 (N_1779,In_3516,In_3703);
xnor U1780 (N_1780,In_2225,In_1630);
nor U1781 (N_1781,In_4969,In_765);
xor U1782 (N_1782,In_2588,In_4951);
nand U1783 (N_1783,In_2591,In_2851);
or U1784 (N_1784,In_4907,In_3680);
or U1785 (N_1785,In_3243,In_1081);
and U1786 (N_1786,In_1580,In_1875);
nor U1787 (N_1787,In_1590,In_2812);
nand U1788 (N_1788,In_300,In_724);
nand U1789 (N_1789,In_3336,In_1869);
or U1790 (N_1790,In_3095,In_330);
or U1791 (N_1791,In_806,In_1588);
nor U1792 (N_1792,In_3449,In_4800);
nand U1793 (N_1793,In_1048,In_1759);
or U1794 (N_1794,In_3998,In_4279);
or U1795 (N_1795,In_3874,In_1113);
or U1796 (N_1796,In_2514,In_1669);
and U1797 (N_1797,In_2294,In_3005);
nor U1798 (N_1798,In_3198,In_4345);
and U1799 (N_1799,In_1573,In_2751);
nor U1800 (N_1800,In_4460,In_4515);
or U1801 (N_1801,In_2532,In_3253);
and U1802 (N_1802,In_2115,In_4406);
and U1803 (N_1803,In_2262,In_4550);
or U1804 (N_1804,In_3239,In_2749);
nor U1805 (N_1805,In_3832,In_2525);
xnor U1806 (N_1806,In_4157,In_4230);
and U1807 (N_1807,In_1301,In_2474);
or U1808 (N_1808,In_2868,In_1311);
or U1809 (N_1809,In_1597,In_4430);
or U1810 (N_1810,In_2300,In_2299);
and U1811 (N_1811,In_3280,In_3863);
xor U1812 (N_1812,In_4142,In_4625);
nand U1813 (N_1813,In_745,In_2863);
and U1814 (N_1814,In_2713,In_305);
and U1815 (N_1815,In_1492,In_1804);
or U1816 (N_1816,In_819,In_529);
or U1817 (N_1817,In_1347,In_3167);
xnor U1818 (N_1818,In_2418,In_2846);
or U1819 (N_1819,In_2694,In_2888);
nand U1820 (N_1820,In_4117,In_4721);
xor U1821 (N_1821,In_2152,In_1465);
xnor U1822 (N_1822,In_1393,In_2552);
nand U1823 (N_1823,In_3278,In_2898);
nand U1824 (N_1824,In_1907,In_831);
nor U1825 (N_1825,In_3592,In_1145);
nand U1826 (N_1826,In_51,In_270);
nor U1827 (N_1827,In_4649,In_902);
xor U1828 (N_1828,In_2935,In_408);
or U1829 (N_1829,In_1344,In_4045);
xor U1830 (N_1830,In_1442,In_613);
and U1831 (N_1831,In_4346,In_4553);
xor U1832 (N_1832,In_2096,In_227);
or U1833 (N_1833,In_3496,In_1665);
or U1834 (N_1834,In_2316,In_3645);
xnor U1835 (N_1835,In_3933,In_2657);
xor U1836 (N_1836,In_375,In_3543);
or U1837 (N_1837,In_1303,In_1656);
and U1838 (N_1838,In_827,In_4380);
xor U1839 (N_1839,In_4644,In_184);
and U1840 (N_1840,In_4571,In_1176);
or U1841 (N_1841,In_4006,In_4964);
nand U1842 (N_1842,In_950,In_4983);
or U1843 (N_1843,In_251,In_3477);
xnor U1844 (N_1844,In_3012,In_2904);
nand U1845 (N_1845,In_2440,In_2046);
xnor U1846 (N_1846,In_713,In_1764);
and U1847 (N_1847,In_3692,In_3270);
xnor U1848 (N_1848,In_135,In_4210);
nor U1849 (N_1849,In_3068,In_2835);
nand U1850 (N_1850,In_3559,In_4190);
and U1851 (N_1851,In_3365,In_648);
and U1852 (N_1852,In_3171,In_4801);
or U1853 (N_1853,In_1232,In_2689);
nor U1854 (N_1854,In_4271,In_692);
nor U1855 (N_1855,In_4363,In_2973);
and U1856 (N_1856,In_3964,In_3900);
and U1857 (N_1857,In_1163,In_3458);
nand U1858 (N_1858,In_1360,In_152);
or U1859 (N_1859,In_598,In_2302);
nand U1860 (N_1860,In_1258,In_2743);
nor U1861 (N_1861,In_4246,In_4544);
and U1862 (N_1862,In_3547,In_1490);
nand U1863 (N_1863,In_2070,In_4353);
or U1864 (N_1864,In_4737,In_4204);
xnor U1865 (N_1865,In_3810,In_506);
nor U1866 (N_1866,In_2206,In_275);
xnor U1867 (N_1867,In_3833,In_2739);
nand U1868 (N_1868,In_4032,In_3576);
xor U1869 (N_1869,In_280,In_2746);
nand U1870 (N_1870,In_352,In_2827);
nand U1871 (N_1871,In_706,In_3918);
xor U1872 (N_1872,In_3382,In_4095);
or U1873 (N_1873,In_158,In_2618);
or U1874 (N_1874,In_2153,In_3999);
xor U1875 (N_1875,In_4836,In_39);
nor U1876 (N_1876,In_4741,In_1458);
nand U1877 (N_1877,In_2197,In_742);
and U1878 (N_1878,In_956,In_539);
nand U1879 (N_1879,In_1502,In_3673);
and U1880 (N_1880,In_575,In_1692);
xnor U1881 (N_1881,In_458,In_3898);
or U1882 (N_1882,In_885,In_3056);
xnor U1883 (N_1883,In_421,In_4302);
nand U1884 (N_1884,In_4321,In_1210);
and U1885 (N_1885,In_1899,In_4568);
and U1886 (N_1886,In_3277,In_4108);
nor U1887 (N_1887,In_1219,In_4146);
or U1888 (N_1888,In_143,In_974);
nor U1889 (N_1889,In_4574,In_1471);
and U1890 (N_1890,In_1015,In_602);
or U1891 (N_1891,In_4707,In_1634);
or U1892 (N_1892,In_1321,In_4523);
nor U1893 (N_1893,In_3251,In_1148);
nand U1894 (N_1894,In_4296,In_3796);
xor U1895 (N_1895,In_2676,In_1004);
xor U1896 (N_1896,In_2807,In_1732);
or U1897 (N_1897,In_1824,In_157);
and U1898 (N_1898,In_4695,In_2417);
nand U1899 (N_1899,In_1383,In_2996);
or U1900 (N_1900,In_2889,In_1177);
or U1901 (N_1901,In_1449,In_499);
nand U1902 (N_1902,In_1690,In_237);
or U1903 (N_1903,In_3378,In_1985);
xnor U1904 (N_1904,In_145,In_2509);
xnor U1905 (N_1905,In_3362,In_292);
nand U1906 (N_1906,In_2196,In_3679);
xor U1907 (N_1907,In_1736,In_3689);
or U1908 (N_1908,In_4205,In_3992);
xor U1909 (N_1909,In_4028,In_1138);
and U1910 (N_1910,In_2786,In_1879);
or U1911 (N_1911,In_2832,In_245);
nor U1912 (N_1912,In_4007,In_2016);
xor U1913 (N_1913,In_4894,In_1281);
nor U1914 (N_1914,In_3062,In_4184);
and U1915 (N_1915,In_1837,In_4119);
and U1916 (N_1916,In_323,In_4638);
or U1917 (N_1917,In_1772,In_3387);
nand U1918 (N_1918,In_48,In_463);
and U1919 (N_1919,In_4203,In_1425);
nor U1920 (N_1920,In_4452,In_2548);
nand U1921 (N_1921,In_4710,In_3925);
nand U1922 (N_1922,In_556,In_3273);
and U1923 (N_1923,In_4808,In_1330);
xor U1924 (N_1924,In_4150,In_4585);
nand U1925 (N_1925,In_2227,In_830);
nand U1926 (N_1926,In_1956,In_4602);
nor U1927 (N_1927,In_791,In_2871);
nand U1928 (N_1928,In_2190,In_1472);
nand U1929 (N_1929,In_965,In_3969);
xnor U1930 (N_1930,In_3617,In_1327);
or U1931 (N_1931,In_951,In_3089);
xnor U1932 (N_1932,In_3480,In_356);
or U1933 (N_1933,In_686,In_4733);
or U1934 (N_1934,In_886,In_1781);
or U1935 (N_1935,In_4266,In_2646);
nor U1936 (N_1936,In_4428,In_298);
xnor U1937 (N_1937,In_4874,In_3570);
nor U1938 (N_1938,In_2559,In_1319);
or U1939 (N_1939,In_1825,In_1629);
nor U1940 (N_1940,In_2837,In_667);
or U1941 (N_1941,In_428,In_4590);
nand U1942 (N_1942,In_4972,In_3720);
nor U1943 (N_1943,In_2593,In_2380);
nor U1944 (N_1944,In_255,In_1146);
nor U1945 (N_1945,In_177,In_4562);
nor U1946 (N_1946,In_471,In_1617);
xor U1947 (N_1947,In_3765,In_1727);
xnor U1948 (N_1948,In_2122,In_627);
nand U1949 (N_1949,In_2138,In_2075);
xnor U1950 (N_1950,In_3890,In_4316);
nand U1951 (N_1951,In_4637,In_2412);
nor U1952 (N_1952,In_653,In_3840);
and U1953 (N_1953,In_2967,In_3838);
and U1954 (N_1954,In_304,In_2524);
nor U1955 (N_1955,In_4796,In_641);
and U1956 (N_1956,In_460,In_4487);
nor U1957 (N_1957,In_4830,In_1243);
nand U1958 (N_1958,In_1276,In_1568);
nor U1959 (N_1959,In_72,In_2124);
xnor U1960 (N_1960,In_4248,In_2637);
and U1961 (N_1961,In_4708,In_4899);
nand U1962 (N_1962,In_3042,In_4738);
xnor U1963 (N_1963,In_1390,In_776);
xnor U1964 (N_1964,In_4825,In_2023);
nand U1965 (N_1965,In_1088,In_967);
nor U1966 (N_1966,In_4165,In_2438);
nor U1967 (N_1967,In_2838,In_695);
and U1968 (N_1968,In_2594,In_2565);
nor U1969 (N_1969,In_896,In_3099);
or U1970 (N_1970,In_4811,In_2790);
xor U1971 (N_1971,In_4736,In_2923);
or U1972 (N_1972,In_4681,In_1480);
xor U1973 (N_1973,In_2422,In_1387);
nand U1974 (N_1974,In_448,In_25);
nand U1975 (N_1975,In_1768,In_4712);
and U1976 (N_1976,In_3026,In_160);
and U1977 (N_1977,In_3967,In_1735);
or U1978 (N_1978,In_1523,In_2537);
xor U1979 (N_1979,In_2805,In_4370);
nand U1980 (N_1980,In_2737,In_4818);
or U1981 (N_1981,In_1503,In_923);
xnor U1982 (N_1982,In_78,In_2960);
nor U1983 (N_1983,In_1461,In_2707);
and U1984 (N_1984,In_3813,In_4491);
and U1985 (N_1985,In_4035,In_3272);
nor U1986 (N_1986,In_3790,In_2263);
and U1987 (N_1987,In_4994,In_2970);
nor U1988 (N_1988,In_4619,In_524);
or U1989 (N_1989,In_2708,In_396);
or U1990 (N_1990,In_4653,In_3488);
or U1991 (N_1991,In_2664,In_903);
nor U1992 (N_1992,In_3359,In_2170);
nand U1993 (N_1993,In_493,In_366);
xor U1994 (N_1994,In_519,In_839);
and U1995 (N_1995,In_2498,In_1316);
nand U1996 (N_1996,In_2920,In_175);
xnor U1997 (N_1997,In_4705,In_3807);
nand U1998 (N_1998,In_2343,In_3398);
nor U1999 (N_1999,In_4453,In_3304);
nor U2000 (N_2000,In_3159,In_49);
nand U2001 (N_2001,In_4537,In_3801);
xnor U2002 (N_2002,In_4076,In_2094);
xor U2003 (N_2003,In_3418,In_4584);
and U2004 (N_2004,In_1904,In_1266);
nor U2005 (N_2005,In_4418,In_743);
or U2006 (N_2006,In_4123,In_2988);
or U2007 (N_2007,In_3166,In_669);
or U2008 (N_2008,In_4086,In_617);
nor U2009 (N_2009,In_795,In_1160);
or U2010 (N_2010,In_725,In_4060);
and U2011 (N_2011,In_3390,In_2787);
xor U2012 (N_2012,In_4996,In_3215);
nand U2013 (N_2013,In_4599,In_2640);
xor U2014 (N_2014,In_2169,In_4129);
nor U2015 (N_2015,In_4471,In_2693);
xor U2016 (N_2016,In_840,In_469);
nand U2017 (N_2017,In_1314,In_4628);
or U2018 (N_2018,In_74,In_220);
nand U2019 (N_2019,In_4153,In_2972);
nand U2020 (N_2020,In_46,In_1298);
xor U2021 (N_2021,In_3571,In_1757);
and U2022 (N_2022,In_2321,In_986);
nand U2023 (N_2023,In_768,In_1065);
or U2024 (N_2024,In_1916,In_4336);
nor U2025 (N_2025,In_55,In_1150);
nor U2026 (N_2026,In_2955,In_1475);
or U2027 (N_2027,In_3061,In_1181);
nand U2028 (N_2028,In_871,In_3127);
or U2029 (N_2029,In_4289,In_870);
and U2030 (N_2030,In_1812,In_3134);
xor U2031 (N_2031,In_4877,In_3622);
or U2032 (N_2032,In_982,In_1143);
nor U2033 (N_2033,In_282,In_97);
nand U2034 (N_2034,In_2545,In_4812);
nand U2035 (N_2035,In_3474,In_1224);
nand U2036 (N_2036,In_1584,In_1774);
nor U2037 (N_2037,In_4971,In_1687);
or U2038 (N_2038,In_2497,In_3809);
or U2039 (N_2039,In_2948,In_434);
nor U2040 (N_2040,In_2834,In_3653);
or U2041 (N_2041,In_2218,In_4820);
or U2042 (N_2042,In_4759,In_3795);
nor U2043 (N_2043,In_957,In_978);
or U2044 (N_2044,In_306,In_454);
xnor U2045 (N_2045,In_195,In_3201);
nand U2046 (N_2046,In_1445,In_26);
xor U2047 (N_2047,In_1591,In_307);
xnor U2048 (N_2048,In_3090,In_1187);
nand U2049 (N_2049,In_1701,In_1710);
and U2050 (N_2050,In_238,In_3531);
or U2051 (N_2051,In_510,In_205);
nand U2052 (N_2052,In_384,In_90);
nor U2053 (N_2053,In_3002,In_3200);
nand U2054 (N_2054,In_3500,In_273);
and U2055 (N_2055,In_2287,In_3651);
or U2056 (N_2056,In_2615,In_972);
and U2057 (N_2057,In_3637,In_77);
nand U2058 (N_2058,In_2192,In_4144);
or U2059 (N_2059,In_1452,In_3745);
xnor U2060 (N_2060,In_4415,In_970);
and U2061 (N_2061,In_1548,In_4967);
nor U2062 (N_2062,In_2285,In_2890);
and U2063 (N_2063,In_399,In_85);
nor U2064 (N_2064,In_4629,In_4124);
xor U2065 (N_2065,In_2128,In_856);
or U2066 (N_2066,In_4444,In_3271);
and U2067 (N_2067,In_3331,In_334);
and U2068 (N_2068,In_2472,In_3084);
or U2069 (N_2069,In_2295,In_4447);
or U2070 (N_2070,In_1464,In_794);
and U2071 (N_2071,In_3721,In_2583);
nand U2072 (N_2072,In_4909,In_3055);
nand U2073 (N_2073,In_4104,In_254);
nand U2074 (N_2074,In_4564,In_3054);
and U2075 (N_2075,In_2873,In_1638);
nand U2076 (N_2076,In_1924,In_1877);
nand U2077 (N_2077,In_4673,In_3993);
xnor U2078 (N_2078,In_3514,In_4004);
nand U2079 (N_2079,In_2191,In_3220);
and U2080 (N_2080,In_63,In_989);
nand U2081 (N_2081,In_2031,In_1640);
or U2082 (N_2082,In_557,In_475);
nor U2083 (N_2083,In_3329,In_681);
nor U2084 (N_2084,In_2060,In_2700);
and U2085 (N_2085,In_720,In_1679);
or U2086 (N_2086,In_2091,In_2397);
nor U2087 (N_2087,In_1159,In_829);
nand U2088 (N_2088,In_1868,In_1011);
or U2089 (N_2089,In_4517,In_1212);
and U2090 (N_2090,In_313,In_1754);
nand U2091 (N_2091,In_1125,In_2740);
and U2092 (N_2092,In_920,In_4099);
nor U2093 (N_2093,In_1129,In_2083);
xnor U2094 (N_2094,In_1097,In_3715);
nand U2095 (N_2095,In_2398,In_4461);
xor U2096 (N_2096,In_864,In_2215);
nand U2097 (N_2097,In_1308,In_4309);
and U2098 (N_2098,In_4424,In_4306);
and U2099 (N_2099,In_516,In_2769);
or U2100 (N_2100,In_502,In_3349);
or U2101 (N_2101,In_4328,In_1201);
or U2102 (N_2102,In_825,In_3453);
or U2103 (N_2103,In_3861,In_3296);
or U2104 (N_2104,In_3517,In_1653);
xor U2105 (N_2105,In_2120,In_3770);
nand U2106 (N_2106,In_1905,In_2587);
nor U2107 (N_2107,In_976,In_2275);
nand U2108 (N_2108,In_2068,In_4411);
and U2109 (N_2109,In_1815,In_1706);
or U2110 (N_2110,In_1431,In_3845);
or U2111 (N_2111,In_1374,In_3439);
or U2112 (N_2112,In_4200,In_4872);
nand U2113 (N_2113,In_3618,In_1974);
or U2114 (N_2114,In_414,In_1300);
nand U2115 (N_2115,In_140,In_3232);
nand U2116 (N_2116,In_919,In_3415);
nor U2117 (N_2117,In_2389,In_3945);
xor U2118 (N_2118,In_977,In_1405);
nor U2119 (N_2119,In_4546,In_4548);
nor U2120 (N_2120,In_3491,In_3830);
nand U2121 (N_2121,In_4932,In_3499);
and U2122 (N_2122,In_2269,In_2180);
xnor U2123 (N_2123,In_3966,In_1170);
or U2124 (N_2124,In_2716,In_2544);
xnor U2125 (N_2125,In_4212,In_2181);
nor U2126 (N_2126,In_1356,In_3078);
xor U2127 (N_2127,In_1814,In_3073);
xor U2128 (N_2128,In_3348,In_1560);
and U2129 (N_2129,In_3785,In_3497);
nand U2130 (N_2130,In_1226,In_4456);
xnor U2131 (N_2131,In_2513,In_786);
and U2132 (N_2132,In_3305,In_3117);
xor U2133 (N_2133,In_2344,In_2008);
nor U2134 (N_2134,In_1891,In_761);
and U2135 (N_2135,In_2446,In_595);
nand U2136 (N_2136,In_4431,In_4275);
or U2137 (N_2137,In_3740,In_2308);
nor U2138 (N_2138,In_4170,In_851);
and U2139 (N_2139,In_2543,In_3341);
or U2140 (N_2140,In_2995,In_3700);
and U2141 (N_2141,In_2240,In_3729);
or U2142 (N_2142,In_4938,In_377);
xnor U2143 (N_2143,In_1746,In_390);
or U2144 (N_2144,In_4307,In_1981);
and U2145 (N_2145,In_3672,In_2073);
xnor U2146 (N_2146,In_4090,In_3153);
nor U2147 (N_2147,In_2985,In_154);
nand U2148 (N_2148,In_1976,In_2419);
nand U2149 (N_2149,In_2258,In_2503);
xor U2150 (N_2150,In_3937,In_2870);
nand U2151 (N_2151,In_1421,In_4255);
and U2152 (N_2152,In_2456,In_120);
nor U2153 (N_2153,In_3238,In_554);
xnor U2154 (N_2154,In_253,In_3065);
nor U2155 (N_2155,In_1032,In_1407);
nor U2156 (N_2156,In_3182,In_4472);
nor U2157 (N_2157,In_2050,In_2978);
xnor U2158 (N_2158,In_1323,In_3839);
or U2159 (N_2159,In_2666,In_299);
nor U2160 (N_2160,In_2819,In_4856);
nor U2161 (N_2161,In_4978,In_4784);
nor U2162 (N_2162,In_1010,In_1969);
and U2163 (N_2163,In_726,In_2742);
xor U2164 (N_2164,In_222,In_3425);
nor U2165 (N_2165,In_4078,In_4270);
or U2166 (N_2166,In_3996,In_111);
xnor U2167 (N_2167,In_1095,In_2997);
and U2168 (N_2168,In_638,In_4335);
nand U2169 (N_2169,In_571,In_2149);
nor U2170 (N_2170,In_4730,In_427);
and U2171 (N_2171,In_3001,In_2069);
nor U2172 (N_2172,In_1832,In_969);
nand U2173 (N_2173,In_2767,In_1694);
or U2174 (N_2174,In_291,In_2475);
and U2175 (N_2175,In_2358,In_263);
nor U2176 (N_2176,In_1058,In_2044);
or U2177 (N_2177,In_2089,In_4604);
or U2178 (N_2178,In_2480,In_4777);
and U2179 (N_2179,In_4304,In_6);
or U2180 (N_2180,In_4906,In_4178);
nor U2181 (N_2181,In_1719,In_2061);
nand U2182 (N_2182,In_1793,In_2535);
nand U2183 (N_2183,In_4679,In_984);
nor U2184 (N_2184,In_4014,In_1897);
or U2185 (N_2185,In_1919,In_3784);
and U2186 (N_2186,In_917,In_762);
xor U2187 (N_2187,In_1414,In_2580);
nand U2188 (N_2188,In_4339,In_4709);
or U2189 (N_2189,In_548,In_309);
xnor U2190 (N_2190,In_877,In_2915);
and U2191 (N_2191,In_91,In_1624);
and U2192 (N_2192,In_1200,In_3887);
xnor U2193 (N_2193,In_3776,In_379);
or U2194 (N_2194,In_2145,In_3364);
nand U2195 (N_2195,In_1147,In_4926);
or U2196 (N_2196,In_2045,In_1485);
nand U2197 (N_2197,In_1778,In_1659);
or U2198 (N_2198,In_118,In_468);
or U2199 (N_2199,In_4068,In_165);
xnor U2200 (N_2200,In_93,In_3669);
xnor U2201 (N_2201,In_114,In_252);
xnor U2202 (N_2202,In_2671,In_1539);
and U2203 (N_2203,In_2844,In_2627);
nor U2204 (N_2204,In_2387,In_1017);
xnor U2205 (N_2205,In_1575,In_723);
xor U2206 (N_2206,In_82,In_3916);
xor U2207 (N_2207,In_1910,In_2178);
nor U2208 (N_2208,In_213,In_898);
nand U2209 (N_2209,In_566,In_1783);
or U2210 (N_2210,In_490,In_4186);
and U2211 (N_2211,In_915,In_1454);
or U2212 (N_2212,In_3256,In_4831);
and U2213 (N_2213,In_3152,In_751);
nor U2214 (N_2214,In_2783,In_1328);
nor U2215 (N_2215,In_2773,In_348);
nor U2216 (N_2216,In_2104,In_3045);
and U2217 (N_2217,In_394,In_3983);
and U2218 (N_2218,In_2927,In_597);
and U2219 (N_2219,In_4793,In_4841);
and U2220 (N_2220,In_3697,In_2653);
nand U2221 (N_2221,In_559,In_1608);
or U2222 (N_2222,In_2928,In_2989);
or U2223 (N_2223,In_451,In_3774);
nand U2224 (N_2224,In_1108,In_924);
or U2225 (N_2225,In_2909,In_2974);
or U2226 (N_2226,In_150,In_4871);
or U2227 (N_2227,In_4356,In_1784);
or U2228 (N_2228,In_431,In_3131);
nand U2229 (N_2229,In_2893,In_1864);
xor U2230 (N_2230,In_4873,In_1761);
or U2231 (N_2231,In_1914,In_192);
nand U2232 (N_2232,In_1029,In_3881);
nand U2233 (N_2233,In_3036,In_405);
xor U2234 (N_2234,In_2937,In_4858);
or U2235 (N_2235,In_3958,In_2938);
and U2236 (N_2236,In_929,In_1069);
nor U2237 (N_2237,In_2347,In_1972);
or U2238 (N_2238,In_3757,In_1459);
and U2239 (N_2239,In_1001,In_3437);
nand U2240 (N_2240,In_4109,In_179);
nand U2241 (N_2241,In_3388,In_4397);
xnor U2242 (N_2242,In_2858,In_2656);
or U2243 (N_2243,In_1377,In_1416);
or U2244 (N_2244,In_4624,In_1111);
nor U2245 (N_2245,In_4847,In_4410);
or U2246 (N_2246,In_2842,In_2166);
nand U2247 (N_2247,In_569,In_1267);
nor U2248 (N_2248,In_789,In_362);
nor U2249 (N_2249,In_206,In_1340);
or U2250 (N_2250,In_4503,In_1466);
and U2251 (N_2251,In_3974,In_2345);
xor U2252 (N_2252,In_2526,In_649);
nor U2253 (N_2253,In_632,In_4048);
nand U2254 (N_2254,In_4939,In_3345);
nand U2255 (N_2255,In_625,In_4241);
xnor U2256 (N_2256,In_209,In_1676);
nor U2257 (N_2257,In_3242,In_4505);
nor U2258 (N_2258,In_714,In_4228);
xor U2259 (N_2259,In_3856,In_3490);
nor U2260 (N_2260,In_87,In_2578);
nand U2261 (N_2261,In_3112,In_172);
or U2262 (N_2262,In_3512,In_295);
or U2263 (N_2263,In_560,In_2789);
nor U2264 (N_2264,In_4384,In_3294);
xor U2265 (N_2265,In_1755,In_4764);
and U2266 (N_2266,In_1718,In_264);
and U2267 (N_2267,In_271,In_319);
and U2268 (N_2268,In_809,In_2372);
or U2269 (N_2269,In_521,In_3315);
or U2270 (N_2270,In_2958,In_3168);
or U2271 (N_2271,In_2434,In_1886);
nor U2272 (N_2272,In_3316,In_337);
or U2273 (N_2273,In_1487,In_2603);
and U2274 (N_2274,In_4280,In_3698);
nor U2275 (N_2275,In_4337,In_1934);
and U2276 (N_2276,In_4285,In_2423);
or U2277 (N_2277,In_2198,In_3608);
nand U2278 (N_2278,In_494,In_4701);
and U2279 (N_2279,In_2809,In_98);
nand U2280 (N_2280,In_2736,In_3230);
nand U2281 (N_2281,In_4860,In_1616);
nor U2282 (N_2282,In_1221,In_4572);
nand U2283 (N_2283,In_2107,In_1262);
xnor U2284 (N_2284,In_3255,In_1332);
or U2285 (N_2285,In_2622,In_1898);
and U2286 (N_2286,In_1611,In_2520);
and U2287 (N_2287,In_4386,In_1808);
and U2288 (N_2288,In_2267,In_3483);
xor U2289 (N_2289,In_4282,In_696);
nand U2290 (N_2290,In_922,In_4331);
nand U2291 (N_2291,In_2758,In_121);
nor U2292 (N_2292,In_204,In_2310);
or U2293 (N_2293,In_1903,In_1544);
xor U2294 (N_2294,In_3738,In_4313);
xor U2295 (N_2295,In_1434,In_558);
xnor U2296 (N_2296,In_3283,In_4185);
nor U2297 (N_2297,In_1353,In_3229);
or U2298 (N_2298,In_3621,In_2981);
or U2299 (N_2299,In_1297,In_3154);
nand U2300 (N_2300,In_1980,In_4842);
xor U2301 (N_2301,In_2628,In_3886);
nand U2302 (N_2302,In_1883,In_860);
xor U2303 (N_2303,In_3684,In_2711);
or U2304 (N_2304,In_3310,In_1403);
and U2305 (N_2305,In_4580,In_2887);
nand U2306 (N_2306,In_4844,In_1291);
or U2307 (N_2307,In_1870,In_2202);
and U2308 (N_2308,In_4177,In_4554);
and U2309 (N_2309,In_3528,In_2430);
nand U2310 (N_2310,In_2112,In_2463);
nor U2311 (N_2311,In_1531,In_616);
nand U2312 (N_2312,In_3188,In_2451);
or U2313 (N_2313,In_4100,In_92);
or U2314 (N_2314,In_2940,In_1780);
nor U2315 (N_2315,In_4851,In_4581);
or U2316 (N_2316,In_4074,In_592);
or U2317 (N_2317,In_2612,In_4999);
nand U2318 (N_2318,In_2511,In_1871);
and U2319 (N_2319,In_3931,In_1117);
xor U2320 (N_2320,In_4070,In_501);
xor U2321 (N_2321,In_1023,In_813);
xnor U2322 (N_2322,In_3299,In_537);
or U2323 (N_2323,In_4483,In_1455);
xnor U2324 (N_2324,In_2346,In_2126);
nor U2325 (N_2325,In_4804,In_1453);
or U2326 (N_2326,In_2015,In_3427);
or U2327 (N_2327,In_430,In_1581);
and U2328 (N_2328,In_3855,In_1322);
xor U2329 (N_2329,In_3145,In_1527);
nor U2330 (N_2330,In_1075,In_324);
nor U2331 (N_2331,In_1637,In_2386);
xor U2332 (N_2332,In_3836,In_640);
nor U2333 (N_2333,In_3141,In_3748);
nand U2334 (N_2334,In_370,In_311);
or U2335 (N_2335,In_2244,In_4058);
nor U2336 (N_2336,In_3741,In_1047);
nand U2337 (N_2337,In_2542,In_3246);
xnor U2338 (N_2338,In_3252,In_1098);
or U2339 (N_2339,In_3069,In_3884);
and U2340 (N_2340,In_4946,In_16);
nor U2341 (N_2341,In_1182,In_429);
nor U2342 (N_2342,In_2782,In_3101);
xnor U2343 (N_2343,In_4062,In_2907);
nand U2344 (N_2344,In_4749,In_1411);
or U2345 (N_2345,In_422,In_3549);
xor U2346 (N_2346,In_2305,In_303);
xnor U2347 (N_2347,In_2802,In_660);
xnor U2348 (N_2348,In_788,In_3164);
nor U2349 (N_2349,In_3852,In_3120);
nor U2350 (N_2350,In_4506,In_4661);
xnor U2351 (N_2351,In_1229,In_3513);
nand U2352 (N_2352,In_2760,In_4538);
xnor U2353 (N_2353,In_4898,In_4446);
nor U2354 (N_2354,In_2551,In_1193);
xnor U2355 (N_2355,In_4258,In_1952);
or U2356 (N_2356,In_1073,In_3896);
nand U2357 (N_2357,In_3116,In_4886);
and U2358 (N_2358,In_105,In_1829);
nand U2359 (N_2359,In_1593,In_1396);
and U2360 (N_2360,In_4767,In_3654);
or U2361 (N_2361,In_4214,In_804);
or U2362 (N_2362,In_849,In_3438);
xnor U2363 (N_2363,In_4250,In_3236);
xnor U2364 (N_2364,In_961,In_4216);
nor U2365 (N_2365,In_4989,In_3902);
nor U2366 (N_2366,In_3656,In_1412);
and U2367 (N_2367,In_1521,In_1491);
or U2368 (N_2368,In_4689,In_1155);
nand U2369 (N_2369,In_2478,In_3102);
xor U2370 (N_2370,In_4848,In_3023);
and U2371 (N_2371,In_3169,In_1418);
or U2372 (N_2372,In_2336,In_2298);
nor U2373 (N_2373,In_4609,In_4043);
nand U2374 (N_2374,In_130,In_515);
or U2375 (N_2375,In_2282,In_425);
nor U2376 (N_2376,In_3658,In_225);
and U2377 (N_2377,In_4044,In_117);
or U2378 (N_2378,In_3432,In_3290);
nor U2379 (N_2379,In_3473,In_2273);
xor U2380 (N_2380,In_999,In_4451);
and U2381 (N_2381,In_848,In_550);
and U2382 (N_2382,In_1978,In_2505);
nor U2383 (N_2383,In_1522,In_535);
nor U2384 (N_2384,In_2470,In_4595);
xnor U2385 (N_2385,In_3057,In_4355);
and U2386 (N_2386,In_3286,In_2051);
or U2387 (N_2387,In_3546,In_3352);
or U2388 (N_2388,In_3610,In_4719);
xor U2389 (N_2389,In_3524,In_2781);
and U2390 (N_2390,In_1183,In_2062);
nand U2391 (N_2391,In_666,In_4982);
or U2392 (N_2392,In_149,In_1494);
and U2393 (N_2393,In_1102,In_2999);
xor U2394 (N_2394,In_426,In_1479);
nor U2395 (N_2395,In_4276,In_4752);
and U2396 (N_2396,In_3053,In_4743);
or U2397 (N_2397,In_2453,In_1235);
xnor U2398 (N_2398,In_2536,In_3155);
or U2399 (N_2399,In_799,In_996);
and U2400 (N_2400,In_3379,In_3118);
xor U2401 (N_2401,In_4189,In_1776);
xor U2402 (N_2402,In_2814,In_718);
xnor U2403 (N_2403,In_3557,In_456);
nand U2404 (N_2404,In_2550,In_3734);
xor U2405 (N_2405,In_4476,In_3343);
nor U2406 (N_2406,In_3643,In_4691);
nand U2407 (N_2407,In_3664,In_1101);
and U2408 (N_2408,In_3596,In_450);
or U2409 (N_2409,In_4756,In_1335);
and U2410 (N_2410,In_1365,In_4312);
nand U2411 (N_2411,In_3080,In_2441);
nor U2412 (N_2412,In_4533,In_3321);
nand U2413 (N_2413,In_3410,In_2420);
xnor U2414 (N_2414,In_2039,In_147);
nand U2415 (N_2415,In_1989,In_581);
or U2416 (N_2416,In_3493,In_1587);
or U2417 (N_2417,In_1255,In_4504);
and U2418 (N_2418,In_3174,In_2204);
nand U2419 (N_2419,In_2735,In_2733);
nand U2420 (N_2420,In_2110,In_4611);
nor U2421 (N_2421,In_3950,In_2271);
nor U2422 (N_2422,In_1817,In_296);
nor U2423 (N_2423,In_580,In_2222);
nor U2424 (N_2424,In_30,In_737);
and U2425 (N_2425,In_3351,In_1105);
xor U2426 (N_2426,In_861,In_3556);
nor U2427 (N_2427,In_948,In_1135);
or U2428 (N_2428,In_4717,In_162);
or U2429 (N_2429,In_4440,In_2705);
and U2430 (N_2430,In_4371,In_783);
xnor U2431 (N_2431,In_2491,In_1997);
nor U2432 (N_2432,In_3172,In_2431);
nor U2433 (N_2433,In_3938,In_178);
xor U2434 (N_2434,In_3475,In_4693);
nor U2435 (N_2435,In_3553,In_4091);
or U2436 (N_2436,In_4732,In_4351);
or U2437 (N_2437,In_141,In_2818);
nand U2438 (N_2438,In_181,In_2547);
nand U2439 (N_2439,In_3346,In_4988);
and U2440 (N_2440,In_310,In_449);
nand U2441 (N_2441,In_2721,In_4098);
nand U2442 (N_2442,In_3254,In_1662);
and U2443 (N_2443,In_508,In_4173);
nand U2444 (N_2444,In_1529,In_2649);
and U2445 (N_2445,In_2232,In_2217);
or U2446 (N_2446,In_3266,In_127);
or U2447 (N_2447,In_2266,In_2261);
nor U2448 (N_2448,In_3939,In_1633);
nand U2449 (N_2449,In_3312,In_3842);
xnor U2450 (N_2450,In_1188,In_1054);
and U2451 (N_2451,In_2659,In_2246);
and U2452 (N_2452,In_3817,In_3082);
nor U2453 (N_2453,In_359,In_459);
and U2454 (N_2454,In_3297,In_685);
or U2455 (N_2455,In_3249,In_985);
or U2456 (N_2456,In_1400,In_4645);
xnor U2457 (N_2457,In_4050,In_168);
nand U2458 (N_2458,In_909,In_4002);
or U2459 (N_2459,In_846,In_491);
xor U2460 (N_2460,In_3930,In_3914);
and U2461 (N_2461,In_4507,In_1705);
or U2462 (N_2462,In_8,In_3870);
and U2463 (N_2463,In_3904,In_3088);
or U2464 (N_2464,In_3311,In_3910);
nand U2465 (N_2465,In_4556,In_4211);
or U2466 (N_2466,In_4433,In_2706);
and U2467 (N_2467,In_2755,In_2477);
nand U2468 (N_2468,In_3585,In_4107);
xnor U2469 (N_2469,In_467,In_2859);
and U2470 (N_2470,In_2770,In_4636);
nor U2471 (N_2471,In_1404,In_3536);
nor U2472 (N_2472,In_1739,In_2619);
nor U2473 (N_2473,In_443,In_4575);
and U2474 (N_2474,In_615,In_1202);
and U2475 (N_2475,In_4238,In_3194);
xor U2476 (N_2476,In_4516,In_101);
and U2477 (N_2477,In_208,In_4790);
nor U2478 (N_2478,In_2764,In_3772);
nand U2479 (N_2479,In_4713,In_4023);
nor U2480 (N_2480,In_3826,In_4508);
nor U2481 (N_2481,In_2762,In_4439);
xnor U2482 (N_2482,In_277,In_4175);
or U2483 (N_2483,In_1052,In_2754);
xor U2484 (N_2484,In_4139,In_446);
and U2485 (N_2485,In_278,In_2406);
xor U2486 (N_2486,In_2054,In_897);
and U2487 (N_2487,In_612,In_1993);
nor U2488 (N_2488,In_2766,In_1798);
nand U2489 (N_2489,In_4416,In_1935);
xor U2490 (N_2490,In_4130,In_3822);
nor U2491 (N_2491,In_3927,In_3739);
xor U2492 (N_2492,In_1722,In_3446);
nor U2493 (N_2493,In_2936,In_2820);
nand U2494 (N_2494,In_4403,In_712);
and U2495 (N_2495,In_3106,In_736);
xnor U2496 (N_2496,In_3077,In_2484);
nand U2497 (N_2497,In_4151,In_385);
and U2498 (N_2498,In_802,In_1984);
nand U2499 (N_2499,In_536,In_2900);
nor U2500 (N_2500,In_1359,In_1278);
nor U2501 (N_2501,In_3848,In_3139);
nor U2502 (N_2502,In_3528,In_4811);
nand U2503 (N_2503,In_2919,In_4305);
nor U2504 (N_2504,In_1233,In_3707);
nand U2505 (N_2505,In_4188,In_4779);
nor U2506 (N_2506,In_2836,In_4869);
and U2507 (N_2507,In_1425,In_245);
nor U2508 (N_2508,In_717,In_4822);
and U2509 (N_2509,In_3122,In_2196);
xnor U2510 (N_2510,In_4058,In_2952);
or U2511 (N_2511,In_2765,In_1765);
nor U2512 (N_2512,In_1158,In_2121);
and U2513 (N_2513,In_2551,In_1864);
or U2514 (N_2514,In_1810,In_240);
and U2515 (N_2515,In_4323,In_1834);
nor U2516 (N_2516,In_3313,In_490);
nor U2517 (N_2517,In_2783,In_4913);
and U2518 (N_2518,In_2025,In_2983);
xor U2519 (N_2519,In_2413,In_3553);
and U2520 (N_2520,In_2172,In_4605);
nand U2521 (N_2521,In_580,In_1505);
or U2522 (N_2522,In_4648,In_1122);
nand U2523 (N_2523,In_3144,In_3154);
or U2524 (N_2524,In_2512,In_4278);
xnor U2525 (N_2525,In_4975,In_3103);
nor U2526 (N_2526,In_2972,In_1605);
nor U2527 (N_2527,In_569,In_4231);
nor U2528 (N_2528,In_917,In_1211);
and U2529 (N_2529,In_593,In_1907);
or U2530 (N_2530,In_2505,In_1114);
nand U2531 (N_2531,In_2807,In_2239);
nand U2532 (N_2532,In_1189,In_1623);
and U2533 (N_2533,In_4220,In_3558);
nand U2534 (N_2534,In_1762,In_636);
nand U2535 (N_2535,In_1683,In_4702);
nand U2536 (N_2536,In_3215,In_1828);
nor U2537 (N_2537,In_749,In_541);
nor U2538 (N_2538,In_2353,In_4458);
nor U2539 (N_2539,In_592,In_858);
or U2540 (N_2540,In_1205,In_1368);
nand U2541 (N_2541,In_2205,In_4218);
nor U2542 (N_2542,In_3245,In_3976);
and U2543 (N_2543,In_918,In_2811);
or U2544 (N_2544,In_4814,In_30);
and U2545 (N_2545,In_1721,In_1694);
nor U2546 (N_2546,In_3276,In_249);
and U2547 (N_2547,In_4326,In_2618);
and U2548 (N_2548,In_4031,In_1652);
or U2549 (N_2549,In_3252,In_4992);
nand U2550 (N_2550,In_645,In_1135);
nor U2551 (N_2551,In_3562,In_2676);
nand U2552 (N_2552,In_4293,In_97);
or U2553 (N_2553,In_3019,In_104);
nor U2554 (N_2554,In_1221,In_1860);
and U2555 (N_2555,In_4492,In_3311);
or U2556 (N_2556,In_4871,In_2573);
xor U2557 (N_2557,In_3429,In_712);
or U2558 (N_2558,In_4691,In_2820);
xor U2559 (N_2559,In_3163,In_895);
xor U2560 (N_2560,In_3761,In_825);
xnor U2561 (N_2561,In_1539,In_2187);
nor U2562 (N_2562,In_1700,In_3690);
and U2563 (N_2563,In_499,In_4799);
nand U2564 (N_2564,In_3446,In_245);
and U2565 (N_2565,In_1344,In_30);
and U2566 (N_2566,In_4749,In_3189);
and U2567 (N_2567,In_1422,In_4038);
and U2568 (N_2568,In_4297,In_1274);
and U2569 (N_2569,In_2739,In_752);
nor U2570 (N_2570,In_1115,In_170);
or U2571 (N_2571,In_11,In_2590);
or U2572 (N_2572,In_2273,In_4812);
nand U2573 (N_2573,In_1753,In_3033);
xor U2574 (N_2574,In_893,In_509);
xnor U2575 (N_2575,In_3909,In_340);
nand U2576 (N_2576,In_3370,In_405);
nand U2577 (N_2577,In_2558,In_1163);
or U2578 (N_2578,In_450,In_3763);
and U2579 (N_2579,In_4503,In_3592);
and U2580 (N_2580,In_369,In_519);
nor U2581 (N_2581,In_48,In_459);
nor U2582 (N_2582,In_4096,In_2504);
nor U2583 (N_2583,In_3817,In_2360);
nand U2584 (N_2584,In_4174,In_730);
xnor U2585 (N_2585,In_3388,In_3406);
nor U2586 (N_2586,In_3249,In_4500);
nor U2587 (N_2587,In_2617,In_1864);
nand U2588 (N_2588,In_2859,In_2730);
nor U2589 (N_2589,In_3443,In_871);
nor U2590 (N_2590,In_4450,In_760);
xnor U2591 (N_2591,In_3727,In_3149);
nor U2592 (N_2592,In_2300,In_3737);
and U2593 (N_2593,In_2379,In_1854);
xor U2594 (N_2594,In_1392,In_600);
or U2595 (N_2595,In_4134,In_3287);
nor U2596 (N_2596,In_920,In_4653);
xor U2597 (N_2597,In_1510,In_3698);
xnor U2598 (N_2598,In_3811,In_2266);
nand U2599 (N_2599,In_208,In_399);
nand U2600 (N_2600,In_1792,In_2427);
nand U2601 (N_2601,In_2531,In_2206);
or U2602 (N_2602,In_2548,In_2697);
or U2603 (N_2603,In_3704,In_1258);
nor U2604 (N_2604,In_1781,In_4012);
nor U2605 (N_2605,In_255,In_1667);
and U2606 (N_2606,In_1191,In_98);
and U2607 (N_2607,In_3493,In_1078);
or U2608 (N_2608,In_4295,In_1934);
nand U2609 (N_2609,In_4286,In_1138);
nor U2610 (N_2610,In_1427,In_3746);
nor U2611 (N_2611,In_4289,In_1181);
xor U2612 (N_2612,In_4633,In_1604);
or U2613 (N_2613,In_3132,In_163);
nor U2614 (N_2614,In_4024,In_3018);
nor U2615 (N_2615,In_2700,In_3413);
nand U2616 (N_2616,In_2684,In_2217);
and U2617 (N_2617,In_3043,In_3911);
nor U2618 (N_2618,In_45,In_4779);
nor U2619 (N_2619,In_2022,In_2175);
xnor U2620 (N_2620,In_3873,In_3150);
or U2621 (N_2621,In_2210,In_2332);
nor U2622 (N_2622,In_3217,In_649);
or U2623 (N_2623,In_604,In_2102);
nor U2624 (N_2624,In_3073,In_4592);
or U2625 (N_2625,In_1134,In_944);
nor U2626 (N_2626,In_3066,In_464);
or U2627 (N_2627,In_3115,In_2598);
nand U2628 (N_2628,In_2949,In_3236);
and U2629 (N_2629,In_3797,In_422);
and U2630 (N_2630,In_1698,In_4192);
xor U2631 (N_2631,In_4173,In_1404);
nand U2632 (N_2632,In_3559,In_2086);
nor U2633 (N_2633,In_3180,In_3779);
or U2634 (N_2634,In_1962,In_857);
nand U2635 (N_2635,In_4998,In_4094);
and U2636 (N_2636,In_2511,In_1860);
or U2637 (N_2637,In_2617,In_3013);
nand U2638 (N_2638,In_2599,In_4749);
nand U2639 (N_2639,In_4298,In_4937);
nor U2640 (N_2640,In_106,In_4050);
or U2641 (N_2641,In_3779,In_3968);
xnor U2642 (N_2642,In_2451,In_2050);
and U2643 (N_2643,In_3542,In_1414);
nor U2644 (N_2644,In_634,In_2615);
nand U2645 (N_2645,In_3767,In_3312);
nand U2646 (N_2646,In_1908,In_368);
and U2647 (N_2647,In_3846,In_586);
or U2648 (N_2648,In_2947,In_4089);
or U2649 (N_2649,In_488,In_1086);
or U2650 (N_2650,In_3575,In_4573);
and U2651 (N_2651,In_4187,In_4457);
nor U2652 (N_2652,In_1081,In_4692);
xor U2653 (N_2653,In_3890,In_375);
nand U2654 (N_2654,In_4341,In_465);
nor U2655 (N_2655,In_1466,In_3124);
and U2656 (N_2656,In_3369,In_40);
nand U2657 (N_2657,In_3189,In_2022);
xnor U2658 (N_2658,In_2977,In_4804);
xor U2659 (N_2659,In_1203,In_611);
nand U2660 (N_2660,In_2925,In_1470);
nor U2661 (N_2661,In_3239,In_3662);
or U2662 (N_2662,In_1238,In_1943);
and U2663 (N_2663,In_1533,In_4796);
xor U2664 (N_2664,In_1495,In_2061);
nor U2665 (N_2665,In_1031,In_2390);
and U2666 (N_2666,In_2341,In_1956);
nand U2667 (N_2667,In_2489,In_915);
and U2668 (N_2668,In_3827,In_804);
or U2669 (N_2669,In_3552,In_3469);
or U2670 (N_2670,In_3733,In_1795);
and U2671 (N_2671,In_391,In_4612);
xnor U2672 (N_2672,In_3090,In_1493);
or U2673 (N_2673,In_4947,In_1493);
or U2674 (N_2674,In_3076,In_4955);
and U2675 (N_2675,In_4893,In_1023);
xor U2676 (N_2676,In_1108,In_3266);
nor U2677 (N_2677,In_3665,In_2833);
or U2678 (N_2678,In_3628,In_3670);
and U2679 (N_2679,In_4043,In_3301);
nand U2680 (N_2680,In_4171,In_4213);
nand U2681 (N_2681,In_790,In_2628);
xnor U2682 (N_2682,In_1714,In_3574);
or U2683 (N_2683,In_566,In_3820);
and U2684 (N_2684,In_3351,In_2111);
or U2685 (N_2685,In_3516,In_4177);
and U2686 (N_2686,In_1952,In_2139);
xnor U2687 (N_2687,In_4639,In_989);
nand U2688 (N_2688,In_1766,In_3895);
nand U2689 (N_2689,In_1091,In_2800);
nand U2690 (N_2690,In_4625,In_4841);
and U2691 (N_2691,In_3164,In_1005);
and U2692 (N_2692,In_1304,In_4698);
nor U2693 (N_2693,In_4353,In_3073);
nand U2694 (N_2694,In_4277,In_589);
nand U2695 (N_2695,In_2481,In_2290);
nor U2696 (N_2696,In_2944,In_292);
nand U2697 (N_2697,In_635,In_250);
xnor U2698 (N_2698,In_4250,In_2681);
xnor U2699 (N_2699,In_4752,In_3411);
or U2700 (N_2700,In_4499,In_3745);
nor U2701 (N_2701,In_4289,In_2704);
nand U2702 (N_2702,In_4177,In_2381);
xnor U2703 (N_2703,In_3432,In_1135);
nor U2704 (N_2704,In_2893,In_3035);
or U2705 (N_2705,In_4305,In_3990);
nand U2706 (N_2706,In_4997,In_397);
and U2707 (N_2707,In_1380,In_3021);
xnor U2708 (N_2708,In_150,In_2042);
nor U2709 (N_2709,In_3767,In_1268);
nand U2710 (N_2710,In_4928,In_1429);
nand U2711 (N_2711,In_2596,In_2046);
nand U2712 (N_2712,In_442,In_3199);
and U2713 (N_2713,In_3372,In_2583);
or U2714 (N_2714,In_3397,In_1824);
and U2715 (N_2715,In_4025,In_3297);
nand U2716 (N_2716,In_1457,In_3961);
and U2717 (N_2717,In_47,In_288);
xor U2718 (N_2718,In_829,In_4678);
and U2719 (N_2719,In_2062,In_4611);
xnor U2720 (N_2720,In_2108,In_3263);
and U2721 (N_2721,In_3393,In_967);
nand U2722 (N_2722,In_3872,In_4749);
or U2723 (N_2723,In_919,In_4514);
and U2724 (N_2724,In_332,In_4841);
nor U2725 (N_2725,In_208,In_2796);
and U2726 (N_2726,In_1745,In_546);
nand U2727 (N_2727,In_4426,In_1857);
nand U2728 (N_2728,In_4626,In_4395);
or U2729 (N_2729,In_1346,In_2738);
nand U2730 (N_2730,In_3059,In_1262);
nand U2731 (N_2731,In_2605,In_4907);
nand U2732 (N_2732,In_854,In_320);
xor U2733 (N_2733,In_2083,In_1488);
and U2734 (N_2734,In_2587,In_43);
nand U2735 (N_2735,In_4194,In_4698);
xor U2736 (N_2736,In_3886,In_4969);
nor U2737 (N_2737,In_2222,In_605);
or U2738 (N_2738,In_1405,In_792);
xnor U2739 (N_2739,In_3677,In_2508);
nor U2740 (N_2740,In_2889,In_1094);
nor U2741 (N_2741,In_2,In_1110);
or U2742 (N_2742,In_2605,In_1319);
and U2743 (N_2743,In_971,In_45);
or U2744 (N_2744,In_948,In_4835);
xor U2745 (N_2745,In_1065,In_4846);
nor U2746 (N_2746,In_4160,In_4148);
or U2747 (N_2747,In_3847,In_941);
xor U2748 (N_2748,In_465,In_3860);
xor U2749 (N_2749,In_3144,In_4947);
and U2750 (N_2750,In_4733,In_1300);
or U2751 (N_2751,In_271,In_176);
xnor U2752 (N_2752,In_2362,In_2544);
nand U2753 (N_2753,In_3135,In_3571);
nand U2754 (N_2754,In_4755,In_3644);
and U2755 (N_2755,In_2261,In_367);
or U2756 (N_2756,In_2125,In_587);
nand U2757 (N_2757,In_4457,In_4568);
nand U2758 (N_2758,In_3959,In_1182);
nor U2759 (N_2759,In_854,In_1504);
xor U2760 (N_2760,In_17,In_3835);
nor U2761 (N_2761,In_2824,In_299);
and U2762 (N_2762,In_3115,In_219);
xnor U2763 (N_2763,In_3477,In_37);
and U2764 (N_2764,In_4584,In_2095);
nand U2765 (N_2765,In_4607,In_1592);
nand U2766 (N_2766,In_1431,In_4930);
nand U2767 (N_2767,In_4469,In_3483);
or U2768 (N_2768,In_2696,In_2708);
xor U2769 (N_2769,In_279,In_1760);
xor U2770 (N_2770,In_3672,In_2721);
or U2771 (N_2771,In_1426,In_604);
and U2772 (N_2772,In_137,In_1726);
and U2773 (N_2773,In_3585,In_2427);
nor U2774 (N_2774,In_994,In_435);
nor U2775 (N_2775,In_1907,In_1820);
nand U2776 (N_2776,In_4516,In_3060);
or U2777 (N_2777,In_3396,In_3459);
nor U2778 (N_2778,In_2387,In_1944);
or U2779 (N_2779,In_202,In_666);
nand U2780 (N_2780,In_803,In_4772);
or U2781 (N_2781,In_2194,In_4956);
xor U2782 (N_2782,In_835,In_3811);
nor U2783 (N_2783,In_2017,In_4455);
and U2784 (N_2784,In_4213,In_4974);
nand U2785 (N_2785,In_611,In_3550);
xnor U2786 (N_2786,In_328,In_4321);
or U2787 (N_2787,In_595,In_1887);
or U2788 (N_2788,In_4966,In_4644);
xor U2789 (N_2789,In_4340,In_421);
nor U2790 (N_2790,In_520,In_4046);
and U2791 (N_2791,In_1725,In_3881);
nand U2792 (N_2792,In_1087,In_367);
nand U2793 (N_2793,In_3971,In_3798);
or U2794 (N_2794,In_2539,In_2795);
or U2795 (N_2795,In_2012,In_3076);
xnor U2796 (N_2796,In_400,In_2207);
nand U2797 (N_2797,In_4927,In_3304);
xnor U2798 (N_2798,In_3959,In_4414);
nor U2799 (N_2799,In_358,In_52);
and U2800 (N_2800,In_1782,In_51);
nand U2801 (N_2801,In_4172,In_3299);
nand U2802 (N_2802,In_3641,In_969);
and U2803 (N_2803,In_1665,In_3073);
nor U2804 (N_2804,In_4418,In_801);
xor U2805 (N_2805,In_4941,In_4323);
nand U2806 (N_2806,In_3887,In_1278);
and U2807 (N_2807,In_250,In_1553);
nand U2808 (N_2808,In_3197,In_3031);
and U2809 (N_2809,In_908,In_4316);
xor U2810 (N_2810,In_2347,In_4209);
and U2811 (N_2811,In_4306,In_4126);
nor U2812 (N_2812,In_1483,In_4863);
nor U2813 (N_2813,In_937,In_2667);
and U2814 (N_2814,In_1538,In_1272);
and U2815 (N_2815,In_1027,In_3426);
nand U2816 (N_2816,In_2667,In_687);
nor U2817 (N_2817,In_616,In_222);
or U2818 (N_2818,In_385,In_1704);
and U2819 (N_2819,In_492,In_2239);
nand U2820 (N_2820,In_2195,In_3480);
xnor U2821 (N_2821,In_1744,In_4619);
nand U2822 (N_2822,In_2923,In_3274);
nand U2823 (N_2823,In_2789,In_1261);
and U2824 (N_2824,In_1884,In_3337);
nand U2825 (N_2825,In_1286,In_482);
nor U2826 (N_2826,In_3644,In_1731);
nor U2827 (N_2827,In_4540,In_2284);
nor U2828 (N_2828,In_2432,In_1954);
xor U2829 (N_2829,In_2751,In_2618);
or U2830 (N_2830,In_541,In_4262);
nand U2831 (N_2831,In_1993,In_1073);
and U2832 (N_2832,In_1815,In_1909);
and U2833 (N_2833,In_2531,In_1897);
and U2834 (N_2834,In_2799,In_758);
nor U2835 (N_2835,In_365,In_754);
nand U2836 (N_2836,In_3467,In_2597);
and U2837 (N_2837,In_355,In_447);
nor U2838 (N_2838,In_836,In_2377);
and U2839 (N_2839,In_1915,In_320);
or U2840 (N_2840,In_676,In_2106);
nor U2841 (N_2841,In_4084,In_1407);
nor U2842 (N_2842,In_2878,In_1785);
nand U2843 (N_2843,In_1969,In_270);
nor U2844 (N_2844,In_1092,In_4153);
and U2845 (N_2845,In_1933,In_828);
or U2846 (N_2846,In_4016,In_3326);
nor U2847 (N_2847,In_4668,In_4989);
nor U2848 (N_2848,In_3905,In_4835);
nand U2849 (N_2849,In_4217,In_158);
and U2850 (N_2850,In_4197,In_2490);
nand U2851 (N_2851,In_3671,In_380);
xor U2852 (N_2852,In_3758,In_1667);
and U2853 (N_2853,In_3554,In_2915);
nor U2854 (N_2854,In_3359,In_4741);
nand U2855 (N_2855,In_2721,In_1557);
nor U2856 (N_2856,In_351,In_3081);
nor U2857 (N_2857,In_3278,In_3988);
xnor U2858 (N_2858,In_4534,In_4940);
and U2859 (N_2859,In_2916,In_135);
or U2860 (N_2860,In_1582,In_4279);
nand U2861 (N_2861,In_419,In_2324);
or U2862 (N_2862,In_176,In_4851);
and U2863 (N_2863,In_3841,In_2657);
and U2864 (N_2864,In_1202,In_2734);
nor U2865 (N_2865,In_3050,In_4691);
nor U2866 (N_2866,In_805,In_2861);
and U2867 (N_2867,In_637,In_1254);
nand U2868 (N_2868,In_2012,In_2097);
or U2869 (N_2869,In_1665,In_4544);
and U2870 (N_2870,In_2472,In_3355);
nand U2871 (N_2871,In_972,In_4458);
nor U2872 (N_2872,In_803,In_2433);
nand U2873 (N_2873,In_4264,In_3215);
or U2874 (N_2874,In_2588,In_2074);
nand U2875 (N_2875,In_3699,In_1237);
xnor U2876 (N_2876,In_3966,In_3913);
nor U2877 (N_2877,In_4899,In_95);
nor U2878 (N_2878,In_2829,In_1334);
nor U2879 (N_2879,In_4705,In_2166);
nand U2880 (N_2880,In_3994,In_3832);
nand U2881 (N_2881,In_1707,In_4441);
or U2882 (N_2882,In_3652,In_2084);
nor U2883 (N_2883,In_1884,In_3358);
or U2884 (N_2884,In_3180,In_3829);
or U2885 (N_2885,In_3417,In_2112);
or U2886 (N_2886,In_1251,In_1770);
and U2887 (N_2887,In_3704,In_4844);
xor U2888 (N_2888,In_4468,In_4751);
nand U2889 (N_2889,In_4660,In_636);
and U2890 (N_2890,In_3276,In_4247);
or U2891 (N_2891,In_794,In_4082);
or U2892 (N_2892,In_3919,In_797);
xor U2893 (N_2893,In_483,In_2051);
nand U2894 (N_2894,In_4508,In_954);
xor U2895 (N_2895,In_2467,In_2621);
nor U2896 (N_2896,In_4526,In_3010);
or U2897 (N_2897,In_1651,In_543);
xnor U2898 (N_2898,In_432,In_4177);
nor U2899 (N_2899,In_3462,In_1991);
and U2900 (N_2900,In_3214,In_4295);
nor U2901 (N_2901,In_3498,In_1180);
nand U2902 (N_2902,In_684,In_3482);
or U2903 (N_2903,In_968,In_1750);
nand U2904 (N_2904,In_691,In_4988);
and U2905 (N_2905,In_4457,In_4031);
nor U2906 (N_2906,In_1907,In_4962);
xnor U2907 (N_2907,In_395,In_2444);
nor U2908 (N_2908,In_2403,In_3915);
and U2909 (N_2909,In_560,In_735);
nor U2910 (N_2910,In_3091,In_4428);
and U2911 (N_2911,In_3266,In_149);
xor U2912 (N_2912,In_1148,In_3010);
nor U2913 (N_2913,In_4042,In_2884);
nor U2914 (N_2914,In_3552,In_3492);
xnor U2915 (N_2915,In_107,In_3591);
and U2916 (N_2916,In_2024,In_1132);
nand U2917 (N_2917,In_1694,In_4707);
nor U2918 (N_2918,In_2053,In_1983);
nand U2919 (N_2919,In_4105,In_3266);
nand U2920 (N_2920,In_3266,In_3168);
or U2921 (N_2921,In_4635,In_176);
nor U2922 (N_2922,In_2589,In_1029);
and U2923 (N_2923,In_3521,In_2627);
nand U2924 (N_2924,In_4455,In_943);
nand U2925 (N_2925,In_245,In_2370);
or U2926 (N_2926,In_2142,In_1353);
and U2927 (N_2927,In_4373,In_2028);
nor U2928 (N_2928,In_1266,In_2802);
or U2929 (N_2929,In_983,In_511);
nand U2930 (N_2930,In_3077,In_3431);
nand U2931 (N_2931,In_4818,In_3484);
xor U2932 (N_2932,In_2870,In_4740);
nand U2933 (N_2933,In_484,In_316);
xnor U2934 (N_2934,In_3181,In_4171);
nand U2935 (N_2935,In_3320,In_4792);
nand U2936 (N_2936,In_1308,In_2466);
and U2937 (N_2937,In_2765,In_744);
nand U2938 (N_2938,In_4792,In_2311);
nor U2939 (N_2939,In_1840,In_1132);
nor U2940 (N_2940,In_3358,In_565);
nand U2941 (N_2941,In_2764,In_1568);
nor U2942 (N_2942,In_4229,In_2543);
or U2943 (N_2943,In_3686,In_1063);
nand U2944 (N_2944,In_640,In_3854);
nor U2945 (N_2945,In_1439,In_2853);
nand U2946 (N_2946,In_3702,In_164);
nand U2947 (N_2947,In_2498,In_4492);
nand U2948 (N_2948,In_2508,In_2481);
or U2949 (N_2949,In_4690,In_3333);
or U2950 (N_2950,In_1435,In_4867);
or U2951 (N_2951,In_676,In_3065);
xor U2952 (N_2952,In_3402,In_4714);
nand U2953 (N_2953,In_666,In_2598);
xor U2954 (N_2954,In_2020,In_3531);
xor U2955 (N_2955,In_4143,In_435);
and U2956 (N_2956,In_2727,In_1637);
nor U2957 (N_2957,In_4401,In_4200);
and U2958 (N_2958,In_2813,In_2414);
xnor U2959 (N_2959,In_2796,In_1961);
and U2960 (N_2960,In_1204,In_2577);
nor U2961 (N_2961,In_328,In_4493);
and U2962 (N_2962,In_2625,In_4267);
xnor U2963 (N_2963,In_855,In_488);
and U2964 (N_2964,In_4034,In_1401);
or U2965 (N_2965,In_2362,In_3171);
and U2966 (N_2966,In_2238,In_1331);
or U2967 (N_2967,In_3233,In_2184);
xnor U2968 (N_2968,In_1087,In_3781);
nand U2969 (N_2969,In_1611,In_4975);
nand U2970 (N_2970,In_4473,In_870);
nor U2971 (N_2971,In_3685,In_3978);
xnor U2972 (N_2972,In_31,In_807);
nand U2973 (N_2973,In_289,In_1918);
xnor U2974 (N_2974,In_392,In_4388);
nand U2975 (N_2975,In_1548,In_362);
and U2976 (N_2976,In_1152,In_612);
nand U2977 (N_2977,In_4547,In_1292);
xnor U2978 (N_2978,In_2309,In_1336);
nand U2979 (N_2979,In_330,In_4276);
or U2980 (N_2980,In_2541,In_2788);
xor U2981 (N_2981,In_1209,In_3226);
and U2982 (N_2982,In_4680,In_4357);
and U2983 (N_2983,In_3360,In_994);
nand U2984 (N_2984,In_3031,In_4245);
nand U2985 (N_2985,In_1478,In_4235);
nand U2986 (N_2986,In_2962,In_2904);
xnor U2987 (N_2987,In_2708,In_1125);
nand U2988 (N_2988,In_994,In_4681);
or U2989 (N_2989,In_839,In_4039);
or U2990 (N_2990,In_3544,In_216);
xor U2991 (N_2991,In_1949,In_347);
and U2992 (N_2992,In_1879,In_4406);
nor U2993 (N_2993,In_4878,In_3416);
nor U2994 (N_2994,In_905,In_3959);
and U2995 (N_2995,In_1454,In_4786);
nand U2996 (N_2996,In_3642,In_2871);
xnor U2997 (N_2997,In_2912,In_4768);
xnor U2998 (N_2998,In_1028,In_4226);
xnor U2999 (N_2999,In_868,In_576);
or U3000 (N_3000,In_4158,In_2322);
nand U3001 (N_3001,In_1443,In_1607);
or U3002 (N_3002,In_3735,In_558);
nand U3003 (N_3003,In_1651,In_585);
nor U3004 (N_3004,In_2785,In_3300);
and U3005 (N_3005,In_246,In_1490);
nand U3006 (N_3006,In_719,In_1250);
xnor U3007 (N_3007,In_3297,In_4772);
nor U3008 (N_3008,In_3171,In_4868);
or U3009 (N_3009,In_346,In_3913);
nor U3010 (N_3010,In_195,In_133);
and U3011 (N_3011,In_4715,In_4275);
nand U3012 (N_3012,In_3574,In_3198);
nand U3013 (N_3013,In_2791,In_1044);
xor U3014 (N_3014,In_1253,In_4826);
and U3015 (N_3015,In_2785,In_2583);
or U3016 (N_3016,In_3748,In_378);
nor U3017 (N_3017,In_1673,In_1423);
nor U3018 (N_3018,In_171,In_2238);
or U3019 (N_3019,In_1496,In_936);
nand U3020 (N_3020,In_2553,In_2750);
nand U3021 (N_3021,In_2356,In_3653);
xnor U3022 (N_3022,In_4225,In_219);
nor U3023 (N_3023,In_2824,In_1187);
and U3024 (N_3024,In_251,In_1907);
xnor U3025 (N_3025,In_853,In_4989);
or U3026 (N_3026,In_79,In_3031);
nor U3027 (N_3027,In_2927,In_23);
and U3028 (N_3028,In_1281,In_2536);
and U3029 (N_3029,In_1710,In_586);
nand U3030 (N_3030,In_4711,In_360);
nand U3031 (N_3031,In_50,In_1112);
or U3032 (N_3032,In_3516,In_147);
xor U3033 (N_3033,In_496,In_3395);
nand U3034 (N_3034,In_4160,In_3044);
or U3035 (N_3035,In_2761,In_4691);
or U3036 (N_3036,In_4739,In_216);
xnor U3037 (N_3037,In_165,In_2286);
and U3038 (N_3038,In_1222,In_2592);
and U3039 (N_3039,In_4907,In_3076);
or U3040 (N_3040,In_896,In_4508);
or U3041 (N_3041,In_3025,In_45);
nand U3042 (N_3042,In_957,In_2616);
and U3043 (N_3043,In_2905,In_480);
and U3044 (N_3044,In_2516,In_4160);
xor U3045 (N_3045,In_3455,In_1148);
and U3046 (N_3046,In_1718,In_1153);
nor U3047 (N_3047,In_3535,In_126);
and U3048 (N_3048,In_219,In_1971);
xor U3049 (N_3049,In_2681,In_3992);
and U3050 (N_3050,In_3409,In_670);
nor U3051 (N_3051,In_1954,In_2654);
xnor U3052 (N_3052,In_3014,In_1195);
nor U3053 (N_3053,In_532,In_3447);
nor U3054 (N_3054,In_4935,In_3409);
and U3055 (N_3055,In_2841,In_1187);
and U3056 (N_3056,In_357,In_3038);
xnor U3057 (N_3057,In_4089,In_3134);
nor U3058 (N_3058,In_1041,In_3929);
or U3059 (N_3059,In_1857,In_3406);
and U3060 (N_3060,In_1969,In_379);
nand U3061 (N_3061,In_4831,In_3162);
and U3062 (N_3062,In_791,In_482);
nor U3063 (N_3063,In_1776,In_756);
nor U3064 (N_3064,In_2940,In_621);
xor U3065 (N_3065,In_3379,In_4128);
nor U3066 (N_3066,In_4552,In_156);
or U3067 (N_3067,In_4017,In_2564);
nor U3068 (N_3068,In_962,In_928);
xor U3069 (N_3069,In_1036,In_3416);
xor U3070 (N_3070,In_4232,In_1268);
and U3071 (N_3071,In_193,In_3487);
and U3072 (N_3072,In_3520,In_3948);
or U3073 (N_3073,In_2356,In_2343);
nand U3074 (N_3074,In_2764,In_3021);
nand U3075 (N_3075,In_1606,In_4975);
nand U3076 (N_3076,In_1929,In_2707);
nor U3077 (N_3077,In_882,In_4288);
and U3078 (N_3078,In_3263,In_4236);
nand U3079 (N_3079,In_3817,In_2847);
and U3080 (N_3080,In_4547,In_1672);
nand U3081 (N_3081,In_3802,In_3206);
xnor U3082 (N_3082,In_3013,In_1329);
nor U3083 (N_3083,In_540,In_4542);
nand U3084 (N_3084,In_3794,In_1461);
nor U3085 (N_3085,In_1158,In_3820);
or U3086 (N_3086,In_2368,In_1999);
xor U3087 (N_3087,In_2875,In_1270);
nor U3088 (N_3088,In_3997,In_139);
nand U3089 (N_3089,In_1129,In_596);
xor U3090 (N_3090,In_3867,In_4461);
and U3091 (N_3091,In_3689,In_3367);
and U3092 (N_3092,In_4528,In_2978);
xor U3093 (N_3093,In_97,In_2354);
or U3094 (N_3094,In_1523,In_1791);
nand U3095 (N_3095,In_2104,In_483);
and U3096 (N_3096,In_1034,In_2145);
nor U3097 (N_3097,In_64,In_3695);
and U3098 (N_3098,In_4578,In_2183);
xnor U3099 (N_3099,In_414,In_2091);
nand U3100 (N_3100,In_2583,In_79);
nand U3101 (N_3101,In_2895,In_1851);
nand U3102 (N_3102,In_2222,In_2061);
and U3103 (N_3103,In_2065,In_2806);
nor U3104 (N_3104,In_735,In_2790);
or U3105 (N_3105,In_972,In_3934);
nor U3106 (N_3106,In_4472,In_2202);
and U3107 (N_3107,In_4822,In_3377);
nand U3108 (N_3108,In_2403,In_1463);
or U3109 (N_3109,In_4350,In_72);
xor U3110 (N_3110,In_801,In_4039);
nor U3111 (N_3111,In_1614,In_1055);
and U3112 (N_3112,In_976,In_4022);
or U3113 (N_3113,In_2849,In_3070);
xnor U3114 (N_3114,In_2459,In_1280);
nor U3115 (N_3115,In_3545,In_233);
xnor U3116 (N_3116,In_3492,In_4693);
xor U3117 (N_3117,In_4087,In_278);
or U3118 (N_3118,In_2647,In_2689);
xor U3119 (N_3119,In_2826,In_747);
and U3120 (N_3120,In_1749,In_2139);
nand U3121 (N_3121,In_1750,In_2574);
nand U3122 (N_3122,In_295,In_2736);
xor U3123 (N_3123,In_2508,In_2609);
xor U3124 (N_3124,In_621,In_1375);
nand U3125 (N_3125,In_1416,In_2269);
and U3126 (N_3126,In_1458,In_577);
nand U3127 (N_3127,In_2128,In_4562);
or U3128 (N_3128,In_4043,In_921);
nor U3129 (N_3129,In_1011,In_628);
xnor U3130 (N_3130,In_2458,In_984);
nor U3131 (N_3131,In_3821,In_610);
nand U3132 (N_3132,In_344,In_1435);
nand U3133 (N_3133,In_4168,In_4322);
and U3134 (N_3134,In_2306,In_1674);
or U3135 (N_3135,In_1411,In_305);
xnor U3136 (N_3136,In_1879,In_3308);
nand U3137 (N_3137,In_1500,In_1971);
nor U3138 (N_3138,In_1756,In_3886);
nand U3139 (N_3139,In_1170,In_242);
or U3140 (N_3140,In_1888,In_2721);
or U3141 (N_3141,In_3581,In_4127);
nand U3142 (N_3142,In_1344,In_4062);
xnor U3143 (N_3143,In_4088,In_904);
xor U3144 (N_3144,In_1244,In_1822);
and U3145 (N_3145,In_1667,In_727);
and U3146 (N_3146,In_4290,In_1194);
and U3147 (N_3147,In_727,In_3648);
xnor U3148 (N_3148,In_4450,In_4394);
xnor U3149 (N_3149,In_392,In_2519);
xnor U3150 (N_3150,In_1816,In_3977);
xor U3151 (N_3151,In_2750,In_1502);
nand U3152 (N_3152,In_3366,In_3892);
xor U3153 (N_3153,In_1888,In_4418);
and U3154 (N_3154,In_1327,In_4165);
and U3155 (N_3155,In_1448,In_392);
or U3156 (N_3156,In_4789,In_3055);
xor U3157 (N_3157,In_1294,In_1238);
or U3158 (N_3158,In_4849,In_3108);
or U3159 (N_3159,In_1885,In_4489);
and U3160 (N_3160,In_4761,In_3915);
or U3161 (N_3161,In_3200,In_2303);
xor U3162 (N_3162,In_3746,In_284);
and U3163 (N_3163,In_3236,In_4980);
xnor U3164 (N_3164,In_254,In_4741);
or U3165 (N_3165,In_2336,In_2220);
nand U3166 (N_3166,In_2719,In_4807);
or U3167 (N_3167,In_2726,In_3484);
xor U3168 (N_3168,In_2005,In_2935);
or U3169 (N_3169,In_4731,In_1792);
and U3170 (N_3170,In_1455,In_3555);
xor U3171 (N_3171,In_4995,In_1706);
and U3172 (N_3172,In_2245,In_3624);
or U3173 (N_3173,In_2482,In_4452);
and U3174 (N_3174,In_1375,In_471);
nand U3175 (N_3175,In_3196,In_2141);
nor U3176 (N_3176,In_49,In_4950);
and U3177 (N_3177,In_3360,In_4181);
nand U3178 (N_3178,In_2985,In_3584);
nand U3179 (N_3179,In_2749,In_2543);
nand U3180 (N_3180,In_4653,In_4075);
xor U3181 (N_3181,In_2419,In_1344);
xnor U3182 (N_3182,In_4487,In_569);
xnor U3183 (N_3183,In_519,In_4048);
and U3184 (N_3184,In_2968,In_3773);
nor U3185 (N_3185,In_4123,In_3453);
nor U3186 (N_3186,In_595,In_4549);
xnor U3187 (N_3187,In_2077,In_4218);
or U3188 (N_3188,In_1188,In_1329);
xnor U3189 (N_3189,In_3657,In_2396);
xor U3190 (N_3190,In_3169,In_1144);
nor U3191 (N_3191,In_47,In_3485);
xor U3192 (N_3192,In_3513,In_1462);
or U3193 (N_3193,In_2238,In_2318);
xnor U3194 (N_3194,In_1153,In_3205);
xor U3195 (N_3195,In_3110,In_3885);
or U3196 (N_3196,In_184,In_1577);
xor U3197 (N_3197,In_1923,In_4446);
nand U3198 (N_3198,In_948,In_2105);
xor U3199 (N_3199,In_1434,In_4326);
nand U3200 (N_3200,In_335,In_1961);
nand U3201 (N_3201,In_3401,In_3540);
xor U3202 (N_3202,In_3031,In_491);
xnor U3203 (N_3203,In_1357,In_4747);
nor U3204 (N_3204,In_4515,In_157);
nand U3205 (N_3205,In_1691,In_3293);
xnor U3206 (N_3206,In_4001,In_2217);
and U3207 (N_3207,In_1330,In_3550);
or U3208 (N_3208,In_4335,In_3555);
or U3209 (N_3209,In_4176,In_4566);
nand U3210 (N_3210,In_2147,In_4325);
and U3211 (N_3211,In_2956,In_821);
or U3212 (N_3212,In_4500,In_1496);
and U3213 (N_3213,In_2730,In_3308);
nand U3214 (N_3214,In_2795,In_2873);
xnor U3215 (N_3215,In_4483,In_3017);
xor U3216 (N_3216,In_2929,In_1513);
nand U3217 (N_3217,In_962,In_2737);
nor U3218 (N_3218,In_4525,In_2817);
and U3219 (N_3219,In_1137,In_4830);
nand U3220 (N_3220,In_496,In_4512);
xor U3221 (N_3221,In_2288,In_3936);
nand U3222 (N_3222,In_2622,In_120);
and U3223 (N_3223,In_3011,In_2807);
or U3224 (N_3224,In_4237,In_4756);
nor U3225 (N_3225,In_4117,In_907);
or U3226 (N_3226,In_457,In_3262);
and U3227 (N_3227,In_3478,In_2048);
xor U3228 (N_3228,In_1375,In_819);
nand U3229 (N_3229,In_1283,In_1980);
nor U3230 (N_3230,In_2243,In_4620);
or U3231 (N_3231,In_3040,In_963);
nand U3232 (N_3232,In_3044,In_4335);
nand U3233 (N_3233,In_4214,In_3780);
nor U3234 (N_3234,In_1730,In_1427);
xor U3235 (N_3235,In_4554,In_1025);
nand U3236 (N_3236,In_3140,In_4261);
nor U3237 (N_3237,In_4437,In_2161);
nor U3238 (N_3238,In_4542,In_3079);
xor U3239 (N_3239,In_2562,In_2642);
nand U3240 (N_3240,In_2033,In_4006);
and U3241 (N_3241,In_4587,In_4838);
xor U3242 (N_3242,In_2331,In_2340);
nand U3243 (N_3243,In_3131,In_4509);
nand U3244 (N_3244,In_3311,In_1304);
nor U3245 (N_3245,In_4417,In_4241);
or U3246 (N_3246,In_4503,In_2437);
nor U3247 (N_3247,In_1982,In_2977);
or U3248 (N_3248,In_1905,In_2325);
or U3249 (N_3249,In_3892,In_720);
nand U3250 (N_3250,In_4151,In_3809);
nand U3251 (N_3251,In_1089,In_4874);
nor U3252 (N_3252,In_4370,In_1242);
nor U3253 (N_3253,In_3799,In_4501);
nor U3254 (N_3254,In_4982,In_2071);
and U3255 (N_3255,In_2982,In_1744);
xor U3256 (N_3256,In_3899,In_2535);
xnor U3257 (N_3257,In_983,In_3664);
and U3258 (N_3258,In_2612,In_2273);
nand U3259 (N_3259,In_4005,In_1627);
and U3260 (N_3260,In_689,In_1869);
or U3261 (N_3261,In_1117,In_2700);
xor U3262 (N_3262,In_2276,In_4712);
or U3263 (N_3263,In_1860,In_1604);
or U3264 (N_3264,In_3009,In_2201);
or U3265 (N_3265,In_2803,In_1320);
and U3266 (N_3266,In_4560,In_3950);
or U3267 (N_3267,In_3609,In_1831);
xor U3268 (N_3268,In_1525,In_2672);
nand U3269 (N_3269,In_4223,In_3493);
xor U3270 (N_3270,In_156,In_604);
and U3271 (N_3271,In_4695,In_2624);
or U3272 (N_3272,In_3603,In_1766);
nor U3273 (N_3273,In_3279,In_4889);
xnor U3274 (N_3274,In_670,In_4384);
nor U3275 (N_3275,In_3825,In_3447);
or U3276 (N_3276,In_4291,In_4904);
and U3277 (N_3277,In_4302,In_2159);
and U3278 (N_3278,In_1304,In_2950);
or U3279 (N_3279,In_4647,In_2898);
nor U3280 (N_3280,In_4341,In_302);
nand U3281 (N_3281,In_3486,In_2233);
xor U3282 (N_3282,In_1824,In_277);
and U3283 (N_3283,In_1019,In_2225);
xor U3284 (N_3284,In_1118,In_4929);
or U3285 (N_3285,In_1277,In_2746);
or U3286 (N_3286,In_1049,In_3125);
or U3287 (N_3287,In_3001,In_40);
nor U3288 (N_3288,In_3231,In_663);
or U3289 (N_3289,In_4283,In_926);
xor U3290 (N_3290,In_2902,In_4847);
or U3291 (N_3291,In_4438,In_415);
and U3292 (N_3292,In_4116,In_1864);
and U3293 (N_3293,In_2756,In_1029);
or U3294 (N_3294,In_1267,In_3695);
xnor U3295 (N_3295,In_757,In_2396);
or U3296 (N_3296,In_3645,In_1309);
and U3297 (N_3297,In_262,In_717);
nor U3298 (N_3298,In_2036,In_1546);
and U3299 (N_3299,In_1484,In_2466);
nor U3300 (N_3300,In_4115,In_717);
or U3301 (N_3301,In_4236,In_360);
and U3302 (N_3302,In_4387,In_89);
nor U3303 (N_3303,In_1563,In_4621);
or U3304 (N_3304,In_3635,In_504);
nor U3305 (N_3305,In_3833,In_3526);
nand U3306 (N_3306,In_2488,In_4313);
nor U3307 (N_3307,In_3279,In_4950);
xor U3308 (N_3308,In_4801,In_1488);
nand U3309 (N_3309,In_50,In_4443);
and U3310 (N_3310,In_4829,In_807);
or U3311 (N_3311,In_822,In_1538);
nand U3312 (N_3312,In_4858,In_1632);
and U3313 (N_3313,In_2262,In_3930);
nand U3314 (N_3314,In_256,In_2136);
xnor U3315 (N_3315,In_3674,In_172);
nand U3316 (N_3316,In_624,In_660);
nand U3317 (N_3317,In_448,In_2431);
xnor U3318 (N_3318,In_21,In_3122);
nor U3319 (N_3319,In_1497,In_1770);
and U3320 (N_3320,In_4186,In_4621);
and U3321 (N_3321,In_1791,In_120);
nor U3322 (N_3322,In_4834,In_1810);
and U3323 (N_3323,In_1376,In_2811);
nor U3324 (N_3324,In_3096,In_754);
or U3325 (N_3325,In_3344,In_901);
or U3326 (N_3326,In_1483,In_1773);
nor U3327 (N_3327,In_2086,In_3761);
or U3328 (N_3328,In_1314,In_508);
and U3329 (N_3329,In_3503,In_470);
and U3330 (N_3330,In_3191,In_2833);
and U3331 (N_3331,In_3907,In_1881);
xnor U3332 (N_3332,In_4423,In_49);
xor U3333 (N_3333,In_3375,In_2788);
nor U3334 (N_3334,In_1014,In_940);
xor U3335 (N_3335,In_156,In_2489);
and U3336 (N_3336,In_3738,In_1248);
or U3337 (N_3337,In_456,In_381);
xnor U3338 (N_3338,In_95,In_4321);
xnor U3339 (N_3339,In_2886,In_1713);
xor U3340 (N_3340,In_4909,In_1247);
or U3341 (N_3341,In_1279,In_397);
nor U3342 (N_3342,In_3970,In_1807);
nor U3343 (N_3343,In_870,In_1489);
or U3344 (N_3344,In_2666,In_4704);
or U3345 (N_3345,In_333,In_1534);
nand U3346 (N_3346,In_4735,In_1748);
nand U3347 (N_3347,In_1244,In_1280);
and U3348 (N_3348,In_2880,In_1656);
nor U3349 (N_3349,In_2363,In_4425);
and U3350 (N_3350,In_808,In_210);
nor U3351 (N_3351,In_4679,In_4548);
and U3352 (N_3352,In_1427,In_2010);
nor U3353 (N_3353,In_77,In_570);
nor U3354 (N_3354,In_4841,In_1110);
and U3355 (N_3355,In_1920,In_2307);
nor U3356 (N_3356,In_487,In_1261);
nor U3357 (N_3357,In_2303,In_743);
nor U3358 (N_3358,In_913,In_3384);
or U3359 (N_3359,In_2006,In_4664);
nand U3360 (N_3360,In_4518,In_744);
and U3361 (N_3361,In_4212,In_4767);
or U3362 (N_3362,In_3656,In_869);
nand U3363 (N_3363,In_3710,In_749);
or U3364 (N_3364,In_2322,In_4862);
xor U3365 (N_3365,In_139,In_1162);
nor U3366 (N_3366,In_480,In_2871);
and U3367 (N_3367,In_4882,In_3494);
and U3368 (N_3368,In_338,In_1676);
nand U3369 (N_3369,In_1380,In_613);
or U3370 (N_3370,In_4293,In_1948);
and U3371 (N_3371,In_1384,In_3909);
nor U3372 (N_3372,In_1466,In_4189);
or U3373 (N_3373,In_3373,In_824);
xor U3374 (N_3374,In_3160,In_2711);
and U3375 (N_3375,In_1626,In_3);
nor U3376 (N_3376,In_757,In_633);
and U3377 (N_3377,In_293,In_3945);
or U3378 (N_3378,In_2976,In_158);
and U3379 (N_3379,In_3318,In_979);
nand U3380 (N_3380,In_698,In_642);
and U3381 (N_3381,In_4259,In_2862);
and U3382 (N_3382,In_516,In_327);
and U3383 (N_3383,In_4283,In_1571);
or U3384 (N_3384,In_576,In_1046);
nor U3385 (N_3385,In_3770,In_1222);
or U3386 (N_3386,In_2213,In_2865);
nor U3387 (N_3387,In_2984,In_1330);
nor U3388 (N_3388,In_1057,In_4190);
and U3389 (N_3389,In_2939,In_4612);
xor U3390 (N_3390,In_3947,In_1061);
and U3391 (N_3391,In_2666,In_570);
or U3392 (N_3392,In_3815,In_1014);
nor U3393 (N_3393,In_703,In_2009);
nand U3394 (N_3394,In_4299,In_3597);
nand U3395 (N_3395,In_4940,In_1510);
nor U3396 (N_3396,In_1225,In_1321);
nand U3397 (N_3397,In_2485,In_929);
and U3398 (N_3398,In_892,In_574);
nand U3399 (N_3399,In_2942,In_4667);
xnor U3400 (N_3400,In_3256,In_2754);
nor U3401 (N_3401,In_2248,In_3638);
nor U3402 (N_3402,In_612,In_1368);
or U3403 (N_3403,In_1422,In_3463);
xor U3404 (N_3404,In_3980,In_475);
xor U3405 (N_3405,In_1442,In_2424);
xor U3406 (N_3406,In_533,In_2976);
xnor U3407 (N_3407,In_1078,In_2094);
or U3408 (N_3408,In_4045,In_2489);
and U3409 (N_3409,In_9,In_975);
and U3410 (N_3410,In_1722,In_2318);
nor U3411 (N_3411,In_1947,In_4313);
nand U3412 (N_3412,In_1160,In_3028);
xnor U3413 (N_3413,In_4293,In_313);
xor U3414 (N_3414,In_2222,In_4020);
xor U3415 (N_3415,In_2728,In_3020);
or U3416 (N_3416,In_1042,In_3555);
nand U3417 (N_3417,In_3185,In_2397);
and U3418 (N_3418,In_81,In_4621);
and U3419 (N_3419,In_168,In_1345);
nand U3420 (N_3420,In_1050,In_192);
nand U3421 (N_3421,In_418,In_1143);
nor U3422 (N_3422,In_1183,In_4582);
nand U3423 (N_3423,In_4067,In_3002);
nor U3424 (N_3424,In_1489,In_2240);
xnor U3425 (N_3425,In_30,In_2549);
nand U3426 (N_3426,In_3290,In_4239);
or U3427 (N_3427,In_34,In_3265);
and U3428 (N_3428,In_1808,In_2170);
nor U3429 (N_3429,In_2781,In_628);
and U3430 (N_3430,In_4012,In_2221);
and U3431 (N_3431,In_3525,In_2441);
and U3432 (N_3432,In_1162,In_2216);
nor U3433 (N_3433,In_189,In_3375);
nor U3434 (N_3434,In_1452,In_4001);
xor U3435 (N_3435,In_627,In_4496);
and U3436 (N_3436,In_880,In_2909);
nand U3437 (N_3437,In_4097,In_3925);
nor U3438 (N_3438,In_468,In_2092);
nor U3439 (N_3439,In_4956,In_1728);
or U3440 (N_3440,In_2802,In_1652);
nor U3441 (N_3441,In_4290,In_3441);
nand U3442 (N_3442,In_2993,In_2906);
xnor U3443 (N_3443,In_4741,In_1723);
nor U3444 (N_3444,In_4401,In_1187);
xnor U3445 (N_3445,In_2678,In_89);
xor U3446 (N_3446,In_2165,In_3732);
or U3447 (N_3447,In_3191,In_1065);
or U3448 (N_3448,In_3667,In_1131);
and U3449 (N_3449,In_4734,In_4410);
xor U3450 (N_3450,In_517,In_4292);
xor U3451 (N_3451,In_4272,In_205);
nor U3452 (N_3452,In_4614,In_3211);
xor U3453 (N_3453,In_1019,In_389);
xor U3454 (N_3454,In_4300,In_1903);
nand U3455 (N_3455,In_2177,In_2899);
and U3456 (N_3456,In_2241,In_475);
and U3457 (N_3457,In_721,In_1446);
and U3458 (N_3458,In_1100,In_4826);
nand U3459 (N_3459,In_3933,In_462);
and U3460 (N_3460,In_3774,In_4362);
nor U3461 (N_3461,In_3789,In_2509);
nand U3462 (N_3462,In_4668,In_2692);
or U3463 (N_3463,In_4941,In_3389);
nand U3464 (N_3464,In_3649,In_708);
xor U3465 (N_3465,In_4120,In_2593);
or U3466 (N_3466,In_2434,In_4087);
xnor U3467 (N_3467,In_2949,In_1723);
and U3468 (N_3468,In_2359,In_3312);
nand U3469 (N_3469,In_422,In_4418);
xnor U3470 (N_3470,In_127,In_4375);
nand U3471 (N_3471,In_131,In_1730);
nand U3472 (N_3472,In_4676,In_1401);
and U3473 (N_3473,In_4485,In_809);
and U3474 (N_3474,In_1709,In_2579);
and U3475 (N_3475,In_619,In_4171);
or U3476 (N_3476,In_1853,In_1474);
nor U3477 (N_3477,In_90,In_2819);
and U3478 (N_3478,In_1775,In_1328);
or U3479 (N_3479,In_1894,In_3812);
nand U3480 (N_3480,In_1109,In_4899);
nor U3481 (N_3481,In_1224,In_1158);
and U3482 (N_3482,In_3612,In_4550);
xnor U3483 (N_3483,In_2336,In_4939);
or U3484 (N_3484,In_3689,In_1062);
nand U3485 (N_3485,In_2727,In_1794);
and U3486 (N_3486,In_2362,In_2990);
nand U3487 (N_3487,In_1550,In_1477);
and U3488 (N_3488,In_1384,In_2399);
nor U3489 (N_3489,In_3834,In_2917);
nand U3490 (N_3490,In_1170,In_4819);
nor U3491 (N_3491,In_2661,In_4855);
xor U3492 (N_3492,In_3960,In_3865);
xor U3493 (N_3493,In_1229,In_4378);
nor U3494 (N_3494,In_4872,In_637);
xnor U3495 (N_3495,In_1430,In_48);
xor U3496 (N_3496,In_106,In_207);
and U3497 (N_3497,In_858,In_659);
nor U3498 (N_3498,In_4024,In_2291);
nor U3499 (N_3499,In_1682,In_4574);
nand U3500 (N_3500,In_3111,In_4543);
xor U3501 (N_3501,In_4736,In_3206);
xor U3502 (N_3502,In_86,In_3129);
xor U3503 (N_3503,In_4023,In_1054);
and U3504 (N_3504,In_4188,In_4359);
or U3505 (N_3505,In_2335,In_3502);
xnor U3506 (N_3506,In_3810,In_4647);
nor U3507 (N_3507,In_3032,In_1935);
xor U3508 (N_3508,In_3894,In_1884);
xnor U3509 (N_3509,In_990,In_808);
or U3510 (N_3510,In_2598,In_25);
and U3511 (N_3511,In_2110,In_4923);
or U3512 (N_3512,In_61,In_2670);
or U3513 (N_3513,In_733,In_80);
or U3514 (N_3514,In_1329,In_443);
nand U3515 (N_3515,In_4723,In_2443);
xor U3516 (N_3516,In_12,In_627);
xor U3517 (N_3517,In_4621,In_4983);
xnor U3518 (N_3518,In_3391,In_1222);
and U3519 (N_3519,In_3784,In_2001);
xor U3520 (N_3520,In_1554,In_2114);
and U3521 (N_3521,In_1956,In_1235);
nor U3522 (N_3522,In_1317,In_2007);
nand U3523 (N_3523,In_4735,In_536);
and U3524 (N_3524,In_2819,In_3325);
or U3525 (N_3525,In_3369,In_934);
nor U3526 (N_3526,In_1253,In_2544);
or U3527 (N_3527,In_2396,In_3671);
and U3528 (N_3528,In_917,In_2759);
xor U3529 (N_3529,In_731,In_4645);
nor U3530 (N_3530,In_485,In_3372);
or U3531 (N_3531,In_644,In_1020);
xor U3532 (N_3532,In_1498,In_2219);
nand U3533 (N_3533,In_2426,In_478);
nand U3534 (N_3534,In_3739,In_2072);
nand U3535 (N_3535,In_196,In_4332);
or U3536 (N_3536,In_1427,In_2505);
nand U3537 (N_3537,In_2323,In_1186);
nor U3538 (N_3538,In_3872,In_1924);
nand U3539 (N_3539,In_4108,In_3942);
nand U3540 (N_3540,In_3311,In_928);
and U3541 (N_3541,In_1103,In_3912);
nor U3542 (N_3542,In_3118,In_1538);
nand U3543 (N_3543,In_1215,In_316);
nand U3544 (N_3544,In_618,In_3218);
xnor U3545 (N_3545,In_2366,In_2401);
nor U3546 (N_3546,In_4891,In_1089);
and U3547 (N_3547,In_4821,In_242);
xor U3548 (N_3548,In_1490,In_704);
nand U3549 (N_3549,In_2545,In_2303);
nand U3550 (N_3550,In_1855,In_1889);
nor U3551 (N_3551,In_4916,In_2809);
nor U3552 (N_3552,In_3002,In_2385);
and U3553 (N_3553,In_2737,In_486);
xnor U3554 (N_3554,In_1299,In_3074);
nand U3555 (N_3555,In_3414,In_4054);
or U3556 (N_3556,In_4503,In_1378);
and U3557 (N_3557,In_3145,In_2232);
nor U3558 (N_3558,In_3413,In_1524);
nand U3559 (N_3559,In_974,In_170);
or U3560 (N_3560,In_4901,In_4855);
or U3561 (N_3561,In_1085,In_1127);
or U3562 (N_3562,In_1362,In_1747);
nand U3563 (N_3563,In_3977,In_4749);
nand U3564 (N_3564,In_1812,In_4787);
or U3565 (N_3565,In_4180,In_3439);
and U3566 (N_3566,In_4628,In_2496);
or U3567 (N_3567,In_4704,In_441);
xor U3568 (N_3568,In_1973,In_3891);
or U3569 (N_3569,In_2660,In_1481);
xnor U3570 (N_3570,In_934,In_652);
xor U3571 (N_3571,In_3984,In_1111);
or U3572 (N_3572,In_3003,In_563);
xnor U3573 (N_3573,In_2280,In_3204);
nor U3574 (N_3574,In_2062,In_4519);
xnor U3575 (N_3575,In_4645,In_4696);
nand U3576 (N_3576,In_2022,In_3504);
xnor U3577 (N_3577,In_2961,In_84);
or U3578 (N_3578,In_3538,In_3362);
or U3579 (N_3579,In_1331,In_2926);
and U3580 (N_3580,In_3603,In_267);
or U3581 (N_3581,In_2785,In_3114);
xnor U3582 (N_3582,In_2357,In_3317);
xor U3583 (N_3583,In_3578,In_3623);
and U3584 (N_3584,In_2640,In_2741);
or U3585 (N_3585,In_3151,In_3834);
nor U3586 (N_3586,In_4718,In_4461);
and U3587 (N_3587,In_1293,In_3651);
or U3588 (N_3588,In_3227,In_1757);
and U3589 (N_3589,In_4995,In_2592);
or U3590 (N_3590,In_4325,In_1181);
and U3591 (N_3591,In_1139,In_3267);
nor U3592 (N_3592,In_676,In_2314);
or U3593 (N_3593,In_4668,In_1322);
or U3594 (N_3594,In_1090,In_1033);
nor U3595 (N_3595,In_2385,In_3646);
xor U3596 (N_3596,In_4464,In_953);
nand U3597 (N_3597,In_4392,In_1411);
and U3598 (N_3598,In_3297,In_1082);
xor U3599 (N_3599,In_3855,In_2379);
xnor U3600 (N_3600,In_4701,In_3917);
nor U3601 (N_3601,In_3346,In_125);
xor U3602 (N_3602,In_4128,In_474);
xnor U3603 (N_3603,In_1156,In_2063);
and U3604 (N_3604,In_1883,In_939);
nor U3605 (N_3605,In_1293,In_682);
xnor U3606 (N_3606,In_4991,In_3665);
and U3607 (N_3607,In_4448,In_2276);
and U3608 (N_3608,In_3921,In_612);
xnor U3609 (N_3609,In_1232,In_4299);
or U3610 (N_3610,In_495,In_1871);
nor U3611 (N_3611,In_4306,In_2152);
xnor U3612 (N_3612,In_3951,In_983);
xnor U3613 (N_3613,In_337,In_2494);
or U3614 (N_3614,In_337,In_1420);
and U3615 (N_3615,In_4994,In_332);
nand U3616 (N_3616,In_2576,In_1076);
xnor U3617 (N_3617,In_4506,In_4233);
and U3618 (N_3618,In_3200,In_4695);
nand U3619 (N_3619,In_1637,In_23);
and U3620 (N_3620,In_1037,In_1539);
nand U3621 (N_3621,In_1704,In_197);
or U3622 (N_3622,In_4897,In_2135);
nand U3623 (N_3623,In_4590,In_520);
or U3624 (N_3624,In_4141,In_2363);
xnor U3625 (N_3625,In_1381,In_235);
or U3626 (N_3626,In_1919,In_2119);
nand U3627 (N_3627,In_459,In_4805);
nand U3628 (N_3628,In_1633,In_438);
or U3629 (N_3629,In_3995,In_3996);
nand U3630 (N_3630,In_1208,In_3269);
or U3631 (N_3631,In_4257,In_4132);
nor U3632 (N_3632,In_4116,In_1691);
xor U3633 (N_3633,In_1489,In_647);
and U3634 (N_3634,In_2414,In_1223);
and U3635 (N_3635,In_3889,In_1368);
nor U3636 (N_3636,In_896,In_793);
nand U3637 (N_3637,In_1566,In_4881);
and U3638 (N_3638,In_1076,In_1);
and U3639 (N_3639,In_378,In_749);
xnor U3640 (N_3640,In_1709,In_1878);
or U3641 (N_3641,In_3283,In_3384);
or U3642 (N_3642,In_1470,In_112);
and U3643 (N_3643,In_3808,In_2105);
nor U3644 (N_3644,In_628,In_3163);
nor U3645 (N_3645,In_4214,In_1473);
xor U3646 (N_3646,In_657,In_209);
or U3647 (N_3647,In_3454,In_4735);
xor U3648 (N_3648,In_603,In_3002);
or U3649 (N_3649,In_1936,In_4945);
xor U3650 (N_3650,In_439,In_2441);
nand U3651 (N_3651,In_4810,In_181);
nor U3652 (N_3652,In_3104,In_406);
and U3653 (N_3653,In_1980,In_1907);
or U3654 (N_3654,In_1586,In_932);
xor U3655 (N_3655,In_2819,In_2447);
nand U3656 (N_3656,In_1432,In_2931);
or U3657 (N_3657,In_1470,In_4057);
nand U3658 (N_3658,In_756,In_2280);
nand U3659 (N_3659,In_3695,In_1796);
nor U3660 (N_3660,In_4633,In_2553);
or U3661 (N_3661,In_4514,In_4136);
and U3662 (N_3662,In_2163,In_2956);
or U3663 (N_3663,In_450,In_2016);
or U3664 (N_3664,In_773,In_1924);
or U3665 (N_3665,In_2679,In_247);
nand U3666 (N_3666,In_3259,In_3940);
or U3667 (N_3667,In_357,In_1055);
or U3668 (N_3668,In_3640,In_1667);
nor U3669 (N_3669,In_2171,In_2113);
or U3670 (N_3670,In_1801,In_3489);
nand U3671 (N_3671,In_3301,In_4067);
and U3672 (N_3672,In_4510,In_2837);
xnor U3673 (N_3673,In_801,In_3716);
xor U3674 (N_3674,In_2420,In_3964);
or U3675 (N_3675,In_906,In_1371);
nand U3676 (N_3676,In_4022,In_4814);
nand U3677 (N_3677,In_2497,In_4972);
xor U3678 (N_3678,In_2228,In_4859);
xor U3679 (N_3679,In_1907,In_360);
or U3680 (N_3680,In_476,In_167);
and U3681 (N_3681,In_3060,In_4443);
nor U3682 (N_3682,In_1331,In_1113);
or U3683 (N_3683,In_3489,In_3022);
nor U3684 (N_3684,In_1839,In_3301);
nor U3685 (N_3685,In_85,In_3162);
xor U3686 (N_3686,In_2111,In_4920);
or U3687 (N_3687,In_690,In_205);
nand U3688 (N_3688,In_4167,In_2076);
and U3689 (N_3689,In_1288,In_3929);
xnor U3690 (N_3690,In_3346,In_2958);
nand U3691 (N_3691,In_4770,In_40);
xor U3692 (N_3692,In_2263,In_1025);
nand U3693 (N_3693,In_4471,In_4460);
or U3694 (N_3694,In_2767,In_4236);
or U3695 (N_3695,In_1431,In_1525);
or U3696 (N_3696,In_3724,In_2431);
or U3697 (N_3697,In_1052,In_2921);
and U3698 (N_3698,In_4298,In_4388);
nor U3699 (N_3699,In_1749,In_1980);
nand U3700 (N_3700,In_851,In_3403);
or U3701 (N_3701,In_3136,In_3340);
or U3702 (N_3702,In_3309,In_1319);
or U3703 (N_3703,In_2061,In_2072);
nand U3704 (N_3704,In_4349,In_523);
nand U3705 (N_3705,In_1423,In_2857);
nor U3706 (N_3706,In_1814,In_1813);
and U3707 (N_3707,In_1346,In_315);
nor U3708 (N_3708,In_2540,In_31);
nand U3709 (N_3709,In_1817,In_3513);
or U3710 (N_3710,In_3539,In_4013);
nor U3711 (N_3711,In_3365,In_2496);
nor U3712 (N_3712,In_1653,In_2139);
and U3713 (N_3713,In_2444,In_1787);
nand U3714 (N_3714,In_3686,In_347);
and U3715 (N_3715,In_1848,In_2380);
nand U3716 (N_3716,In_1739,In_3550);
nand U3717 (N_3717,In_396,In_2899);
and U3718 (N_3718,In_1102,In_3774);
nand U3719 (N_3719,In_523,In_2297);
or U3720 (N_3720,In_4123,In_1515);
and U3721 (N_3721,In_6,In_48);
nor U3722 (N_3722,In_4563,In_247);
or U3723 (N_3723,In_3736,In_1291);
or U3724 (N_3724,In_1599,In_2875);
nor U3725 (N_3725,In_384,In_1132);
and U3726 (N_3726,In_3303,In_131);
and U3727 (N_3727,In_4352,In_4900);
xnor U3728 (N_3728,In_2542,In_4365);
and U3729 (N_3729,In_852,In_81);
or U3730 (N_3730,In_2749,In_3637);
nand U3731 (N_3731,In_4607,In_817);
nor U3732 (N_3732,In_2219,In_3662);
or U3733 (N_3733,In_1099,In_4598);
nand U3734 (N_3734,In_4133,In_4985);
xor U3735 (N_3735,In_4890,In_2798);
nor U3736 (N_3736,In_1315,In_4487);
xor U3737 (N_3737,In_4350,In_4798);
and U3738 (N_3738,In_2417,In_2028);
nand U3739 (N_3739,In_1282,In_2392);
nor U3740 (N_3740,In_911,In_4424);
nor U3741 (N_3741,In_159,In_2740);
or U3742 (N_3742,In_4662,In_3861);
nand U3743 (N_3743,In_3711,In_4904);
xnor U3744 (N_3744,In_3413,In_4366);
nor U3745 (N_3745,In_3698,In_2204);
nor U3746 (N_3746,In_2041,In_3998);
nor U3747 (N_3747,In_1894,In_784);
nand U3748 (N_3748,In_3773,In_3899);
xor U3749 (N_3749,In_1120,In_3360);
nor U3750 (N_3750,In_218,In_2009);
nor U3751 (N_3751,In_2138,In_1578);
or U3752 (N_3752,In_2474,In_2832);
or U3753 (N_3753,In_859,In_3685);
or U3754 (N_3754,In_2877,In_1358);
and U3755 (N_3755,In_3241,In_4079);
nand U3756 (N_3756,In_1277,In_4959);
xor U3757 (N_3757,In_4875,In_4347);
and U3758 (N_3758,In_2064,In_3563);
xor U3759 (N_3759,In_3075,In_295);
xor U3760 (N_3760,In_1049,In_3799);
or U3761 (N_3761,In_3784,In_3345);
and U3762 (N_3762,In_1656,In_4726);
or U3763 (N_3763,In_2148,In_3006);
or U3764 (N_3764,In_29,In_2563);
nor U3765 (N_3765,In_1104,In_510);
and U3766 (N_3766,In_2109,In_434);
and U3767 (N_3767,In_3558,In_4298);
xor U3768 (N_3768,In_4347,In_2713);
or U3769 (N_3769,In_112,In_908);
and U3770 (N_3770,In_3193,In_3618);
nor U3771 (N_3771,In_3975,In_4967);
or U3772 (N_3772,In_3695,In_4168);
nor U3773 (N_3773,In_86,In_2652);
nand U3774 (N_3774,In_3344,In_3067);
nand U3775 (N_3775,In_4762,In_4837);
or U3776 (N_3776,In_1491,In_2060);
nand U3777 (N_3777,In_825,In_963);
nor U3778 (N_3778,In_3595,In_1921);
nor U3779 (N_3779,In_4493,In_3530);
or U3780 (N_3780,In_2860,In_538);
and U3781 (N_3781,In_2044,In_761);
xnor U3782 (N_3782,In_3138,In_409);
nor U3783 (N_3783,In_4957,In_2199);
xnor U3784 (N_3784,In_3838,In_3390);
or U3785 (N_3785,In_4780,In_2519);
or U3786 (N_3786,In_323,In_875);
nor U3787 (N_3787,In_4289,In_1935);
nand U3788 (N_3788,In_525,In_2943);
or U3789 (N_3789,In_4680,In_4117);
xor U3790 (N_3790,In_4593,In_4647);
xor U3791 (N_3791,In_4540,In_3944);
xnor U3792 (N_3792,In_349,In_4789);
nand U3793 (N_3793,In_484,In_2137);
and U3794 (N_3794,In_4788,In_1890);
and U3795 (N_3795,In_4173,In_2031);
nor U3796 (N_3796,In_1179,In_1779);
xnor U3797 (N_3797,In_415,In_1841);
xor U3798 (N_3798,In_351,In_1895);
nor U3799 (N_3799,In_495,In_4606);
or U3800 (N_3800,In_3753,In_2435);
nor U3801 (N_3801,In_2991,In_4056);
nor U3802 (N_3802,In_1695,In_1683);
nand U3803 (N_3803,In_3203,In_1825);
nor U3804 (N_3804,In_810,In_1121);
or U3805 (N_3805,In_216,In_1378);
and U3806 (N_3806,In_384,In_85);
nor U3807 (N_3807,In_2223,In_599);
xnor U3808 (N_3808,In_2638,In_1169);
nand U3809 (N_3809,In_2321,In_3518);
nor U3810 (N_3810,In_3037,In_35);
xnor U3811 (N_3811,In_2496,In_528);
nand U3812 (N_3812,In_3337,In_4622);
nand U3813 (N_3813,In_659,In_187);
xor U3814 (N_3814,In_1097,In_1541);
and U3815 (N_3815,In_4758,In_1202);
xor U3816 (N_3816,In_2044,In_1047);
nor U3817 (N_3817,In_2475,In_2486);
nor U3818 (N_3818,In_1980,In_3354);
nor U3819 (N_3819,In_3027,In_911);
nand U3820 (N_3820,In_4115,In_2920);
nor U3821 (N_3821,In_3655,In_578);
and U3822 (N_3822,In_2617,In_3846);
and U3823 (N_3823,In_806,In_2092);
nor U3824 (N_3824,In_337,In_2538);
xnor U3825 (N_3825,In_75,In_1314);
or U3826 (N_3826,In_1516,In_2350);
and U3827 (N_3827,In_1730,In_712);
nor U3828 (N_3828,In_3788,In_2128);
nor U3829 (N_3829,In_1252,In_2239);
xor U3830 (N_3830,In_1736,In_2251);
xnor U3831 (N_3831,In_287,In_3601);
or U3832 (N_3832,In_4117,In_2004);
nor U3833 (N_3833,In_4834,In_2682);
nor U3834 (N_3834,In_2262,In_1119);
nand U3835 (N_3835,In_2908,In_2199);
nor U3836 (N_3836,In_3777,In_4439);
nand U3837 (N_3837,In_2776,In_32);
nor U3838 (N_3838,In_537,In_1245);
nor U3839 (N_3839,In_1032,In_4421);
and U3840 (N_3840,In_1062,In_4116);
xnor U3841 (N_3841,In_2273,In_1750);
nand U3842 (N_3842,In_3993,In_1589);
nor U3843 (N_3843,In_1930,In_2700);
xor U3844 (N_3844,In_579,In_3292);
and U3845 (N_3845,In_3285,In_1778);
or U3846 (N_3846,In_1410,In_2992);
and U3847 (N_3847,In_3974,In_2446);
nand U3848 (N_3848,In_3545,In_2602);
xor U3849 (N_3849,In_226,In_976);
or U3850 (N_3850,In_1665,In_2585);
or U3851 (N_3851,In_4725,In_718);
xor U3852 (N_3852,In_4194,In_3021);
nor U3853 (N_3853,In_4126,In_1663);
and U3854 (N_3854,In_318,In_2391);
and U3855 (N_3855,In_4078,In_2689);
or U3856 (N_3856,In_3959,In_3884);
nor U3857 (N_3857,In_4029,In_3132);
nand U3858 (N_3858,In_1557,In_140);
nor U3859 (N_3859,In_4429,In_2991);
and U3860 (N_3860,In_2434,In_1955);
nor U3861 (N_3861,In_4040,In_3587);
xor U3862 (N_3862,In_4636,In_1063);
or U3863 (N_3863,In_3802,In_2865);
or U3864 (N_3864,In_340,In_4228);
xor U3865 (N_3865,In_4551,In_1579);
or U3866 (N_3866,In_4465,In_1139);
nand U3867 (N_3867,In_376,In_240);
nor U3868 (N_3868,In_1719,In_640);
nand U3869 (N_3869,In_3709,In_1331);
nand U3870 (N_3870,In_4188,In_45);
or U3871 (N_3871,In_2188,In_2806);
nand U3872 (N_3872,In_2864,In_2107);
nor U3873 (N_3873,In_2526,In_4464);
xnor U3874 (N_3874,In_2731,In_1313);
and U3875 (N_3875,In_2300,In_4650);
or U3876 (N_3876,In_775,In_3752);
xnor U3877 (N_3877,In_1343,In_1361);
and U3878 (N_3878,In_3203,In_2507);
nand U3879 (N_3879,In_3045,In_2559);
nand U3880 (N_3880,In_385,In_4560);
nand U3881 (N_3881,In_999,In_4671);
xnor U3882 (N_3882,In_1549,In_1281);
and U3883 (N_3883,In_1643,In_435);
and U3884 (N_3884,In_2830,In_3433);
xor U3885 (N_3885,In_1703,In_4031);
nand U3886 (N_3886,In_4908,In_2972);
and U3887 (N_3887,In_2578,In_3619);
xnor U3888 (N_3888,In_4926,In_1030);
and U3889 (N_3889,In_4426,In_967);
xnor U3890 (N_3890,In_4112,In_3250);
nor U3891 (N_3891,In_4625,In_3642);
xnor U3892 (N_3892,In_315,In_4719);
and U3893 (N_3893,In_3207,In_4562);
nand U3894 (N_3894,In_4711,In_3809);
or U3895 (N_3895,In_3460,In_4110);
nor U3896 (N_3896,In_4789,In_3241);
nand U3897 (N_3897,In_341,In_4316);
nor U3898 (N_3898,In_3301,In_2473);
nand U3899 (N_3899,In_58,In_4586);
xnor U3900 (N_3900,In_4854,In_4524);
and U3901 (N_3901,In_4071,In_55);
and U3902 (N_3902,In_4509,In_3746);
and U3903 (N_3903,In_907,In_309);
or U3904 (N_3904,In_4803,In_4580);
and U3905 (N_3905,In_904,In_2562);
nor U3906 (N_3906,In_1982,In_966);
nor U3907 (N_3907,In_4556,In_297);
nand U3908 (N_3908,In_2398,In_4704);
xnor U3909 (N_3909,In_1667,In_4182);
or U3910 (N_3910,In_4370,In_3341);
or U3911 (N_3911,In_2556,In_4146);
nand U3912 (N_3912,In_2364,In_4541);
and U3913 (N_3913,In_831,In_291);
and U3914 (N_3914,In_1660,In_3890);
and U3915 (N_3915,In_2451,In_3964);
and U3916 (N_3916,In_4206,In_1458);
and U3917 (N_3917,In_4203,In_4780);
xnor U3918 (N_3918,In_4981,In_1652);
nor U3919 (N_3919,In_3966,In_4891);
xor U3920 (N_3920,In_4981,In_2940);
xor U3921 (N_3921,In_435,In_2050);
nand U3922 (N_3922,In_3684,In_3751);
nand U3923 (N_3923,In_4389,In_4139);
nand U3924 (N_3924,In_1911,In_4578);
nand U3925 (N_3925,In_2175,In_4204);
nand U3926 (N_3926,In_4129,In_3104);
and U3927 (N_3927,In_1864,In_2767);
nor U3928 (N_3928,In_2492,In_1378);
or U3929 (N_3929,In_3448,In_3360);
or U3930 (N_3930,In_3481,In_1703);
or U3931 (N_3931,In_1963,In_3074);
or U3932 (N_3932,In_4676,In_2904);
xor U3933 (N_3933,In_296,In_4904);
xor U3934 (N_3934,In_3892,In_272);
xor U3935 (N_3935,In_962,In_1252);
or U3936 (N_3936,In_550,In_2009);
and U3937 (N_3937,In_724,In_903);
nor U3938 (N_3938,In_4214,In_1169);
xor U3939 (N_3939,In_887,In_1371);
xnor U3940 (N_3940,In_1108,In_1796);
and U3941 (N_3941,In_1996,In_2174);
or U3942 (N_3942,In_1189,In_1143);
xor U3943 (N_3943,In_339,In_2366);
nand U3944 (N_3944,In_997,In_3870);
nor U3945 (N_3945,In_793,In_2033);
nand U3946 (N_3946,In_2530,In_3077);
nor U3947 (N_3947,In_4742,In_2214);
nand U3948 (N_3948,In_2200,In_889);
xor U3949 (N_3949,In_4882,In_2356);
xor U3950 (N_3950,In_1432,In_3726);
nand U3951 (N_3951,In_4268,In_4123);
and U3952 (N_3952,In_732,In_2103);
nand U3953 (N_3953,In_3017,In_2910);
nor U3954 (N_3954,In_3223,In_1540);
and U3955 (N_3955,In_1366,In_2422);
nor U3956 (N_3956,In_2144,In_4563);
nand U3957 (N_3957,In_3745,In_421);
nand U3958 (N_3958,In_1840,In_4038);
nor U3959 (N_3959,In_2696,In_3062);
xor U3960 (N_3960,In_2212,In_1182);
and U3961 (N_3961,In_3656,In_3584);
nor U3962 (N_3962,In_796,In_3906);
xnor U3963 (N_3963,In_913,In_3707);
xnor U3964 (N_3964,In_4139,In_2190);
and U3965 (N_3965,In_1577,In_398);
nor U3966 (N_3966,In_4855,In_4532);
nor U3967 (N_3967,In_1971,In_1032);
xnor U3968 (N_3968,In_3925,In_2959);
nor U3969 (N_3969,In_39,In_1644);
nand U3970 (N_3970,In_4218,In_1526);
and U3971 (N_3971,In_3646,In_4415);
nand U3972 (N_3972,In_1858,In_414);
and U3973 (N_3973,In_1611,In_4124);
nor U3974 (N_3974,In_2388,In_1847);
nor U3975 (N_3975,In_654,In_1562);
or U3976 (N_3976,In_392,In_4396);
and U3977 (N_3977,In_3399,In_1926);
or U3978 (N_3978,In_3498,In_1753);
nand U3979 (N_3979,In_696,In_2419);
or U3980 (N_3980,In_1909,In_1218);
nor U3981 (N_3981,In_1693,In_103);
or U3982 (N_3982,In_2742,In_3231);
and U3983 (N_3983,In_1027,In_2583);
nor U3984 (N_3984,In_2931,In_1120);
or U3985 (N_3985,In_733,In_190);
nor U3986 (N_3986,In_247,In_2422);
xnor U3987 (N_3987,In_3492,In_3838);
nand U3988 (N_3988,In_768,In_2004);
and U3989 (N_3989,In_717,In_54);
and U3990 (N_3990,In_4733,In_92);
nor U3991 (N_3991,In_1703,In_3031);
and U3992 (N_3992,In_1033,In_3278);
nor U3993 (N_3993,In_1104,In_623);
xnor U3994 (N_3994,In_3514,In_775);
xor U3995 (N_3995,In_461,In_4980);
nor U3996 (N_3996,In_2517,In_2682);
or U3997 (N_3997,In_1514,In_3419);
nand U3998 (N_3998,In_1242,In_238);
nand U3999 (N_3999,In_3168,In_3876);
or U4000 (N_4000,In_967,In_2203);
xor U4001 (N_4001,In_4404,In_2253);
nor U4002 (N_4002,In_1952,In_4801);
and U4003 (N_4003,In_1832,In_3469);
or U4004 (N_4004,In_302,In_3281);
nor U4005 (N_4005,In_4085,In_3792);
and U4006 (N_4006,In_773,In_1489);
or U4007 (N_4007,In_4199,In_2407);
xor U4008 (N_4008,In_4152,In_279);
or U4009 (N_4009,In_773,In_498);
nand U4010 (N_4010,In_306,In_705);
or U4011 (N_4011,In_1725,In_1213);
and U4012 (N_4012,In_4589,In_2737);
nand U4013 (N_4013,In_3403,In_1127);
nor U4014 (N_4014,In_4256,In_2873);
nor U4015 (N_4015,In_844,In_2005);
nand U4016 (N_4016,In_3441,In_1328);
or U4017 (N_4017,In_207,In_3775);
nand U4018 (N_4018,In_1809,In_3499);
xor U4019 (N_4019,In_3911,In_1417);
or U4020 (N_4020,In_1611,In_1030);
nor U4021 (N_4021,In_1300,In_66);
nand U4022 (N_4022,In_4616,In_1660);
nand U4023 (N_4023,In_2868,In_1171);
nand U4024 (N_4024,In_2301,In_2262);
or U4025 (N_4025,In_1540,In_2712);
or U4026 (N_4026,In_2398,In_1747);
xor U4027 (N_4027,In_4244,In_4401);
and U4028 (N_4028,In_3961,In_1406);
nor U4029 (N_4029,In_3434,In_2538);
xnor U4030 (N_4030,In_1048,In_3718);
nor U4031 (N_4031,In_1039,In_485);
nand U4032 (N_4032,In_1379,In_774);
and U4033 (N_4033,In_3707,In_320);
and U4034 (N_4034,In_2322,In_1915);
nor U4035 (N_4035,In_2314,In_2939);
xnor U4036 (N_4036,In_2749,In_886);
or U4037 (N_4037,In_4843,In_410);
and U4038 (N_4038,In_4665,In_4852);
nor U4039 (N_4039,In_4444,In_3631);
or U4040 (N_4040,In_3198,In_892);
or U4041 (N_4041,In_3492,In_2091);
and U4042 (N_4042,In_3011,In_1070);
and U4043 (N_4043,In_239,In_3919);
nor U4044 (N_4044,In_3574,In_2712);
xnor U4045 (N_4045,In_262,In_1150);
xnor U4046 (N_4046,In_2603,In_3845);
nor U4047 (N_4047,In_2871,In_3268);
and U4048 (N_4048,In_587,In_1544);
nand U4049 (N_4049,In_1363,In_4206);
and U4050 (N_4050,In_482,In_1101);
nand U4051 (N_4051,In_871,In_3759);
nand U4052 (N_4052,In_1466,In_616);
nor U4053 (N_4053,In_306,In_3526);
and U4054 (N_4054,In_3393,In_449);
or U4055 (N_4055,In_707,In_2944);
or U4056 (N_4056,In_1891,In_3253);
xnor U4057 (N_4057,In_3627,In_205);
nor U4058 (N_4058,In_3297,In_633);
nor U4059 (N_4059,In_2458,In_1499);
nor U4060 (N_4060,In_1821,In_4720);
nor U4061 (N_4061,In_3393,In_4384);
or U4062 (N_4062,In_328,In_697);
or U4063 (N_4063,In_1118,In_48);
nand U4064 (N_4064,In_1598,In_4485);
and U4065 (N_4065,In_3732,In_3583);
nand U4066 (N_4066,In_945,In_4220);
or U4067 (N_4067,In_243,In_3672);
or U4068 (N_4068,In_4767,In_4116);
nand U4069 (N_4069,In_3192,In_4923);
and U4070 (N_4070,In_2484,In_605);
xnor U4071 (N_4071,In_4508,In_1346);
nor U4072 (N_4072,In_3341,In_3757);
or U4073 (N_4073,In_3606,In_4158);
or U4074 (N_4074,In_4593,In_1838);
and U4075 (N_4075,In_4347,In_1046);
nand U4076 (N_4076,In_3586,In_4716);
xnor U4077 (N_4077,In_3518,In_2354);
and U4078 (N_4078,In_2640,In_4482);
and U4079 (N_4079,In_907,In_3370);
nor U4080 (N_4080,In_2410,In_4695);
or U4081 (N_4081,In_2199,In_4028);
xor U4082 (N_4082,In_1738,In_2787);
or U4083 (N_4083,In_4594,In_4743);
or U4084 (N_4084,In_866,In_1926);
and U4085 (N_4085,In_1808,In_187);
or U4086 (N_4086,In_448,In_4369);
nor U4087 (N_4087,In_406,In_4026);
xor U4088 (N_4088,In_695,In_4506);
xor U4089 (N_4089,In_29,In_628);
or U4090 (N_4090,In_265,In_3102);
and U4091 (N_4091,In_2031,In_224);
nor U4092 (N_4092,In_4873,In_4993);
xor U4093 (N_4093,In_1520,In_3689);
nand U4094 (N_4094,In_840,In_3087);
and U4095 (N_4095,In_2972,In_2223);
xnor U4096 (N_4096,In_936,In_4051);
nand U4097 (N_4097,In_2541,In_1291);
xor U4098 (N_4098,In_2913,In_2750);
and U4099 (N_4099,In_2150,In_3347);
or U4100 (N_4100,In_4476,In_490);
nor U4101 (N_4101,In_243,In_3864);
and U4102 (N_4102,In_4165,In_54);
nand U4103 (N_4103,In_3157,In_2574);
xor U4104 (N_4104,In_4489,In_1470);
and U4105 (N_4105,In_2245,In_3280);
or U4106 (N_4106,In_509,In_2029);
nand U4107 (N_4107,In_1636,In_2283);
xor U4108 (N_4108,In_4403,In_2046);
xnor U4109 (N_4109,In_3061,In_228);
and U4110 (N_4110,In_3614,In_3606);
nor U4111 (N_4111,In_4808,In_1408);
nand U4112 (N_4112,In_2860,In_1376);
nor U4113 (N_4113,In_3,In_2312);
nor U4114 (N_4114,In_890,In_4477);
or U4115 (N_4115,In_3321,In_3419);
nand U4116 (N_4116,In_3901,In_4937);
or U4117 (N_4117,In_4078,In_582);
or U4118 (N_4118,In_2407,In_2506);
or U4119 (N_4119,In_311,In_2531);
or U4120 (N_4120,In_158,In_772);
nor U4121 (N_4121,In_4115,In_3006);
and U4122 (N_4122,In_780,In_1973);
or U4123 (N_4123,In_3369,In_4762);
nand U4124 (N_4124,In_1577,In_2631);
nand U4125 (N_4125,In_4588,In_2948);
xor U4126 (N_4126,In_4949,In_634);
and U4127 (N_4127,In_537,In_298);
nor U4128 (N_4128,In_4106,In_3017);
xnor U4129 (N_4129,In_3138,In_3156);
or U4130 (N_4130,In_1115,In_4674);
nor U4131 (N_4131,In_2789,In_4098);
or U4132 (N_4132,In_4771,In_649);
and U4133 (N_4133,In_2101,In_4555);
or U4134 (N_4134,In_916,In_4623);
and U4135 (N_4135,In_1507,In_1319);
and U4136 (N_4136,In_3117,In_930);
nor U4137 (N_4137,In_3779,In_3672);
nand U4138 (N_4138,In_1102,In_80);
xor U4139 (N_4139,In_2679,In_3392);
and U4140 (N_4140,In_801,In_2903);
xnor U4141 (N_4141,In_4426,In_4338);
or U4142 (N_4142,In_347,In_17);
and U4143 (N_4143,In_4540,In_261);
and U4144 (N_4144,In_1582,In_3329);
or U4145 (N_4145,In_2610,In_2263);
xor U4146 (N_4146,In_2215,In_4892);
xor U4147 (N_4147,In_4211,In_4571);
xnor U4148 (N_4148,In_413,In_431);
and U4149 (N_4149,In_3503,In_1844);
and U4150 (N_4150,In_4318,In_4989);
or U4151 (N_4151,In_1446,In_2859);
nand U4152 (N_4152,In_2171,In_2967);
nand U4153 (N_4153,In_1450,In_4947);
nand U4154 (N_4154,In_1273,In_1485);
and U4155 (N_4155,In_3530,In_3706);
nor U4156 (N_4156,In_3938,In_1095);
nor U4157 (N_4157,In_3615,In_1389);
nor U4158 (N_4158,In_2587,In_1252);
xor U4159 (N_4159,In_4652,In_3115);
and U4160 (N_4160,In_2026,In_501);
nand U4161 (N_4161,In_4614,In_4462);
nand U4162 (N_4162,In_632,In_4330);
nand U4163 (N_4163,In_3739,In_3792);
and U4164 (N_4164,In_515,In_585);
nand U4165 (N_4165,In_3721,In_2884);
or U4166 (N_4166,In_1090,In_646);
nand U4167 (N_4167,In_1231,In_3782);
or U4168 (N_4168,In_1338,In_3655);
xor U4169 (N_4169,In_1130,In_1713);
xor U4170 (N_4170,In_2613,In_886);
nor U4171 (N_4171,In_1443,In_881);
nor U4172 (N_4172,In_1277,In_2774);
nor U4173 (N_4173,In_836,In_48);
or U4174 (N_4174,In_3949,In_2061);
and U4175 (N_4175,In_1433,In_1241);
or U4176 (N_4176,In_1270,In_3262);
nand U4177 (N_4177,In_1807,In_401);
nand U4178 (N_4178,In_3340,In_3292);
nand U4179 (N_4179,In_360,In_4688);
nand U4180 (N_4180,In_552,In_2245);
nand U4181 (N_4181,In_4753,In_2275);
nor U4182 (N_4182,In_624,In_3285);
xnor U4183 (N_4183,In_3447,In_4768);
xor U4184 (N_4184,In_4734,In_143);
nand U4185 (N_4185,In_527,In_2616);
nor U4186 (N_4186,In_2227,In_4372);
or U4187 (N_4187,In_1254,In_561);
and U4188 (N_4188,In_2272,In_399);
nand U4189 (N_4189,In_665,In_1341);
nand U4190 (N_4190,In_3917,In_3402);
and U4191 (N_4191,In_32,In_4616);
and U4192 (N_4192,In_2151,In_1645);
nor U4193 (N_4193,In_4407,In_1444);
xor U4194 (N_4194,In_1338,In_4627);
or U4195 (N_4195,In_2562,In_2878);
and U4196 (N_4196,In_4605,In_2077);
and U4197 (N_4197,In_4960,In_2463);
nand U4198 (N_4198,In_3284,In_423);
nor U4199 (N_4199,In_329,In_3828);
and U4200 (N_4200,In_2788,In_3661);
xor U4201 (N_4201,In_873,In_4317);
nor U4202 (N_4202,In_1262,In_4390);
nor U4203 (N_4203,In_2955,In_1410);
and U4204 (N_4204,In_1448,In_3591);
nor U4205 (N_4205,In_3234,In_4533);
or U4206 (N_4206,In_2129,In_2255);
nand U4207 (N_4207,In_4238,In_371);
xnor U4208 (N_4208,In_2986,In_2842);
or U4209 (N_4209,In_1514,In_2110);
nand U4210 (N_4210,In_3224,In_738);
and U4211 (N_4211,In_800,In_4617);
xor U4212 (N_4212,In_135,In_2772);
nand U4213 (N_4213,In_2530,In_4559);
and U4214 (N_4214,In_3536,In_2331);
or U4215 (N_4215,In_733,In_3299);
nor U4216 (N_4216,In_4113,In_4537);
nand U4217 (N_4217,In_3795,In_3810);
nor U4218 (N_4218,In_1852,In_3238);
or U4219 (N_4219,In_2191,In_4279);
and U4220 (N_4220,In_549,In_2337);
and U4221 (N_4221,In_767,In_2321);
and U4222 (N_4222,In_1377,In_2869);
nand U4223 (N_4223,In_408,In_245);
nor U4224 (N_4224,In_3237,In_4138);
nor U4225 (N_4225,In_4625,In_2454);
nand U4226 (N_4226,In_2390,In_1425);
nor U4227 (N_4227,In_3297,In_1207);
xor U4228 (N_4228,In_1666,In_3620);
nor U4229 (N_4229,In_3118,In_528);
nor U4230 (N_4230,In_4097,In_2602);
nor U4231 (N_4231,In_1891,In_3080);
nor U4232 (N_4232,In_2693,In_1707);
nor U4233 (N_4233,In_560,In_4634);
and U4234 (N_4234,In_2936,In_679);
xnor U4235 (N_4235,In_4701,In_4529);
and U4236 (N_4236,In_1844,In_4522);
and U4237 (N_4237,In_3276,In_3288);
nand U4238 (N_4238,In_2671,In_3750);
xnor U4239 (N_4239,In_4469,In_2551);
or U4240 (N_4240,In_1398,In_2747);
nor U4241 (N_4241,In_2627,In_3494);
nor U4242 (N_4242,In_1445,In_2399);
and U4243 (N_4243,In_4725,In_4429);
or U4244 (N_4244,In_2998,In_3072);
nand U4245 (N_4245,In_3934,In_4150);
nand U4246 (N_4246,In_1537,In_4530);
nand U4247 (N_4247,In_630,In_2911);
nand U4248 (N_4248,In_533,In_2630);
and U4249 (N_4249,In_3089,In_2179);
or U4250 (N_4250,In_3383,In_4540);
and U4251 (N_4251,In_4544,In_3592);
nand U4252 (N_4252,In_2448,In_2708);
nor U4253 (N_4253,In_1077,In_1253);
or U4254 (N_4254,In_3254,In_2792);
xnor U4255 (N_4255,In_1997,In_4144);
xnor U4256 (N_4256,In_4950,In_4398);
or U4257 (N_4257,In_1098,In_4342);
or U4258 (N_4258,In_175,In_700);
and U4259 (N_4259,In_3396,In_73);
nand U4260 (N_4260,In_192,In_3589);
or U4261 (N_4261,In_2420,In_3312);
and U4262 (N_4262,In_4131,In_2237);
or U4263 (N_4263,In_951,In_1751);
nor U4264 (N_4264,In_1998,In_719);
nor U4265 (N_4265,In_609,In_4935);
xor U4266 (N_4266,In_4333,In_491);
or U4267 (N_4267,In_3783,In_2947);
xnor U4268 (N_4268,In_2345,In_1216);
or U4269 (N_4269,In_425,In_982);
or U4270 (N_4270,In_2309,In_1352);
nand U4271 (N_4271,In_604,In_4128);
nand U4272 (N_4272,In_4779,In_1618);
or U4273 (N_4273,In_4036,In_4302);
nor U4274 (N_4274,In_3283,In_601);
nand U4275 (N_4275,In_3022,In_2238);
and U4276 (N_4276,In_4493,In_858);
nor U4277 (N_4277,In_3666,In_4640);
and U4278 (N_4278,In_435,In_982);
nor U4279 (N_4279,In_1320,In_1122);
nor U4280 (N_4280,In_4792,In_1833);
xor U4281 (N_4281,In_147,In_4170);
or U4282 (N_4282,In_964,In_2763);
or U4283 (N_4283,In_1065,In_119);
and U4284 (N_4284,In_2092,In_3413);
and U4285 (N_4285,In_1521,In_4820);
nor U4286 (N_4286,In_985,In_1748);
xnor U4287 (N_4287,In_4708,In_1877);
and U4288 (N_4288,In_2259,In_947);
nand U4289 (N_4289,In_2752,In_1944);
and U4290 (N_4290,In_2184,In_3016);
nand U4291 (N_4291,In_441,In_459);
or U4292 (N_4292,In_1548,In_2530);
xor U4293 (N_4293,In_3448,In_3590);
nand U4294 (N_4294,In_488,In_3043);
nand U4295 (N_4295,In_4537,In_4232);
and U4296 (N_4296,In_3743,In_2085);
or U4297 (N_4297,In_2574,In_4911);
and U4298 (N_4298,In_876,In_101);
nand U4299 (N_4299,In_1068,In_4947);
or U4300 (N_4300,In_1061,In_4572);
nand U4301 (N_4301,In_483,In_2603);
or U4302 (N_4302,In_774,In_4180);
nand U4303 (N_4303,In_3436,In_3003);
and U4304 (N_4304,In_2680,In_765);
or U4305 (N_4305,In_1889,In_1234);
and U4306 (N_4306,In_934,In_1734);
or U4307 (N_4307,In_4324,In_1325);
or U4308 (N_4308,In_1550,In_613);
and U4309 (N_4309,In_1095,In_344);
xnor U4310 (N_4310,In_1265,In_1718);
nor U4311 (N_4311,In_2260,In_1093);
nor U4312 (N_4312,In_4830,In_268);
nand U4313 (N_4313,In_70,In_4925);
nor U4314 (N_4314,In_3365,In_2879);
nor U4315 (N_4315,In_1540,In_3065);
nor U4316 (N_4316,In_3834,In_4304);
nand U4317 (N_4317,In_2186,In_3167);
and U4318 (N_4318,In_1346,In_1994);
xor U4319 (N_4319,In_4888,In_3495);
or U4320 (N_4320,In_3129,In_2997);
nand U4321 (N_4321,In_4232,In_4525);
and U4322 (N_4322,In_2467,In_1);
nor U4323 (N_4323,In_3694,In_4628);
nor U4324 (N_4324,In_4928,In_2931);
or U4325 (N_4325,In_4274,In_111);
nor U4326 (N_4326,In_4942,In_4776);
or U4327 (N_4327,In_3064,In_3935);
and U4328 (N_4328,In_2935,In_2898);
xor U4329 (N_4329,In_3161,In_4607);
and U4330 (N_4330,In_4335,In_4658);
nor U4331 (N_4331,In_3521,In_1437);
and U4332 (N_4332,In_2843,In_3730);
and U4333 (N_4333,In_4976,In_1082);
nand U4334 (N_4334,In_2147,In_541);
nor U4335 (N_4335,In_1467,In_2154);
and U4336 (N_4336,In_810,In_3181);
and U4337 (N_4337,In_1392,In_419);
and U4338 (N_4338,In_2857,In_1062);
nor U4339 (N_4339,In_2747,In_3146);
or U4340 (N_4340,In_4965,In_2277);
xnor U4341 (N_4341,In_1215,In_4526);
xor U4342 (N_4342,In_4377,In_1747);
nand U4343 (N_4343,In_446,In_40);
xnor U4344 (N_4344,In_1788,In_3557);
and U4345 (N_4345,In_3329,In_754);
or U4346 (N_4346,In_1989,In_2180);
and U4347 (N_4347,In_1058,In_1245);
and U4348 (N_4348,In_680,In_297);
nand U4349 (N_4349,In_1466,In_4981);
nand U4350 (N_4350,In_3832,In_4449);
xor U4351 (N_4351,In_501,In_4807);
and U4352 (N_4352,In_1235,In_4047);
or U4353 (N_4353,In_212,In_4002);
and U4354 (N_4354,In_1448,In_1203);
xor U4355 (N_4355,In_4588,In_4109);
nand U4356 (N_4356,In_1414,In_4143);
and U4357 (N_4357,In_3831,In_2363);
xor U4358 (N_4358,In_4766,In_2772);
nor U4359 (N_4359,In_3571,In_1495);
nand U4360 (N_4360,In_4280,In_454);
xor U4361 (N_4361,In_1245,In_2306);
and U4362 (N_4362,In_3800,In_2157);
nand U4363 (N_4363,In_1365,In_3498);
xnor U4364 (N_4364,In_3964,In_918);
xor U4365 (N_4365,In_2268,In_3611);
xnor U4366 (N_4366,In_562,In_2977);
and U4367 (N_4367,In_4943,In_2559);
xnor U4368 (N_4368,In_2351,In_4873);
or U4369 (N_4369,In_4018,In_1416);
or U4370 (N_4370,In_2598,In_1627);
or U4371 (N_4371,In_4439,In_4842);
xor U4372 (N_4372,In_3312,In_2016);
nand U4373 (N_4373,In_3682,In_430);
and U4374 (N_4374,In_1715,In_3924);
xor U4375 (N_4375,In_4022,In_4495);
or U4376 (N_4376,In_703,In_4180);
nor U4377 (N_4377,In_2327,In_1771);
nor U4378 (N_4378,In_4624,In_4060);
nand U4379 (N_4379,In_3441,In_3669);
xor U4380 (N_4380,In_3335,In_4388);
xor U4381 (N_4381,In_1246,In_163);
and U4382 (N_4382,In_3797,In_3248);
nor U4383 (N_4383,In_1409,In_4107);
nand U4384 (N_4384,In_4930,In_3481);
and U4385 (N_4385,In_3143,In_245);
or U4386 (N_4386,In_666,In_2055);
xnor U4387 (N_4387,In_71,In_4895);
nor U4388 (N_4388,In_3196,In_4069);
xor U4389 (N_4389,In_3251,In_3970);
xnor U4390 (N_4390,In_99,In_3995);
nand U4391 (N_4391,In_930,In_2692);
nand U4392 (N_4392,In_1930,In_1124);
nor U4393 (N_4393,In_3882,In_4154);
xnor U4394 (N_4394,In_4964,In_2623);
or U4395 (N_4395,In_4004,In_3620);
xnor U4396 (N_4396,In_4863,In_4854);
xnor U4397 (N_4397,In_3468,In_4711);
xor U4398 (N_4398,In_1760,In_2242);
xnor U4399 (N_4399,In_3801,In_2741);
or U4400 (N_4400,In_2780,In_2974);
or U4401 (N_4401,In_2243,In_1053);
or U4402 (N_4402,In_1663,In_3167);
or U4403 (N_4403,In_1099,In_1569);
nor U4404 (N_4404,In_4460,In_1731);
and U4405 (N_4405,In_1000,In_209);
nor U4406 (N_4406,In_496,In_3568);
nor U4407 (N_4407,In_3673,In_4353);
and U4408 (N_4408,In_1542,In_2698);
nand U4409 (N_4409,In_2251,In_1194);
or U4410 (N_4410,In_2633,In_3738);
nor U4411 (N_4411,In_2018,In_1635);
xnor U4412 (N_4412,In_235,In_2120);
nand U4413 (N_4413,In_1254,In_2301);
nor U4414 (N_4414,In_2125,In_748);
or U4415 (N_4415,In_4836,In_174);
or U4416 (N_4416,In_1240,In_1012);
nand U4417 (N_4417,In_776,In_3652);
nand U4418 (N_4418,In_1640,In_4690);
xnor U4419 (N_4419,In_2764,In_3628);
nand U4420 (N_4420,In_2775,In_4152);
or U4421 (N_4421,In_2380,In_1788);
xor U4422 (N_4422,In_3139,In_4996);
xor U4423 (N_4423,In_226,In_942);
nand U4424 (N_4424,In_3441,In_4731);
nor U4425 (N_4425,In_3360,In_415);
xnor U4426 (N_4426,In_2478,In_2837);
nand U4427 (N_4427,In_4616,In_1031);
xnor U4428 (N_4428,In_4927,In_3612);
nand U4429 (N_4429,In_3531,In_1425);
or U4430 (N_4430,In_1727,In_2492);
and U4431 (N_4431,In_3707,In_3164);
xor U4432 (N_4432,In_1284,In_954);
or U4433 (N_4433,In_1339,In_3353);
nor U4434 (N_4434,In_363,In_2415);
or U4435 (N_4435,In_3952,In_2348);
and U4436 (N_4436,In_413,In_1980);
xnor U4437 (N_4437,In_4369,In_3905);
and U4438 (N_4438,In_4749,In_605);
xor U4439 (N_4439,In_4936,In_1712);
nand U4440 (N_4440,In_2157,In_2416);
nor U4441 (N_4441,In_2443,In_3656);
xnor U4442 (N_4442,In_651,In_997);
nor U4443 (N_4443,In_4305,In_958);
or U4444 (N_4444,In_1890,In_105);
nand U4445 (N_4445,In_1758,In_2949);
nor U4446 (N_4446,In_4869,In_4779);
nor U4447 (N_4447,In_2297,In_2205);
nand U4448 (N_4448,In_4483,In_1045);
or U4449 (N_4449,In_196,In_3135);
or U4450 (N_4450,In_3953,In_3133);
nand U4451 (N_4451,In_3235,In_4546);
or U4452 (N_4452,In_2970,In_1496);
or U4453 (N_4453,In_3200,In_1599);
or U4454 (N_4454,In_2020,In_1438);
nor U4455 (N_4455,In_434,In_117);
nor U4456 (N_4456,In_249,In_1943);
and U4457 (N_4457,In_1640,In_1618);
and U4458 (N_4458,In_2143,In_3877);
or U4459 (N_4459,In_4110,In_2201);
and U4460 (N_4460,In_153,In_2945);
nor U4461 (N_4461,In_2584,In_2240);
nand U4462 (N_4462,In_2338,In_4848);
nand U4463 (N_4463,In_1377,In_2707);
xor U4464 (N_4464,In_1697,In_3246);
or U4465 (N_4465,In_3521,In_2983);
or U4466 (N_4466,In_4640,In_4692);
nand U4467 (N_4467,In_2852,In_3261);
and U4468 (N_4468,In_2326,In_101);
and U4469 (N_4469,In_4361,In_4133);
nand U4470 (N_4470,In_4063,In_93);
nand U4471 (N_4471,In_4715,In_4798);
and U4472 (N_4472,In_1222,In_3639);
nor U4473 (N_4473,In_4399,In_3917);
or U4474 (N_4474,In_2908,In_2409);
nand U4475 (N_4475,In_3263,In_4430);
xnor U4476 (N_4476,In_1565,In_4464);
xor U4477 (N_4477,In_4458,In_2811);
xnor U4478 (N_4478,In_2576,In_3925);
nand U4479 (N_4479,In_3512,In_1101);
and U4480 (N_4480,In_3464,In_2053);
or U4481 (N_4481,In_2055,In_601);
and U4482 (N_4482,In_1260,In_4144);
xnor U4483 (N_4483,In_412,In_4352);
xor U4484 (N_4484,In_130,In_823);
or U4485 (N_4485,In_2627,In_713);
or U4486 (N_4486,In_1794,In_4832);
nor U4487 (N_4487,In_2584,In_3266);
nor U4488 (N_4488,In_3918,In_4318);
xnor U4489 (N_4489,In_4932,In_2245);
nand U4490 (N_4490,In_2666,In_1852);
xor U4491 (N_4491,In_1703,In_3901);
nand U4492 (N_4492,In_4992,In_1139);
nand U4493 (N_4493,In_3984,In_2691);
nor U4494 (N_4494,In_4489,In_1795);
or U4495 (N_4495,In_3178,In_4335);
nor U4496 (N_4496,In_1896,In_1942);
and U4497 (N_4497,In_1955,In_4574);
and U4498 (N_4498,In_1502,In_3348);
nand U4499 (N_4499,In_4140,In_4238);
nor U4500 (N_4500,In_352,In_4716);
nor U4501 (N_4501,In_3136,In_4756);
and U4502 (N_4502,In_285,In_131);
nor U4503 (N_4503,In_3713,In_204);
nand U4504 (N_4504,In_3357,In_1456);
and U4505 (N_4505,In_1308,In_3619);
and U4506 (N_4506,In_742,In_4067);
nor U4507 (N_4507,In_3033,In_3174);
xnor U4508 (N_4508,In_4395,In_366);
xnor U4509 (N_4509,In_3297,In_3537);
nor U4510 (N_4510,In_1299,In_2306);
or U4511 (N_4511,In_3087,In_2231);
and U4512 (N_4512,In_659,In_836);
nand U4513 (N_4513,In_2600,In_3545);
xor U4514 (N_4514,In_4402,In_4304);
or U4515 (N_4515,In_2337,In_2360);
nor U4516 (N_4516,In_1164,In_581);
nor U4517 (N_4517,In_2329,In_3172);
xor U4518 (N_4518,In_4480,In_176);
xnor U4519 (N_4519,In_1645,In_3995);
xor U4520 (N_4520,In_3785,In_199);
xnor U4521 (N_4521,In_4003,In_840);
xor U4522 (N_4522,In_3469,In_4383);
xnor U4523 (N_4523,In_1776,In_4905);
or U4524 (N_4524,In_2663,In_2427);
or U4525 (N_4525,In_4904,In_992);
nor U4526 (N_4526,In_3351,In_2954);
or U4527 (N_4527,In_1304,In_878);
and U4528 (N_4528,In_4952,In_4540);
or U4529 (N_4529,In_2082,In_2655);
and U4530 (N_4530,In_420,In_3832);
nor U4531 (N_4531,In_2344,In_708);
nor U4532 (N_4532,In_3156,In_3358);
xor U4533 (N_4533,In_1602,In_2198);
nor U4534 (N_4534,In_1400,In_1725);
and U4535 (N_4535,In_1018,In_57);
and U4536 (N_4536,In_4858,In_1635);
xor U4537 (N_4537,In_3557,In_3843);
xor U4538 (N_4538,In_4426,In_400);
and U4539 (N_4539,In_3611,In_3268);
or U4540 (N_4540,In_405,In_82);
and U4541 (N_4541,In_4517,In_1385);
nor U4542 (N_4542,In_4490,In_2407);
or U4543 (N_4543,In_1628,In_4534);
and U4544 (N_4544,In_168,In_2);
or U4545 (N_4545,In_2506,In_4040);
nand U4546 (N_4546,In_4322,In_4127);
nand U4547 (N_4547,In_3807,In_387);
nor U4548 (N_4548,In_4185,In_4924);
xnor U4549 (N_4549,In_3656,In_4937);
and U4550 (N_4550,In_4540,In_3057);
or U4551 (N_4551,In_2728,In_4470);
or U4552 (N_4552,In_1546,In_761);
nor U4553 (N_4553,In_4521,In_1917);
nand U4554 (N_4554,In_784,In_3247);
or U4555 (N_4555,In_615,In_1460);
or U4556 (N_4556,In_4671,In_3598);
or U4557 (N_4557,In_2427,In_3543);
nand U4558 (N_4558,In_2444,In_570);
or U4559 (N_4559,In_4665,In_3496);
nor U4560 (N_4560,In_2357,In_3671);
nor U4561 (N_4561,In_4654,In_1403);
xor U4562 (N_4562,In_3936,In_4350);
or U4563 (N_4563,In_2764,In_2478);
and U4564 (N_4564,In_2820,In_2109);
and U4565 (N_4565,In_1259,In_1613);
nor U4566 (N_4566,In_4474,In_4310);
nand U4567 (N_4567,In_2942,In_1900);
and U4568 (N_4568,In_2779,In_1093);
nor U4569 (N_4569,In_600,In_4937);
nor U4570 (N_4570,In_4211,In_1544);
nand U4571 (N_4571,In_1560,In_4541);
nor U4572 (N_4572,In_1490,In_1746);
nand U4573 (N_4573,In_4276,In_530);
nand U4574 (N_4574,In_1634,In_885);
or U4575 (N_4575,In_4000,In_226);
or U4576 (N_4576,In_1398,In_1319);
or U4577 (N_4577,In_2963,In_3548);
or U4578 (N_4578,In_2991,In_1583);
nor U4579 (N_4579,In_335,In_62);
xnor U4580 (N_4580,In_3408,In_1926);
nand U4581 (N_4581,In_3329,In_2945);
nor U4582 (N_4582,In_4213,In_1750);
or U4583 (N_4583,In_3150,In_4888);
nand U4584 (N_4584,In_3621,In_4259);
nor U4585 (N_4585,In_4803,In_3759);
xnor U4586 (N_4586,In_897,In_781);
and U4587 (N_4587,In_2496,In_2955);
and U4588 (N_4588,In_1453,In_20);
or U4589 (N_4589,In_2205,In_4286);
or U4590 (N_4590,In_860,In_4158);
xnor U4591 (N_4591,In_4945,In_1882);
xnor U4592 (N_4592,In_21,In_2656);
and U4593 (N_4593,In_3381,In_1335);
or U4594 (N_4594,In_1625,In_4602);
xnor U4595 (N_4595,In_404,In_3357);
xnor U4596 (N_4596,In_2503,In_831);
or U4597 (N_4597,In_3087,In_1112);
nor U4598 (N_4598,In_3709,In_1733);
and U4599 (N_4599,In_2938,In_3467);
xor U4600 (N_4600,In_4542,In_4853);
and U4601 (N_4601,In_929,In_412);
nor U4602 (N_4602,In_2983,In_3927);
and U4603 (N_4603,In_4418,In_4866);
nor U4604 (N_4604,In_2441,In_701);
nor U4605 (N_4605,In_2423,In_3641);
and U4606 (N_4606,In_2667,In_4527);
and U4607 (N_4607,In_4069,In_3555);
nor U4608 (N_4608,In_1741,In_3951);
nor U4609 (N_4609,In_4229,In_2365);
nor U4610 (N_4610,In_178,In_2155);
xnor U4611 (N_4611,In_4447,In_4233);
and U4612 (N_4612,In_438,In_1430);
or U4613 (N_4613,In_4470,In_4528);
or U4614 (N_4614,In_4039,In_1137);
and U4615 (N_4615,In_3525,In_4702);
nand U4616 (N_4616,In_2753,In_3049);
or U4617 (N_4617,In_4095,In_2604);
nor U4618 (N_4618,In_2044,In_2792);
and U4619 (N_4619,In_3793,In_1315);
nor U4620 (N_4620,In_4042,In_1716);
xnor U4621 (N_4621,In_4480,In_532);
xnor U4622 (N_4622,In_2123,In_1173);
xnor U4623 (N_4623,In_4265,In_2983);
nand U4624 (N_4624,In_2439,In_584);
and U4625 (N_4625,In_3203,In_670);
nand U4626 (N_4626,In_1997,In_3585);
xor U4627 (N_4627,In_3632,In_4783);
and U4628 (N_4628,In_4048,In_3585);
xor U4629 (N_4629,In_4331,In_4178);
nand U4630 (N_4630,In_352,In_4243);
or U4631 (N_4631,In_4474,In_1729);
xnor U4632 (N_4632,In_3735,In_2503);
xnor U4633 (N_4633,In_335,In_4841);
or U4634 (N_4634,In_3068,In_1420);
or U4635 (N_4635,In_4755,In_3885);
nor U4636 (N_4636,In_1167,In_4989);
or U4637 (N_4637,In_1766,In_1343);
nor U4638 (N_4638,In_1835,In_3421);
or U4639 (N_4639,In_174,In_2397);
or U4640 (N_4640,In_1122,In_4624);
nor U4641 (N_4641,In_1856,In_72);
xor U4642 (N_4642,In_4096,In_4793);
or U4643 (N_4643,In_3203,In_4676);
xor U4644 (N_4644,In_642,In_4505);
and U4645 (N_4645,In_3598,In_2042);
nor U4646 (N_4646,In_2036,In_3867);
or U4647 (N_4647,In_2424,In_2901);
nor U4648 (N_4648,In_1973,In_3771);
and U4649 (N_4649,In_1753,In_3232);
and U4650 (N_4650,In_61,In_4833);
and U4651 (N_4651,In_3753,In_1093);
and U4652 (N_4652,In_2706,In_434);
nor U4653 (N_4653,In_1527,In_2862);
xnor U4654 (N_4654,In_2161,In_353);
or U4655 (N_4655,In_14,In_3399);
and U4656 (N_4656,In_4688,In_1264);
nand U4657 (N_4657,In_3605,In_4473);
or U4658 (N_4658,In_721,In_853);
or U4659 (N_4659,In_1428,In_87);
nand U4660 (N_4660,In_56,In_569);
nand U4661 (N_4661,In_4894,In_3174);
and U4662 (N_4662,In_3380,In_790);
nor U4663 (N_4663,In_275,In_4193);
or U4664 (N_4664,In_867,In_4561);
xnor U4665 (N_4665,In_905,In_4754);
and U4666 (N_4666,In_800,In_1074);
or U4667 (N_4667,In_637,In_4759);
nor U4668 (N_4668,In_2404,In_3520);
and U4669 (N_4669,In_4325,In_1076);
nand U4670 (N_4670,In_3978,In_2593);
and U4671 (N_4671,In_1688,In_2308);
xnor U4672 (N_4672,In_2394,In_1329);
or U4673 (N_4673,In_1071,In_4863);
or U4674 (N_4674,In_3432,In_2932);
nor U4675 (N_4675,In_3668,In_2414);
or U4676 (N_4676,In_824,In_606);
and U4677 (N_4677,In_3203,In_2542);
or U4678 (N_4678,In_3347,In_3053);
nor U4679 (N_4679,In_2523,In_3328);
nor U4680 (N_4680,In_2158,In_2065);
and U4681 (N_4681,In_3600,In_859);
nand U4682 (N_4682,In_4786,In_3237);
nand U4683 (N_4683,In_3698,In_2262);
nand U4684 (N_4684,In_552,In_499);
nand U4685 (N_4685,In_4422,In_4048);
nand U4686 (N_4686,In_2499,In_410);
and U4687 (N_4687,In_256,In_4246);
or U4688 (N_4688,In_1294,In_2915);
nand U4689 (N_4689,In_3260,In_307);
xnor U4690 (N_4690,In_2586,In_760);
and U4691 (N_4691,In_2981,In_3014);
or U4692 (N_4692,In_1739,In_2169);
nand U4693 (N_4693,In_3798,In_4728);
or U4694 (N_4694,In_3852,In_4645);
xnor U4695 (N_4695,In_778,In_297);
and U4696 (N_4696,In_3609,In_1162);
nor U4697 (N_4697,In_438,In_1007);
xnor U4698 (N_4698,In_417,In_2415);
xor U4699 (N_4699,In_4065,In_1528);
and U4700 (N_4700,In_1672,In_1338);
or U4701 (N_4701,In_131,In_3621);
xor U4702 (N_4702,In_4037,In_2221);
xnor U4703 (N_4703,In_1587,In_2153);
or U4704 (N_4704,In_791,In_4982);
xor U4705 (N_4705,In_615,In_4500);
nor U4706 (N_4706,In_4120,In_278);
and U4707 (N_4707,In_4643,In_1955);
nand U4708 (N_4708,In_2214,In_2029);
xnor U4709 (N_4709,In_2512,In_3678);
xnor U4710 (N_4710,In_1531,In_479);
and U4711 (N_4711,In_4226,In_2656);
xnor U4712 (N_4712,In_2284,In_878);
xor U4713 (N_4713,In_3442,In_2571);
xor U4714 (N_4714,In_519,In_2764);
or U4715 (N_4715,In_3747,In_1029);
and U4716 (N_4716,In_981,In_1527);
nand U4717 (N_4717,In_2343,In_4037);
and U4718 (N_4718,In_4297,In_2010);
and U4719 (N_4719,In_729,In_2266);
and U4720 (N_4720,In_4556,In_4869);
or U4721 (N_4721,In_4149,In_2663);
or U4722 (N_4722,In_3172,In_2000);
nand U4723 (N_4723,In_114,In_3249);
or U4724 (N_4724,In_1536,In_1992);
xnor U4725 (N_4725,In_387,In_4139);
or U4726 (N_4726,In_722,In_3381);
xnor U4727 (N_4727,In_1569,In_4104);
xnor U4728 (N_4728,In_1801,In_3175);
nand U4729 (N_4729,In_2833,In_2345);
nor U4730 (N_4730,In_1193,In_87);
nor U4731 (N_4731,In_2590,In_4509);
xor U4732 (N_4732,In_46,In_4994);
or U4733 (N_4733,In_4307,In_721);
or U4734 (N_4734,In_2701,In_3298);
nor U4735 (N_4735,In_263,In_3306);
xnor U4736 (N_4736,In_3776,In_4931);
xor U4737 (N_4737,In_2734,In_688);
xnor U4738 (N_4738,In_1652,In_648);
nor U4739 (N_4739,In_531,In_2260);
nand U4740 (N_4740,In_1489,In_4537);
nor U4741 (N_4741,In_3445,In_1423);
nor U4742 (N_4742,In_2966,In_1800);
nand U4743 (N_4743,In_2334,In_3860);
and U4744 (N_4744,In_4035,In_1991);
nor U4745 (N_4745,In_2818,In_2826);
nor U4746 (N_4746,In_1196,In_1302);
xor U4747 (N_4747,In_3179,In_2300);
and U4748 (N_4748,In_1113,In_2127);
xor U4749 (N_4749,In_1584,In_3718);
nand U4750 (N_4750,In_3807,In_2905);
or U4751 (N_4751,In_4121,In_3192);
xnor U4752 (N_4752,In_3824,In_687);
nand U4753 (N_4753,In_717,In_3495);
or U4754 (N_4754,In_1488,In_631);
nor U4755 (N_4755,In_3048,In_3956);
nor U4756 (N_4756,In_4819,In_2892);
nand U4757 (N_4757,In_3862,In_2127);
nor U4758 (N_4758,In_1546,In_4709);
xnor U4759 (N_4759,In_2800,In_3470);
or U4760 (N_4760,In_2640,In_3160);
nor U4761 (N_4761,In_2485,In_2599);
xnor U4762 (N_4762,In_2666,In_4200);
xnor U4763 (N_4763,In_3267,In_2602);
nor U4764 (N_4764,In_826,In_2915);
or U4765 (N_4765,In_161,In_2385);
xnor U4766 (N_4766,In_985,In_1670);
xor U4767 (N_4767,In_4936,In_608);
nor U4768 (N_4768,In_2205,In_1172);
and U4769 (N_4769,In_2314,In_608);
nand U4770 (N_4770,In_4555,In_2987);
nor U4771 (N_4771,In_246,In_4900);
or U4772 (N_4772,In_2532,In_2979);
nor U4773 (N_4773,In_2396,In_1660);
nor U4774 (N_4774,In_795,In_4729);
xnor U4775 (N_4775,In_4512,In_2389);
xor U4776 (N_4776,In_3098,In_4593);
xnor U4777 (N_4777,In_1002,In_1018);
or U4778 (N_4778,In_2811,In_3953);
nand U4779 (N_4779,In_1008,In_765);
nand U4780 (N_4780,In_9,In_1348);
xor U4781 (N_4781,In_370,In_2244);
xnor U4782 (N_4782,In_75,In_1896);
nor U4783 (N_4783,In_586,In_4989);
and U4784 (N_4784,In_2478,In_483);
nand U4785 (N_4785,In_1555,In_2236);
xnor U4786 (N_4786,In_1350,In_2677);
xor U4787 (N_4787,In_1454,In_4066);
or U4788 (N_4788,In_3535,In_4601);
and U4789 (N_4789,In_1889,In_2756);
nor U4790 (N_4790,In_1365,In_3716);
nor U4791 (N_4791,In_2306,In_172);
nand U4792 (N_4792,In_4607,In_2782);
nor U4793 (N_4793,In_727,In_1286);
nor U4794 (N_4794,In_3324,In_2099);
nand U4795 (N_4795,In_4928,In_737);
or U4796 (N_4796,In_359,In_3779);
and U4797 (N_4797,In_2625,In_4376);
and U4798 (N_4798,In_2383,In_2860);
and U4799 (N_4799,In_3867,In_3949);
nor U4800 (N_4800,In_2308,In_3694);
and U4801 (N_4801,In_4181,In_2101);
nor U4802 (N_4802,In_3904,In_1274);
or U4803 (N_4803,In_2716,In_4144);
or U4804 (N_4804,In_1307,In_67);
or U4805 (N_4805,In_3754,In_1434);
and U4806 (N_4806,In_2089,In_2351);
or U4807 (N_4807,In_1744,In_100);
or U4808 (N_4808,In_1398,In_1884);
and U4809 (N_4809,In_3178,In_3672);
xor U4810 (N_4810,In_1903,In_4156);
nand U4811 (N_4811,In_173,In_2086);
or U4812 (N_4812,In_4044,In_4883);
nor U4813 (N_4813,In_4365,In_3955);
or U4814 (N_4814,In_2878,In_2152);
nand U4815 (N_4815,In_603,In_2356);
xnor U4816 (N_4816,In_2170,In_2477);
and U4817 (N_4817,In_4047,In_1149);
or U4818 (N_4818,In_3520,In_775);
xor U4819 (N_4819,In_3936,In_1535);
xor U4820 (N_4820,In_3494,In_2909);
and U4821 (N_4821,In_2773,In_378);
xor U4822 (N_4822,In_828,In_3860);
or U4823 (N_4823,In_1118,In_2176);
nand U4824 (N_4824,In_1077,In_1687);
xnor U4825 (N_4825,In_1725,In_1394);
xnor U4826 (N_4826,In_266,In_2530);
and U4827 (N_4827,In_2366,In_649);
nand U4828 (N_4828,In_705,In_1212);
and U4829 (N_4829,In_3450,In_4870);
and U4830 (N_4830,In_3691,In_445);
nand U4831 (N_4831,In_1427,In_1538);
nand U4832 (N_4832,In_3973,In_2132);
or U4833 (N_4833,In_1843,In_4963);
and U4834 (N_4834,In_4803,In_3405);
and U4835 (N_4835,In_1399,In_4558);
nor U4836 (N_4836,In_2931,In_4721);
xnor U4837 (N_4837,In_4686,In_851);
and U4838 (N_4838,In_3618,In_2585);
xor U4839 (N_4839,In_2802,In_4072);
or U4840 (N_4840,In_3347,In_1018);
nor U4841 (N_4841,In_337,In_2647);
xnor U4842 (N_4842,In_138,In_1089);
and U4843 (N_4843,In_368,In_1613);
and U4844 (N_4844,In_4170,In_2031);
and U4845 (N_4845,In_801,In_1121);
or U4846 (N_4846,In_32,In_3383);
nor U4847 (N_4847,In_2165,In_4284);
or U4848 (N_4848,In_4598,In_4402);
nand U4849 (N_4849,In_1175,In_4517);
xnor U4850 (N_4850,In_2813,In_4086);
or U4851 (N_4851,In_1430,In_2285);
or U4852 (N_4852,In_2904,In_4821);
nand U4853 (N_4853,In_2279,In_1367);
or U4854 (N_4854,In_3530,In_312);
or U4855 (N_4855,In_257,In_967);
or U4856 (N_4856,In_2546,In_817);
nand U4857 (N_4857,In_4975,In_740);
and U4858 (N_4858,In_3067,In_2738);
xor U4859 (N_4859,In_869,In_3432);
nor U4860 (N_4860,In_3568,In_3286);
and U4861 (N_4861,In_348,In_1969);
nand U4862 (N_4862,In_4468,In_1141);
and U4863 (N_4863,In_766,In_2165);
or U4864 (N_4864,In_3076,In_2640);
nand U4865 (N_4865,In_979,In_2416);
nor U4866 (N_4866,In_4254,In_2976);
xnor U4867 (N_4867,In_2648,In_1326);
nor U4868 (N_4868,In_1498,In_3641);
and U4869 (N_4869,In_651,In_850);
or U4870 (N_4870,In_1390,In_3485);
and U4871 (N_4871,In_1862,In_3775);
and U4872 (N_4872,In_1805,In_1968);
nand U4873 (N_4873,In_3808,In_906);
nor U4874 (N_4874,In_636,In_4322);
nand U4875 (N_4875,In_1399,In_198);
and U4876 (N_4876,In_2201,In_2076);
and U4877 (N_4877,In_819,In_1275);
nor U4878 (N_4878,In_1936,In_3963);
xor U4879 (N_4879,In_3502,In_1180);
or U4880 (N_4880,In_4858,In_2401);
nor U4881 (N_4881,In_4003,In_3915);
or U4882 (N_4882,In_18,In_1968);
nor U4883 (N_4883,In_1871,In_1935);
nor U4884 (N_4884,In_3550,In_4621);
nor U4885 (N_4885,In_2076,In_3727);
xnor U4886 (N_4886,In_1420,In_4869);
and U4887 (N_4887,In_4749,In_4982);
and U4888 (N_4888,In_1808,In_1869);
or U4889 (N_4889,In_2383,In_3120);
xnor U4890 (N_4890,In_1496,In_2412);
or U4891 (N_4891,In_325,In_2666);
or U4892 (N_4892,In_20,In_3758);
or U4893 (N_4893,In_729,In_315);
xnor U4894 (N_4894,In_4618,In_2839);
xnor U4895 (N_4895,In_4851,In_4535);
nand U4896 (N_4896,In_2612,In_1732);
or U4897 (N_4897,In_4216,In_3555);
and U4898 (N_4898,In_3114,In_3698);
nand U4899 (N_4899,In_4892,In_199);
nor U4900 (N_4900,In_2242,In_855);
and U4901 (N_4901,In_4510,In_1428);
xor U4902 (N_4902,In_2562,In_1859);
xor U4903 (N_4903,In_1203,In_2714);
and U4904 (N_4904,In_2405,In_1045);
nand U4905 (N_4905,In_4141,In_4368);
xnor U4906 (N_4906,In_3515,In_3024);
nor U4907 (N_4907,In_1980,In_2951);
xor U4908 (N_4908,In_79,In_2741);
or U4909 (N_4909,In_4022,In_3991);
or U4910 (N_4910,In_2672,In_4785);
xnor U4911 (N_4911,In_2618,In_1372);
nor U4912 (N_4912,In_1389,In_1099);
and U4913 (N_4913,In_3584,In_1316);
and U4914 (N_4914,In_1327,In_4107);
xor U4915 (N_4915,In_2240,In_3758);
xor U4916 (N_4916,In_2262,In_2991);
nor U4917 (N_4917,In_1491,In_328);
nand U4918 (N_4918,In_4188,In_4222);
or U4919 (N_4919,In_3506,In_3546);
xnor U4920 (N_4920,In_676,In_1190);
xnor U4921 (N_4921,In_3888,In_2759);
nor U4922 (N_4922,In_2734,In_2617);
or U4923 (N_4923,In_416,In_812);
nand U4924 (N_4924,In_3850,In_2807);
and U4925 (N_4925,In_1091,In_3043);
and U4926 (N_4926,In_2035,In_3226);
xor U4927 (N_4927,In_2508,In_3600);
nand U4928 (N_4928,In_1582,In_313);
xor U4929 (N_4929,In_4879,In_1282);
nor U4930 (N_4930,In_4936,In_2002);
nor U4931 (N_4931,In_4674,In_1723);
or U4932 (N_4932,In_3091,In_4345);
or U4933 (N_4933,In_3206,In_2499);
xor U4934 (N_4934,In_2851,In_2069);
nand U4935 (N_4935,In_4070,In_158);
or U4936 (N_4936,In_2314,In_1376);
and U4937 (N_4937,In_1795,In_4304);
xnor U4938 (N_4938,In_668,In_3869);
nand U4939 (N_4939,In_1427,In_91);
nor U4940 (N_4940,In_3313,In_801);
and U4941 (N_4941,In_4602,In_1780);
nor U4942 (N_4942,In_3018,In_1812);
nor U4943 (N_4943,In_4215,In_2398);
nor U4944 (N_4944,In_4288,In_1171);
or U4945 (N_4945,In_1107,In_1856);
or U4946 (N_4946,In_611,In_1840);
or U4947 (N_4947,In_1239,In_1087);
or U4948 (N_4948,In_917,In_541);
nor U4949 (N_4949,In_3566,In_1373);
or U4950 (N_4950,In_4332,In_4521);
and U4951 (N_4951,In_811,In_3186);
and U4952 (N_4952,In_3739,In_2905);
nand U4953 (N_4953,In_3598,In_3744);
nand U4954 (N_4954,In_1516,In_4033);
nor U4955 (N_4955,In_4404,In_295);
and U4956 (N_4956,In_4925,In_1024);
nand U4957 (N_4957,In_4657,In_2666);
or U4958 (N_4958,In_4154,In_2484);
nand U4959 (N_4959,In_3277,In_2182);
nor U4960 (N_4960,In_2952,In_2828);
nor U4961 (N_4961,In_1246,In_1774);
xnor U4962 (N_4962,In_2481,In_298);
nand U4963 (N_4963,In_4151,In_2987);
nor U4964 (N_4964,In_2184,In_3543);
or U4965 (N_4965,In_2562,In_3196);
or U4966 (N_4966,In_699,In_4118);
or U4967 (N_4967,In_2821,In_4896);
nor U4968 (N_4968,In_29,In_4990);
xor U4969 (N_4969,In_3020,In_3330);
nand U4970 (N_4970,In_4619,In_1752);
and U4971 (N_4971,In_4252,In_4373);
nor U4972 (N_4972,In_2762,In_4877);
and U4973 (N_4973,In_4992,In_563);
nor U4974 (N_4974,In_4175,In_4716);
nor U4975 (N_4975,In_2801,In_4076);
or U4976 (N_4976,In_1813,In_4389);
and U4977 (N_4977,In_310,In_1673);
nor U4978 (N_4978,In_3167,In_4266);
and U4979 (N_4979,In_3982,In_4794);
xnor U4980 (N_4980,In_4654,In_2303);
or U4981 (N_4981,In_302,In_2426);
nand U4982 (N_4982,In_1331,In_501);
or U4983 (N_4983,In_364,In_1730);
xnor U4984 (N_4984,In_2830,In_2413);
xor U4985 (N_4985,In_2431,In_2450);
and U4986 (N_4986,In_2758,In_4097);
or U4987 (N_4987,In_2436,In_2382);
and U4988 (N_4988,In_2716,In_2725);
nor U4989 (N_4989,In_4381,In_4047);
or U4990 (N_4990,In_3130,In_3270);
and U4991 (N_4991,In_3158,In_1155);
and U4992 (N_4992,In_2809,In_46);
and U4993 (N_4993,In_21,In_1410);
and U4994 (N_4994,In_850,In_1266);
nor U4995 (N_4995,In_4350,In_4920);
xor U4996 (N_4996,In_854,In_241);
xnor U4997 (N_4997,In_4959,In_2602);
or U4998 (N_4998,In_3210,In_3339);
nor U4999 (N_4999,In_2091,In_2503);
nor U5000 (N_5000,N_557,N_4173);
and U5001 (N_5001,N_1036,N_4707);
and U5002 (N_5002,N_865,N_4519);
xor U5003 (N_5003,N_24,N_818);
and U5004 (N_5004,N_4191,N_4846);
xor U5005 (N_5005,N_1331,N_4367);
nor U5006 (N_5006,N_3668,N_4652);
xor U5007 (N_5007,N_2155,N_1689);
xor U5008 (N_5008,N_3531,N_3122);
xnor U5009 (N_5009,N_2527,N_711);
or U5010 (N_5010,N_4650,N_3840);
nor U5011 (N_5011,N_4006,N_2048);
or U5012 (N_5012,N_2588,N_433);
nand U5013 (N_5013,N_4831,N_2000);
nand U5014 (N_5014,N_2774,N_184);
or U5015 (N_5015,N_498,N_61);
nor U5016 (N_5016,N_2376,N_802);
or U5017 (N_5017,N_1122,N_3113);
and U5018 (N_5018,N_3574,N_4234);
or U5019 (N_5019,N_3292,N_97);
or U5020 (N_5020,N_2154,N_218);
nand U5021 (N_5021,N_3946,N_3036);
and U5022 (N_5022,N_3791,N_1991);
and U5023 (N_5023,N_4794,N_4828);
or U5024 (N_5024,N_2882,N_1186);
or U5025 (N_5025,N_4597,N_1014);
nand U5026 (N_5026,N_4911,N_155);
xnor U5027 (N_5027,N_1451,N_3844);
nand U5028 (N_5028,N_4710,N_1504);
xor U5029 (N_5029,N_568,N_243);
nand U5030 (N_5030,N_3646,N_2615);
nor U5031 (N_5031,N_3331,N_2476);
and U5032 (N_5032,N_3701,N_2685);
xnor U5033 (N_5033,N_1264,N_1402);
nand U5034 (N_5034,N_3078,N_2092);
or U5035 (N_5035,N_4452,N_3811);
and U5036 (N_5036,N_4678,N_1116);
nor U5037 (N_5037,N_2178,N_1432);
or U5038 (N_5038,N_3814,N_2958);
nor U5039 (N_5039,N_2282,N_308);
or U5040 (N_5040,N_4222,N_3517);
xor U5041 (N_5041,N_4808,N_1230);
xnor U5042 (N_5042,N_245,N_593);
nor U5043 (N_5043,N_3854,N_3730);
or U5044 (N_5044,N_1425,N_266);
xor U5045 (N_5045,N_448,N_2466);
and U5046 (N_5046,N_1956,N_2254);
nand U5047 (N_5047,N_803,N_3971);
xnor U5048 (N_5048,N_378,N_4844);
nand U5049 (N_5049,N_2937,N_3549);
nor U5050 (N_5050,N_2801,N_3733);
and U5051 (N_5051,N_3296,N_3841);
and U5052 (N_5052,N_123,N_3679);
nor U5053 (N_5053,N_4259,N_4186);
xnor U5054 (N_5054,N_4172,N_2131);
nand U5055 (N_5055,N_586,N_1157);
xnor U5056 (N_5056,N_3399,N_1865);
and U5057 (N_5057,N_1517,N_875);
nor U5058 (N_5058,N_4915,N_2911);
and U5059 (N_5059,N_3110,N_496);
or U5060 (N_5060,N_4796,N_1180);
and U5061 (N_5061,N_4506,N_1453);
nor U5062 (N_5062,N_2499,N_4639);
nor U5063 (N_5063,N_473,N_2324);
xnor U5064 (N_5064,N_44,N_4033);
xnor U5065 (N_5065,N_856,N_4139);
nor U5066 (N_5066,N_1009,N_2360);
or U5067 (N_5067,N_828,N_3072);
nand U5068 (N_5068,N_1165,N_1692);
xnor U5069 (N_5069,N_3105,N_951);
or U5070 (N_5070,N_2136,N_3261);
xnor U5071 (N_5071,N_2301,N_1054);
nand U5072 (N_5072,N_3372,N_3076);
and U5073 (N_5073,N_1346,N_2142);
xor U5074 (N_5074,N_1761,N_3433);
xor U5075 (N_5075,N_1738,N_4963);
xor U5076 (N_5076,N_186,N_1273);
xnor U5077 (N_5077,N_2627,N_3691);
nand U5078 (N_5078,N_1840,N_1442);
nand U5079 (N_5079,N_3928,N_590);
and U5080 (N_5080,N_4739,N_4572);
nand U5081 (N_5081,N_1536,N_3907);
or U5082 (N_5082,N_4392,N_4932);
nor U5083 (N_5083,N_2590,N_1998);
nor U5084 (N_5084,N_1469,N_3991);
nor U5085 (N_5085,N_4228,N_2143);
xor U5086 (N_5086,N_3916,N_2658);
nor U5087 (N_5087,N_617,N_258);
or U5088 (N_5088,N_63,N_4495);
nor U5089 (N_5089,N_2032,N_226);
xor U5090 (N_5090,N_4985,N_3100);
xnor U5091 (N_5091,N_69,N_214);
nand U5092 (N_5092,N_1281,N_2646);
or U5093 (N_5093,N_2029,N_1155);
and U5094 (N_5094,N_2806,N_2374);
and U5095 (N_5095,N_1721,N_11);
or U5096 (N_5096,N_2846,N_3579);
and U5097 (N_5097,N_3282,N_4558);
xor U5098 (N_5098,N_4056,N_2756);
xnor U5099 (N_5099,N_3852,N_4032);
nor U5100 (N_5100,N_492,N_4196);
and U5101 (N_5101,N_3856,N_2043);
nor U5102 (N_5102,N_765,N_2200);
nand U5103 (N_5103,N_925,N_2830);
or U5104 (N_5104,N_2117,N_3047);
and U5105 (N_5105,N_4069,N_4353);
xor U5106 (N_5106,N_390,N_4675);
nand U5107 (N_5107,N_3809,N_1246);
nand U5108 (N_5108,N_1891,N_897);
and U5109 (N_5109,N_2183,N_2746);
xnor U5110 (N_5110,N_962,N_3103);
or U5111 (N_5111,N_3529,N_3826);
nand U5112 (N_5112,N_2648,N_1508);
nor U5113 (N_5113,N_2837,N_4670);
or U5114 (N_5114,N_4833,N_4061);
or U5115 (N_5115,N_1610,N_4178);
and U5116 (N_5116,N_1354,N_3473);
nand U5117 (N_5117,N_540,N_228);
nand U5118 (N_5118,N_4630,N_639);
nand U5119 (N_5119,N_2322,N_4555);
xor U5120 (N_5120,N_681,N_432);
nand U5121 (N_5121,N_1522,N_1377);
or U5122 (N_5122,N_2221,N_49);
and U5123 (N_5123,N_2034,N_1214);
nand U5124 (N_5124,N_505,N_3761);
nand U5125 (N_5125,N_1086,N_440);
xnor U5126 (N_5126,N_3125,N_1845);
nor U5127 (N_5127,N_3664,N_2577);
nor U5128 (N_5128,N_1183,N_2464);
or U5129 (N_5129,N_3242,N_2011);
nor U5130 (N_5130,N_107,N_230);
nand U5131 (N_5131,N_2775,N_934);
or U5132 (N_5132,N_121,N_1660);
xor U5133 (N_5133,N_2369,N_1549);
nand U5134 (N_5134,N_3756,N_1724);
xor U5135 (N_5135,N_2457,N_3917);
and U5136 (N_5136,N_4237,N_1128);
and U5137 (N_5137,N_2037,N_3158);
xor U5138 (N_5138,N_647,N_4637);
xor U5139 (N_5139,N_1756,N_2656);
or U5140 (N_5140,N_3894,N_4066);
nand U5141 (N_5141,N_2299,N_1555);
or U5142 (N_5142,N_2579,N_2556);
nand U5143 (N_5143,N_1781,N_457);
nand U5144 (N_5144,N_1048,N_1518);
xor U5145 (N_5145,N_1437,N_212);
and U5146 (N_5146,N_4854,N_796);
nand U5147 (N_5147,N_4102,N_4216);
xor U5148 (N_5148,N_221,N_2537);
or U5149 (N_5149,N_4753,N_1663);
and U5150 (N_5150,N_4593,N_1494);
xnor U5151 (N_5151,N_874,N_1050);
or U5152 (N_5152,N_452,N_3133);
nand U5153 (N_5153,N_4377,N_1816);
xnor U5154 (N_5154,N_78,N_2286);
or U5155 (N_5155,N_2562,N_2731);
and U5156 (N_5156,N_3313,N_3526);
and U5157 (N_5157,N_4774,N_156);
xor U5158 (N_5158,N_4357,N_3054);
xor U5159 (N_5159,N_4004,N_2148);
and U5160 (N_5160,N_4984,N_750);
nand U5161 (N_5161,N_2285,N_915);
nor U5162 (N_5162,N_2269,N_2581);
xnor U5163 (N_5163,N_2817,N_958);
nor U5164 (N_5164,N_1237,N_4460);
and U5165 (N_5165,N_4053,N_2245);
and U5166 (N_5166,N_628,N_3019);
or U5167 (N_5167,N_889,N_4028);
nand U5168 (N_5168,N_1232,N_598);
xor U5169 (N_5169,N_2660,N_734);
or U5170 (N_5170,N_1154,N_3376);
or U5171 (N_5171,N_4897,N_2015);
xor U5172 (N_5172,N_3532,N_3775);
nor U5173 (N_5173,N_858,N_3120);
or U5174 (N_5174,N_3497,N_1872);
nand U5175 (N_5175,N_137,N_592);
nand U5176 (N_5176,N_139,N_3471);
nand U5177 (N_5177,N_20,N_3798);
and U5178 (N_5178,N_4559,N_1678);
xor U5179 (N_5179,N_2554,N_3937);
nand U5180 (N_5180,N_2293,N_3196);
nand U5181 (N_5181,N_887,N_892);
nand U5182 (N_5182,N_3487,N_2314);
or U5183 (N_5183,N_251,N_1153);
or U5184 (N_5184,N_4628,N_1315);
nand U5185 (N_5185,N_607,N_3430);
nor U5186 (N_5186,N_4626,N_2838);
nor U5187 (N_5187,N_622,N_4777);
nand U5188 (N_5188,N_4496,N_1791);
xnor U5189 (N_5189,N_2758,N_1250);
and U5190 (N_5190,N_2544,N_3350);
nor U5191 (N_5191,N_2676,N_4594);
xnor U5192 (N_5192,N_1184,N_344);
xnor U5193 (N_5193,N_2983,N_3274);
or U5194 (N_5194,N_1045,N_1297);
and U5195 (N_5195,N_2428,N_2697);
xor U5196 (N_5196,N_166,N_1851);
nor U5197 (N_5197,N_4978,N_3851);
or U5198 (N_5198,N_4328,N_1160);
and U5199 (N_5199,N_3651,N_443);
nand U5200 (N_5200,N_4581,N_3454);
xnor U5201 (N_5201,N_2036,N_4604);
xnor U5202 (N_5202,N_1406,N_806);
nor U5203 (N_5203,N_2971,N_649);
and U5204 (N_5204,N_688,N_4406);
xnor U5205 (N_5205,N_1140,N_3882);
nand U5206 (N_5206,N_3432,N_1106);
or U5207 (N_5207,N_4603,N_2062);
and U5208 (N_5208,N_1899,N_1994);
and U5209 (N_5209,N_3106,N_2042);
nor U5210 (N_5210,N_2999,N_745);
nor U5211 (N_5211,N_1340,N_1194);
nand U5212 (N_5212,N_2759,N_4679);
nor U5213 (N_5213,N_3692,N_3822);
and U5214 (N_5214,N_1490,N_4202);
xnor U5215 (N_5215,N_2768,N_1105);
nor U5216 (N_5216,N_4624,N_4394);
and U5217 (N_5217,N_4454,N_2194);
and U5218 (N_5218,N_3051,N_3484);
nand U5219 (N_5219,N_3897,N_1870);
or U5220 (N_5220,N_4941,N_1362);
or U5221 (N_5221,N_4755,N_4413);
and U5222 (N_5222,N_4945,N_3802);
xnor U5223 (N_5223,N_1475,N_4812);
nand U5224 (N_5224,N_2952,N_4779);
and U5225 (N_5225,N_4068,N_2994);
xor U5226 (N_5226,N_2171,N_1668);
xor U5227 (N_5227,N_4302,N_2152);
nor U5228 (N_5228,N_846,N_778);
nor U5229 (N_5229,N_1553,N_4712);
nor U5230 (N_5230,N_4161,N_4760);
xor U5231 (N_5231,N_1719,N_2953);
xnor U5232 (N_5232,N_3860,N_793);
and U5233 (N_5233,N_1152,N_859);
nor U5234 (N_5234,N_198,N_1304);
nand U5235 (N_5235,N_2808,N_2001);
xnor U5236 (N_5236,N_888,N_585);
or U5237 (N_5237,N_89,N_1570);
nand U5238 (N_5238,N_2553,N_4967);
nor U5239 (N_5239,N_1016,N_2928);
nor U5240 (N_5240,N_4525,N_2929);
or U5241 (N_5241,N_736,N_286);
or U5242 (N_5242,N_197,N_4065);
nor U5243 (N_5243,N_4784,N_2392);
or U5244 (N_5244,N_4240,N_4210);
and U5245 (N_5245,N_1733,N_2265);
and U5246 (N_5246,N_1608,N_3002);
nor U5247 (N_5247,N_1546,N_3688);
and U5248 (N_5248,N_3396,N_4926);
nor U5249 (N_5249,N_1267,N_3348);
and U5250 (N_5250,N_1287,N_4343);
nand U5251 (N_5251,N_114,N_2606);
xnor U5252 (N_5252,N_972,N_3309);
nand U5253 (N_5253,N_1101,N_3778);
or U5254 (N_5254,N_2234,N_1953);
or U5255 (N_5255,N_471,N_784);
xor U5256 (N_5256,N_1768,N_444);
xor U5257 (N_5257,N_2365,N_968);
and U5258 (N_5258,N_2184,N_808);
and U5259 (N_5259,N_4633,N_461);
xnor U5260 (N_5260,N_4117,N_3429);
xor U5261 (N_5261,N_4332,N_2176);
nor U5262 (N_5262,N_562,N_1276);
nor U5263 (N_5263,N_578,N_2654);
nand U5264 (N_5264,N_1228,N_405);
xnor U5265 (N_5265,N_836,N_1333);
nor U5266 (N_5266,N_2302,N_2290);
and U5267 (N_5267,N_4175,N_4366);
or U5268 (N_5268,N_129,N_3575);
or U5269 (N_5269,N_2294,N_2744);
and U5270 (N_5270,N_1725,N_1713);
nor U5271 (N_5271,N_1334,N_1229);
and U5272 (N_5272,N_484,N_2752);
nor U5273 (N_5273,N_1973,N_4934);
xnor U5274 (N_5274,N_4313,N_1759);
xnor U5275 (N_5275,N_322,N_325);
nand U5276 (N_5276,N_975,N_795);
nor U5277 (N_5277,N_4584,N_1142);
and U5278 (N_5278,N_3335,N_2270);
xor U5279 (N_5279,N_1130,N_4194);
nor U5280 (N_5280,N_3792,N_3546);
or U5281 (N_5281,N_3315,N_3390);
nand U5282 (N_5282,N_2595,N_3751);
nand U5283 (N_5283,N_4310,N_2437);
nor U5284 (N_5284,N_559,N_4334);
nand U5285 (N_5285,N_1671,N_4086);
and U5286 (N_5286,N_1762,N_4998);
nor U5287 (N_5287,N_3255,N_4308);
xor U5288 (N_5288,N_294,N_3003);
or U5289 (N_5289,N_1951,N_3431);
xor U5290 (N_5290,N_2803,N_296);
nor U5291 (N_5291,N_2671,N_4950);
nor U5292 (N_5292,N_662,N_12);
xor U5293 (N_5293,N_4537,N_2607);
and U5294 (N_5294,N_3655,N_2120);
nor U5295 (N_5295,N_3702,N_1804);
nand U5296 (N_5296,N_928,N_1465);
nor U5297 (N_5297,N_3489,N_192);
and U5298 (N_5298,N_4108,N_922);
nor U5299 (N_5299,N_756,N_3164);
nand U5300 (N_5300,N_2690,N_3850);
xnor U5301 (N_5301,N_4255,N_1092);
nor U5302 (N_5302,N_2106,N_3147);
and U5303 (N_5303,N_1578,N_4213);
or U5304 (N_5304,N_3708,N_74);
and U5305 (N_5305,N_2565,N_2071);
nand U5306 (N_5306,N_1649,N_2777);
xnor U5307 (N_5307,N_2046,N_1421);
and U5308 (N_5308,N_2504,N_4094);
nor U5309 (N_5309,N_2339,N_395);
nor U5310 (N_5310,N_935,N_2101);
and U5311 (N_5311,N_4365,N_4641);
nor U5312 (N_5312,N_1676,N_1712);
nor U5313 (N_5313,N_2632,N_3115);
nor U5314 (N_5314,N_281,N_1974);
xnor U5315 (N_5315,N_954,N_4686);
or U5316 (N_5316,N_2764,N_664);
xnor U5317 (N_5317,N_914,N_1029);
and U5318 (N_5318,N_4577,N_389);
and U5319 (N_5319,N_1163,N_3556);
or U5320 (N_5320,N_2251,N_1193);
xnor U5321 (N_5321,N_35,N_4824);
nor U5322 (N_5322,N_3742,N_4080);
nor U5323 (N_5323,N_1710,N_2028);
nand U5324 (N_5324,N_4456,N_4329);
xnor U5325 (N_5325,N_345,N_3808);
or U5326 (N_5326,N_3447,N_1384);
xnor U5327 (N_5327,N_1038,N_3890);
or U5328 (N_5328,N_2433,N_1103);
xor U5329 (N_5329,N_1790,N_2730);
or U5330 (N_5330,N_2485,N_1877);
or U5331 (N_5331,N_826,N_3915);
and U5332 (N_5332,N_709,N_2385);
xnor U5333 (N_5333,N_2968,N_3270);
xor U5334 (N_5334,N_1200,N_430);
nand U5335 (N_5335,N_4426,N_3082);
xnor U5336 (N_5336,N_4793,N_886);
nor U5337 (N_5337,N_2298,N_321);
and U5338 (N_5338,N_1270,N_1728);
and U5339 (N_5339,N_257,N_1802);
or U5340 (N_5340,N_3061,N_3838);
nand U5341 (N_5341,N_4852,N_53);
or U5342 (N_5342,N_323,N_4867);
or U5343 (N_5343,N_1904,N_4813);
nor U5344 (N_5344,N_3176,N_2833);
or U5345 (N_5345,N_1351,N_3200);
xnor U5346 (N_5346,N_3277,N_4242);
nor U5347 (N_5347,N_1013,N_4600);
and U5348 (N_5348,N_1976,N_3983);
and U5349 (N_5349,N_392,N_1484);
and U5350 (N_5350,N_819,N_3703);
and U5351 (N_5351,N_1338,N_1814);
nor U5352 (N_5352,N_3178,N_1133);
and U5353 (N_5353,N_1164,N_2111);
nor U5354 (N_5354,N_1793,N_4997);
and U5355 (N_5355,N_2422,N_2508);
nand U5356 (N_5356,N_4326,N_3717);
xnor U5357 (N_5357,N_737,N_4295);
and U5358 (N_5358,N_632,N_39);
and U5359 (N_5359,N_3059,N_2289);
or U5360 (N_5360,N_2068,N_271);
nor U5361 (N_5361,N_1758,N_1558);
nand U5362 (N_5362,N_4049,N_3161);
or U5363 (N_5363,N_964,N_526);
or U5364 (N_5364,N_1702,N_490);
nor U5365 (N_5365,N_1380,N_3616);
nor U5366 (N_5366,N_2674,N_2076);
or U5367 (N_5367,N_3220,N_1970);
and U5368 (N_5368,N_3140,N_4084);
and U5369 (N_5369,N_1896,N_996);
and U5370 (N_5370,N_554,N_1808);
nor U5371 (N_5371,N_4076,N_1107);
and U5372 (N_5372,N_1809,N_1403);
nand U5373 (N_5373,N_1718,N_363);
and U5374 (N_5374,N_4912,N_3262);
xnor U5375 (N_5375,N_678,N_4817);
and U5376 (N_5376,N_986,N_2924);
or U5377 (N_5377,N_4333,N_1881);
nand U5378 (N_5378,N_3423,N_700);
xnor U5379 (N_5379,N_3344,N_3338);
or U5380 (N_5380,N_1329,N_413);
xnor U5381 (N_5381,N_1039,N_726);
nand U5382 (N_5382,N_2257,N_994);
nand U5383 (N_5383,N_515,N_614);
and U5384 (N_5384,N_725,N_4567);
nor U5385 (N_5385,N_2021,N_1084);
and U5386 (N_5386,N_2198,N_3229);
or U5387 (N_5387,N_147,N_3409);
or U5388 (N_5388,N_3896,N_288);
xnor U5389 (N_5389,N_1188,N_1168);
nor U5390 (N_5390,N_4657,N_2467);
or U5391 (N_5391,N_175,N_630);
and U5392 (N_5392,N_2356,N_3857);
and U5393 (N_5393,N_2005,N_3038);
nand U5394 (N_5394,N_3479,N_1875);
nand U5395 (N_5395,N_3676,N_2945);
nor U5396 (N_5396,N_1630,N_2018);
or U5397 (N_5397,N_3768,N_1044);
nand U5398 (N_5398,N_2341,N_1387);
nor U5399 (N_5399,N_182,N_3011);
xnor U5400 (N_5400,N_656,N_264);
xor U5401 (N_5401,N_4580,N_2491);
nor U5402 (N_5402,N_2506,N_2677);
nand U5403 (N_5403,N_1674,N_1028);
nor U5404 (N_5404,N_3823,N_1428);
or U5405 (N_5405,N_3018,N_982);
nor U5406 (N_5406,N_984,N_3921);
nor U5407 (N_5407,N_4721,N_4974);
or U5408 (N_5408,N_2226,N_3134);
or U5409 (N_5409,N_1765,N_4251);
and U5410 (N_5410,N_2920,N_355);
nor U5411 (N_5411,N_2943,N_4008);
and U5412 (N_5412,N_724,N_46);
and U5413 (N_5413,N_2426,N_4457);
and U5414 (N_5414,N_3264,N_3341);
nor U5415 (N_5415,N_879,N_838);
xnor U5416 (N_5416,N_1633,N_2168);
nor U5417 (N_5417,N_2698,N_1041);
xnor U5418 (N_5418,N_3652,N_4160);
nor U5419 (N_5419,N_4671,N_2104);
xor U5420 (N_5420,N_4583,N_4491);
or U5421 (N_5421,N_1182,N_4350);
nor U5422 (N_5422,N_1817,N_822);
nor U5423 (N_5423,N_3619,N_1089);
nor U5424 (N_5424,N_3478,N_967);
and U5425 (N_5425,N_259,N_2342);
xor U5426 (N_5426,N_219,N_2840);
nand U5427 (N_5427,N_2240,N_4680);
and U5428 (N_5428,N_1146,N_2586);
xor U5429 (N_5429,N_1900,N_2686);
or U5430 (N_5430,N_1008,N_4398);
and U5431 (N_5431,N_1627,N_4101);
and U5432 (N_5432,N_612,N_3293);
nand U5433 (N_5433,N_2798,N_616);
nor U5434 (N_5434,N_2088,N_2242);
or U5435 (N_5435,N_2644,N_1025);
nand U5436 (N_5436,N_1093,N_4223);
nand U5437 (N_5437,N_3040,N_343);
nand U5438 (N_5438,N_2860,N_3572);
and U5439 (N_5439,N_4247,N_2220);
or U5440 (N_5440,N_3360,N_3905);
and U5441 (N_5441,N_2057,N_4800);
nand U5442 (N_5442,N_3771,N_1265);
xor U5443 (N_5443,N_2721,N_3174);
and U5444 (N_5444,N_4384,N_2963);
nor U5445 (N_5445,N_2058,N_844);
and U5446 (N_5446,N_2310,N_3425);
and U5447 (N_5447,N_1280,N_375);
xnor U5448 (N_5448,N_4149,N_3680);
and U5449 (N_5449,N_3254,N_3669);
xor U5450 (N_5450,N_2053,N_661);
and U5451 (N_5451,N_3908,N_3126);
nor U5452 (N_5452,N_2597,N_476);
and U5453 (N_5453,N_1680,N_866);
nand U5454 (N_5454,N_1564,N_4942);
nor U5455 (N_5455,N_401,N_164);
or U5456 (N_5456,N_4248,N_791);
or U5457 (N_5457,N_545,N_451);
nor U5458 (N_5458,N_165,N_1511);
or U5459 (N_5459,N_1082,N_1400);
and U5460 (N_5460,N_4241,N_170);
and U5461 (N_5461,N_349,N_1113);
xnor U5462 (N_5462,N_172,N_2002);
nand U5463 (N_5463,N_2996,N_3820);
nor U5464 (N_5464,N_2091,N_87);
or U5465 (N_5465,N_2509,N_683);
nand U5466 (N_5466,N_648,N_4304);
or U5467 (N_5467,N_2657,N_3749);
and U5468 (N_5468,N_4522,N_775);
nand U5469 (N_5469,N_3551,N_85);
xor U5470 (N_5470,N_2720,N_2533);
or U5471 (N_5471,N_1496,N_3149);
xnor U5472 (N_5472,N_328,N_3193);
or U5473 (N_5473,N_2349,N_3605);
or U5474 (N_5474,N_1004,N_4072);
nor U5475 (N_5475,N_733,N_4528);
nand U5476 (N_5476,N_453,N_2571);
nand U5477 (N_5477,N_287,N_2742);
nor U5478 (N_5478,N_3525,N_3389);
xnor U5479 (N_5479,N_297,N_830);
and U5480 (N_5480,N_3678,N_1063);
nor U5481 (N_5481,N_3855,N_3900);
or U5482 (N_5482,N_3408,N_1109);
or U5483 (N_5483,N_14,N_1433);
nor U5484 (N_5484,N_4609,N_410);
and U5485 (N_5485,N_4427,N_3635);
nor U5486 (N_5486,N_1796,N_442);
or U5487 (N_5487,N_2747,N_3570);
nor U5488 (N_5488,N_2733,N_1512);
or U5489 (N_5489,N_3878,N_4669);
nand U5490 (N_5490,N_331,N_3281);
or U5491 (N_5491,N_4940,N_3179);
xnor U5492 (N_5492,N_2253,N_1788);
nand U5493 (N_5493,N_4981,N_977);
or U5494 (N_5494,N_2214,N_2839);
nand U5495 (N_5495,N_2275,N_4245);
nor U5496 (N_5496,N_1283,N_702);
nand U5497 (N_5497,N_4435,N_4048);
xor U5498 (N_5498,N_2141,N_2007);
xnor U5499 (N_5499,N_193,N_1730);
xnor U5500 (N_5500,N_3827,N_3612);
nor U5501 (N_5501,N_4441,N_2603);
nor U5502 (N_5502,N_961,N_907);
and U5503 (N_5503,N_2703,N_398);
nor U5504 (N_5504,N_1571,N_3436);
nand U5505 (N_5505,N_4147,N_3405);
or U5506 (N_5506,N_3464,N_521);
nor U5507 (N_5507,N_4047,N_240);
nor U5508 (N_5508,N_4836,N_1701);
or U5509 (N_5509,N_2244,N_3580);
xor U5510 (N_5510,N_1631,N_1523);
xor U5511 (N_5511,N_23,N_3114);
nor U5512 (N_5512,N_2395,N_1860);
nor U5513 (N_5513,N_3083,N_4075);
or U5514 (N_5514,N_1381,N_4214);
and U5515 (N_5515,N_4132,N_2804);
nor U5516 (N_5516,N_130,N_2982);
nand U5517 (N_5517,N_783,N_4005);
or U5518 (N_5518,N_311,N_761);
or U5519 (N_5519,N_1059,N_4839);
or U5520 (N_5520,N_4937,N_1061);
nor U5521 (N_5521,N_852,N_3163);
nor U5522 (N_5522,N_3636,N_2815);
or U5523 (N_5523,N_4122,N_2233);
or U5524 (N_5524,N_2948,N_2998);
nor U5525 (N_5525,N_1149,N_1108);
xor U5526 (N_5526,N_1736,N_1621);
xnor U5527 (N_5527,N_3729,N_3986);
or U5528 (N_5528,N_1753,N_4258);
or U5529 (N_5529,N_2450,N_1669);
or U5530 (N_5530,N_1260,N_905);
nand U5531 (N_5531,N_4416,N_3911);
or U5532 (N_5532,N_1841,N_1873);
and U5533 (N_5533,N_3225,N_3108);
and U5534 (N_5534,N_1483,N_4688);
or U5535 (N_5535,N_4995,N_3839);
and U5536 (N_5536,N_1205,N_707);
xor U5537 (N_5537,N_1887,N_2065);
xor U5538 (N_5538,N_3153,N_3034);
xnor U5539 (N_5539,N_3039,N_909);
and U5540 (N_5540,N_1474,N_2085);
xnor U5541 (N_5541,N_3523,N_4762);
or U5542 (N_5542,N_4772,N_3403);
and U5543 (N_5543,N_4003,N_4936);
nand U5544 (N_5544,N_1330,N_1986);
nand U5545 (N_5545,N_2633,N_1480);
or U5546 (N_5546,N_2067,N_3428);
nand U5547 (N_5547,N_890,N_2723);
nand U5548 (N_5548,N_4913,N_619);
or U5549 (N_5549,N_3177,N_3444);
or U5550 (N_5550,N_2981,N_3961);
and U5551 (N_5551,N_1749,N_183);
nand U5552 (N_5552,N_753,N_1445);
and U5553 (N_5553,N_3799,N_1407);
nand U5554 (N_5554,N_3330,N_4693);
or U5555 (N_5555,N_4757,N_849);
nand U5556 (N_5556,N_1468,N_4025);
or U5557 (N_5557,N_2386,N_2858);
or U5558 (N_5558,N_3861,N_4014);
nor U5559 (N_5559,N_4918,N_1923);
nand U5560 (N_5560,N_3610,N_387);
and U5561 (N_5561,N_1415,N_2879);
and U5562 (N_5562,N_2600,N_3303);
xor U5563 (N_5563,N_4756,N_4702);
nor U5564 (N_5564,N_3868,N_2122);
or U5565 (N_5565,N_3272,N_1497);
nor U5566 (N_5566,N_4070,N_3557);
nand U5567 (N_5567,N_1467,N_729);
nand U5568 (N_5568,N_232,N_369);
xor U5569 (N_5569,N_4159,N_2113);
nor U5570 (N_5570,N_877,N_3145);
nand U5571 (N_5571,N_2532,N_673);
nor U5572 (N_5572,N_2884,N_3629);
xor U5573 (N_5573,N_2225,N_1812);
nand U5574 (N_5574,N_2914,N_507);
xor U5575 (N_5575,N_1509,N_4919);
xnor U5576 (N_5576,N_4616,N_2139);
and U5577 (N_5577,N_3043,N_2619);
nor U5578 (N_5578,N_1015,N_2522);
and U5579 (N_5579,N_3789,N_2664);
nor U5580 (N_5580,N_695,N_3323);
and U5581 (N_5581,N_1889,N_2510);
and U5582 (N_5582,N_2083,N_1217);
nor U5583 (N_5583,N_4349,N_2714);
xor U5584 (N_5584,N_4021,N_936);
or U5585 (N_5585,N_1653,N_4602);
or U5586 (N_5586,N_4103,N_4994);
and U5587 (N_5587,N_3481,N_2695);
nand U5588 (N_5588,N_4461,N_2003);
xnor U5589 (N_5589,N_2126,N_4436);
nor U5590 (N_5590,N_3477,N_4440);
nand U5591 (N_5591,N_2947,N_1294);
and U5592 (N_5592,N_4582,N_1269);
and U5593 (N_5593,N_1062,N_4424);
nand U5594 (N_5594,N_3804,N_1962);
or U5595 (N_5595,N_3046,N_4564);
or U5596 (N_5596,N_4335,N_1477);
nor U5597 (N_5597,N_885,N_4783);
or U5598 (N_5598,N_845,N_3682);
nand U5599 (N_5599,N_863,N_2827);
or U5600 (N_5600,N_2099,N_3859);
or U5601 (N_5601,N_3661,N_4683);
or U5602 (N_5602,N_2757,N_589);
and U5603 (N_5603,N_4039,N_1458);
and U5604 (N_5604,N_1204,N_3965);
or U5605 (N_5605,N_1798,N_3324);
nor U5606 (N_5606,N_1622,N_4002);
and U5607 (N_5607,N_1492,N_3097);
and U5608 (N_5608,N_2792,N_2398);
or U5609 (N_5609,N_3263,N_1832);
or U5610 (N_5610,N_3332,N_2439);
nand U5611 (N_5611,N_1410,N_1639);
and U5612 (N_5612,N_333,N_1049);
nor U5613 (N_5613,N_3988,N_1784);
and U5614 (N_5614,N_3662,N_524);
xor U5615 (N_5615,N_2363,N_4162);
and U5616 (N_5616,N_923,N_4619);
and U5617 (N_5617,N_626,N_1472);
xor U5618 (N_5618,N_210,N_3440);
xnor U5619 (N_5619,N_1939,N_2078);
xnor U5620 (N_5620,N_4960,N_3006);
or U5621 (N_5621,N_3964,N_629);
or U5622 (N_5622,N_4991,N_1505);
and U5623 (N_5623,N_4078,N_4381);
and U5624 (N_5624,N_4548,N_1573);
xor U5625 (N_5625,N_4553,N_3116);
nand U5626 (N_5626,N_1166,N_1042);
and U5627 (N_5627,N_1958,N_640);
nor U5628 (N_5628,N_3345,N_916);
nor U5629 (N_5629,N_1828,N_161);
nor U5630 (N_5630,N_2688,N_1618);
nand U5631 (N_5631,N_2252,N_1769);
and U5632 (N_5632,N_2224,N_2138);
and U5633 (N_5633,N_3929,N_2334);
nor U5634 (N_5634,N_2539,N_3902);
or U5635 (N_5635,N_535,N_680);
nor U5636 (N_5636,N_3626,N_2869);
or U5637 (N_5637,N_4481,N_205);
nand U5638 (N_5638,N_2754,N_2631);
nand U5639 (N_5639,N_920,N_4488);
nor U5640 (N_5640,N_4588,N_1734);
xor U5641 (N_5641,N_2572,N_4442);
and U5642 (N_5642,N_3977,N_3973);
xor U5643 (N_5643,N_4336,N_1423);
xnor U5644 (N_5644,N_3025,N_4914);
nor U5645 (N_5645,N_2772,N_1539);
nand U5646 (N_5646,N_4674,N_2854);
and U5647 (N_5647,N_1302,N_2035);
nand U5648 (N_5648,N_2812,N_4818);
nor U5649 (N_5649,N_13,N_2512);
or U5650 (N_5650,N_279,N_974);
and U5651 (N_5651,N_1871,N_1772);
nor U5652 (N_5652,N_3638,N_3797);
nand U5653 (N_5653,N_215,N_1901);
and U5654 (N_5654,N_2760,N_4989);
xor U5655 (N_5655,N_4471,N_5);
nand U5656 (N_5656,N_1957,N_1910);
xnor U5657 (N_5657,N_1760,N_2347);
and U5658 (N_5658,N_2022,N_3815);
or U5659 (N_5659,N_4585,N_4087);
xor U5660 (N_5660,N_1905,N_2526);
or U5661 (N_5661,N_2816,N_382);
nor U5662 (N_5662,N_4309,N_2584);
and U5663 (N_5663,N_3275,N_4575);
xnor U5664 (N_5664,N_227,N_3284);
nor U5665 (N_5665,N_1336,N_1352);
nand U5666 (N_5666,N_1700,N_4699);
nand U5667 (N_5667,N_893,N_3130);
nand U5668 (N_5668,N_4150,N_4177);
nand U5669 (N_5669,N_6,N_832);
or U5670 (N_5670,N_815,N_1847);
nand U5671 (N_5671,N_261,N_2704);
nand U5672 (N_5672,N_1616,N_2327);
and U5673 (N_5673,N_4661,N_523);
xnor U5674 (N_5674,N_1548,N_3892);
or U5675 (N_5675,N_4330,N_4348);
xor U5676 (N_5676,N_3832,N_584);
and U5677 (N_5677,N_4323,N_2326);
or U5678 (N_5678,N_1394,N_3603);
nor U5679 (N_5679,N_4133,N_4835);
or U5680 (N_5680,N_327,N_2672);
and U5681 (N_5681,N_2895,N_4822);
or U5682 (N_5682,N_133,N_2623);
xnor U5683 (N_5683,N_4797,N_380);
nor U5684 (N_5684,N_4673,N_3456);
xor U5685 (N_5685,N_1358,N_2173);
nand U5686 (N_5686,N_549,N_4853);
xor U5687 (N_5687,N_2505,N_4763);
nand U5688 (N_5688,N_4340,N_1906);
xnor U5689 (N_5689,N_3598,N_103);
and U5690 (N_5690,N_2019,N_2832);
nand U5691 (N_5691,N_843,N_1742);
and U5692 (N_5692,N_3269,N_2370);
and U5693 (N_5693,N_1501,N_4395);
or U5694 (N_5694,N_4279,N_1882);
xnor U5695 (N_5695,N_4944,N_2559);
and U5696 (N_5696,N_2206,N_1586);
nor U5697 (N_5697,N_4776,N_2033);
and U5698 (N_5698,N_4676,N_4487);
xor U5699 (N_5699,N_1977,N_347);
or U5700 (N_5700,N_3364,N_2305);
xnor U5701 (N_5701,N_4141,N_1322);
nor U5702 (N_5702,N_1594,N_4608);
and U5703 (N_5703,N_2594,N_581);
xnor U5704 (N_5704,N_701,N_262);
nand U5705 (N_5705,N_1810,N_1919);
nand U5706 (N_5706,N_1173,N_3805);
xnor U5707 (N_5707,N_2933,N_1638);
xor U5708 (N_5708,N_1568,N_1739);
or U5709 (N_5709,N_1069,N_4019);
and U5710 (N_5710,N_1215,N_77);
xnor U5711 (N_5711,N_3930,N_1341);
nand U5712 (N_5712,N_2045,N_2044);
nand U5713 (N_5713,N_465,N_706);
nor U5714 (N_5714,N_3187,N_3418);
and U5715 (N_5715,N_4502,N_313);
and U5716 (N_5716,N_927,N_4894);
nor U5717 (N_5717,N_1481,N_1975);
or U5718 (N_5718,N_2972,N_4081);
and U5719 (N_5719,N_950,N_3352);
and U5720 (N_5720,N_2566,N_1751);
xor U5721 (N_5721,N_3813,N_1470);
and U5722 (N_5722,N_1514,N_2484);
nand U5723 (N_5723,N_4654,N_3340);
xor U5724 (N_5724,N_1988,N_1567);
xnor U5725 (N_5725,N_931,N_2075);
or U5726 (N_5726,N_4857,N_134);
nand U5727 (N_5727,N_4771,N_563);
or U5728 (N_5728,N_3342,N_666);
nor U5729 (N_5729,N_4337,N_3217);
nor U5730 (N_5730,N_4238,N_4034);
nor U5731 (N_5731,N_1181,N_786);
nor U5732 (N_5732,N_4475,N_1783);
and U5733 (N_5733,N_4317,N_4727);
or U5734 (N_5734,N_3234,N_3351);
nor U5735 (N_5735,N_213,N_2103);
nor U5736 (N_5736,N_2247,N_878);
and U5737 (N_5737,N_394,N_1210);
nor U5738 (N_5738,N_2828,N_4042);
nor U5739 (N_5739,N_3087,N_3942);
nand U5740 (N_5740,N_3210,N_2014);
xor U5741 (N_5741,N_4751,N_4352);
nor U5742 (N_5742,N_4870,N_4606);
nor U5743 (N_5743,N_68,N_1880);
nor U5744 (N_5744,N_3439,N_3258);
xor U5745 (N_5745,N_1827,N_4546);
or U5746 (N_5746,N_1544,N_1370);
nand U5747 (N_5747,N_4832,N_3978);
nand U5748 (N_5748,N_3188,N_995);
nand U5749 (N_5749,N_1818,N_2824);
or U5750 (N_5750,N_1767,N_663);
nor U5751 (N_5751,N_3144,N_4050);
or U5752 (N_5752,N_4468,N_4244);
nor U5753 (N_5753,N_3452,N_1000);
nor U5754 (N_5754,N_4315,N_2406);
nand U5755 (N_5755,N_3643,N_4773);
xor U5756 (N_5756,N_60,N_3035);
nor U5757 (N_5757,N_4470,N_3185);
and U5758 (N_5758,N_4390,N_3673);
or U5759 (N_5759,N_4736,N_997);
nand U5760 (N_5760,N_1686,N_145);
and U5761 (N_5761,N_117,N_4570);
or U5762 (N_5762,N_1617,N_4542);
xor U5763 (N_5763,N_4166,N_3166);
nor U5764 (N_5764,N_1386,N_386);
nor U5765 (N_5765,N_1968,N_787);
and U5766 (N_5766,N_4379,N_906);
or U5767 (N_5767,N_1876,N_263);
or U5768 (N_5768,N_1677,N_4096);
nand U5769 (N_5769,N_2930,N_3068);
nand U5770 (N_5770,N_3694,N_2343);
nor U5771 (N_5771,N_3491,N_1489);
nand U5772 (N_5772,N_4855,N_3972);
nor U5773 (N_5773,N_3128,N_3091);
xnor U5774 (N_5774,N_4955,N_472);
nand U5775 (N_5775,N_2931,N_3312);
nand U5776 (N_5776,N_4987,N_3760);
nor U5777 (N_5777,N_2694,N_2668);
or U5778 (N_5778,N_2535,N_2552);
nand U5779 (N_5779,N_1158,N_3180);
nand U5780 (N_5780,N_1572,N_1615);
or U5781 (N_5781,N_4587,N_1197);
xor U5782 (N_5782,N_1950,N_3622);
nand U5783 (N_5783,N_4283,N_3448);
nor U5784 (N_5784,N_2222,N_2417);
or U5785 (N_5785,N_1455,N_536);
nand U5786 (N_5786,N_1757,N_167);
nand U5787 (N_5787,N_3710,N_3573);
nor U5788 (N_5788,N_1850,N_4562);
or U5789 (N_5789,N_759,N_4882);
nor U5790 (N_5790,N_603,N_3918);
nand U5791 (N_5791,N_2427,N_2098);
xor U5792 (N_5792,N_1826,N_2430);
or U5793 (N_5793,N_2908,N_1611);
and U5794 (N_5794,N_30,N_2902);
xor U5795 (N_5795,N_40,N_4477);
and U5796 (N_5796,N_4499,N_2236);
nand U5797 (N_5797,N_2330,N_1797);
nor U5798 (N_5798,N_19,N_3830);
or U5799 (N_5799,N_190,N_3457);
xor U5800 (N_5800,N_2538,N_3232);
and U5801 (N_5801,N_2229,N_4717);
nor U5802 (N_5802,N_3548,N_3739);
nor U5803 (N_5803,N_307,N_2250);
nor U5804 (N_5804,N_2217,N_3438);
nor U5805 (N_5805,N_2487,N_3631);
nand U5806 (N_5806,N_15,N_4199);
and U5807 (N_5807,N_2010,N_2307);
xor U5808 (N_5808,N_1820,N_3512);
nor U5809 (N_5809,N_357,N_2789);
or U5810 (N_5810,N_1782,N_776);
xor U5811 (N_5811,N_3948,N_1345);
and U5812 (N_5812,N_1506,N_2276);
xnor U5813 (N_5813,N_1174,N_2555);
nor U5814 (N_5814,N_3831,N_1949);
xor U5815 (N_5815,N_4925,N_3578);
nor U5816 (N_5816,N_4909,N_2950);
and U5817 (N_5817,N_1679,N_1556);
or U5818 (N_5818,N_642,N_4734);
xor U5819 (N_5819,N_1427,N_1414);
and U5820 (N_5820,N_949,N_1777);
or U5821 (N_5821,N_3211,N_2446);
or U5822 (N_5822,N_3520,N_1211);
nor U5823 (N_5823,N_1419,N_3154);
nor U5824 (N_5824,N_1159,N_4549);
nand U5825 (N_5825,N_1516,N_106);
and U5826 (N_5826,N_1792,N_81);
xor U5827 (N_5827,N_2818,N_4803);
nand U5828 (N_5828,N_1533,N_4207);
xor U5829 (N_5829,N_3544,N_1030);
nand U5830 (N_5830,N_4666,N_1268);
nand U5831 (N_5831,N_4264,N_3092);
and U5832 (N_5832,N_4962,N_2192);
or U5833 (N_5833,N_3783,N_54);
nor U5834 (N_5834,N_4689,N_4089);
and U5835 (N_5835,N_3647,N_3283);
nand U5836 (N_5836,N_4623,N_2258);
nor U5837 (N_5837,N_1922,N_1390);
nand U5838 (N_5838,N_3996,N_1207);
xor U5839 (N_5839,N_1227,N_4467);
nand U5840 (N_5840,N_3848,N_1112);
nor U5841 (N_5841,N_2156,N_2604);
nor U5842 (N_5842,N_336,N_834);
nand U5843 (N_5843,N_2241,N_4363);
nand U5844 (N_5844,N_3417,N_1459);
xor U5845 (N_5845,N_3697,N_3496);
xor U5846 (N_5846,N_2311,N_1837);
nor U5847 (N_5847,N_1614,N_613);
xor U5848 (N_5848,N_4770,N_1347);
nor U5849 (N_5849,N_1503,N_4910);
or U5850 (N_5850,N_4312,N_3715);
nand U5851 (N_5851,N_2608,N_1684);
xor U5852 (N_5852,N_4151,N_4625);
or U5853 (N_5853,N_1737,N_98);
nor U5854 (N_5854,N_1085,N_4507);
or U5855 (N_5855,N_973,N_391);
or U5856 (N_5856,N_1253,N_2593);
and U5857 (N_5857,N_4599,N_4119);
nand U5858 (N_5858,N_3773,N_3609);
nand U5859 (N_5859,N_2905,N_963);
or U5860 (N_5860,N_952,N_2069);
nor U5861 (N_5861,N_824,N_422);
and U5862 (N_5862,N_3334,N_4785);
and U5863 (N_5863,N_4827,N_2502);
and U5864 (N_5864,N_4814,N_500);
nand U5865 (N_5865,N_570,N_2536);
and U5866 (N_5866,N_3474,N_3536);
xor U5867 (N_5867,N_506,N_2170);
nor U5868 (N_5868,N_4374,N_2112);
and U5869 (N_5869,N_154,N_2149);
nor U5870 (N_5870,N_3155,N_1697);
xnor U5871 (N_5871,N_3297,N_4908);
xor U5872 (N_5872,N_1127,N_1895);
nand U5873 (N_5873,N_110,N_4115);
or U5874 (N_5874,N_55,N_4620);
and U5875 (N_5875,N_4646,N_2199);
nor U5876 (N_5876,N_3592,N_871);
nor U5877 (N_5877,N_4540,N_933);
xor U5878 (N_5878,N_2191,N_4866);
and U5879 (N_5879,N_2712,N_1732);
or U5880 (N_5880,N_4359,N_3480);
nor U5881 (N_5881,N_246,N_1396);
nor U5882 (N_5882,N_3310,N_3984);
xor U5883 (N_5883,N_2959,N_4498);
and U5884 (N_5884,N_4062,N_1);
or U5885 (N_5885,N_3563,N_1708);
and U5886 (N_5886,N_4841,N_517);
xnor U5887 (N_5887,N_4948,N_1431);
nand U5888 (N_5888,N_195,N_3793);
nor U5889 (N_5889,N_4124,N_3062);
nand U5890 (N_5890,N_811,N_4165);
nand U5891 (N_5891,N_3325,N_4863);
nor U5892 (N_5892,N_2647,N_4215);
and U5893 (N_5893,N_2891,N_2684);
and U5894 (N_5894,N_1731,N_2472);
nor U5895 (N_5895,N_1424,N_1744);
or U5896 (N_5896,N_3042,N_2115);
or U5897 (N_5897,N_3182,N_2709);
xor U5898 (N_5898,N_2637,N_1011);
nand U5899 (N_5899,N_2743,N_4226);
xnor U5900 (N_5900,N_3649,N_3004);
nor U5901 (N_5901,N_250,N_2197);
nor U5902 (N_5902,N_2970,N_2162);
or U5903 (N_5903,N_2412,N_741);
nand U5904 (N_5904,N_1766,N_1695);
and U5905 (N_5905,N_1046,N_4322);
nand U5906 (N_5906,N_4750,N_379);
nor U5907 (N_5907,N_487,N_2873);
or U5908 (N_5908,N_3732,N_329);
nand U5909 (N_5909,N_1981,N_3367);
and U5910 (N_5910,N_728,N_3414);
xnor U5911 (N_5911,N_1435,N_857);
nor U5912 (N_5912,N_3306,N_2926);
nor U5913 (N_5913,N_2049,N_3181);
nand U5914 (N_5914,N_917,N_4276);
nor U5915 (N_5915,N_436,N_2380);
and U5916 (N_5916,N_4380,N_1972);
or U5917 (N_5917,N_3540,N_2006);
and U5918 (N_5918,N_2008,N_2788);
nor U5919 (N_5919,N_3607,N_2889);
nor U5920 (N_5920,N_708,N_1226);
and U5921 (N_5921,N_4903,N_3932);
or U5922 (N_5922,N_2421,N_3402);
nor U5923 (N_5923,N_3898,N_418);
or U5924 (N_5924,N_1743,N_419);
nand U5925 (N_5925,N_4074,N_4692);
xnor U5926 (N_5926,N_3800,N_872);
xor U5927 (N_5927,N_4726,N_3589);
or U5928 (N_5928,N_2316,N_774);
and U5929 (N_5929,N_2403,N_3564);
xor U5930 (N_5930,N_4085,N_1935);
nand U5931 (N_5931,N_1078,N_3194);
nand U5932 (N_5932,N_3267,N_1420);
nand U5933 (N_5933,N_1928,N_122);
nand U5934 (N_5934,N_751,N_1787);
and U5935 (N_5935,N_131,N_2488);
xor U5936 (N_5936,N_577,N_3190);
xnor U5937 (N_5937,N_1110,N_4057);
and U5938 (N_5938,N_2345,N_346);
and U5939 (N_5939,N_1067,N_3041);
xnor U5940 (N_5940,N_4167,N_1554);
xnor U5941 (N_5941,N_4209,N_2462);
xor U5942 (N_5942,N_1694,N_2040);
nor U5943 (N_5943,N_4146,N_3770);
and U5944 (N_5944,N_3201,N_1825);
nand U5945 (N_5945,N_4968,N_4052);
or U5946 (N_5946,N_1717,N_2628);
or U5947 (N_5947,N_4752,N_4425);
nand U5948 (N_5948,N_4060,N_1239);
nand U5949 (N_5949,N_4429,N_3659);
nor U5950 (N_5950,N_2469,N_3245);
nor U5951 (N_5951,N_4786,N_2292);
nand U5952 (N_5952,N_2665,N_3801);
nand U5953 (N_5953,N_4382,N_1286);
nand U5954 (N_5954,N_2093,N_2780);
nand U5955 (N_5955,N_426,N_3118);
and U5956 (N_5956,N_851,N_3974);
nor U5957 (N_5957,N_804,N_2012);
or U5958 (N_5958,N_3660,N_4883);
or U5959 (N_5959,N_2503,N_2303);
nor U5960 (N_5960,N_4345,N_3666);
nor U5961 (N_5961,N_3391,N_3127);
and U5962 (N_5962,N_4408,N_1399);
and U5963 (N_5963,N_1959,N_1852);
or U5964 (N_5964,N_2492,N_4082);
nand U5965 (N_5965,N_2906,N_72);
nand U5966 (N_5966,N_2471,N_359);
xnor U5967 (N_5967,N_1911,N_142);
or U5968 (N_5968,N_533,N_2157);
and U5969 (N_5969,N_3321,N_3316);
xnor U5970 (N_5970,N_3533,N_3080);
nand U5971 (N_5971,N_2119,N_2901);
and U5972 (N_5972,N_1206,N_2262);
and U5973 (N_5973,N_2315,N_4969);
nor U5974 (N_5974,N_2907,N_3818);
xnor U5975 (N_5975,N_4607,N_4865);
xnor U5976 (N_5976,N_850,N_861);
nor U5977 (N_5977,N_2892,N_4996);
or U5978 (N_5978,N_1866,N_3542);
xnor U5979 (N_5979,N_3959,N_1599);
xor U5980 (N_5980,N_3371,N_1491);
xnor U5981 (N_5981,N_1350,N_3713);
nor U5982 (N_5982,N_943,N_3681);
nor U5983 (N_5983,N_2867,N_2651);
or U5984 (N_5984,N_4116,N_4531);
nand U5985 (N_5985,N_3449,N_674);
or U5986 (N_5986,N_3023,N_489);
nor U5987 (N_5987,N_3075,N_3960);
or U5988 (N_5988,N_4318,N_4282);
xor U5989 (N_5989,N_1969,N_2267);
xor U5990 (N_5990,N_3248,N_4051);
and U5991 (N_5991,N_687,N_894);
nand U5992 (N_5992,N_2397,N_1869);
and U5993 (N_5993,N_764,N_1813);
and U5994 (N_5994,N_1931,N_1774);
or U5995 (N_5995,N_4206,N_4598);
xnor U5996 (N_5996,N_4230,N_2762);
and U5997 (N_5997,N_3990,N_2284);
xor U5998 (N_5998,N_4437,N_3952);
xnor U5999 (N_5999,N_2587,N_4965);
and U6000 (N_6000,N_1833,N_2463);
and U6001 (N_6001,N_3876,N_1299);
nor U6002 (N_6002,N_4046,N_2494);
nand U6003 (N_6003,N_1685,N_276);
nor U6004 (N_6004,N_2209,N_2496);
and U6005 (N_6005,N_1829,N_2611);
nor U6006 (N_6006,N_488,N_602);
or U6007 (N_6007,N_1655,N_2211);
and U6008 (N_6008,N_4685,N_4221);
and U6009 (N_6009,N_4513,N_2849);
xnor U6010 (N_6010,N_4677,N_1897);
nand U6011 (N_6011,N_2480,N_3286);
nor U6012 (N_6012,N_4530,N_1007);
xor U6013 (N_6013,N_2483,N_265);
nand U6014 (N_6014,N_4509,N_4362);
nand U6015 (N_6015,N_300,N_1047);
and U6016 (N_6016,N_3628,N_4538);
or U6017 (N_6017,N_3238,N_573);
and U6018 (N_6018,N_4232,N_2204);
nand U6019 (N_6019,N_4725,N_740);
nor U6020 (N_6020,N_1926,N_1830);
xnor U6021 (N_6021,N_2456,N_1416);
or U6022 (N_6022,N_2728,N_2216);
nand U6023 (N_6023,N_3690,N_4645);
or U6024 (N_6024,N_3535,N_4949);
and U6025 (N_6025,N_16,N_4231);
or U6026 (N_6026,N_966,N_2338);
nor U6027 (N_6027,N_284,N_2771);
or U6028 (N_6028,N_3380,N_310);
or U6029 (N_6029,N_3369,N_236);
xnor U6030 (N_6030,N_2373,N_3828);
nand U6031 (N_6031,N_2350,N_2084);
xor U6032 (N_6032,N_1507,N_1510);
xor U6033 (N_6033,N_4389,N_3785);
nor U6034 (N_6034,N_1404,N_2897);
nor U6035 (N_6035,N_2378,N_754);
or U6036 (N_6036,N_1914,N_1017);
xor U6037 (N_6037,N_1275,N_1918);
xnor U6038 (N_6038,N_3927,N_368);
xor U6039 (N_6039,N_2560,N_17);
or U6040 (N_6040,N_2108,N_1378);
nor U6041 (N_6041,N_1740,N_4111);
and U6042 (N_6042,N_4975,N_2087);
or U6043 (N_6043,N_2451,N_4983);
nor U6044 (N_6044,N_3381,N_2814);
xnor U6045 (N_6045,N_4711,N_1393);
and U6046 (N_6046,N_4142,N_999);
xnor U6047 (N_6047,N_314,N_3081);
nor U6048 (N_6048,N_2235,N_4700);
nand U6049 (N_6049,N_722,N_3606);
or U6050 (N_6050,N_2734,N_1290);
and U6051 (N_6051,N_3304,N_2279);
or U6052 (N_6052,N_4480,N_2642);
and U6053 (N_6053,N_1907,N_651);
xor U6054 (N_6054,N_2853,N_3466);
and U6055 (N_6055,N_1095,N_3096);
xnor U6056 (N_6056,N_4720,N_393);
or U6057 (N_6057,N_1690,N_3098);
xor U6058 (N_6058,N_3485,N_3554);
nand U6059 (N_6059,N_4140,N_4512);
or U6060 (N_6060,N_1902,N_486);
nor U6061 (N_6061,N_1999,N_4174);
or U6062 (N_6062,N_1208,N_3333);
xnor U6063 (N_6063,N_2102,N_4899);
nor U6064 (N_6064,N_3862,N_324);
nand U6065 (N_6065,N_2582,N_278);
and U6066 (N_6066,N_2352,N_2601);
nand U6067 (N_6067,N_4289,N_3849);
and U6068 (N_6068,N_316,N_1530);
nor U6069 (N_6069,N_2741,N_1650);
nand U6070 (N_6070,N_4261,N_638);
and U6071 (N_6071,N_4730,N_3494);
and U6072 (N_6072,N_2249,N_2570);
and U6073 (N_6073,N_1831,N_3975);
nor U6074 (N_6074,N_2617,N_3784);
nand U6075 (N_6075,N_196,N_56);
xor U6076 (N_6076,N_2161,N_870);
xor U6077 (N_6077,N_115,N_4973);
and U6078 (N_6078,N_3853,N_4500);
nand U6079 (N_6079,N_2181,N_978);
xnor U6080 (N_6080,N_285,N_773);
nand U6081 (N_6081,N_686,N_1703);
or U6082 (N_6082,N_2189,N_1482);
and U6083 (N_6083,N_2361,N_2576);
nand U6084 (N_6084,N_116,N_2459);
nor U6085 (N_6085,N_4433,N_4270);
and U6086 (N_6086,N_1715,N_3737);
nand U6087 (N_6087,N_1243,N_2266);
or U6088 (N_6088,N_4268,N_1937);
xor U6089 (N_6089,N_677,N_2016);
xnor U6090 (N_6090,N_3596,N_1526);
and U6091 (N_6091,N_2569,N_2915);
nor U6092 (N_6092,N_2243,N_2864);
nor U6093 (N_6093,N_862,N_407);
or U6094 (N_6094,N_454,N_2313);
nand U6095 (N_6095,N_356,N_28);
or U6096 (N_6096,N_1222,N_4446);
nor U6097 (N_6097,N_2652,N_4494);
nand U6098 (N_6098,N_3671,N_4378);
nor U6099 (N_6099,N_3642,N_2271);
or U6100 (N_6100,N_3538,N_3980);
nor U6101 (N_6101,N_4419,N_339);
and U6102 (N_6102,N_4552,N_2137);
nor U6103 (N_6103,N_4288,N_2561);
nand U6104 (N_6104,N_384,N_3);
and U6105 (N_6105,N_229,N_4492);
nand U6106 (N_6106,N_1196,N_2531);
nand U6107 (N_6107,N_82,N_1920);
xor U6108 (N_6108,N_1342,N_727);
nor U6109 (N_6109,N_148,N_367);
nor U6110 (N_6110,N_953,N_2936);
and U6111 (N_6111,N_1328,N_3287);
nand U6112 (N_6112,N_2309,N_1199);
and U6113 (N_6113,N_199,N_3198);
nor U6114 (N_6114,N_29,N_2724);
or U6115 (N_6115,N_3204,N_1537);
nor U6116 (N_6116,N_2726,N_4595);
nand U6117 (N_6117,N_1723,N_1261);
and U6118 (N_6118,N_1051,N_4183);
nand U6119 (N_6119,N_3550,N_2977);
and U6120 (N_6120,N_3320,N_3318);
or U6121 (N_6121,N_4892,N_235);
or U6122 (N_6122,N_3522,N_2614);
xnor U6123 (N_6123,N_4099,N_3486);
or U6124 (N_6124,N_4106,N_3621);
xor U6125 (N_6125,N_597,N_3233);
and U6126 (N_6126,N_1461,N_4956);
and U6127 (N_6127,N_1426,N_2669);
xor U6128 (N_6128,N_2419,N_1943);
and U6129 (N_6129,N_691,N_2169);
nor U6130 (N_6130,N_3780,N_1980);
or U6131 (N_6131,N_1141,N_2662);
nor U6132 (N_6132,N_2910,N_508);
nor U6133 (N_6133,N_2185,N_2052);
and U6134 (N_6134,N_2423,N_2813);
nor U6135 (N_6135,N_2434,N_2272);
nor U6136 (N_6136,N_3891,N_976);
and U6137 (N_6137,N_2739,N_4529);
or U6138 (N_6138,N_2399,N_721);
or U6139 (N_6139,N_1248,N_1037);
xnor U6140 (N_6140,N_3562,N_720);
and U6141 (N_6141,N_4407,N_153);
or U6142 (N_6142,N_1285,N_2799);
xnor U6143 (N_6143,N_3374,N_3510);
nor U6144 (N_6144,N_2086,N_1316);
or U6145 (N_6145,N_3314,N_4163);
xor U6146 (N_6146,N_2918,N_3723);
and U6147 (N_6147,N_2766,N_217);
and U6148 (N_6148,N_204,N_3375);
nand U6149 (N_6149,N_2215,N_4601);
nand U6150 (N_6150,N_2585,N_241);
or U6151 (N_6151,N_4009,N_3615);
nor U6152 (N_6152,N_1659,N_4071);
and U6153 (N_6153,N_3027,N_2878);
nand U6154 (N_6154,N_3397,N_779);
nand U6155 (N_6155,N_3384,N_3104);
and U6156 (N_6156,N_2969,N_4490);
and U6157 (N_6157,N_3625,N_4029);
nor U6158 (N_6158,N_4267,N_4935);
xnor U6159 (N_6159,N_2418,N_4667);
or U6160 (N_6160,N_1538,N_2900);
nor U6161 (N_6161,N_1683,N_4023);
nand U6162 (N_6162,N_3301,N_1696);
nor U6163 (N_6163,N_2212,N_1349);
and U6164 (N_6164,N_3872,N_247);
and U6165 (N_6165,N_544,N_2549);
and U6166 (N_6166,N_4256,N_4463);
nor U6167 (N_6167,N_1309,N_2455);
nor U6168 (N_6168,N_3591,N_1704);
nor U6169 (N_6169,N_2454,N_4861);
xor U6170 (N_6170,N_4517,N_2541);
or U6171 (N_6171,N_4153,N_3280);
xnor U6172 (N_6172,N_1598,N_2641);
or U6173 (N_6173,N_3171,N_3593);
nand U6174 (N_6174,N_548,N_4791);
nand U6175 (N_6175,N_3191,N_940);
and U6176 (N_6176,N_1666,N_2118);
nor U6177 (N_6177,N_817,N_3093);
and U6178 (N_6178,N_414,N_1187);
xnor U6179 (N_6179,N_634,N_3604);
and U6180 (N_6180,N_2404,N_1241);
nand U6181 (N_6181,N_2366,N_2885);
or U6182 (N_6182,N_4521,N_938);
nor U6183 (N_6183,N_3790,N_3307);
nand U6184 (N_6184,N_4778,N_3720);
and U6185 (N_6185,N_234,N_1031);
xnor U6186 (N_6186,N_1589,N_644);
and U6187 (N_6187,N_2921,N_574);
and U6188 (N_6188,N_4649,N_3936);
nor U6189 (N_6189,N_1376,N_2004);
and U6190 (N_6190,N_439,N_99);
nand U6191 (N_6191,N_2966,N_4249);
nor U6192 (N_6192,N_2797,N_2308);
and U6193 (N_6193,N_1520,N_2534);
nor U6194 (N_6194,N_2382,N_1306);
nand U6195 (N_6195,N_4274,N_3246);
nand U6196 (N_6196,N_3005,N_1185);
nor U6197 (N_6197,N_4574,N_174);
or U6198 (N_6198,N_1323,N_2708);
and U6199 (N_6199,N_1498,N_2995);
or U6200 (N_6200,N_4354,N_4455);
xor U6201 (N_6201,N_2218,N_2109);
and U6202 (N_6202,N_3945,N_37);
and U6203 (N_6203,N_3914,N_2328);
and U6204 (N_6204,N_4532,N_2865);
nor U6205 (N_6205,N_3385,N_2940);
xor U6206 (N_6206,N_4660,N_3968);
and U6207 (N_6207,N_22,N_2655);
or U6208 (N_6208,N_411,N_2643);
xor U6209 (N_6209,N_2107,N_1835);
xor U6210 (N_6210,N_3235,N_342);
xor U6211 (N_6211,N_330,N_2055);
nor U6212 (N_6212,N_2700,N_4383);
xnor U6213 (N_6213,N_109,N_4044);
nor U6214 (N_6214,N_2128,N_3803);
nor U6215 (N_6215,N_4795,N_1529);
nand U6216 (N_6216,N_206,N_3585);
nor U6217 (N_6217,N_558,N_427);
or U6218 (N_6218,N_2785,N_1308);
xor U6219 (N_6219,N_3530,N_4181);
nand U6220 (N_6220,N_4358,N_4466);
and U6221 (N_6221,N_3387,N_3634);
and U6222 (N_6222,N_4372,N_2375);
or U6223 (N_6223,N_1440,N_1010);
nand U6224 (N_6224,N_1858,N_2530);
nand U6225 (N_6225,N_4902,N_67);
nand U6226 (N_6226,N_2898,N_25);
nand U6227 (N_6227,N_3215,N_4758);
and U6228 (N_6228,N_146,N_4527);
nand U6229 (N_6229,N_2097,N_3252);
and U6230 (N_6230,N_1240,N_4735);
nor U6231 (N_6231,N_1780,N_4107);
nor U6232 (N_6232,N_3955,N_1531);
nand U6233 (N_6233,N_3146,N_1576);
or U6234 (N_6234,N_4007,N_3349);
or U6235 (N_6235,N_3725,N_315);
nor U6236 (N_6236,N_3712,N_1764);
or U6237 (N_6237,N_530,N_1888);
or U6238 (N_6238,N_3141,N_1946);
nand U6239 (N_6239,N_93,N_1605);
or U6240 (N_6240,N_2634,N_4420);
xnor U6241 (N_6241,N_1317,N_3271);
and U6242 (N_6242,N_3227,N_3998);
and U6243 (N_6243,N_3317,N_4493);
nor U6244 (N_6244,N_2160,N_152);
nand U6245 (N_6245,N_80,N_1681);
nand U6246 (N_6246,N_2629,N_34);
or U6247 (N_6247,N_1258,N_3969);
or U6248 (N_6248,N_3677,N_1672);
xor U6249 (N_6249,N_1314,N_4120);
nand U6250 (N_6250,N_4198,N_2866);
and U6251 (N_6251,N_3620,N_2689);
or U6252 (N_6252,N_3796,N_4091);
and U6253 (N_6253,N_3222,N_1081);
or U6254 (N_6254,N_509,N_2364);
nand U6255 (N_6255,N_4713,N_4401);
or U6256 (N_6256,N_854,N_2135);
xor U6257 (N_6257,N_4728,N_2304);
nand U6258 (N_6258,N_3435,N_1862);
xnor U6259 (N_6259,N_713,N_1849);
nor U6260 (N_6260,N_2548,N_157);
and U6261 (N_6261,N_2405,N_1454);
xor U6262 (N_6262,N_2486,N_1190);
xor U6263 (N_6263,N_4211,N_3687);
xor U6264 (N_6264,N_520,N_3020);
and U6265 (N_6265,N_646,N_4432);
nand U6266 (N_6266,N_3685,N_4482);
nand U6267 (N_6267,N_1123,N_546);
and U6268 (N_6268,N_2127,N_842);
nor U6269 (N_6269,N_481,N_4451);
or U6270 (N_6270,N_32,N_692);
xor U6271 (N_6271,N_2602,N_868);
or U6272 (N_6272,N_827,N_659);
xor U6273 (N_6273,N_27,N_2066);
xnor U6274 (N_6274,N_304,N_1534);
xor U6275 (N_6275,N_2123,N_2431);
and U6276 (N_6276,N_3762,N_306);
or U6277 (N_6277,N_2517,N_2845);
and U6278 (N_6278,N_553,N_4990);
or U6279 (N_6279,N_3000,N_86);
or U6280 (N_6280,N_4980,N_3993);
or U6281 (N_6281,N_1486,N_3488);
or U6282 (N_6282,N_2150,N_1288);
and U6283 (N_6283,N_4360,N_4874);
and U6284 (N_6284,N_3709,N_891);
or U6285 (N_6285,N_4200,N_4339);
nand U6286 (N_6286,N_3705,N_1263);
and U6287 (N_6287,N_3901,N_2452);
xor U6288 (N_6288,N_47,N_4403);
nor U6289 (N_6289,N_2384,N_768);
and U6290 (N_6290,N_1637,N_1040);
and U6291 (N_6291,N_4281,N_643);
xnor U6292 (N_6292,N_1295,N_3395);
or U6293 (N_6293,N_2273,N_1997);
nor U6294 (N_6294,N_2962,N_3693);
and U6295 (N_6295,N_2186,N_1192);
or U6296 (N_6296,N_4741,N_1625);
nor U6297 (N_6297,N_270,N_3135);
xnor U6298 (N_6298,N_2913,N_1763);
and U6299 (N_6299,N_3518,N_1409);
or U6300 (N_6300,N_3825,N_3016);
nand U6301 (N_6301,N_3997,N_1857);
nor U6302 (N_6302,N_3904,N_4030);
xor U6303 (N_6303,N_1026,N_4239);
xnor U6304 (N_6304,N_3223,N_2072);
nand U6305 (N_6305,N_1581,N_4877);
nor U6306 (N_6306,N_4405,N_3451);
or U6307 (N_6307,N_4860,N_4010);
xnor U6308 (N_6308,N_3460,N_3925);
and U6309 (N_6309,N_3458,N_901);
nand U6310 (N_6310,N_3305,N_965);
xnor U6311 (N_6311,N_1178,N_3139);
or U6312 (N_6312,N_3858,N_4135);
xnor U6313 (N_6313,N_3590,N_4781);
and U6314 (N_6314,N_1244,N_3641);
and U6315 (N_6315,N_618,N_2666);
or U6316 (N_6316,N_1667,N_3741);
nor U6317 (N_6317,N_3152,N_3650);
or U6318 (N_6318,N_3875,N_1541);
or U6319 (N_6319,N_2715,N_3724);
or U6320 (N_6320,N_3788,N_3358);
or U6321 (N_6321,N_2794,N_1408);
nor U6322 (N_6322,N_1170,N_2991);
nand U6323 (N_6323,N_4438,N_1412);
nand U6324 (N_6324,N_4026,N_1064);
nand U6325 (N_6325,N_4843,N_477);
nand U6326 (N_6326,N_3150,N_3055);
xor U6327 (N_6327,N_1446,N_4484);
xor U6328 (N_6328,N_3728,N_4338);
nand U6329 (N_6329,N_1853,N_73);
nor U6330 (N_6330,N_4618,N_4826);
or U6331 (N_6331,N_1601,N_1597);
xnor U6332 (N_6332,N_3119,N_318);
or U6333 (N_6333,N_4536,N_4287);
nand U6334 (N_6334,N_2489,N_431);
nand U6335 (N_6335,N_4154,N_971);
xor U6336 (N_6336,N_1664,N_853);
xor U6337 (N_6337,N_4905,N_4535);
and U6338 (N_6338,N_623,N_1422);
and U6339 (N_6339,N_3013,N_1234);
xnor U6340 (N_6340,N_1139,N_1099);
nand U6341 (N_6341,N_946,N_4638);
nor U6342 (N_6342,N_503,N_2856);
and U6343 (N_6343,N_1993,N_4040);
nand U6344 (N_6344,N_2793,N_4804);
xor U6345 (N_6345,N_2205,N_290);
and U6346 (N_6346,N_4331,N_3101);
or U6347 (N_6347,N_676,N_1005);
nor U6348 (N_6348,N_3714,N_1515);
and U6349 (N_6349,N_4399,N_3388);
and U6350 (N_6350,N_1272,N_4344);
or U6351 (N_6351,N_4881,N_839);
and U6352 (N_6352,N_360,N_4889);
nand U6353 (N_6353,N_1971,N_4706);
xor U6354 (N_6354,N_1565,N_3151);
nand U6355 (N_6355,N_3377,N_1052);
xnor U6356 (N_6356,N_3654,N_2903);
or U6357 (N_6357,N_2732,N_4143);
nor U6358 (N_6358,N_4848,N_7);
nand U6359 (N_6359,N_4449,N_1819);
nand U6360 (N_6360,N_4714,N_2835);
and U6361 (N_6361,N_350,N_2023);
or U6362 (N_6362,N_1055,N_657);
nor U6363 (N_6363,N_3810,N_399);
xor U6364 (N_6364,N_1444,N_3219);
nand U6365 (N_6365,N_4842,N_4578);
nand U6366 (N_6366,N_807,N_1952);
or U6367 (N_6367,N_792,N_3887);
or U6368 (N_6368,N_4464,N_2821);
nor U6369 (N_6369,N_4629,N_2401);
and U6370 (N_6370,N_1353,N_785);
or U6371 (N_6371,N_3157,N_3266);
xor U6372 (N_6372,N_3595,N_2259);
xor U6373 (N_6373,N_1002,N_4621);
xor U6374 (N_6374,N_4422,N_3545);
xnor U6375 (N_6375,N_4327,N_4168);
or U6376 (N_6376,N_1388,N_4524);
or U6377 (N_6377,N_119,N_1135);
and U6378 (N_6378,N_2325,N_3472);
and U6379 (N_6379,N_2745,N_2410);
and U6380 (N_6380,N_4001,N_3434);
or U6381 (N_6381,N_3294,N_3290);
and U6382 (N_6382,N_3386,N_4229);
or U6383 (N_6383,N_3731,N_3608);
xor U6384 (N_6384,N_2622,N_1488);
nand U6385 (N_6385,N_2230,N_2077);
nand U6386 (N_6386,N_1282,N_4187);
and U6387 (N_6387,N_4591,N_3365);
and U6388 (N_6388,N_527,N_4045);
and U6389 (N_6389,N_3776,N_1856);
or U6390 (N_6390,N_637,N_4090);
and U6391 (N_6391,N_3407,N_679);
or U6392 (N_6392,N_160,N_3981);
xnor U6393 (N_6393,N_1385,N_3461);
nor U6394 (N_6394,N_758,N_2518);
nand U6395 (N_6395,N_1557,N_3674);
nand U6396 (N_6396,N_3249,N_2473);
xor U6397 (N_6397,N_3363,N_1032);
nor U6398 (N_6398,N_3273,N_370);
or U6399 (N_6399,N_3909,N_45);
nand U6400 (N_6400,N_420,N_3985);
nor U6401 (N_6401,N_2841,N_140);
nor U6402 (N_6402,N_4850,N_956);
and U6403 (N_6403,N_1628,N_4114);
nor U6404 (N_6404,N_3056,N_1027);
or U6405 (N_6405,N_1982,N_2064);
and U6406 (N_6406,N_1584,N_789);
nor U6407 (N_6407,N_238,N_1596);
or U6408 (N_6408,N_2089,N_2524);
nor U6409 (N_6409,N_4439,N_3302);
nand U6410 (N_6410,N_3329,N_209);
or U6411 (N_6411,N_3627,N_641);
or U6412 (N_6412,N_2295,N_3587);
and U6413 (N_6413,N_2624,N_4554);
xor U6414 (N_6414,N_4724,N_1729);
or U6415 (N_6415,N_3109,N_1355);
or U6416 (N_6416,N_1098,N_2979);
nand U6417 (N_6417,N_1513,N_1120);
or U6418 (N_6418,N_1448,N_3230);
and U6419 (N_6419,N_2782,N_4088);
and U6420 (N_6420,N_4749,N_882);
nand U6421 (N_6421,N_4539,N_1635);
nand U6422 (N_6422,N_1438,N_4612);
nand U6423 (N_6423,N_2146,N_4503);
nor U6424 (N_6424,N_2859,N_514);
and U6425 (N_6425,N_3186,N_3049);
and U6426 (N_6426,N_64,N_1592);
or U6427 (N_6427,N_4568,N_3437);
or U6428 (N_6428,N_2013,N_3247);
and U6429 (N_6429,N_159,N_531);
and U6430 (N_6430,N_1124,N_3366);
xor U6431 (N_6431,N_2415,N_3560);
and U6432 (N_6432,N_4418,N_1096);
and U6433 (N_6433,N_3944,N_2986);
nor U6434 (N_6434,N_4930,N_299);
nand U6435 (N_6435,N_1613,N_4971);
xnor U6436 (N_6436,N_4518,N_652);
xor U6437 (N_6437,N_594,N_269);
nand U6438 (N_6438,N_1574,N_2147);
nand U6439 (N_6439,N_2132,N_3524);
and U6440 (N_6440,N_4462,N_1838);
nor U6441 (N_6441,N_409,N_207);
and U6442 (N_6442,N_4489,N_2965);
nor U6443 (N_6443,N_3028,N_4012);
xnor U6444 (N_6444,N_2941,N_1652);
or U6445 (N_6445,N_3168,N_1874);
or U6446 (N_6446,N_2121,N_1162);
xnor U6447 (N_6447,N_2394,N_41);
or U6448 (N_6448,N_3136,N_685);
and U6449 (N_6449,N_2883,N_1878);
xnor U6450 (N_6450,N_3470,N_1577);
and U6451 (N_6451,N_1941,N_1151);
or U6452 (N_6452,N_2182,N_3957);
xor U6453 (N_6453,N_903,N_1365);
nor U6454 (N_6454,N_3566,N_1111);
xnor U6455 (N_6455,N_317,N_4476);
nor U6456 (N_6456,N_1499,N_2288);
or U6457 (N_6457,N_4825,N_1471);
xor U6458 (N_6458,N_3117,N_1449);
and U6459 (N_6459,N_437,N_1603);
or U6460 (N_6460,N_75,N_3754);
nand U6461 (N_6461,N_1665,N_3401);
xnor U6462 (N_6462,N_4077,N_2151);
xor U6463 (N_6463,N_2389,N_1855);
nand U6464 (N_6464,N_4893,N_3053);
or U6465 (N_6465,N_816,N_4668);
or U6466 (N_6466,N_1478,N_4789);
and U6467 (N_6467,N_3555,N_930);
and U6468 (N_6468,N_1343,N_4504);
and U6469 (N_6469,N_1839,N_1293);
or U6470 (N_6470,N_665,N_719);
nor U6471 (N_6471,N_3700,N_1255);
nand U6472 (N_6472,N_396,N_1266);
or U6473 (N_6473,N_3237,N_4719);
xor U6474 (N_6474,N_1335,N_2056);
xor U6475 (N_6475,N_3033,N_3683);
and U6476 (N_6476,N_2667,N_3599);
xor U6477 (N_6477,N_4376,N_4954);
and U6478 (N_6478,N_1479,N_2609);
xor U6479 (N_6479,N_3172,N_4931);
nand U6480 (N_6480,N_883,N_141);
nand U6481 (N_6481,N_3411,N_1836);
xor U6482 (N_6482,N_441,N_898);
nor U6483 (N_6483,N_1908,N_2371);
or U6484 (N_6484,N_2942,N_4192);
nor U6485 (N_6485,N_539,N_2054);
or U6486 (N_6486,N_1779,N_2348);
nor U6487 (N_6487,N_579,N_3509);
nor U6488 (N_6488,N_3624,N_4479);
nor U6489 (N_6489,N_1500,N_425);
or U6490 (N_6490,N_1954,N_2210);
nand U6491 (N_6491,N_2519,N_564);
nor U6492 (N_6492,N_2767,N_1235);
nand U6493 (N_6493,N_4823,N_1456);
xor U6494 (N_6494,N_3319,N_1561);
nand U6495 (N_6495,N_447,N_1118);
nor U6496 (N_6496,N_66,N_2458);
or U6497 (N_6497,N_4816,N_3837);
nor U6498 (N_6498,N_1021,N_1366);
nand U6499 (N_6499,N_600,N_4592);
nor U6500 (N_6500,N_3031,N_3966);
or U6501 (N_6501,N_4286,N_2442);
xor U6502 (N_6502,N_3213,N_960);
nor U6503 (N_6503,N_4453,N_1485);
and U6504 (N_6504,N_4257,N_2516);
nand U6505 (N_6505,N_3750,N_3167);
xnor U6506 (N_6506,N_542,N_58);
nor U6507 (N_6507,N_163,N_3727);
and U6508 (N_6508,N_1065,N_3632);
xnor U6509 (N_6509,N_4856,N_4273);
nand U6510 (N_6510,N_128,N_3913);
or U6511 (N_6511,N_1585,N_3354);
xor U6512 (N_6512,N_4806,N_4020);
and U6513 (N_6513,N_1167,N_4158);
nand U6514 (N_6514,N_4563,N_1198);
and U6515 (N_6515,N_2987,N_2213);
nor U6516 (N_6516,N_3528,N_606);
nand U6517 (N_6517,N_2336,N_3010);
nand U6518 (N_6518,N_2640,N_3322);
xor U6519 (N_6519,N_2949,N_1148);
nor U6520 (N_6520,N_2447,N_400);
xor U6521 (N_6521,N_2673,N_1332);
and U6522 (N_6522,N_1369,N_2274);
xor U6523 (N_6523,N_1057,N_1893);
nand U6524 (N_6524,N_4285,N_4888);
xor U6525 (N_6525,N_1291,N_2896);
and U6526 (N_6526,N_538,N_2461);
xnor U6527 (N_6527,N_113,N_2737);
and U6528 (N_6528,N_1452,N_2145);
nand U6529 (N_6529,N_2144,N_4260);
and U6530 (N_6530,N_474,N_2187);
or U6531 (N_6531,N_4121,N_742);
and U6532 (N_6532,N_3442,N_2625);
or U6533 (N_6533,N_424,N_1588);
nor U6534 (N_6534,N_749,N_2738);
xor U6535 (N_6535,N_908,N_4320);
xor U6536 (N_6536,N_4277,N_1436);
nand U6537 (N_6537,N_1795,N_1087);
and U6538 (N_6538,N_2026,N_4556);
or U6539 (N_6539,N_31,N_4356);
xor U6540 (N_6540,N_4787,N_3787);
nor U6541 (N_6541,N_3633,N_4361);
nor U6542 (N_6542,N_608,N_3665);
nor U6543 (N_6543,N_3842,N_4617);
xnor U6544 (N_6544,N_3553,N_373);
nand U6545 (N_6545,N_4747,N_3156);
nand U6546 (N_6546,N_3923,N_1034);
or U6547 (N_6547,N_3834,N_4126);
or U6548 (N_6548,N_3137,N_2984);
nand U6549 (N_6549,N_3954,N_4737);
nand U6550 (N_6550,N_274,N_3565);
xnor U6551 (N_6551,N_1176,N_1279);
xor U6552 (N_6552,N_1805,N_3888);
xnor U6553 (N_6553,N_4868,N_365);
and U6554 (N_6554,N_4272,N_794);
nor U6555 (N_6555,N_4297,N_3240);
nor U6556 (N_6556,N_1771,N_1654);
nor U6557 (N_6557,N_3836,N_3300);
nand U6558 (N_6558,N_3567,N_4799);
xnor U6559 (N_6559,N_3999,N_3919);
nand U6560 (N_6560,N_338,N_560);
or U6561 (N_6561,N_4917,N_2281);
and U6562 (N_6562,N_256,N_120);
nand U6563 (N_6563,N_4551,N_2515);
or U6564 (N_6564,N_2193,N_3427);
nand U6565 (N_6565,N_50,N_1657);
and U6566 (N_6566,N_693,N_4840);
nand U6567 (N_6567,N_3597,N_3716);
and U6568 (N_6568,N_2990,N_456);
xnor U6569 (N_6569,N_1629,N_3879);
and U6570 (N_6570,N_926,N_4988);
xor U6571 (N_6571,N_519,N_860);
and U6572 (N_6572,N_660,N_4474);
nor U6573 (N_6573,N_3368,N_3617);
nand U6574 (N_6574,N_932,N_1203);
nand U6575 (N_6575,N_1136,N_2501);
nand U6576 (N_6576,N_3236,N_2362);
nor U6577 (N_6577,N_4858,N_1936);
nor U6578 (N_6578,N_301,N_3940);
nor U6579 (N_6579,N_3623,N_2596);
nor U6580 (N_6580,N_2114,N_3873);
or U6581 (N_6581,N_3050,N_4233);
nand U6582 (N_6582,N_2944,N_550);
or U6583 (N_6583,N_4647,N_3052);
and U6584 (N_6584,N_216,N_3807);
xnor U6585 (N_6585,N_3931,N_3953);
nor U6586 (N_6586,N_4644,N_2323);
nor U6587 (N_6587,N_4184,N_671);
nand U6588 (N_6588,N_684,N_348);
xor U6589 (N_6589,N_4691,N_624);
xor U6590 (N_6590,N_2843,N_1821);
nor U6591 (N_6591,N_1886,N_3212);
and U6592 (N_6592,N_4896,N_2735);
and U6593 (N_6593,N_2976,N_2228);
and U6594 (N_6594,N_4743,N_4134);
or U6595 (N_6595,N_576,N_3007);
or U6596 (N_6596,N_2823,N_3507);
nor U6597 (N_6597,N_127,N_2201);
or U6598 (N_6598,N_3920,N_941);
xor U6599 (N_6599,N_2960,N_2863);
xnor U6600 (N_6600,N_2073,N_406);
nor U6601 (N_6601,N_670,N_993);
and U6602 (N_6602,N_497,N_1100);
xnor U6603 (N_6603,N_4347,N_1356);
and U6604 (N_6604,N_2635,N_3752);
xnor U6605 (N_6605,N_2679,N_2894);
nand U6606 (N_6606,N_1898,N_1413);
nand U6607 (N_6607,N_493,N_1675);
nand U6608 (N_6608,N_1129,N_541);
nand U6609 (N_6609,N_4643,N_3216);
and U6610 (N_6610,N_3327,N_1242);
nor U6611 (N_6611,N_2725,N_18);
and U6612 (N_6612,N_1225,N_2888);
and U6613 (N_6613,N_3285,N_2202);
xnor U6614 (N_6614,N_3400,N_1012);
nand U6615 (N_6615,N_1320,N_4547);
xor U6616 (N_6616,N_3718,N_1075);
nor U6617 (N_6617,N_260,N_3085);
nor U6618 (N_6618,N_4152,N_3064);
and U6619 (N_6619,N_38,N_4622);
and U6620 (N_6620,N_1716,N_4129);
nor U6621 (N_6621,N_2227,N_1535);
xor U6622 (N_6622,N_3543,N_4092);
nor U6623 (N_6623,N_2344,N_4112);
or U6624 (N_6624,N_132,N_96);
and U6625 (N_6625,N_2020,N_2523);
nor U6626 (N_6626,N_864,N_2682);
xor U6627 (N_6627,N_3356,N_3067);
or U6628 (N_6628,N_2332,N_781);
or U6629 (N_6629,N_4924,N_428);
xnor U6630 (N_6630,N_1619,N_2390);
nor U6631 (N_6631,N_4838,N_2105);
nand U6632 (N_6632,N_3379,N_3173);
or U6633 (N_6633,N_4939,N_460);
nand U6634 (N_6634,N_2520,N_143);
xnor U6635 (N_6635,N_2545,N_1262);
nand U6636 (N_6636,N_3355,N_267);
nand U6637 (N_6637,N_3759,N_831);
xnor U6638 (N_6638,N_3278,N_138);
nand U6639 (N_6639,N_4560,N_4798);
nor U6640 (N_6640,N_3410,N_4387);
xnor U6641 (N_6641,N_2751,N_1575);
and U6642 (N_6642,N_3416,N_2819);
nand U6643 (N_6643,N_1961,N_4732);
nand U6644 (N_6644,N_766,N_2232);
and U6645 (N_6645,N_4397,N_254);
and U6646 (N_6646,N_1693,N_21);
or U6647 (N_6647,N_353,N_1430);
xor U6648 (N_6648,N_4986,N_3208);
nand U6649 (N_6649,N_4642,N_181);
and U6650 (N_6650,N_3648,N_2681);
xnor U6651 (N_6651,N_672,N_2649);
nand U6652 (N_6652,N_2887,N_4871);
or U6653 (N_6653,N_2787,N_1251);
and U6654 (N_6654,N_3253,N_1080);
or U6655 (N_6655,N_4819,N_1606);
xor U6656 (N_6656,N_3169,N_2164);
and U6657 (N_6657,N_4195,N_2529);
nor U6658 (N_6658,N_3406,N_2291);
and U6659 (N_6659,N_2237,N_4508);
xor U6660 (N_6660,N_704,N_2497);
or U6661 (N_6661,N_1429,N_1223);
or U6662 (N_6662,N_150,N_2420);
xor U6663 (N_6663,N_3124,N_2822);
nor U6664 (N_6664,N_985,N_2783);
or U6665 (N_6665,N_4105,N_1462);
xor U6666 (N_6666,N_1843,N_4946);
nor U6667 (N_6667,N_3476,N_2935);
nor U6668 (N_6668,N_4631,N_4579);
or U6669 (N_6669,N_2955,N_211);
xnor U6670 (N_6670,N_3505,N_3847);
nor U6671 (N_6671,N_3373,N_615);
nand U6672 (N_6672,N_482,N_4252);
and U6673 (N_6673,N_4219,N_2811);
nor U6674 (N_6674,N_2753,N_717);
xor U6675 (N_6675,N_2650,N_543);
or U6676 (N_6676,N_4801,N_1861);
nor U6677 (N_6677,N_1327,N_3588);
xnor U6678 (N_6678,N_1379,N_177);
nor U6679 (N_6679,N_595,N_3095);
and U6680 (N_6680,N_1018,N_2);
nand U6681 (N_6681,N_1389,N_690);
nand U6682 (N_6682,N_571,N_755);
or U6683 (N_6683,N_1220,N_4130);
nand U6684 (N_6684,N_88,N_188);
nand U6685 (N_6685,N_1543,N_4767);
or U6686 (N_6686,N_3743,N_4761);
and U6687 (N_6687,N_1254,N_2358);
nor U6688 (N_6688,N_463,N_3060);
nand U6689 (N_6689,N_1542,N_823);
and U6690 (N_6690,N_3107,N_518);
nor U6691 (N_6691,N_194,N_2583);
nand U6692 (N_6692,N_4658,N_2511);
or U6693 (N_6693,N_1126,N_760);
nor U6694 (N_6694,N_735,N_1540);
and U6695 (N_6695,N_3601,N_4890);
and U6696 (N_6696,N_1623,N_135);
or U6697 (N_6697,N_92,N_4185);
and U6698 (N_6698,N_3298,N_2750);
nor U6699 (N_6699,N_3736,N_1439);
xnor U6700 (N_6700,N_769,N_4766);
xor U6701 (N_6701,N_4156,N_3170);
nand U6702 (N_6702,N_3895,N_4723);
nand U6703 (N_6703,N_445,N_694);
nor U6704 (N_6704,N_2256,N_2177);
and U6705 (N_6705,N_162,N_4298);
or U6706 (N_6706,N_3547,N_2479);
and U6707 (N_6707,N_2557,N_2612);
nor U6708 (N_6708,N_3308,N_2761);
nand U6709 (N_6709,N_944,N_4409);
xor U6710 (N_6710,N_1966,N_3353);
xor U6711 (N_6711,N_2705,N_2124);
nand U6712 (N_6712,N_4400,N_744);
nand U6713 (N_6713,N_4929,N_625);
xor U6714 (N_6714,N_2263,N_3251);
nand U6715 (N_6715,N_2683,N_3939);
or U6716 (N_6716,N_1303,N_4922);
and U6717 (N_6717,N_2424,N_334);
or U6718 (N_6718,N_2061,N_2030);
xnor U6719 (N_6719,N_2796,N_1019);
nand U6720 (N_6720,N_3378,N_732);
nor U6721 (N_6721,N_2208,N_547);
and U6722 (N_6722,N_3260,N_2831);
nor U6723 (N_6723,N_3014,N_1213);
or U6724 (N_6724,N_4225,N_104);
xor U6725 (N_6725,N_3949,N_4873);
and U6726 (N_6726,N_2133,N_2934);
nor U6727 (N_6727,N_1912,N_1447);
and U6728 (N_6728,N_780,N_788);
nor U6729 (N_6729,N_4829,N_4180);
nand U6730 (N_6730,N_2166,N_748);
or U6731 (N_6731,N_1600,N_1256);
or U6732 (N_6732,N_847,N_459);
xnor U6733 (N_6733,N_1643,N_2765);
and U6734 (N_6734,N_650,N_2255);
xnor U6735 (N_6735,N_2551,N_3586);
nand U6736 (N_6736,N_1277,N_2904);
and U6737 (N_6737,N_4709,N_3658);
nand U6738 (N_6738,N_469,N_4058);
nor U6739 (N_6739,N_446,N_3935);
nor U6740 (N_6740,N_2528,N_3045);
nor U6741 (N_6741,N_2498,N_4690);
xor U6742 (N_6742,N_621,N_2407);
xnor U6743 (N_6743,N_1296,N_2748);
and U6744 (N_6744,N_714,N_2474);
nand U6745 (N_6745,N_2478,N_36);
or U6746 (N_6746,N_746,N_2321);
or U6747 (N_6747,N_2095,N_83);
and U6748 (N_6748,N_295,N_991);
or U6749 (N_6749,N_798,N_3256);
xnor U6750 (N_6750,N_4275,N_947);
nor U6751 (N_6751,N_4431,N_2050);
and U6752 (N_6752,N_1175,N_2540);
xor U6753 (N_6753,N_4027,N_989);
nor U6754 (N_6754,N_2713,N_1863);
or U6755 (N_6755,N_2079,N_821);
or U6756 (N_6756,N_4782,N_1868);
nand U6757 (N_6757,N_4314,N_939);
nor U6758 (N_6758,N_3870,N_556);
or U6759 (N_6759,N_1963,N_4729);
xnor U6760 (N_6760,N_3582,N_203);
xnor U6761 (N_6761,N_825,N_4351);
and U6762 (N_6762,N_412,N_782);
nor U6763 (N_6763,N_2763,N_3490);
nor U6764 (N_6764,N_1464,N_3199);
nand U6765 (N_6765,N_710,N_3877);
nand U6766 (N_6766,N_248,N_1097);
or U6767 (N_6767,N_4884,N_125);
and U6768 (N_6768,N_4953,N_2180);
and U6769 (N_6769,N_1058,N_959);
and U6770 (N_6770,N_4742,N_987);
nor U6771 (N_6771,N_2460,N_3558);
xnor U6772 (N_6772,N_3467,N_3519);
xnor U6773 (N_6773,N_4136,N_2575);
or U6774 (N_6774,N_580,N_4684);
and U6775 (N_6775,N_3001,N_2736);
nor U6776 (N_6776,N_743,N_1658);
nand U6777 (N_6777,N_4373,N_2939);
or U6778 (N_6778,N_4635,N_4662);
and U6779 (N_6779,N_3672,N_158);
and U6780 (N_6780,N_2547,N_3214);
xnor U6781 (N_6781,N_812,N_4972);
nor U6782 (N_6782,N_1620,N_2699);
xnor U6783 (N_6783,N_4687,N_319);
or U6784 (N_6784,N_4118,N_242);
or U6785 (N_6785,N_2219,N_1364);
and U6786 (N_6786,N_1927,N_1074);
and U6787 (N_6787,N_1775,N_4388);
xor U6788 (N_6788,N_3938,N_1373);
and U6789 (N_6789,N_2844,N_3499);
and U6790 (N_6790,N_3816,N_4024);
nand U6791 (N_6791,N_480,N_1357);
nand U6792 (N_6792,N_2440,N_2179);
nor U6793 (N_6793,N_1803,N_4201);
xor U6794 (N_6794,N_738,N_4611);
and U6795 (N_6795,N_4697,N_1815);
and U6796 (N_6796,N_3462,N_667);
nand U6797 (N_6797,N_1741,N_4759);
or U6798 (N_6798,N_1091,N_3581);
xnor U6799 (N_6799,N_4810,N_599);
and U6800 (N_6800,N_340,N_1903);
nor U6801 (N_6801,N_1418,N_231);
nor U6802 (N_6802,N_620,N_532);
and U6803 (N_6803,N_1043,N_3951);
xor U6804 (N_6804,N_1711,N_4615);
nor U6805 (N_6805,N_1892,N_4901);
nor U6806 (N_6806,N_2558,N_1551);
xnor U6807 (N_6807,N_33,N_797);
nand U6808 (N_6808,N_4459,N_1150);
xor U6809 (N_6809,N_2875,N_4465);
nand U6810 (N_6810,N_2130,N_1391);
nand U6811 (N_6811,N_561,N_458);
and U6812 (N_6812,N_3295,N_3412);
nor U6813 (N_6813,N_4613,N_3393);
nor U6814 (N_6814,N_3032,N_4263);
or U6815 (N_6815,N_4895,N_255);
xnor U6816 (N_6816,N_3767,N_3910);
nand U6817 (N_6817,N_2770,N_2432);
nor U6818 (N_6818,N_4704,N_1359);
and U6819 (N_6819,N_2702,N_3552);
nand U6820 (N_6820,N_1524,N_4718);
or U6821 (N_6821,N_3746,N_341);
xor U6822 (N_6822,N_3195,N_1319);
xnor U6823 (N_6823,N_4188,N_4510);
nor U6824 (N_6824,N_3239,N_2810);
and U6825 (N_6825,N_1989,N_3912);
nand U6826 (N_6826,N_2372,N_3684);
xnor U6827 (N_6827,N_4243,N_3276);
xor U6828 (N_6828,N_2946,N_377);
nand U6829 (N_6829,N_3074,N_2444);
and U6830 (N_6830,N_4300,N_3475);
nor U6831 (N_6831,N_611,N_1249);
nand U6832 (N_6832,N_2009,N_2876);
nor U6833 (N_6833,N_376,N_1709);
and U6834 (N_6834,N_988,N_1368);
nand U6835 (N_6835,N_2381,N_873);
and U6836 (N_6836,N_4038,N_1001);
nand U6837 (N_6837,N_3289,N_4501);
or U6838 (N_6838,N_3311,N_4421);
or U6839 (N_6839,N_4627,N_2850);
and U6840 (N_6840,N_3459,N_4217);
or U6841 (N_6841,N_3863,N_3772);
nor U6842 (N_6842,N_2776,N_3527);
and U6843 (N_6843,N_1367,N_3982);
and U6844 (N_6844,N_1727,N_4634);
xor U6845 (N_6845,N_1257,N_2477);
nand U6846 (N_6846,N_2190,N_2956);
and U6847 (N_6847,N_136,N_2791);
xnor U6848 (N_6848,N_4208,N_4170);
and U6849 (N_6849,N_2964,N_587);
nor U6850 (N_6850,N_2041,N_4079);
nand U6851 (N_6851,N_4656,N_2335);
xnor U6852 (N_6852,N_767,N_4342);
nand U6853 (N_6853,N_79,N_2567);
xor U6854 (N_6854,N_381,N_4951);
xor U6855 (N_6855,N_4851,N_3192);
nand U6856 (N_6856,N_2306,N_4961);
nand U6857 (N_6857,N_42,N_3602);
nor U6858 (N_6858,N_3670,N_3614);
nand U6859 (N_6859,N_2842,N_1770);
and U6860 (N_6860,N_3539,N_4976);
nor U6861 (N_6861,N_1645,N_4095);
xor U6862 (N_6862,N_305,N_332);
or U6863 (N_6863,N_9,N_335);
or U6864 (N_6864,N_2165,N_4450);
nand U6865 (N_6865,N_3571,N_2807);
xor U6866 (N_6866,N_4415,N_937);
nor U6867 (N_6867,N_3189,N_43);
and U6868 (N_6868,N_2377,N_1940);
or U6869 (N_6869,N_631,N_1073);
xor U6870 (N_6870,N_4271,N_2134);
nand U6871 (N_6871,N_1372,N_1955);
and U6872 (N_6872,N_4543,N_712);
nand U6873 (N_6873,N_3469,N_1119);
and U6874 (N_6874,N_1132,N_2388);
nor U6875 (N_6875,N_2059,N_403);
nor U6876 (N_6876,N_178,N_3420);
xor U6877 (N_6877,N_1773,N_2513);
xnor U6878 (N_6878,N_801,N_945);
nand U6879 (N_6879,N_2687,N_4483);
nor U6880 (N_6880,N_4169,N_1305);
xor U6881 (N_6881,N_3656,N_2993);
nand U6882 (N_6882,N_485,N_3989);
and U6883 (N_6883,N_601,N_3735);
or U6884 (N_6884,N_3833,N_1944);
nor U6885 (N_6885,N_4790,N_4959);
or U6886 (N_6886,N_4113,N_990);
xnor U6887 (N_6887,N_4640,N_3129);
or U6888 (N_6888,N_1348,N_4947);
xor U6889 (N_6889,N_149,N_2296);
nor U6890 (N_6890,N_4371,N_4788);
xor U6891 (N_6891,N_3979,N_494);
nand U6892 (N_6892,N_1965,N_2481);
and U6893 (N_6893,N_2621,N_3148);
nor U6894 (N_6894,N_4341,N_3819);
or U6895 (N_6895,N_3058,N_1842);
and U6896 (N_6896,N_2453,N_1337);
and U6897 (N_6897,N_2988,N_911);
and U6898 (N_6898,N_3483,N_3326);
or U6899 (N_6899,N_2663,N_537);
xnor U6900 (N_6900,N_3132,N_2400);
or U6901 (N_6901,N_4299,N_1547);
xnor U6902 (N_6902,N_118,N_4516);
or U6903 (N_6903,N_3657,N_3521);
nand U6904 (N_6904,N_4316,N_187);
or U6905 (N_6905,N_272,N_2300);
xnor U6906 (N_6906,N_4733,N_4375);
nor U6907 (N_6907,N_3576,N_3515);
or U6908 (N_6908,N_1662,N_3044);
and U6909 (N_6909,N_65,N_4293);
xnor U6910 (N_6910,N_4703,N_4458);
nand U6911 (N_6911,N_510,N_4093);
or U6912 (N_6912,N_1822,N_501);
nand U6913 (N_6913,N_1006,N_3734);
and U6914 (N_6914,N_4927,N_402);
nand U6915 (N_6915,N_3506,N_2967);
and U6916 (N_6916,N_2264,N_144);
or U6917 (N_6917,N_4659,N_1985);
nand U6918 (N_6918,N_4682,N_4125);
or U6919 (N_6919,N_70,N_2196);
nor U6920 (N_6920,N_948,N_1705);
nand U6921 (N_6921,N_4632,N_1307);
xnor U6922 (N_6922,N_1473,N_4386);
xor U6923 (N_6923,N_4064,N_4876);
or U6924 (N_6924,N_1990,N_277);
nor U6925 (N_6925,N_57,N_1673);
xnor U6926 (N_6926,N_1236,N_841);
and U6927 (N_6927,N_1823,N_4864);
xor U6928 (N_6928,N_3121,N_1114);
xor U6929 (N_6929,N_4966,N_1125);
nor U6930 (N_6930,N_2391,N_3453);
nor U6931 (N_6931,N_2368,N_1060);
nor U6932 (N_6932,N_4278,N_689);
xnor U6933 (N_6933,N_2630,N_4655);
xor U6934 (N_6934,N_1624,N_168);
nand U6935 (N_6935,N_4486,N_4869);
xor U6936 (N_6936,N_3343,N_3777);
nand U6937 (N_6937,N_2283,N_2938);
or U6938 (N_6938,N_3958,N_435);
and U6939 (N_6939,N_3987,N_4414);
and U6940 (N_6940,N_4862,N_813);
nor U6941 (N_6941,N_3202,N_4220);
nand U6942 (N_6942,N_4879,N_4768);
xor U6943 (N_6943,N_4218,N_1224);
nand U6944 (N_6944,N_2090,N_337);
and U6945 (N_6945,N_1651,N_3413);
nand U6946 (N_6946,N_3337,N_3398);
and U6947 (N_6947,N_2094,N_2475);
or U6948 (N_6948,N_1807,N_4875);
xnor U6949 (N_6949,N_2379,N_2116);
or U6950 (N_6950,N_3541,N_2613);
nor U6951 (N_6951,N_1115,N_653);
and U6952 (N_6952,N_268,N_1383);
xor U6953 (N_6953,N_2874,N_575);
nand U6954 (N_6954,N_2800,N_551);
nand U6955 (N_6955,N_201,N_2919);
nand U6956 (N_6956,N_225,N_3956);
and U6957 (N_6957,N_249,N_1691);
nor U6958 (N_6958,N_4769,N_1519);
nand U6959 (N_6959,N_1201,N_108);
nor U6960 (N_6960,N_696,N_233);
or U6961 (N_6961,N_3009,N_1930);
xnor U6962 (N_6962,N_4891,N_1318);
or U6963 (N_6963,N_2580,N_3899);
xnor U6964 (N_6964,N_529,N_2435);
nand U6965 (N_6965,N_2618,N_3183);
nand U6966 (N_6966,N_4197,N_3537);
nor U6967 (N_6967,N_2927,N_1071);
or U6968 (N_6968,N_3758,N_1967);
xnor U6969 (N_6969,N_1785,N_2025);
and U6970 (N_6970,N_2493,N_4834);
nand U6971 (N_6971,N_809,N_3089);
nand U6972 (N_6972,N_1247,N_4880);
nor U6973 (N_6973,N_675,N_2393);
nor U6974 (N_6974,N_3738,N_4815);
and U6975 (N_6975,N_528,N_312);
xor U6976 (N_6976,N_3102,N_2031);
nand U6977 (N_6977,N_2868,N_4715);
nor U6978 (N_6978,N_2546,N_924);
nor U6979 (N_6979,N_3745,N_2848);
nor U6980 (N_6980,N_1147,N_1646);
or U6981 (N_6981,N_4775,N_1077);
and U6982 (N_6982,N_499,N_2992);
or U6983 (N_6983,N_478,N_1102);
nand U6984 (N_6984,N_4952,N_4393);
and U6985 (N_6985,N_3131,N_566);
and U6986 (N_6986,N_2238,N_669);
and U6987 (N_6987,N_3206,N_2465);
or U6988 (N_6988,N_1397,N_3933);
nor U6989 (N_6989,N_3441,N_4571);
or U6990 (N_6990,N_1925,N_4738);
nor U6991 (N_6991,N_1641,N_2387);
or U6992 (N_6992,N_275,N_4305);
or U6993 (N_6993,N_3740,N_3559);
xnor U6994 (N_6994,N_2359,N_3600);
nor U6995 (N_6995,N_252,N_1867);
nor U6996 (N_6996,N_1023,N_1284);
nor U6997 (N_6997,N_2261,N_4227);
or U6998 (N_6998,N_3726,N_3947);
or U6999 (N_6999,N_3584,N_1104);
xor U7000 (N_7000,N_635,N_3782);
xnor U7001 (N_7001,N_1648,N_4041);
nor U7002 (N_7002,N_3719,N_3383);
nor U7003 (N_7003,N_555,N_3976);
and U7004 (N_7004,N_1755,N_2855);
xnor U7005 (N_7005,N_3008,N_3707);
or U7006 (N_7006,N_942,N_534);
xor U7007 (N_7007,N_4754,N_552);
and U7008 (N_7008,N_51,N_3503);
nor U7009 (N_7009,N_2693,N_3867);
and U7010 (N_7010,N_4098,N_1221);
xor U7011 (N_7011,N_283,N_896);
xor U7012 (N_7012,N_105,N_1859);
nor U7013 (N_7013,N_569,N_124);
and U7014 (N_7014,N_1466,N_2639);
and U7015 (N_7015,N_3017,N_3970);
or U7016 (N_7016,N_1595,N_1854);
and U7017 (N_7017,N_4970,N_1884);
and U7018 (N_7018,N_4740,N_3864);
nand U7019 (N_7019,N_3244,N_470);
nand U7020 (N_7020,N_1566,N_4698);
nand U7021 (N_7021,N_3138,N_3165);
nor U7022 (N_7022,N_3048,N_2769);
and U7023 (N_7023,N_4557,N_1921);
xnor U7024 (N_7024,N_3637,N_1527);
xnor U7025 (N_7025,N_3207,N_4933);
or U7026 (N_7026,N_4900,N_4610);
and U7027 (N_7027,N_3817,N_2414);
and U7028 (N_7028,N_1848,N_1344);
and U7029 (N_7029,N_880,N_3231);
nand U7030 (N_7030,N_1212,N_3569);
nand U7031 (N_7031,N_1964,N_4428);
xor U7032 (N_7032,N_2039,N_2710);
nand U7033 (N_7033,N_1325,N_1722);
nand U7034 (N_7034,N_1156,N_1750);
or U7035 (N_7035,N_2346,N_423);
and U7036 (N_7036,N_4694,N_1401);
xor U7037 (N_7037,N_3394,N_3094);
nand U7038 (N_7038,N_3962,N_3753);
nor U7039 (N_7039,N_3445,N_1144);
and U7040 (N_7040,N_59,N_4402);
xor U7041 (N_7041,N_1879,N_4015);
nor U7042 (N_7042,N_2277,N_4977);
nand U7043 (N_7043,N_4265,N_326);
or U7044 (N_7044,N_1083,N_2616);
nor U7045 (N_7045,N_3012,N_2922);
nor U7046 (N_7046,N_4016,N_3455);
and U7047 (N_7047,N_4224,N_2722);
nor U7048 (N_7048,N_1634,N_2989);
xnor U7049 (N_7049,N_3577,N_3347);
xnor U7050 (N_7050,N_1076,N_4821);
nand U7051 (N_7051,N_2675,N_3769);
nor U7052 (N_7052,N_3865,N_1642);
nand U7053 (N_7053,N_2482,N_4292);
nor U7054 (N_7054,N_2495,N_1844);
nand U7055 (N_7055,N_4515,N_1706);
xor U7056 (N_7056,N_1450,N_1559);
or U7057 (N_7057,N_869,N_2129);
or U7058 (N_7058,N_4792,N_1924);
or U7059 (N_7059,N_4128,N_1552);
nor U7060 (N_7060,N_1602,N_4845);
xor U7061 (N_7061,N_1714,N_2974);
nand U7062 (N_7062,N_2260,N_3653);
nor U7063 (N_7063,N_91,N_1521);
and U7064 (N_7064,N_1582,N_723);
nor U7065 (N_7065,N_3197,N_4059);
nor U7066 (N_7066,N_3675,N_52);
nor U7067 (N_7067,N_71,N_3450);
nand U7068 (N_7068,N_3994,N_1580);
xnor U7069 (N_7069,N_2727,N_2287);
nor U7070 (N_7070,N_4212,N_2396);
nor U7071 (N_7071,N_4764,N_1747);
or U7072 (N_7072,N_835,N_101);
nand U7073 (N_7073,N_3795,N_3328);
or U7074 (N_7074,N_2784,N_3594);
nand U7075 (N_7075,N_2985,N_3021);
nand U7076 (N_7076,N_1172,N_3493);
or U7077 (N_7077,N_2163,N_2975);
nand U7078 (N_7078,N_1068,N_2951);
or U7079 (N_7079,N_4534,N_191);
nor U7080 (N_7080,N_1090,N_4849);
xnor U7081 (N_7081,N_3763,N_4746);
nand U7082 (N_7082,N_491,N_1894);
and U7083 (N_7083,N_3779,N_829);
nand U7084 (N_7084,N_2096,N_4807);
nand U7085 (N_7085,N_282,N_1398);
nor U7086 (N_7086,N_4923,N_1885);
nand U7087 (N_7087,N_2153,N_2925);
nor U7088 (N_7088,N_3689,N_2172);
xnor U7089 (N_7089,N_4802,N_2802);
nand U7090 (N_7090,N_3583,N_1947);
and U7091 (N_7091,N_4999,N_352);
xor U7092 (N_7092,N_3880,N_1441);
xor U7093 (N_7093,N_2779,N_1171);
or U7094 (N_7094,N_4104,N_2980);
xor U7095 (N_7095,N_2795,N_2997);
nand U7096 (N_7096,N_4485,N_4636);
nand U7097 (N_7097,N_4904,N_2351);
nor U7098 (N_7098,N_3279,N_2319);
and U7099 (N_7099,N_4368,N_4569);
xnor U7100 (N_7100,N_3057,N_3443);
nor U7101 (N_7101,N_3618,N_1656);
xnor U7102 (N_7102,N_3963,N_1312);
xnor U7103 (N_7103,N_1363,N_2636);
and U7104 (N_7104,N_3226,N_1929);
nor U7105 (N_7105,N_2857,N_2954);
nor U7106 (N_7106,N_4370,N_4);
nand U7107 (N_7107,N_3640,N_2525);
xnor U7108 (N_7108,N_1864,N_1495);
or U7109 (N_7109,N_3079,N_2599);
or U7110 (N_7110,N_2329,N_881);
nor U7111 (N_7111,N_3869,N_3568);
nor U7112 (N_7112,N_1252,N_1933);
or U7113 (N_7113,N_3922,N_111);
nor U7114 (N_7114,N_4189,N_3291);
nor U7115 (N_7115,N_1216,N_1395);
nand U7116 (N_7116,N_2195,N_2568);
or U7117 (N_7117,N_4396,N_244);
and U7118 (N_7118,N_4885,N_3243);
and U7119 (N_7119,N_1292,N_567);
and U7120 (N_7120,N_2239,N_2659);
or U7121 (N_7121,N_2063,N_1487);
and U7122 (N_7122,N_3069,N_1245);
xnor U7123 (N_7123,N_189,N_1218);
or U7124 (N_7124,N_2175,N_362);
or U7125 (N_7125,N_3883,N_2696);
nor U7126 (N_7126,N_220,N_495);
and U7127 (N_7127,N_1644,N_4958);
nand U7128 (N_7128,N_1411,N_3561);
nand U7129 (N_7129,N_4235,N_388);
xnor U7130 (N_7130,N_2923,N_2578);
nor U7131 (N_7131,N_2825,N_2448);
or U7132 (N_7132,N_705,N_4545);
xor U7133 (N_7133,N_4964,N_468);
nor U7134 (N_7134,N_1800,N_4269);
and U7135 (N_7135,N_2449,N_361);
nand U7136 (N_7136,N_3339,N_2862);
and U7137 (N_7137,N_4859,N_3361);
or U7138 (N_7138,N_4055,N_4590);
nor U7139 (N_7139,N_4830,N_1324);
xnor U7140 (N_7140,N_202,N_655);
nand U7141 (N_7141,N_4511,N_4820);
or U7142 (N_7142,N_4236,N_2438);
xnor U7143 (N_7143,N_1640,N_4280);
xnor U7144 (N_7144,N_1463,N_3359);
nand U7145 (N_7145,N_3288,N_1545);
and U7146 (N_7146,N_3885,N_3024);
nor U7147 (N_7147,N_2158,N_4036);
and U7148 (N_7148,N_516,N_2297);
nor U7149 (N_7149,N_3630,N_1890);
xnor U7150 (N_7150,N_2550,N_981);
xor U7151 (N_7151,N_2051,N_1079);
nor U7152 (N_7152,N_415,N_429);
nand U7153 (N_7153,N_3209,N_4144);
nand U7154 (N_7154,N_918,N_449);
and U7155 (N_7155,N_790,N_610);
xor U7156 (N_7156,N_3721,N_3063);
xor U7157 (N_7157,N_102,N_3934);
and U7158 (N_7158,N_2573,N_1278);
nor U7159 (N_7159,N_1326,N_1361);
or U7160 (N_7160,N_604,N_3698);
xor U7161 (N_7161,N_2331,N_4653);
or U7162 (N_7162,N_2847,N_2716);
xor U7163 (N_7163,N_2829,N_1321);
nor U7164 (N_7164,N_4205,N_4445);
xnor U7165 (N_7165,N_3065,N_3482);
nand U7166 (N_7166,N_455,N_94);
or U7167 (N_7167,N_1983,N_3175);
nor U7168 (N_7168,N_4073,N_302);
xor U7169 (N_7169,N_4526,N_3786);
nand U7170 (N_7170,N_4765,N_1066);
nand U7171 (N_7171,N_1647,N_1995);
nand U7172 (N_7172,N_76,N_900);
nor U7173 (N_7173,N_2820,N_3224);
and U7174 (N_7174,N_4648,N_291);
nand U7175 (N_7175,N_1460,N_1938);
or U7176 (N_7176,N_1088,N_4681);
nand U7177 (N_7177,N_1984,N_4022);
nor U7178 (N_7178,N_3513,N_180);
or U7179 (N_7179,N_3755,N_2047);
and U7180 (N_7180,N_4921,N_763);
xor U7181 (N_7181,N_4031,N_1024);
or U7182 (N_7182,N_992,N_3382);
xor U7183 (N_7183,N_3265,N_4296);
nand U7184 (N_7184,N_416,N_4017);
and U7185 (N_7185,N_2383,N_698);
nand U7186 (N_7186,N_876,N_833);
nand U7187 (N_7187,N_2826,N_3511);
xor U7188 (N_7188,N_504,N_777);
and U7189 (N_7189,N_1735,N_633);
or U7190 (N_7190,N_799,N_3812);
and U7191 (N_7191,N_4100,N_3821);
and U7192 (N_7192,N_4369,N_3704);
xnor U7193 (N_7193,N_1072,N_3203);
and U7194 (N_7194,N_3722,N_1138);
nor U7195 (N_7195,N_1300,N_4018);
nand U7196 (N_7196,N_3084,N_3843);
nand U7197 (N_7197,N_273,N_1748);
or U7198 (N_7198,N_3516,N_4391);
nand U7199 (N_7199,N_3611,N_4097);
xnor U7200 (N_7200,N_1209,N_3835);
nand U7201 (N_7201,N_2574,N_772);
and U7202 (N_7202,N_1688,N_983);
and U7203 (N_7203,N_4696,N_95);
or U7204 (N_7204,N_2881,N_1682);
nand U7205 (N_7205,N_4469,N_4672);
xnor U7206 (N_7206,N_1915,N_3824);
nor U7207 (N_7207,N_2445,N_970);
or U7208 (N_7208,N_366,N_814);
nand U7209 (N_7209,N_895,N_3268);
nor U7210 (N_7210,N_1754,N_3143);
xnor U7211 (N_7211,N_4447,N_2337);
nand U7212 (N_7212,N_4520,N_3706);
nand U7213 (N_7213,N_840,N_2620);
xor U7214 (N_7214,N_3534,N_3257);
xor U7215 (N_7215,N_3299,N_4346);
nor U7216 (N_7216,N_3881,N_4722);
nor U7217 (N_7217,N_820,N_4992);
and U7218 (N_7218,N_4878,N_770);
nand U7219 (N_7219,N_1786,N_1550);
and U7220 (N_7220,N_4179,N_884);
nor U7221 (N_7221,N_3967,N_3159);
and U7222 (N_7222,N_2514,N_4364);
and U7223 (N_7223,N_4928,N_3066);
xor U7224 (N_7224,N_1752,N_1310);
xnor U7225 (N_7225,N_3711,N_2207);
nor U7226 (N_7226,N_2961,N_1801);
nand U7227 (N_7227,N_1374,N_4497);
and U7228 (N_7228,N_292,N_2081);
or U7229 (N_7229,N_2416,N_1934);
and U7230 (N_7230,N_1960,N_3906);
nor U7231 (N_7231,N_3613,N_1799);
xor U7232 (N_7232,N_2231,N_3415);
and U7233 (N_7233,N_208,N_4780);
or U7234 (N_7234,N_1231,N_2707);
or U7235 (N_7235,N_1371,N_3744);
and U7236 (N_7236,N_4872,N_1339);
nand U7237 (N_7237,N_4550,N_4083);
and U7238 (N_7238,N_1776,N_752);
and U7239 (N_7239,N_1360,N_2354);
xnor U7240 (N_7240,N_919,N_2645);
nor U7241 (N_7241,N_1707,N_654);
or U7242 (N_7242,N_2125,N_4505);
nand U7243 (N_7243,N_4614,N_4979);
nand U7244 (N_7244,N_3419,N_4294);
or U7245 (N_7245,N_2680,N_475);
nand U7246 (N_7246,N_2278,N_1301);
and U7247 (N_7247,N_4847,N_4541);
and U7248 (N_7248,N_1233,N_2425);
xnor U7249 (N_7249,N_3765,N_2203);
nor U7250 (N_7250,N_1978,N_2598);
nor U7251 (N_7251,N_358,N_0);
xnor U7252 (N_7252,N_224,N_4701);
and U7253 (N_7253,N_4837,N_605);
nor U7254 (N_7254,N_2355,N_253);
nand U7255 (N_7255,N_2188,N_4182);
xnor U7256 (N_7256,N_3468,N_2507);
or U7257 (N_7257,N_2872,N_2778);
and U7258 (N_7258,N_1131,N_1313);
xor U7259 (N_7259,N_4254,N_2443);
nand U7260 (N_7260,N_4155,N_2542);
xor U7261 (N_7261,N_1612,N_3943);
xor U7262 (N_7262,N_2159,N_565);
xor U7263 (N_7263,N_1434,N_1591);
nor U7264 (N_7264,N_4982,N_438);
nand U7265 (N_7265,N_1687,N_4596);
nand U7266 (N_7266,N_699,N_4037);
or U7267 (N_7267,N_4907,N_8);
nand U7268 (N_7268,N_3886,N_3926);
nor U7269 (N_7269,N_682,N_3015);
or U7270 (N_7270,N_1532,N_3446);
nand U7271 (N_7271,N_4266,N_1726);
nand U7272 (N_7272,N_4067,N_525);
and U7273 (N_7273,N_2413,N_4190);
and U7274 (N_7274,N_572,N_2786);
nand U7275 (N_7275,N_1916,N_1834);
xnor U7276 (N_7276,N_4589,N_837);
nand U7277 (N_7277,N_2706,N_955);
or U7278 (N_7278,N_2436,N_2402);
or U7279 (N_7279,N_645,N_1169);
xor U7280 (N_7280,N_1745,N_3644);
or U7281 (N_7281,N_26,N_351);
nand U7282 (N_7282,N_4748,N_2701);
and U7283 (N_7283,N_3846,N_3421);
nor U7284 (N_7284,N_4434,N_2834);
xnor U7285 (N_7285,N_3774,N_3022);
and U7286 (N_7286,N_4430,N_588);
and U7287 (N_7287,N_4290,N_2973);
nand U7288 (N_7288,N_757,N_4311);
and U7289 (N_7289,N_1493,N_2038);
xnor U7290 (N_7290,N_1161,N_169);
nor U7291 (N_7291,N_2409,N_2809);
and U7292 (N_7292,N_3866,N_1274);
or U7293 (N_7293,N_222,N_762);
xnor U7294 (N_7294,N_2500,N_2740);
or U7295 (N_7295,N_4137,N_4301);
xor U7296 (N_7296,N_3070,N_1562);
xnor U7297 (N_7297,N_3893,N_4533);
or U7298 (N_7298,N_2718,N_2521);
nand U7299 (N_7299,N_354,N_1117);
nand U7300 (N_7300,N_1003,N_921);
and U7301 (N_7301,N_185,N_3903);
xnor U7302 (N_7302,N_4478,N_3757);
and U7303 (N_7303,N_4035,N_4561);
nand U7304 (N_7304,N_4306,N_3241);
and U7305 (N_7305,N_303,N_3508);
nand U7306 (N_7306,N_1699,N_2670);
and U7307 (N_7307,N_2978,N_4744);
or U7308 (N_7308,N_1996,N_3463);
nor U7309 (N_7309,N_371,N_1202);
and U7310 (N_7310,N_1609,N_1056);
xnor U7311 (N_7311,N_4448,N_90);
or U7312 (N_7312,N_4321,N_731);
xnor U7313 (N_7313,N_1579,N_1382);
nand U7314 (N_7314,N_913,N_3465);
and U7315 (N_7315,N_372,N_3501);
nand U7316 (N_7316,N_4665,N_3259);
and U7317 (N_7317,N_3766,N_4412);
nand U7318 (N_7318,N_1121,N_4110);
or U7319 (N_7319,N_4811,N_1137);
and U7320 (N_7320,N_1179,N_3995);
xnor U7321 (N_7321,N_4417,N_4157);
nand U7322 (N_7322,N_980,N_2880);
xnor U7323 (N_7323,N_2790,N_1259);
and U7324 (N_7324,N_2877,N_4716);
nand U7325 (N_7325,N_4176,N_3950);
xnor U7326 (N_7326,N_2080,N_668);
nor U7327 (N_7327,N_3370,N_718);
xor U7328 (N_7328,N_1022,N_2605);
and U7329 (N_7329,N_4573,N_4054);
nand U7330 (N_7330,N_1789,N_2932);
nor U7331 (N_7331,N_1948,N_1271);
or U7332 (N_7332,N_1670,N_1392);
nor U7333 (N_7333,N_855,N_998);
xnor U7334 (N_7334,N_309,N_2691);
nand U7335 (N_7335,N_320,N_2589);
and U7336 (N_7336,N_383,N_4605);
xor U7337 (N_7337,N_2912,N_3874);
and U7338 (N_7338,N_4809,N_3184);
or U7339 (N_7339,N_3829,N_3123);
xor U7340 (N_7340,N_3026,N_4411);
and U7341 (N_7341,N_805,N_4566);
and U7342 (N_7342,N_4514,N_1219);
and U7343 (N_7343,N_2692,N_3696);
xnor U7344 (N_7344,N_697,N_2082);
xnor U7345 (N_7345,N_1457,N_1846);
xor U7346 (N_7346,N_716,N_969);
and U7347 (N_7347,N_2353,N_4171);
nand U7348 (N_7348,N_1806,N_2174);
and U7349 (N_7349,N_4886,N_2340);
or U7350 (N_7350,N_2060,N_658);
nor U7351 (N_7351,N_1811,N_3336);
xor U7352 (N_7352,N_4586,N_298);
xnor U7353 (N_7353,N_3667,N_1604);
xnor U7354 (N_7354,N_4284,N_1311);
nor U7355 (N_7355,N_1932,N_3492);
nand U7356 (N_7356,N_929,N_3392);
or U7357 (N_7357,N_4887,N_2638);
nand U7358 (N_7358,N_1528,N_3112);
and U7359 (N_7359,N_2893,N_715);
and U7360 (N_7360,N_2653,N_3794);
nand U7361 (N_7361,N_2167,N_2429);
nor U7362 (N_7362,N_4957,N_636);
nand U7363 (N_7363,N_2755,N_4148);
or U7364 (N_7364,N_2280,N_2661);
xor U7365 (N_7365,N_1883,N_4324);
xor U7366 (N_7366,N_2851,N_2074);
nand U7367 (N_7367,N_1417,N_289);
nand U7368 (N_7368,N_479,N_1070);
xnor U7369 (N_7369,N_3090,N_4805);
xnor U7370 (N_7370,N_1134,N_450);
or U7371 (N_7371,N_3250,N_2223);
nand U7372 (N_7372,N_730,N_582);
nand U7373 (N_7373,N_867,N_4246);
and U7374 (N_7374,N_4663,N_1590);
xnor U7375 (N_7375,N_4444,N_293);
and U7376 (N_7376,N_3205,N_2027);
nor U7377 (N_7377,N_4011,N_1913);
nor U7378 (N_7378,N_3362,N_4938);
and U7379 (N_7379,N_979,N_4325);
nor U7380 (N_7380,N_3695,N_2610);
and U7381 (N_7381,N_3992,N_1824);
and U7382 (N_7382,N_4472,N_771);
nand U7383 (N_7383,N_899,N_2070);
and U7384 (N_7384,N_609,N_3037);
and U7385 (N_7385,N_4708,N_2564);
and U7386 (N_7386,N_1979,N_2024);
nor U7387 (N_7387,N_4253,N_703);
or U7388 (N_7388,N_1238,N_2592);
nand U7389 (N_7389,N_4109,N_583);
nor U7390 (N_7390,N_100,N_4203);
xor U7391 (N_7391,N_483,N_3099);
nor U7392 (N_7392,N_4906,N_4898);
nor U7393 (N_7393,N_464,N_3639);
nor U7394 (N_7394,N_3500,N_2411);
nor U7395 (N_7395,N_1143,N_1476);
nor U7396 (N_7396,N_1794,N_2805);
xor U7397 (N_7397,N_2110,N_3747);
or U7398 (N_7398,N_1632,N_171);
nor U7399 (N_7399,N_4319,N_1035);
xor U7400 (N_7400,N_1942,N_4262);
xor U7401 (N_7401,N_848,N_2773);
and U7402 (N_7402,N_4355,N_4473);
and U7403 (N_7403,N_4138,N_1917);
xnor U7404 (N_7404,N_4404,N_3941);
xnor U7405 (N_7405,N_1636,N_2852);
nand U7406 (N_7406,N_434,N_179);
nor U7407 (N_7407,N_397,N_2246);
xor U7408 (N_7408,N_3111,N_4443);
nor U7409 (N_7409,N_126,N_404);
nand U7410 (N_7410,N_4745,N_3495);
xnor U7411 (N_7411,N_1177,N_3924);
nor U7412 (N_7412,N_3071,N_1607);
xor U7413 (N_7413,N_1569,N_3426);
nand U7414 (N_7414,N_2408,N_237);
nor U7415 (N_7415,N_4307,N_4523);
nand U7416 (N_7416,N_4993,N_3142);
nor U7417 (N_7417,N_4127,N_62);
nor U7418 (N_7418,N_4063,N_4423);
nor U7419 (N_7419,N_3030,N_1626);
and U7420 (N_7420,N_2563,N_3346);
nand U7421 (N_7421,N_1053,N_4123);
xor U7422 (N_7422,N_1502,N_1945);
or U7423 (N_7423,N_957,N_2367);
nor U7424 (N_7424,N_364,N_3699);
and U7425 (N_7425,N_1987,N_3514);
xnor U7426 (N_7426,N_1720,N_3498);
nand U7427 (N_7427,N_3663,N_1992);
nand U7428 (N_7428,N_4544,N_48);
xnor U7429 (N_7429,N_3424,N_2333);
and U7430 (N_7430,N_902,N_3357);
or U7431 (N_7431,N_2248,N_511);
xnor U7432 (N_7432,N_2717,N_3764);
and U7433 (N_7433,N_2871,N_2357);
nand U7434 (N_7434,N_2781,N_4291);
and U7435 (N_7435,N_2886,N_467);
nor U7436 (N_7436,N_912,N_904);
nand U7437 (N_7437,N_4943,N_2719);
and U7438 (N_7438,N_4164,N_2140);
nor U7439 (N_7439,N_1593,N_3073);
nand U7440 (N_7440,N_2836,N_2318);
xor U7441 (N_7441,N_3871,N_3645);
or U7442 (N_7442,N_4145,N_408);
xor U7443 (N_7443,N_1405,N_2916);
and U7444 (N_7444,N_1191,N_1375);
or U7445 (N_7445,N_280,N_151);
or U7446 (N_7446,N_4651,N_3504);
nor U7447 (N_7447,N_84,N_4000);
and U7448 (N_7448,N_1560,N_3686);
or U7449 (N_7449,N_1698,N_374);
and U7450 (N_7450,N_4131,N_910);
nand U7451 (N_7451,N_4385,N_1661);
nand U7452 (N_7452,N_1094,N_1525);
or U7453 (N_7453,N_3422,N_627);
nand U7454 (N_7454,N_4250,N_2861);
xor U7455 (N_7455,N_200,N_3218);
xnor U7456 (N_7456,N_596,N_1145);
nand U7457 (N_7457,N_4576,N_2490);
xor U7458 (N_7458,N_1583,N_239);
nor U7459 (N_7459,N_3502,N_417);
nand U7460 (N_7460,N_3781,N_4193);
or U7461 (N_7461,N_112,N_2917);
xor U7462 (N_7462,N_4731,N_2017);
nor U7463 (N_7463,N_591,N_4303);
nor U7464 (N_7464,N_1746,N_1587);
nor U7465 (N_7465,N_2678,N_4204);
xor U7466 (N_7466,N_513,N_800);
xnor U7467 (N_7467,N_2729,N_4920);
nor U7468 (N_7468,N_1443,N_223);
or U7469 (N_7469,N_10,N_2749);
and U7470 (N_7470,N_2100,N_1909);
xnor U7471 (N_7471,N_512,N_3088);
nand U7472 (N_7472,N_522,N_4664);
nand U7473 (N_7473,N_2870,N_4043);
or U7474 (N_7474,N_3086,N_3806);
nor U7475 (N_7475,N_385,N_1195);
nand U7476 (N_7476,N_739,N_2317);
or U7477 (N_7477,N_1189,N_3162);
or U7478 (N_7478,N_2909,N_2312);
xor U7479 (N_7479,N_1563,N_462);
or U7480 (N_7480,N_3884,N_2890);
and U7481 (N_7481,N_2320,N_3845);
or U7482 (N_7482,N_2591,N_4916);
or U7483 (N_7483,N_466,N_3748);
nand U7484 (N_7484,N_4705,N_1033);
or U7485 (N_7485,N_3221,N_2468);
and U7486 (N_7486,N_2711,N_2268);
xor U7487 (N_7487,N_3404,N_173);
xor U7488 (N_7488,N_421,N_810);
or U7489 (N_7489,N_2957,N_3077);
xor U7490 (N_7490,N_1298,N_2470);
and U7491 (N_7491,N_3228,N_3889);
and U7492 (N_7492,N_1289,N_502);
or U7493 (N_7493,N_176,N_1778);
nand U7494 (N_7494,N_4013,N_1020);
or U7495 (N_7495,N_3029,N_3160);
and U7496 (N_7496,N_4565,N_4410);
xor U7497 (N_7497,N_2543,N_2626);
or U7498 (N_7498,N_4695,N_747);
nor U7499 (N_7499,N_2441,N_2899);
and U7500 (N_7500,N_4901,N_3572);
nor U7501 (N_7501,N_1153,N_2706);
nor U7502 (N_7502,N_1211,N_1472);
and U7503 (N_7503,N_1040,N_2198);
or U7504 (N_7504,N_711,N_2096);
or U7505 (N_7505,N_4923,N_4919);
xnor U7506 (N_7506,N_4238,N_1032);
nand U7507 (N_7507,N_2376,N_941);
or U7508 (N_7508,N_4604,N_2774);
or U7509 (N_7509,N_1586,N_2778);
or U7510 (N_7510,N_1346,N_4445);
xor U7511 (N_7511,N_304,N_481);
nand U7512 (N_7512,N_4611,N_552);
and U7513 (N_7513,N_423,N_1500);
nor U7514 (N_7514,N_1685,N_2009);
nand U7515 (N_7515,N_2950,N_4440);
nor U7516 (N_7516,N_2267,N_3554);
xnor U7517 (N_7517,N_2894,N_1665);
or U7518 (N_7518,N_3234,N_4414);
nor U7519 (N_7519,N_3948,N_2801);
nand U7520 (N_7520,N_1428,N_2055);
nor U7521 (N_7521,N_4944,N_2716);
nor U7522 (N_7522,N_3332,N_1570);
xor U7523 (N_7523,N_414,N_1645);
and U7524 (N_7524,N_2186,N_272);
or U7525 (N_7525,N_543,N_4232);
xor U7526 (N_7526,N_1507,N_4199);
or U7527 (N_7527,N_2959,N_1575);
and U7528 (N_7528,N_4622,N_3102);
or U7529 (N_7529,N_83,N_3281);
and U7530 (N_7530,N_4252,N_1399);
and U7531 (N_7531,N_3000,N_3624);
and U7532 (N_7532,N_4344,N_2494);
nand U7533 (N_7533,N_2341,N_878);
nor U7534 (N_7534,N_2401,N_1203);
nand U7535 (N_7535,N_430,N_1268);
nand U7536 (N_7536,N_4558,N_184);
nor U7537 (N_7537,N_2403,N_837);
and U7538 (N_7538,N_1475,N_1000);
and U7539 (N_7539,N_4241,N_2258);
nand U7540 (N_7540,N_4397,N_3446);
xnor U7541 (N_7541,N_4522,N_1833);
nor U7542 (N_7542,N_4119,N_4104);
and U7543 (N_7543,N_2601,N_737);
nor U7544 (N_7544,N_1661,N_3300);
nand U7545 (N_7545,N_648,N_1769);
and U7546 (N_7546,N_1506,N_2615);
or U7547 (N_7547,N_1813,N_1631);
nand U7548 (N_7548,N_3852,N_2690);
nor U7549 (N_7549,N_1671,N_1621);
and U7550 (N_7550,N_1352,N_4427);
and U7551 (N_7551,N_169,N_3011);
nand U7552 (N_7552,N_1345,N_3877);
or U7553 (N_7553,N_1958,N_2876);
xnor U7554 (N_7554,N_380,N_4009);
xnor U7555 (N_7555,N_4095,N_1972);
xnor U7556 (N_7556,N_3301,N_3019);
nand U7557 (N_7557,N_2668,N_1518);
xor U7558 (N_7558,N_2541,N_3250);
nor U7559 (N_7559,N_3909,N_3143);
xor U7560 (N_7560,N_79,N_143);
and U7561 (N_7561,N_634,N_4458);
or U7562 (N_7562,N_610,N_1480);
nor U7563 (N_7563,N_1610,N_1411);
and U7564 (N_7564,N_3739,N_1769);
nor U7565 (N_7565,N_3984,N_1377);
nand U7566 (N_7566,N_1049,N_3451);
and U7567 (N_7567,N_782,N_862);
xnor U7568 (N_7568,N_2130,N_4022);
nor U7569 (N_7569,N_3054,N_4470);
nor U7570 (N_7570,N_2192,N_4058);
or U7571 (N_7571,N_150,N_283);
nor U7572 (N_7572,N_3505,N_41);
nand U7573 (N_7573,N_182,N_3242);
nand U7574 (N_7574,N_1218,N_585);
and U7575 (N_7575,N_3918,N_938);
xor U7576 (N_7576,N_105,N_102);
nand U7577 (N_7577,N_3769,N_1877);
xor U7578 (N_7578,N_3454,N_3693);
or U7579 (N_7579,N_2925,N_3881);
or U7580 (N_7580,N_4743,N_1562);
nand U7581 (N_7581,N_128,N_1174);
and U7582 (N_7582,N_1541,N_4292);
or U7583 (N_7583,N_3945,N_2163);
nand U7584 (N_7584,N_2789,N_122);
or U7585 (N_7585,N_3052,N_4455);
or U7586 (N_7586,N_564,N_2969);
or U7587 (N_7587,N_1076,N_3793);
and U7588 (N_7588,N_1196,N_3994);
xor U7589 (N_7589,N_3368,N_4408);
nor U7590 (N_7590,N_228,N_4241);
xnor U7591 (N_7591,N_1767,N_4181);
or U7592 (N_7592,N_4784,N_3659);
nor U7593 (N_7593,N_4861,N_4679);
nand U7594 (N_7594,N_4016,N_2917);
nor U7595 (N_7595,N_1890,N_2753);
nand U7596 (N_7596,N_105,N_1373);
and U7597 (N_7597,N_103,N_4206);
xnor U7598 (N_7598,N_4789,N_2460);
and U7599 (N_7599,N_4458,N_1158);
and U7600 (N_7600,N_4905,N_862);
nand U7601 (N_7601,N_3712,N_1407);
or U7602 (N_7602,N_4928,N_1263);
nor U7603 (N_7603,N_3347,N_1501);
nor U7604 (N_7604,N_347,N_4286);
nand U7605 (N_7605,N_1950,N_2589);
nand U7606 (N_7606,N_1597,N_2589);
or U7607 (N_7607,N_1053,N_1504);
xnor U7608 (N_7608,N_1501,N_4839);
nand U7609 (N_7609,N_314,N_2886);
and U7610 (N_7610,N_4488,N_1338);
or U7611 (N_7611,N_1331,N_2619);
or U7612 (N_7612,N_2046,N_3032);
and U7613 (N_7613,N_2045,N_3542);
nor U7614 (N_7614,N_592,N_96);
or U7615 (N_7615,N_1928,N_4866);
nand U7616 (N_7616,N_3552,N_1729);
xnor U7617 (N_7617,N_227,N_1928);
xor U7618 (N_7618,N_2467,N_2749);
and U7619 (N_7619,N_3838,N_4886);
nor U7620 (N_7620,N_4932,N_2033);
nand U7621 (N_7621,N_694,N_812);
and U7622 (N_7622,N_2368,N_585);
xnor U7623 (N_7623,N_1903,N_3793);
or U7624 (N_7624,N_2881,N_689);
xnor U7625 (N_7625,N_621,N_2773);
or U7626 (N_7626,N_4590,N_2446);
nor U7627 (N_7627,N_2181,N_456);
and U7628 (N_7628,N_2733,N_3525);
and U7629 (N_7629,N_4234,N_3146);
or U7630 (N_7630,N_311,N_3720);
and U7631 (N_7631,N_3619,N_241);
xnor U7632 (N_7632,N_4237,N_2982);
or U7633 (N_7633,N_3568,N_1180);
nand U7634 (N_7634,N_1304,N_1267);
nand U7635 (N_7635,N_2892,N_337);
xnor U7636 (N_7636,N_3241,N_3908);
and U7637 (N_7637,N_748,N_475);
nand U7638 (N_7638,N_4542,N_301);
or U7639 (N_7639,N_384,N_4809);
or U7640 (N_7640,N_637,N_2832);
xnor U7641 (N_7641,N_158,N_4461);
nand U7642 (N_7642,N_3041,N_2035);
nor U7643 (N_7643,N_1753,N_3691);
or U7644 (N_7644,N_3101,N_2319);
nor U7645 (N_7645,N_4198,N_1073);
or U7646 (N_7646,N_2129,N_3789);
nand U7647 (N_7647,N_1642,N_659);
or U7648 (N_7648,N_614,N_2447);
and U7649 (N_7649,N_1921,N_4720);
nor U7650 (N_7650,N_3526,N_1523);
xor U7651 (N_7651,N_1391,N_822);
or U7652 (N_7652,N_1056,N_2355);
xnor U7653 (N_7653,N_845,N_387);
nor U7654 (N_7654,N_763,N_3932);
nand U7655 (N_7655,N_52,N_2070);
and U7656 (N_7656,N_1316,N_3854);
or U7657 (N_7657,N_2695,N_2959);
nor U7658 (N_7658,N_3294,N_3613);
nand U7659 (N_7659,N_3746,N_1322);
nand U7660 (N_7660,N_2722,N_927);
or U7661 (N_7661,N_2457,N_1000);
nor U7662 (N_7662,N_2810,N_4424);
and U7663 (N_7663,N_1303,N_790);
or U7664 (N_7664,N_4873,N_1091);
nand U7665 (N_7665,N_703,N_1128);
and U7666 (N_7666,N_3015,N_3129);
nor U7667 (N_7667,N_4998,N_3942);
nor U7668 (N_7668,N_1458,N_2716);
nand U7669 (N_7669,N_4185,N_1793);
and U7670 (N_7670,N_440,N_2477);
nand U7671 (N_7671,N_2073,N_874);
or U7672 (N_7672,N_2784,N_4770);
xor U7673 (N_7673,N_4774,N_4342);
or U7674 (N_7674,N_280,N_4152);
nand U7675 (N_7675,N_3797,N_730);
nor U7676 (N_7676,N_2002,N_4510);
nor U7677 (N_7677,N_2345,N_4405);
or U7678 (N_7678,N_102,N_2906);
and U7679 (N_7679,N_3391,N_703);
or U7680 (N_7680,N_279,N_1626);
and U7681 (N_7681,N_2366,N_4639);
xor U7682 (N_7682,N_1083,N_2408);
nand U7683 (N_7683,N_2331,N_2364);
and U7684 (N_7684,N_2704,N_3931);
xor U7685 (N_7685,N_2048,N_803);
and U7686 (N_7686,N_779,N_2380);
or U7687 (N_7687,N_541,N_3350);
or U7688 (N_7688,N_4936,N_4461);
and U7689 (N_7689,N_955,N_1282);
or U7690 (N_7690,N_1649,N_50);
and U7691 (N_7691,N_2696,N_3531);
nor U7692 (N_7692,N_954,N_503);
xnor U7693 (N_7693,N_513,N_739);
or U7694 (N_7694,N_2642,N_1540);
and U7695 (N_7695,N_4955,N_3712);
or U7696 (N_7696,N_3969,N_4158);
nor U7697 (N_7697,N_4984,N_368);
nand U7698 (N_7698,N_2875,N_134);
xor U7699 (N_7699,N_2933,N_2413);
nand U7700 (N_7700,N_4627,N_3360);
and U7701 (N_7701,N_1854,N_441);
and U7702 (N_7702,N_1278,N_2976);
nand U7703 (N_7703,N_1076,N_2260);
nand U7704 (N_7704,N_645,N_4336);
and U7705 (N_7705,N_3459,N_2713);
or U7706 (N_7706,N_4414,N_4650);
or U7707 (N_7707,N_87,N_3376);
nor U7708 (N_7708,N_1753,N_1796);
nor U7709 (N_7709,N_114,N_1039);
or U7710 (N_7710,N_1762,N_2078);
nand U7711 (N_7711,N_2216,N_2220);
and U7712 (N_7712,N_642,N_4313);
xor U7713 (N_7713,N_481,N_993);
nand U7714 (N_7714,N_444,N_4102);
nor U7715 (N_7715,N_2601,N_2137);
xnor U7716 (N_7716,N_4030,N_4172);
and U7717 (N_7717,N_1382,N_245);
xnor U7718 (N_7718,N_3341,N_828);
nor U7719 (N_7719,N_2922,N_2833);
or U7720 (N_7720,N_98,N_4103);
or U7721 (N_7721,N_4507,N_4614);
nand U7722 (N_7722,N_682,N_2863);
nor U7723 (N_7723,N_3810,N_2115);
nand U7724 (N_7724,N_3173,N_651);
and U7725 (N_7725,N_2821,N_424);
or U7726 (N_7726,N_82,N_4436);
and U7727 (N_7727,N_3629,N_4443);
nor U7728 (N_7728,N_3594,N_467);
or U7729 (N_7729,N_3858,N_4526);
and U7730 (N_7730,N_4183,N_3000);
or U7731 (N_7731,N_227,N_1863);
and U7732 (N_7732,N_4746,N_3097);
nor U7733 (N_7733,N_4238,N_2382);
xnor U7734 (N_7734,N_2297,N_2322);
or U7735 (N_7735,N_1935,N_4343);
xnor U7736 (N_7736,N_493,N_4998);
nand U7737 (N_7737,N_1711,N_2218);
nand U7738 (N_7738,N_292,N_4658);
nor U7739 (N_7739,N_1505,N_1376);
or U7740 (N_7740,N_2025,N_1736);
or U7741 (N_7741,N_4900,N_4964);
nand U7742 (N_7742,N_1873,N_1982);
and U7743 (N_7743,N_1615,N_2647);
xor U7744 (N_7744,N_1352,N_4591);
xor U7745 (N_7745,N_921,N_4171);
or U7746 (N_7746,N_3830,N_1881);
and U7747 (N_7747,N_2742,N_3677);
or U7748 (N_7748,N_3969,N_29);
xnor U7749 (N_7749,N_584,N_3249);
xnor U7750 (N_7750,N_2734,N_3039);
xnor U7751 (N_7751,N_4954,N_1456);
nor U7752 (N_7752,N_1784,N_403);
or U7753 (N_7753,N_4982,N_3744);
nor U7754 (N_7754,N_1472,N_2545);
and U7755 (N_7755,N_3348,N_3434);
xor U7756 (N_7756,N_1914,N_3883);
or U7757 (N_7757,N_3727,N_3435);
nand U7758 (N_7758,N_358,N_2773);
nand U7759 (N_7759,N_642,N_436);
or U7760 (N_7760,N_3496,N_3319);
xnor U7761 (N_7761,N_3851,N_689);
or U7762 (N_7762,N_2485,N_905);
xor U7763 (N_7763,N_1991,N_865);
xor U7764 (N_7764,N_4517,N_687);
or U7765 (N_7765,N_1181,N_255);
nor U7766 (N_7766,N_114,N_632);
or U7767 (N_7767,N_715,N_2292);
or U7768 (N_7768,N_2427,N_3151);
nand U7769 (N_7769,N_3771,N_2450);
nor U7770 (N_7770,N_4821,N_3059);
nand U7771 (N_7771,N_4249,N_393);
and U7772 (N_7772,N_1110,N_3307);
or U7773 (N_7773,N_221,N_1915);
xor U7774 (N_7774,N_2769,N_767);
nor U7775 (N_7775,N_1325,N_3669);
or U7776 (N_7776,N_1174,N_3444);
or U7777 (N_7777,N_883,N_204);
nand U7778 (N_7778,N_2119,N_2883);
nand U7779 (N_7779,N_1451,N_4290);
nor U7780 (N_7780,N_1839,N_4806);
nor U7781 (N_7781,N_489,N_587);
nor U7782 (N_7782,N_2217,N_2894);
xnor U7783 (N_7783,N_172,N_279);
nor U7784 (N_7784,N_506,N_4819);
xor U7785 (N_7785,N_3779,N_1916);
nand U7786 (N_7786,N_2565,N_3032);
nor U7787 (N_7787,N_3323,N_3390);
xnor U7788 (N_7788,N_1426,N_4668);
xor U7789 (N_7789,N_999,N_4026);
nor U7790 (N_7790,N_3557,N_2805);
nand U7791 (N_7791,N_1007,N_2322);
nand U7792 (N_7792,N_1116,N_3728);
and U7793 (N_7793,N_3962,N_2595);
and U7794 (N_7794,N_4939,N_1420);
nor U7795 (N_7795,N_1647,N_210);
xnor U7796 (N_7796,N_4087,N_1120);
or U7797 (N_7797,N_306,N_588);
and U7798 (N_7798,N_671,N_1630);
nand U7799 (N_7799,N_3195,N_186);
xor U7800 (N_7800,N_4062,N_2826);
or U7801 (N_7801,N_1874,N_3110);
nor U7802 (N_7802,N_768,N_3678);
nor U7803 (N_7803,N_3650,N_3787);
nor U7804 (N_7804,N_4632,N_2187);
or U7805 (N_7805,N_1977,N_4488);
or U7806 (N_7806,N_4736,N_766);
nand U7807 (N_7807,N_1239,N_2076);
or U7808 (N_7808,N_1000,N_3591);
xor U7809 (N_7809,N_1764,N_1021);
xnor U7810 (N_7810,N_2889,N_2941);
nor U7811 (N_7811,N_2533,N_381);
nor U7812 (N_7812,N_2277,N_2423);
or U7813 (N_7813,N_4869,N_1021);
and U7814 (N_7814,N_3492,N_2941);
xnor U7815 (N_7815,N_3249,N_3002);
nor U7816 (N_7816,N_1141,N_3620);
or U7817 (N_7817,N_1574,N_1083);
or U7818 (N_7818,N_76,N_2663);
and U7819 (N_7819,N_1297,N_319);
nand U7820 (N_7820,N_2520,N_3377);
nor U7821 (N_7821,N_502,N_3226);
or U7822 (N_7822,N_3526,N_4322);
and U7823 (N_7823,N_4336,N_3950);
and U7824 (N_7824,N_2231,N_1707);
nand U7825 (N_7825,N_1732,N_1481);
or U7826 (N_7826,N_4528,N_106);
xor U7827 (N_7827,N_2789,N_3472);
xnor U7828 (N_7828,N_888,N_4307);
or U7829 (N_7829,N_890,N_1155);
xor U7830 (N_7830,N_4500,N_4411);
nand U7831 (N_7831,N_3907,N_2399);
or U7832 (N_7832,N_2283,N_473);
nor U7833 (N_7833,N_4931,N_4947);
xor U7834 (N_7834,N_2638,N_3388);
nand U7835 (N_7835,N_777,N_3759);
nor U7836 (N_7836,N_4369,N_3813);
xor U7837 (N_7837,N_3574,N_4992);
nand U7838 (N_7838,N_1096,N_2255);
xnor U7839 (N_7839,N_827,N_2109);
and U7840 (N_7840,N_4256,N_1486);
nand U7841 (N_7841,N_4394,N_222);
xor U7842 (N_7842,N_1792,N_218);
nand U7843 (N_7843,N_1869,N_4612);
nand U7844 (N_7844,N_974,N_2567);
or U7845 (N_7845,N_4674,N_3696);
or U7846 (N_7846,N_2977,N_3456);
xnor U7847 (N_7847,N_626,N_1676);
xnor U7848 (N_7848,N_1282,N_2812);
nor U7849 (N_7849,N_2070,N_700);
or U7850 (N_7850,N_3956,N_2662);
or U7851 (N_7851,N_561,N_1972);
or U7852 (N_7852,N_369,N_135);
xnor U7853 (N_7853,N_1843,N_643);
nand U7854 (N_7854,N_152,N_2596);
and U7855 (N_7855,N_2820,N_1909);
and U7856 (N_7856,N_2904,N_3828);
and U7857 (N_7857,N_539,N_4542);
xnor U7858 (N_7858,N_2505,N_3580);
and U7859 (N_7859,N_1303,N_2892);
xnor U7860 (N_7860,N_1225,N_539);
nand U7861 (N_7861,N_712,N_163);
nor U7862 (N_7862,N_4828,N_4267);
and U7863 (N_7863,N_2856,N_2326);
xor U7864 (N_7864,N_2978,N_2951);
and U7865 (N_7865,N_3240,N_1467);
xor U7866 (N_7866,N_120,N_1248);
or U7867 (N_7867,N_438,N_2003);
or U7868 (N_7868,N_1773,N_3587);
nand U7869 (N_7869,N_674,N_4274);
nor U7870 (N_7870,N_4392,N_2452);
nand U7871 (N_7871,N_328,N_1421);
xnor U7872 (N_7872,N_402,N_252);
and U7873 (N_7873,N_1578,N_2494);
nand U7874 (N_7874,N_2055,N_1388);
nand U7875 (N_7875,N_4994,N_683);
or U7876 (N_7876,N_4907,N_2071);
and U7877 (N_7877,N_3248,N_4897);
nand U7878 (N_7878,N_3353,N_1368);
nand U7879 (N_7879,N_3795,N_1764);
nand U7880 (N_7880,N_2568,N_2404);
xor U7881 (N_7881,N_1248,N_1968);
xor U7882 (N_7882,N_1435,N_1930);
or U7883 (N_7883,N_4738,N_4570);
nor U7884 (N_7884,N_239,N_3194);
or U7885 (N_7885,N_3735,N_3534);
xnor U7886 (N_7886,N_856,N_2748);
nor U7887 (N_7887,N_1193,N_4528);
nand U7888 (N_7888,N_2910,N_2789);
or U7889 (N_7889,N_4800,N_2631);
or U7890 (N_7890,N_2182,N_4042);
xor U7891 (N_7891,N_2070,N_3252);
nor U7892 (N_7892,N_3109,N_2966);
or U7893 (N_7893,N_482,N_4733);
xor U7894 (N_7894,N_2941,N_4346);
nor U7895 (N_7895,N_1610,N_929);
xor U7896 (N_7896,N_4891,N_4984);
xnor U7897 (N_7897,N_1039,N_2821);
and U7898 (N_7898,N_1977,N_3898);
xnor U7899 (N_7899,N_2690,N_2190);
or U7900 (N_7900,N_168,N_1754);
xor U7901 (N_7901,N_3783,N_643);
nand U7902 (N_7902,N_1116,N_3579);
nand U7903 (N_7903,N_2292,N_1118);
and U7904 (N_7904,N_2571,N_4357);
or U7905 (N_7905,N_1738,N_2070);
nand U7906 (N_7906,N_4215,N_168);
xnor U7907 (N_7907,N_3026,N_1405);
and U7908 (N_7908,N_4387,N_4394);
or U7909 (N_7909,N_104,N_2693);
nor U7910 (N_7910,N_2318,N_588);
xnor U7911 (N_7911,N_4629,N_454);
and U7912 (N_7912,N_3324,N_4552);
nand U7913 (N_7913,N_458,N_259);
xnor U7914 (N_7914,N_3217,N_3886);
or U7915 (N_7915,N_2585,N_1910);
nor U7916 (N_7916,N_2489,N_4195);
or U7917 (N_7917,N_2084,N_2661);
and U7918 (N_7918,N_1082,N_928);
nand U7919 (N_7919,N_363,N_3334);
xor U7920 (N_7920,N_530,N_337);
nand U7921 (N_7921,N_220,N_1290);
or U7922 (N_7922,N_3048,N_189);
xor U7923 (N_7923,N_972,N_1713);
xor U7924 (N_7924,N_4491,N_2437);
nor U7925 (N_7925,N_3017,N_3061);
nand U7926 (N_7926,N_2908,N_1826);
or U7927 (N_7927,N_1038,N_2939);
xnor U7928 (N_7928,N_3304,N_2492);
or U7929 (N_7929,N_2525,N_1197);
nand U7930 (N_7930,N_2593,N_2520);
nor U7931 (N_7931,N_2678,N_906);
xor U7932 (N_7932,N_4293,N_2530);
or U7933 (N_7933,N_1684,N_1906);
nor U7934 (N_7934,N_3086,N_1125);
or U7935 (N_7935,N_4058,N_2577);
or U7936 (N_7936,N_2153,N_1933);
or U7937 (N_7937,N_4471,N_3295);
xor U7938 (N_7938,N_2405,N_3623);
and U7939 (N_7939,N_1291,N_3580);
and U7940 (N_7940,N_1232,N_4099);
nor U7941 (N_7941,N_1874,N_3362);
xor U7942 (N_7942,N_1791,N_293);
xnor U7943 (N_7943,N_227,N_4453);
or U7944 (N_7944,N_1333,N_943);
nor U7945 (N_7945,N_4081,N_2792);
nor U7946 (N_7946,N_4196,N_644);
or U7947 (N_7947,N_2088,N_752);
nor U7948 (N_7948,N_4416,N_110);
xnor U7949 (N_7949,N_1553,N_3167);
and U7950 (N_7950,N_4415,N_22);
nand U7951 (N_7951,N_1778,N_1882);
nand U7952 (N_7952,N_838,N_2180);
nand U7953 (N_7953,N_3738,N_708);
nor U7954 (N_7954,N_661,N_380);
xnor U7955 (N_7955,N_3422,N_1124);
xor U7956 (N_7956,N_3477,N_3324);
nand U7957 (N_7957,N_139,N_4233);
or U7958 (N_7958,N_1370,N_3142);
nand U7959 (N_7959,N_3302,N_3623);
xor U7960 (N_7960,N_3012,N_3415);
nor U7961 (N_7961,N_785,N_2656);
or U7962 (N_7962,N_993,N_2514);
nand U7963 (N_7963,N_2009,N_3372);
or U7964 (N_7964,N_1503,N_3628);
nor U7965 (N_7965,N_3162,N_135);
and U7966 (N_7966,N_557,N_4186);
or U7967 (N_7967,N_497,N_2976);
and U7968 (N_7968,N_460,N_2786);
or U7969 (N_7969,N_56,N_3932);
and U7970 (N_7970,N_1734,N_1793);
nor U7971 (N_7971,N_3641,N_3747);
and U7972 (N_7972,N_2002,N_630);
nor U7973 (N_7973,N_1784,N_2434);
nor U7974 (N_7974,N_4545,N_3056);
or U7975 (N_7975,N_1233,N_1171);
xor U7976 (N_7976,N_2143,N_2647);
or U7977 (N_7977,N_3252,N_1041);
xnor U7978 (N_7978,N_4851,N_3694);
nand U7979 (N_7979,N_2033,N_4962);
nand U7980 (N_7980,N_4330,N_1025);
xnor U7981 (N_7981,N_3575,N_3615);
or U7982 (N_7982,N_2754,N_1685);
nor U7983 (N_7983,N_2924,N_1435);
and U7984 (N_7984,N_4,N_2655);
xnor U7985 (N_7985,N_3556,N_4236);
or U7986 (N_7986,N_2311,N_1364);
nor U7987 (N_7987,N_796,N_2248);
nand U7988 (N_7988,N_1491,N_3182);
or U7989 (N_7989,N_4523,N_2075);
or U7990 (N_7990,N_4537,N_827);
nor U7991 (N_7991,N_4891,N_349);
nand U7992 (N_7992,N_4550,N_819);
and U7993 (N_7993,N_3478,N_2611);
nor U7994 (N_7994,N_2228,N_1377);
nor U7995 (N_7995,N_1886,N_3141);
xor U7996 (N_7996,N_3155,N_423);
or U7997 (N_7997,N_587,N_3152);
nand U7998 (N_7998,N_4305,N_4021);
nor U7999 (N_7999,N_2900,N_2004);
nand U8000 (N_8000,N_3089,N_3200);
nor U8001 (N_8001,N_166,N_3002);
and U8002 (N_8002,N_2065,N_2273);
nand U8003 (N_8003,N_180,N_2759);
or U8004 (N_8004,N_1562,N_90);
and U8005 (N_8005,N_4206,N_1343);
nor U8006 (N_8006,N_2562,N_4585);
or U8007 (N_8007,N_2975,N_1131);
xor U8008 (N_8008,N_4753,N_1570);
nand U8009 (N_8009,N_475,N_3459);
and U8010 (N_8010,N_1653,N_143);
or U8011 (N_8011,N_2980,N_2185);
nor U8012 (N_8012,N_2517,N_1295);
nand U8013 (N_8013,N_3545,N_4380);
xor U8014 (N_8014,N_2767,N_3641);
and U8015 (N_8015,N_2610,N_4059);
or U8016 (N_8016,N_4916,N_1365);
or U8017 (N_8017,N_4506,N_3819);
nor U8018 (N_8018,N_806,N_3478);
or U8019 (N_8019,N_424,N_3648);
or U8020 (N_8020,N_3011,N_3702);
nand U8021 (N_8021,N_1862,N_410);
nor U8022 (N_8022,N_4010,N_4074);
or U8023 (N_8023,N_3210,N_184);
nor U8024 (N_8024,N_3376,N_659);
nand U8025 (N_8025,N_4941,N_848);
and U8026 (N_8026,N_253,N_2526);
xor U8027 (N_8027,N_2716,N_4288);
nor U8028 (N_8028,N_3330,N_3146);
and U8029 (N_8029,N_3203,N_1082);
nand U8030 (N_8030,N_923,N_2312);
and U8031 (N_8031,N_4324,N_695);
and U8032 (N_8032,N_50,N_4985);
or U8033 (N_8033,N_3131,N_885);
xnor U8034 (N_8034,N_1075,N_3054);
nor U8035 (N_8035,N_2848,N_3261);
and U8036 (N_8036,N_1252,N_4124);
or U8037 (N_8037,N_4278,N_1099);
and U8038 (N_8038,N_4077,N_3085);
nand U8039 (N_8039,N_747,N_2788);
nor U8040 (N_8040,N_2672,N_2044);
nor U8041 (N_8041,N_3760,N_835);
nand U8042 (N_8042,N_4936,N_3136);
nor U8043 (N_8043,N_1465,N_3679);
nand U8044 (N_8044,N_2259,N_865);
and U8045 (N_8045,N_3282,N_1973);
xor U8046 (N_8046,N_713,N_1615);
and U8047 (N_8047,N_257,N_1292);
nand U8048 (N_8048,N_44,N_2621);
or U8049 (N_8049,N_3075,N_1843);
nor U8050 (N_8050,N_2355,N_4606);
and U8051 (N_8051,N_4620,N_3226);
and U8052 (N_8052,N_2415,N_2321);
and U8053 (N_8053,N_4369,N_4497);
nor U8054 (N_8054,N_3298,N_323);
or U8055 (N_8055,N_1273,N_1733);
xnor U8056 (N_8056,N_3669,N_1333);
nand U8057 (N_8057,N_3109,N_1100);
xnor U8058 (N_8058,N_3475,N_2894);
and U8059 (N_8059,N_2887,N_138);
or U8060 (N_8060,N_862,N_920);
nand U8061 (N_8061,N_884,N_1057);
xor U8062 (N_8062,N_2649,N_3332);
nor U8063 (N_8063,N_591,N_374);
nor U8064 (N_8064,N_4402,N_1091);
nor U8065 (N_8065,N_1605,N_4784);
xor U8066 (N_8066,N_3286,N_947);
xor U8067 (N_8067,N_973,N_1575);
or U8068 (N_8068,N_1896,N_4098);
nand U8069 (N_8069,N_318,N_357);
or U8070 (N_8070,N_4960,N_1027);
nand U8071 (N_8071,N_1141,N_2022);
xor U8072 (N_8072,N_709,N_1399);
or U8073 (N_8073,N_3838,N_208);
xnor U8074 (N_8074,N_58,N_372);
nand U8075 (N_8075,N_782,N_3088);
and U8076 (N_8076,N_1481,N_1150);
nand U8077 (N_8077,N_2436,N_3509);
and U8078 (N_8078,N_4698,N_63);
or U8079 (N_8079,N_39,N_3211);
and U8080 (N_8080,N_1694,N_960);
xnor U8081 (N_8081,N_2055,N_3892);
or U8082 (N_8082,N_4749,N_4881);
nor U8083 (N_8083,N_4385,N_1793);
nand U8084 (N_8084,N_3608,N_4722);
nand U8085 (N_8085,N_4314,N_132);
or U8086 (N_8086,N_2331,N_4928);
and U8087 (N_8087,N_4497,N_358);
and U8088 (N_8088,N_2768,N_4030);
nor U8089 (N_8089,N_3790,N_2131);
or U8090 (N_8090,N_3420,N_1565);
and U8091 (N_8091,N_2748,N_3672);
or U8092 (N_8092,N_3555,N_72);
or U8093 (N_8093,N_600,N_1409);
nand U8094 (N_8094,N_471,N_1418);
or U8095 (N_8095,N_3188,N_2071);
or U8096 (N_8096,N_3985,N_2083);
xor U8097 (N_8097,N_4224,N_3134);
xnor U8098 (N_8098,N_2297,N_1255);
nor U8099 (N_8099,N_4330,N_86);
xor U8100 (N_8100,N_4358,N_3928);
or U8101 (N_8101,N_2449,N_4273);
xnor U8102 (N_8102,N_539,N_2728);
and U8103 (N_8103,N_880,N_3393);
xnor U8104 (N_8104,N_4658,N_912);
nor U8105 (N_8105,N_4446,N_1426);
xor U8106 (N_8106,N_464,N_2490);
xor U8107 (N_8107,N_3207,N_4525);
nand U8108 (N_8108,N_131,N_2853);
nand U8109 (N_8109,N_778,N_1575);
nand U8110 (N_8110,N_4907,N_4197);
or U8111 (N_8111,N_4247,N_1385);
nand U8112 (N_8112,N_589,N_2966);
and U8113 (N_8113,N_3057,N_275);
and U8114 (N_8114,N_3836,N_2972);
and U8115 (N_8115,N_4577,N_883);
and U8116 (N_8116,N_650,N_1364);
or U8117 (N_8117,N_748,N_3265);
nor U8118 (N_8118,N_773,N_662);
nor U8119 (N_8119,N_3379,N_4208);
and U8120 (N_8120,N_3877,N_1360);
nor U8121 (N_8121,N_2276,N_400);
xnor U8122 (N_8122,N_4633,N_4820);
nor U8123 (N_8123,N_3301,N_2110);
or U8124 (N_8124,N_4057,N_4799);
nand U8125 (N_8125,N_2125,N_2745);
nand U8126 (N_8126,N_1141,N_2878);
nor U8127 (N_8127,N_4845,N_140);
nor U8128 (N_8128,N_4405,N_1517);
and U8129 (N_8129,N_1785,N_2719);
and U8130 (N_8130,N_4262,N_3649);
nor U8131 (N_8131,N_1075,N_2887);
and U8132 (N_8132,N_4317,N_1659);
nor U8133 (N_8133,N_2772,N_4829);
and U8134 (N_8134,N_494,N_2602);
and U8135 (N_8135,N_2288,N_2518);
xnor U8136 (N_8136,N_161,N_216);
xor U8137 (N_8137,N_2481,N_496);
xor U8138 (N_8138,N_2133,N_2332);
or U8139 (N_8139,N_4661,N_4151);
xor U8140 (N_8140,N_2946,N_4731);
xnor U8141 (N_8141,N_4613,N_4517);
xnor U8142 (N_8142,N_2224,N_2090);
nand U8143 (N_8143,N_1217,N_4149);
nor U8144 (N_8144,N_1428,N_1389);
xnor U8145 (N_8145,N_2124,N_1431);
and U8146 (N_8146,N_3619,N_3865);
or U8147 (N_8147,N_37,N_1427);
and U8148 (N_8148,N_1354,N_533);
and U8149 (N_8149,N_898,N_4702);
xor U8150 (N_8150,N_1618,N_4072);
or U8151 (N_8151,N_2261,N_1209);
xor U8152 (N_8152,N_3440,N_803);
xor U8153 (N_8153,N_946,N_4770);
and U8154 (N_8154,N_3756,N_3513);
and U8155 (N_8155,N_2736,N_3544);
xor U8156 (N_8156,N_3884,N_4463);
nand U8157 (N_8157,N_4460,N_4471);
or U8158 (N_8158,N_4191,N_3045);
or U8159 (N_8159,N_2474,N_20);
xor U8160 (N_8160,N_3243,N_3681);
or U8161 (N_8161,N_3097,N_863);
nand U8162 (N_8162,N_4236,N_2280);
or U8163 (N_8163,N_4374,N_4189);
nand U8164 (N_8164,N_4073,N_3690);
or U8165 (N_8165,N_1613,N_2371);
or U8166 (N_8166,N_3609,N_3151);
or U8167 (N_8167,N_2284,N_1756);
or U8168 (N_8168,N_2961,N_1196);
nor U8169 (N_8169,N_3844,N_3148);
and U8170 (N_8170,N_232,N_4654);
nor U8171 (N_8171,N_1196,N_4349);
nor U8172 (N_8172,N_3908,N_681);
nand U8173 (N_8173,N_4102,N_3996);
or U8174 (N_8174,N_3754,N_3871);
nand U8175 (N_8175,N_4091,N_1862);
and U8176 (N_8176,N_131,N_2325);
and U8177 (N_8177,N_3667,N_2336);
nor U8178 (N_8178,N_632,N_564);
nor U8179 (N_8179,N_3501,N_1961);
and U8180 (N_8180,N_4789,N_689);
xor U8181 (N_8181,N_1585,N_950);
and U8182 (N_8182,N_3412,N_1654);
or U8183 (N_8183,N_86,N_3552);
xnor U8184 (N_8184,N_1969,N_1204);
or U8185 (N_8185,N_2017,N_3414);
nand U8186 (N_8186,N_4007,N_719);
or U8187 (N_8187,N_20,N_1655);
xor U8188 (N_8188,N_4543,N_4833);
nand U8189 (N_8189,N_4075,N_4876);
xor U8190 (N_8190,N_4653,N_3805);
xor U8191 (N_8191,N_4075,N_3393);
nand U8192 (N_8192,N_1007,N_1928);
nand U8193 (N_8193,N_441,N_1842);
xnor U8194 (N_8194,N_4885,N_778);
nand U8195 (N_8195,N_2934,N_3971);
nand U8196 (N_8196,N_3059,N_4505);
nor U8197 (N_8197,N_3885,N_4475);
nand U8198 (N_8198,N_808,N_4499);
or U8199 (N_8199,N_4147,N_3069);
and U8200 (N_8200,N_4051,N_1490);
nor U8201 (N_8201,N_4081,N_3648);
or U8202 (N_8202,N_4473,N_751);
xnor U8203 (N_8203,N_3277,N_297);
nand U8204 (N_8204,N_1950,N_2980);
nor U8205 (N_8205,N_90,N_2617);
nor U8206 (N_8206,N_77,N_1715);
or U8207 (N_8207,N_216,N_664);
nand U8208 (N_8208,N_4488,N_4475);
nor U8209 (N_8209,N_4337,N_1221);
nor U8210 (N_8210,N_985,N_1952);
xor U8211 (N_8211,N_1778,N_3003);
nor U8212 (N_8212,N_3354,N_4070);
and U8213 (N_8213,N_4697,N_2505);
nand U8214 (N_8214,N_1423,N_313);
and U8215 (N_8215,N_213,N_969);
nand U8216 (N_8216,N_3591,N_4780);
nor U8217 (N_8217,N_1913,N_4019);
nor U8218 (N_8218,N_875,N_849);
and U8219 (N_8219,N_3984,N_3444);
nor U8220 (N_8220,N_3314,N_1213);
nand U8221 (N_8221,N_4991,N_2910);
or U8222 (N_8222,N_328,N_1402);
nand U8223 (N_8223,N_4189,N_211);
nand U8224 (N_8224,N_3156,N_3056);
and U8225 (N_8225,N_633,N_916);
xnor U8226 (N_8226,N_4800,N_3468);
xnor U8227 (N_8227,N_2120,N_4849);
xnor U8228 (N_8228,N_888,N_3871);
nor U8229 (N_8229,N_4618,N_3233);
nand U8230 (N_8230,N_1534,N_4267);
and U8231 (N_8231,N_2453,N_3333);
and U8232 (N_8232,N_2142,N_1676);
nor U8233 (N_8233,N_1211,N_1540);
or U8234 (N_8234,N_2142,N_2979);
xnor U8235 (N_8235,N_4873,N_4161);
nor U8236 (N_8236,N_3219,N_3933);
nand U8237 (N_8237,N_985,N_267);
nor U8238 (N_8238,N_1048,N_329);
nand U8239 (N_8239,N_3190,N_1107);
xnor U8240 (N_8240,N_2854,N_3577);
nand U8241 (N_8241,N_2024,N_1342);
nand U8242 (N_8242,N_1321,N_3611);
nand U8243 (N_8243,N_4133,N_164);
xnor U8244 (N_8244,N_2729,N_1230);
nand U8245 (N_8245,N_1680,N_1326);
or U8246 (N_8246,N_4671,N_4175);
or U8247 (N_8247,N_3668,N_168);
xnor U8248 (N_8248,N_4531,N_4144);
xor U8249 (N_8249,N_1575,N_4733);
or U8250 (N_8250,N_3701,N_1776);
xnor U8251 (N_8251,N_1699,N_4567);
nand U8252 (N_8252,N_3057,N_1543);
or U8253 (N_8253,N_2536,N_794);
nand U8254 (N_8254,N_3349,N_730);
and U8255 (N_8255,N_3323,N_2885);
or U8256 (N_8256,N_2563,N_1202);
and U8257 (N_8257,N_4477,N_517);
xnor U8258 (N_8258,N_2488,N_307);
or U8259 (N_8259,N_1535,N_2331);
nor U8260 (N_8260,N_1306,N_580);
or U8261 (N_8261,N_3957,N_4753);
nor U8262 (N_8262,N_1087,N_347);
nand U8263 (N_8263,N_1098,N_694);
xor U8264 (N_8264,N_2553,N_1475);
nor U8265 (N_8265,N_2348,N_2458);
or U8266 (N_8266,N_4927,N_4005);
nand U8267 (N_8267,N_2237,N_4578);
and U8268 (N_8268,N_247,N_3877);
or U8269 (N_8269,N_1824,N_4735);
xnor U8270 (N_8270,N_3067,N_4549);
or U8271 (N_8271,N_3616,N_1416);
or U8272 (N_8272,N_713,N_4600);
and U8273 (N_8273,N_3807,N_4710);
or U8274 (N_8274,N_2123,N_3268);
nor U8275 (N_8275,N_4563,N_4391);
xor U8276 (N_8276,N_1268,N_3401);
nor U8277 (N_8277,N_3855,N_1984);
and U8278 (N_8278,N_4308,N_3105);
or U8279 (N_8279,N_169,N_3619);
or U8280 (N_8280,N_3899,N_1920);
or U8281 (N_8281,N_319,N_3912);
xnor U8282 (N_8282,N_2911,N_4099);
or U8283 (N_8283,N_1555,N_1158);
or U8284 (N_8284,N_1909,N_4332);
or U8285 (N_8285,N_3413,N_1926);
nor U8286 (N_8286,N_1336,N_929);
and U8287 (N_8287,N_307,N_531);
and U8288 (N_8288,N_4093,N_699);
nand U8289 (N_8289,N_1000,N_2170);
nor U8290 (N_8290,N_2107,N_4264);
nand U8291 (N_8291,N_4427,N_3512);
xor U8292 (N_8292,N_2620,N_1248);
nor U8293 (N_8293,N_3850,N_604);
or U8294 (N_8294,N_1994,N_4532);
and U8295 (N_8295,N_1045,N_4175);
nand U8296 (N_8296,N_1435,N_2982);
xor U8297 (N_8297,N_3774,N_3282);
xor U8298 (N_8298,N_4528,N_2661);
and U8299 (N_8299,N_3979,N_313);
nand U8300 (N_8300,N_3875,N_3098);
xnor U8301 (N_8301,N_4801,N_4462);
nor U8302 (N_8302,N_1379,N_1431);
and U8303 (N_8303,N_891,N_1643);
nand U8304 (N_8304,N_1995,N_4322);
or U8305 (N_8305,N_3855,N_3146);
nand U8306 (N_8306,N_2592,N_4212);
nor U8307 (N_8307,N_3377,N_794);
and U8308 (N_8308,N_3032,N_3955);
or U8309 (N_8309,N_89,N_4838);
and U8310 (N_8310,N_4169,N_4714);
nand U8311 (N_8311,N_1949,N_4744);
or U8312 (N_8312,N_1335,N_3844);
nor U8313 (N_8313,N_569,N_4072);
xnor U8314 (N_8314,N_1122,N_3895);
xor U8315 (N_8315,N_539,N_2450);
nand U8316 (N_8316,N_4433,N_1791);
nand U8317 (N_8317,N_3440,N_464);
xor U8318 (N_8318,N_2785,N_2840);
nor U8319 (N_8319,N_2022,N_3873);
nand U8320 (N_8320,N_144,N_3749);
and U8321 (N_8321,N_4622,N_731);
xnor U8322 (N_8322,N_2054,N_4694);
nor U8323 (N_8323,N_982,N_2511);
and U8324 (N_8324,N_3933,N_433);
xnor U8325 (N_8325,N_3348,N_2059);
xnor U8326 (N_8326,N_793,N_4650);
and U8327 (N_8327,N_2062,N_1806);
nor U8328 (N_8328,N_4239,N_2005);
nor U8329 (N_8329,N_781,N_3980);
and U8330 (N_8330,N_2914,N_3309);
nor U8331 (N_8331,N_87,N_3511);
or U8332 (N_8332,N_4248,N_2808);
xnor U8333 (N_8333,N_3439,N_2387);
xor U8334 (N_8334,N_3768,N_4710);
and U8335 (N_8335,N_2479,N_3697);
and U8336 (N_8336,N_1761,N_2160);
or U8337 (N_8337,N_4323,N_2520);
xor U8338 (N_8338,N_2222,N_4436);
and U8339 (N_8339,N_2,N_1162);
xnor U8340 (N_8340,N_128,N_3034);
and U8341 (N_8341,N_4677,N_1285);
or U8342 (N_8342,N_2389,N_2259);
or U8343 (N_8343,N_2640,N_4579);
nand U8344 (N_8344,N_3062,N_3946);
xnor U8345 (N_8345,N_672,N_4536);
or U8346 (N_8346,N_1012,N_4157);
nand U8347 (N_8347,N_4437,N_2995);
nor U8348 (N_8348,N_1627,N_564);
and U8349 (N_8349,N_497,N_4828);
nand U8350 (N_8350,N_2476,N_3526);
and U8351 (N_8351,N_4091,N_3672);
or U8352 (N_8352,N_1139,N_2747);
nand U8353 (N_8353,N_1041,N_2028);
or U8354 (N_8354,N_2075,N_1672);
xor U8355 (N_8355,N_2608,N_1330);
nor U8356 (N_8356,N_136,N_3705);
and U8357 (N_8357,N_1256,N_3528);
nand U8358 (N_8358,N_2100,N_134);
nand U8359 (N_8359,N_1341,N_4144);
xnor U8360 (N_8360,N_1420,N_3048);
or U8361 (N_8361,N_4445,N_4640);
and U8362 (N_8362,N_1122,N_4026);
nand U8363 (N_8363,N_4527,N_4459);
or U8364 (N_8364,N_4023,N_187);
nand U8365 (N_8365,N_2793,N_3855);
nand U8366 (N_8366,N_3703,N_4822);
or U8367 (N_8367,N_4377,N_953);
and U8368 (N_8368,N_1848,N_16);
and U8369 (N_8369,N_2994,N_2125);
or U8370 (N_8370,N_130,N_1010);
nor U8371 (N_8371,N_3302,N_1616);
nor U8372 (N_8372,N_2894,N_8);
and U8373 (N_8373,N_2231,N_1594);
xnor U8374 (N_8374,N_367,N_2830);
and U8375 (N_8375,N_4148,N_4835);
and U8376 (N_8376,N_3168,N_2363);
or U8377 (N_8377,N_3923,N_4582);
or U8378 (N_8378,N_379,N_3844);
and U8379 (N_8379,N_3672,N_560);
xnor U8380 (N_8380,N_4695,N_164);
nor U8381 (N_8381,N_4123,N_3686);
nor U8382 (N_8382,N_3602,N_616);
xnor U8383 (N_8383,N_2877,N_3462);
or U8384 (N_8384,N_1719,N_3286);
and U8385 (N_8385,N_3128,N_2277);
or U8386 (N_8386,N_1792,N_3458);
or U8387 (N_8387,N_3791,N_2608);
xor U8388 (N_8388,N_3099,N_2569);
and U8389 (N_8389,N_2264,N_4940);
or U8390 (N_8390,N_4927,N_1559);
and U8391 (N_8391,N_3017,N_3765);
or U8392 (N_8392,N_708,N_4737);
or U8393 (N_8393,N_3076,N_1979);
nor U8394 (N_8394,N_4266,N_2426);
nor U8395 (N_8395,N_189,N_1626);
and U8396 (N_8396,N_1197,N_3613);
nor U8397 (N_8397,N_128,N_2196);
nor U8398 (N_8398,N_3089,N_590);
nor U8399 (N_8399,N_2291,N_4332);
or U8400 (N_8400,N_3336,N_3096);
xor U8401 (N_8401,N_4270,N_2386);
and U8402 (N_8402,N_1525,N_4249);
or U8403 (N_8403,N_4472,N_1219);
nor U8404 (N_8404,N_3823,N_1295);
and U8405 (N_8405,N_1344,N_2207);
and U8406 (N_8406,N_4135,N_3682);
xor U8407 (N_8407,N_1537,N_4872);
xor U8408 (N_8408,N_2060,N_1225);
and U8409 (N_8409,N_1184,N_4644);
or U8410 (N_8410,N_4769,N_3786);
nand U8411 (N_8411,N_2276,N_1741);
nand U8412 (N_8412,N_4086,N_3869);
or U8413 (N_8413,N_2319,N_1127);
nor U8414 (N_8414,N_317,N_202);
nand U8415 (N_8415,N_3302,N_4750);
xnor U8416 (N_8416,N_563,N_4788);
nor U8417 (N_8417,N_691,N_848);
nor U8418 (N_8418,N_2148,N_3337);
xnor U8419 (N_8419,N_1273,N_3952);
nor U8420 (N_8420,N_2675,N_4000);
xor U8421 (N_8421,N_1514,N_3753);
or U8422 (N_8422,N_2901,N_596);
and U8423 (N_8423,N_3784,N_2053);
nand U8424 (N_8424,N_2655,N_2641);
or U8425 (N_8425,N_185,N_429);
or U8426 (N_8426,N_2095,N_149);
nand U8427 (N_8427,N_440,N_1652);
and U8428 (N_8428,N_3016,N_1387);
and U8429 (N_8429,N_4081,N_548);
xnor U8430 (N_8430,N_3117,N_2370);
or U8431 (N_8431,N_69,N_3736);
nor U8432 (N_8432,N_231,N_3589);
nand U8433 (N_8433,N_703,N_3224);
nor U8434 (N_8434,N_2808,N_2172);
nor U8435 (N_8435,N_4972,N_1488);
nand U8436 (N_8436,N_1095,N_2109);
or U8437 (N_8437,N_1251,N_3758);
nor U8438 (N_8438,N_3524,N_852);
xor U8439 (N_8439,N_357,N_4521);
and U8440 (N_8440,N_3034,N_61);
nor U8441 (N_8441,N_3375,N_408);
xnor U8442 (N_8442,N_141,N_2923);
xor U8443 (N_8443,N_319,N_1465);
nand U8444 (N_8444,N_2914,N_1765);
or U8445 (N_8445,N_4610,N_2008);
xnor U8446 (N_8446,N_808,N_3438);
nand U8447 (N_8447,N_4960,N_2786);
nor U8448 (N_8448,N_568,N_4408);
xnor U8449 (N_8449,N_4451,N_4734);
xnor U8450 (N_8450,N_3872,N_1673);
nand U8451 (N_8451,N_2335,N_3427);
nand U8452 (N_8452,N_1730,N_2872);
nand U8453 (N_8453,N_1304,N_600);
or U8454 (N_8454,N_4806,N_2725);
or U8455 (N_8455,N_4806,N_3560);
xnor U8456 (N_8456,N_2639,N_2419);
and U8457 (N_8457,N_2186,N_737);
and U8458 (N_8458,N_1575,N_3903);
xor U8459 (N_8459,N_4159,N_978);
xor U8460 (N_8460,N_2633,N_1601);
nor U8461 (N_8461,N_3945,N_2693);
or U8462 (N_8462,N_3953,N_1538);
nor U8463 (N_8463,N_937,N_4328);
and U8464 (N_8464,N_2684,N_2183);
or U8465 (N_8465,N_492,N_1452);
nor U8466 (N_8466,N_319,N_2969);
and U8467 (N_8467,N_878,N_2129);
nor U8468 (N_8468,N_4482,N_1339);
or U8469 (N_8469,N_716,N_3380);
nand U8470 (N_8470,N_3816,N_3488);
and U8471 (N_8471,N_4891,N_4930);
xor U8472 (N_8472,N_1790,N_1707);
or U8473 (N_8473,N_1246,N_3559);
or U8474 (N_8474,N_1903,N_2085);
nor U8475 (N_8475,N_1285,N_464);
or U8476 (N_8476,N_212,N_3870);
xnor U8477 (N_8477,N_1346,N_2243);
nor U8478 (N_8478,N_3687,N_4295);
nand U8479 (N_8479,N_2893,N_2005);
nor U8480 (N_8480,N_1218,N_4575);
or U8481 (N_8481,N_3233,N_1771);
or U8482 (N_8482,N_130,N_2649);
and U8483 (N_8483,N_2158,N_4559);
nand U8484 (N_8484,N_1434,N_529);
xnor U8485 (N_8485,N_4819,N_3871);
nor U8486 (N_8486,N_1581,N_504);
nand U8487 (N_8487,N_1282,N_672);
xnor U8488 (N_8488,N_2131,N_3357);
and U8489 (N_8489,N_292,N_4567);
or U8490 (N_8490,N_1876,N_1110);
nand U8491 (N_8491,N_3873,N_2808);
and U8492 (N_8492,N_1057,N_1846);
xor U8493 (N_8493,N_2710,N_2611);
or U8494 (N_8494,N_1199,N_3486);
nand U8495 (N_8495,N_4473,N_4116);
xor U8496 (N_8496,N_3268,N_3846);
and U8497 (N_8497,N_4067,N_4243);
or U8498 (N_8498,N_2972,N_2031);
and U8499 (N_8499,N_4999,N_1089);
nand U8500 (N_8500,N_534,N_3821);
and U8501 (N_8501,N_3423,N_2065);
nand U8502 (N_8502,N_4941,N_1002);
nor U8503 (N_8503,N_2143,N_4328);
nand U8504 (N_8504,N_2303,N_1069);
or U8505 (N_8505,N_3481,N_1576);
and U8506 (N_8506,N_864,N_3326);
nand U8507 (N_8507,N_2781,N_292);
xor U8508 (N_8508,N_169,N_2271);
xor U8509 (N_8509,N_2919,N_4381);
or U8510 (N_8510,N_3343,N_1247);
nor U8511 (N_8511,N_4021,N_3431);
nand U8512 (N_8512,N_2452,N_4547);
nand U8513 (N_8513,N_2597,N_392);
and U8514 (N_8514,N_4372,N_2087);
nor U8515 (N_8515,N_4214,N_3701);
nor U8516 (N_8516,N_4854,N_2930);
xor U8517 (N_8517,N_325,N_2169);
nand U8518 (N_8518,N_133,N_1824);
xor U8519 (N_8519,N_1148,N_528);
and U8520 (N_8520,N_2269,N_3993);
nand U8521 (N_8521,N_2793,N_294);
and U8522 (N_8522,N_3685,N_4617);
or U8523 (N_8523,N_1593,N_1620);
xnor U8524 (N_8524,N_3157,N_3409);
xnor U8525 (N_8525,N_234,N_3248);
nand U8526 (N_8526,N_959,N_4598);
nand U8527 (N_8527,N_3089,N_2300);
or U8528 (N_8528,N_4280,N_2974);
nor U8529 (N_8529,N_1615,N_2965);
or U8530 (N_8530,N_1362,N_1265);
nand U8531 (N_8531,N_4971,N_177);
nand U8532 (N_8532,N_4453,N_1461);
nand U8533 (N_8533,N_3774,N_2227);
nand U8534 (N_8534,N_4291,N_1779);
and U8535 (N_8535,N_959,N_1198);
and U8536 (N_8536,N_4006,N_3942);
xnor U8537 (N_8537,N_539,N_3964);
nand U8538 (N_8538,N_1675,N_3660);
and U8539 (N_8539,N_2789,N_1764);
xnor U8540 (N_8540,N_2854,N_331);
nor U8541 (N_8541,N_4471,N_4806);
nand U8542 (N_8542,N_487,N_462);
nor U8543 (N_8543,N_2582,N_320);
and U8544 (N_8544,N_850,N_4856);
and U8545 (N_8545,N_920,N_2904);
or U8546 (N_8546,N_994,N_2722);
or U8547 (N_8547,N_993,N_1134);
nor U8548 (N_8548,N_2861,N_2270);
or U8549 (N_8549,N_2772,N_4014);
or U8550 (N_8550,N_4781,N_1052);
nor U8551 (N_8551,N_3032,N_240);
and U8552 (N_8552,N_2970,N_4951);
and U8553 (N_8553,N_3647,N_1165);
nor U8554 (N_8554,N_3240,N_4540);
or U8555 (N_8555,N_686,N_1041);
and U8556 (N_8556,N_1976,N_744);
nor U8557 (N_8557,N_2370,N_735);
and U8558 (N_8558,N_3997,N_386);
xor U8559 (N_8559,N_1003,N_449);
or U8560 (N_8560,N_3350,N_1027);
and U8561 (N_8561,N_398,N_4503);
and U8562 (N_8562,N_1497,N_145);
xor U8563 (N_8563,N_1913,N_1592);
nor U8564 (N_8564,N_1148,N_3831);
nor U8565 (N_8565,N_4055,N_4042);
nor U8566 (N_8566,N_4092,N_2041);
nand U8567 (N_8567,N_2725,N_4314);
nand U8568 (N_8568,N_1869,N_1677);
and U8569 (N_8569,N_4085,N_3916);
xor U8570 (N_8570,N_2653,N_2429);
nor U8571 (N_8571,N_551,N_2119);
xor U8572 (N_8572,N_2357,N_3192);
or U8573 (N_8573,N_4771,N_708);
nand U8574 (N_8574,N_3274,N_2527);
nor U8575 (N_8575,N_4690,N_3137);
nor U8576 (N_8576,N_1536,N_1521);
and U8577 (N_8577,N_1976,N_3884);
nor U8578 (N_8578,N_1529,N_4909);
or U8579 (N_8579,N_4937,N_4369);
nor U8580 (N_8580,N_623,N_4035);
nor U8581 (N_8581,N_3390,N_507);
nor U8582 (N_8582,N_3092,N_445);
xnor U8583 (N_8583,N_538,N_1252);
and U8584 (N_8584,N_2093,N_100);
nand U8585 (N_8585,N_237,N_3057);
or U8586 (N_8586,N_2176,N_2341);
nand U8587 (N_8587,N_1533,N_899);
or U8588 (N_8588,N_1953,N_1457);
nor U8589 (N_8589,N_4346,N_4682);
nor U8590 (N_8590,N_3686,N_4415);
or U8591 (N_8591,N_3763,N_2005);
or U8592 (N_8592,N_2402,N_689);
nor U8593 (N_8593,N_2710,N_1889);
xor U8594 (N_8594,N_1288,N_1615);
nand U8595 (N_8595,N_611,N_4472);
nand U8596 (N_8596,N_509,N_1857);
nand U8597 (N_8597,N_2359,N_3425);
nand U8598 (N_8598,N_1251,N_3678);
xnor U8599 (N_8599,N_4287,N_2855);
nand U8600 (N_8600,N_3561,N_3280);
xor U8601 (N_8601,N_4446,N_3315);
xor U8602 (N_8602,N_2383,N_372);
nand U8603 (N_8603,N_4203,N_3621);
or U8604 (N_8604,N_3264,N_4405);
nor U8605 (N_8605,N_2028,N_2221);
nand U8606 (N_8606,N_1909,N_4753);
xor U8607 (N_8607,N_3255,N_1486);
nand U8608 (N_8608,N_1807,N_2102);
and U8609 (N_8609,N_1064,N_4008);
xor U8610 (N_8610,N_2277,N_3909);
and U8611 (N_8611,N_2971,N_408);
xor U8612 (N_8612,N_2344,N_146);
nor U8613 (N_8613,N_4637,N_3198);
nor U8614 (N_8614,N_3802,N_423);
or U8615 (N_8615,N_479,N_11);
and U8616 (N_8616,N_1197,N_3896);
xnor U8617 (N_8617,N_1915,N_2921);
nor U8618 (N_8618,N_4839,N_1564);
nand U8619 (N_8619,N_2525,N_414);
nor U8620 (N_8620,N_4835,N_951);
and U8621 (N_8621,N_488,N_727);
nand U8622 (N_8622,N_1826,N_2472);
or U8623 (N_8623,N_4944,N_3114);
and U8624 (N_8624,N_981,N_4548);
nand U8625 (N_8625,N_4125,N_4445);
and U8626 (N_8626,N_4827,N_4694);
nand U8627 (N_8627,N_2900,N_1368);
or U8628 (N_8628,N_3968,N_3924);
nor U8629 (N_8629,N_3551,N_2664);
or U8630 (N_8630,N_307,N_47);
nor U8631 (N_8631,N_2934,N_2851);
or U8632 (N_8632,N_2652,N_914);
and U8633 (N_8633,N_1558,N_1855);
or U8634 (N_8634,N_2154,N_2911);
nor U8635 (N_8635,N_2332,N_3210);
xor U8636 (N_8636,N_4437,N_967);
or U8637 (N_8637,N_1139,N_583);
nand U8638 (N_8638,N_583,N_3570);
xor U8639 (N_8639,N_4,N_2970);
nor U8640 (N_8640,N_505,N_2334);
xnor U8641 (N_8641,N_1847,N_4680);
nor U8642 (N_8642,N_4931,N_4588);
nand U8643 (N_8643,N_2520,N_4215);
or U8644 (N_8644,N_3098,N_2222);
and U8645 (N_8645,N_1577,N_418);
nor U8646 (N_8646,N_1492,N_1656);
xor U8647 (N_8647,N_1519,N_3722);
xnor U8648 (N_8648,N_2231,N_88);
nor U8649 (N_8649,N_4710,N_1270);
or U8650 (N_8650,N_2165,N_1255);
nand U8651 (N_8651,N_3570,N_364);
nor U8652 (N_8652,N_4223,N_1337);
xor U8653 (N_8653,N_4972,N_3885);
or U8654 (N_8654,N_3045,N_2047);
or U8655 (N_8655,N_2908,N_7);
or U8656 (N_8656,N_3460,N_78);
and U8657 (N_8657,N_4317,N_1587);
and U8658 (N_8658,N_1671,N_1365);
or U8659 (N_8659,N_613,N_3819);
and U8660 (N_8660,N_773,N_904);
or U8661 (N_8661,N_2757,N_3546);
or U8662 (N_8662,N_2617,N_3416);
nor U8663 (N_8663,N_3403,N_1369);
nor U8664 (N_8664,N_2932,N_4111);
or U8665 (N_8665,N_3443,N_1426);
or U8666 (N_8666,N_3342,N_268);
and U8667 (N_8667,N_1225,N_3032);
xnor U8668 (N_8668,N_4646,N_972);
nand U8669 (N_8669,N_4346,N_1437);
nand U8670 (N_8670,N_4922,N_1579);
xor U8671 (N_8671,N_1732,N_904);
xor U8672 (N_8672,N_4493,N_2927);
nor U8673 (N_8673,N_2538,N_980);
nor U8674 (N_8674,N_4018,N_3938);
nor U8675 (N_8675,N_2714,N_1684);
and U8676 (N_8676,N_130,N_3724);
and U8677 (N_8677,N_1796,N_1802);
or U8678 (N_8678,N_4964,N_1862);
nand U8679 (N_8679,N_965,N_3053);
xnor U8680 (N_8680,N_4527,N_1913);
and U8681 (N_8681,N_112,N_1724);
or U8682 (N_8682,N_2330,N_918);
or U8683 (N_8683,N_4186,N_3252);
nand U8684 (N_8684,N_4538,N_4180);
or U8685 (N_8685,N_4915,N_1345);
nand U8686 (N_8686,N_2773,N_4025);
and U8687 (N_8687,N_4245,N_3062);
nand U8688 (N_8688,N_2199,N_4622);
or U8689 (N_8689,N_3440,N_3558);
and U8690 (N_8690,N_136,N_2392);
nand U8691 (N_8691,N_2123,N_1697);
and U8692 (N_8692,N_3618,N_4139);
or U8693 (N_8693,N_3552,N_950);
and U8694 (N_8694,N_4148,N_4837);
xor U8695 (N_8695,N_219,N_1752);
and U8696 (N_8696,N_30,N_1456);
nand U8697 (N_8697,N_637,N_4846);
or U8698 (N_8698,N_4149,N_4241);
xor U8699 (N_8699,N_4695,N_4288);
nand U8700 (N_8700,N_4153,N_3135);
and U8701 (N_8701,N_3762,N_3854);
or U8702 (N_8702,N_1914,N_1128);
nand U8703 (N_8703,N_395,N_3386);
nor U8704 (N_8704,N_3378,N_458);
nor U8705 (N_8705,N_3527,N_3702);
xnor U8706 (N_8706,N_1302,N_3030);
nand U8707 (N_8707,N_3146,N_4122);
xnor U8708 (N_8708,N_3825,N_1242);
nand U8709 (N_8709,N_529,N_4652);
and U8710 (N_8710,N_3732,N_3600);
xnor U8711 (N_8711,N_3561,N_718);
nand U8712 (N_8712,N_4114,N_2420);
and U8713 (N_8713,N_3382,N_1379);
nor U8714 (N_8714,N_4644,N_2328);
and U8715 (N_8715,N_73,N_4482);
and U8716 (N_8716,N_2999,N_2061);
xor U8717 (N_8717,N_4283,N_3047);
and U8718 (N_8718,N_580,N_1233);
nand U8719 (N_8719,N_40,N_3149);
or U8720 (N_8720,N_2321,N_470);
nand U8721 (N_8721,N_2268,N_3434);
and U8722 (N_8722,N_2476,N_296);
xnor U8723 (N_8723,N_3600,N_2951);
nor U8724 (N_8724,N_2481,N_4524);
xor U8725 (N_8725,N_4282,N_12);
nor U8726 (N_8726,N_2407,N_3644);
or U8727 (N_8727,N_1182,N_4338);
nor U8728 (N_8728,N_1496,N_1287);
or U8729 (N_8729,N_4957,N_1642);
nor U8730 (N_8730,N_2665,N_667);
xnor U8731 (N_8731,N_3950,N_3560);
nor U8732 (N_8732,N_3103,N_347);
xor U8733 (N_8733,N_4676,N_2850);
or U8734 (N_8734,N_1509,N_3924);
and U8735 (N_8735,N_2930,N_2793);
or U8736 (N_8736,N_703,N_2036);
nand U8737 (N_8737,N_3374,N_1056);
or U8738 (N_8738,N_36,N_4410);
xnor U8739 (N_8739,N_55,N_4261);
nor U8740 (N_8740,N_1988,N_969);
and U8741 (N_8741,N_3502,N_3904);
nor U8742 (N_8742,N_100,N_3498);
nand U8743 (N_8743,N_2500,N_2086);
nor U8744 (N_8744,N_1267,N_3964);
and U8745 (N_8745,N_1837,N_871);
nand U8746 (N_8746,N_2955,N_81);
or U8747 (N_8747,N_3565,N_1030);
and U8748 (N_8748,N_4029,N_181);
and U8749 (N_8749,N_4869,N_2624);
nand U8750 (N_8750,N_716,N_2918);
nand U8751 (N_8751,N_257,N_1817);
nor U8752 (N_8752,N_484,N_4298);
or U8753 (N_8753,N_2822,N_4779);
xnor U8754 (N_8754,N_2832,N_59);
nand U8755 (N_8755,N_2772,N_872);
nand U8756 (N_8756,N_2786,N_3544);
nand U8757 (N_8757,N_4952,N_1395);
nor U8758 (N_8758,N_3745,N_4727);
or U8759 (N_8759,N_1011,N_697);
xnor U8760 (N_8760,N_2617,N_3557);
and U8761 (N_8761,N_2233,N_1635);
nor U8762 (N_8762,N_4841,N_793);
xnor U8763 (N_8763,N_3940,N_3881);
and U8764 (N_8764,N_4630,N_4007);
nand U8765 (N_8765,N_2116,N_2101);
nand U8766 (N_8766,N_3713,N_700);
nor U8767 (N_8767,N_4918,N_3821);
nand U8768 (N_8768,N_4224,N_4922);
nor U8769 (N_8769,N_4693,N_4567);
nor U8770 (N_8770,N_1944,N_3416);
nor U8771 (N_8771,N_2850,N_2965);
and U8772 (N_8772,N_1781,N_1584);
xor U8773 (N_8773,N_2413,N_2841);
xor U8774 (N_8774,N_2493,N_1357);
or U8775 (N_8775,N_4675,N_3367);
and U8776 (N_8776,N_1586,N_4893);
nand U8777 (N_8777,N_4621,N_2556);
or U8778 (N_8778,N_2554,N_2972);
xnor U8779 (N_8779,N_4082,N_350);
nand U8780 (N_8780,N_1113,N_3797);
and U8781 (N_8781,N_3552,N_4341);
and U8782 (N_8782,N_4801,N_4756);
and U8783 (N_8783,N_4614,N_3388);
and U8784 (N_8784,N_3113,N_314);
nand U8785 (N_8785,N_270,N_3248);
nand U8786 (N_8786,N_29,N_3096);
or U8787 (N_8787,N_3798,N_892);
and U8788 (N_8788,N_3514,N_1483);
and U8789 (N_8789,N_3355,N_2004);
nand U8790 (N_8790,N_4420,N_1906);
xor U8791 (N_8791,N_3823,N_1436);
nand U8792 (N_8792,N_2749,N_1140);
and U8793 (N_8793,N_1734,N_1700);
or U8794 (N_8794,N_1233,N_3359);
and U8795 (N_8795,N_2516,N_3309);
and U8796 (N_8796,N_172,N_2709);
xnor U8797 (N_8797,N_654,N_3520);
and U8798 (N_8798,N_2908,N_2308);
nand U8799 (N_8799,N_222,N_4660);
or U8800 (N_8800,N_596,N_2771);
nor U8801 (N_8801,N_858,N_2480);
nand U8802 (N_8802,N_2031,N_3525);
and U8803 (N_8803,N_1633,N_4859);
or U8804 (N_8804,N_4204,N_4887);
or U8805 (N_8805,N_2773,N_2692);
and U8806 (N_8806,N_2120,N_307);
nand U8807 (N_8807,N_2450,N_427);
and U8808 (N_8808,N_112,N_315);
nand U8809 (N_8809,N_2716,N_4109);
xnor U8810 (N_8810,N_4798,N_156);
xnor U8811 (N_8811,N_3205,N_4723);
xnor U8812 (N_8812,N_3386,N_3706);
nor U8813 (N_8813,N_3274,N_3637);
or U8814 (N_8814,N_1751,N_2141);
or U8815 (N_8815,N_4948,N_2840);
xnor U8816 (N_8816,N_3356,N_4718);
or U8817 (N_8817,N_2514,N_153);
nand U8818 (N_8818,N_3445,N_1636);
nor U8819 (N_8819,N_1489,N_1738);
nor U8820 (N_8820,N_3918,N_825);
nand U8821 (N_8821,N_4217,N_591);
nand U8822 (N_8822,N_1878,N_2100);
and U8823 (N_8823,N_2883,N_4634);
nand U8824 (N_8824,N_4528,N_3131);
nand U8825 (N_8825,N_1875,N_2537);
nor U8826 (N_8826,N_2118,N_1735);
and U8827 (N_8827,N_4894,N_846);
nor U8828 (N_8828,N_4267,N_3216);
xor U8829 (N_8829,N_1100,N_1115);
nor U8830 (N_8830,N_1027,N_48);
nand U8831 (N_8831,N_171,N_4953);
and U8832 (N_8832,N_2398,N_4313);
and U8833 (N_8833,N_3185,N_566);
or U8834 (N_8834,N_4004,N_2070);
nor U8835 (N_8835,N_2905,N_4082);
xor U8836 (N_8836,N_606,N_4911);
xor U8837 (N_8837,N_3687,N_1197);
and U8838 (N_8838,N_2550,N_4376);
nor U8839 (N_8839,N_845,N_3303);
nand U8840 (N_8840,N_4283,N_3115);
and U8841 (N_8841,N_3283,N_581);
nand U8842 (N_8842,N_4686,N_687);
nor U8843 (N_8843,N_3165,N_1561);
xnor U8844 (N_8844,N_4171,N_1595);
and U8845 (N_8845,N_4366,N_2407);
and U8846 (N_8846,N_1503,N_3710);
xnor U8847 (N_8847,N_393,N_3603);
nor U8848 (N_8848,N_2148,N_2510);
xnor U8849 (N_8849,N_1358,N_1259);
xnor U8850 (N_8850,N_3710,N_3542);
or U8851 (N_8851,N_2504,N_2419);
or U8852 (N_8852,N_3655,N_3305);
nand U8853 (N_8853,N_4600,N_3187);
and U8854 (N_8854,N_3109,N_3759);
nand U8855 (N_8855,N_3673,N_141);
nand U8856 (N_8856,N_4999,N_1756);
nand U8857 (N_8857,N_4795,N_1298);
and U8858 (N_8858,N_1281,N_4913);
nand U8859 (N_8859,N_3900,N_1910);
and U8860 (N_8860,N_3361,N_4525);
xnor U8861 (N_8861,N_4997,N_3560);
xor U8862 (N_8862,N_4299,N_4254);
xnor U8863 (N_8863,N_1171,N_99);
nor U8864 (N_8864,N_2573,N_1954);
nand U8865 (N_8865,N_4248,N_3951);
xor U8866 (N_8866,N_4923,N_2486);
xnor U8867 (N_8867,N_1086,N_521);
or U8868 (N_8868,N_1392,N_2050);
or U8869 (N_8869,N_2589,N_373);
nand U8870 (N_8870,N_2139,N_2567);
or U8871 (N_8871,N_4699,N_2724);
nand U8872 (N_8872,N_4540,N_1180);
nand U8873 (N_8873,N_3678,N_356);
nand U8874 (N_8874,N_3941,N_1742);
or U8875 (N_8875,N_4777,N_2958);
nor U8876 (N_8876,N_2642,N_2860);
and U8877 (N_8877,N_1846,N_4371);
or U8878 (N_8878,N_1224,N_3415);
and U8879 (N_8879,N_2990,N_2233);
and U8880 (N_8880,N_2916,N_2694);
nor U8881 (N_8881,N_1656,N_510);
or U8882 (N_8882,N_4937,N_3873);
xor U8883 (N_8883,N_4708,N_3161);
nor U8884 (N_8884,N_1063,N_2399);
nor U8885 (N_8885,N_2990,N_2373);
or U8886 (N_8886,N_3327,N_4704);
nor U8887 (N_8887,N_3014,N_2778);
or U8888 (N_8888,N_4832,N_1834);
and U8889 (N_8889,N_2735,N_4846);
or U8890 (N_8890,N_3791,N_3217);
or U8891 (N_8891,N_59,N_3908);
or U8892 (N_8892,N_1850,N_38);
nor U8893 (N_8893,N_4918,N_488);
xnor U8894 (N_8894,N_2176,N_2535);
xor U8895 (N_8895,N_1256,N_2207);
and U8896 (N_8896,N_1267,N_1153);
nand U8897 (N_8897,N_2819,N_2542);
or U8898 (N_8898,N_831,N_4633);
nor U8899 (N_8899,N_3988,N_4070);
nand U8900 (N_8900,N_3761,N_2023);
and U8901 (N_8901,N_3866,N_3080);
or U8902 (N_8902,N_2753,N_3685);
nor U8903 (N_8903,N_1495,N_725);
nor U8904 (N_8904,N_2374,N_2775);
and U8905 (N_8905,N_940,N_4421);
or U8906 (N_8906,N_4987,N_1156);
or U8907 (N_8907,N_1895,N_3376);
nand U8908 (N_8908,N_4668,N_2460);
and U8909 (N_8909,N_2317,N_2501);
nand U8910 (N_8910,N_2720,N_3196);
xor U8911 (N_8911,N_4025,N_2730);
nor U8912 (N_8912,N_1060,N_513);
nand U8913 (N_8913,N_19,N_3014);
nor U8914 (N_8914,N_1765,N_4807);
and U8915 (N_8915,N_3366,N_4273);
or U8916 (N_8916,N_4314,N_3629);
nand U8917 (N_8917,N_1707,N_4643);
or U8918 (N_8918,N_1034,N_1743);
nand U8919 (N_8919,N_892,N_3635);
and U8920 (N_8920,N_1893,N_2892);
or U8921 (N_8921,N_2090,N_2652);
nor U8922 (N_8922,N_2254,N_716);
xor U8923 (N_8923,N_890,N_1538);
xor U8924 (N_8924,N_1800,N_3645);
or U8925 (N_8925,N_2210,N_2354);
and U8926 (N_8926,N_1273,N_1476);
nand U8927 (N_8927,N_1750,N_1961);
or U8928 (N_8928,N_2439,N_2064);
xnor U8929 (N_8929,N_2292,N_3278);
and U8930 (N_8930,N_4678,N_3836);
or U8931 (N_8931,N_981,N_1376);
and U8932 (N_8932,N_1298,N_1393);
nor U8933 (N_8933,N_4931,N_1239);
or U8934 (N_8934,N_969,N_2934);
and U8935 (N_8935,N_2390,N_1920);
or U8936 (N_8936,N_988,N_2824);
and U8937 (N_8937,N_240,N_2212);
and U8938 (N_8938,N_2238,N_939);
and U8939 (N_8939,N_3801,N_1077);
and U8940 (N_8940,N_3845,N_3921);
nand U8941 (N_8941,N_4492,N_3671);
or U8942 (N_8942,N_3915,N_2177);
or U8943 (N_8943,N_4368,N_4835);
nor U8944 (N_8944,N_4002,N_840);
nand U8945 (N_8945,N_1167,N_4712);
and U8946 (N_8946,N_2581,N_1449);
and U8947 (N_8947,N_4907,N_4225);
or U8948 (N_8948,N_4632,N_3847);
or U8949 (N_8949,N_3734,N_1185);
nor U8950 (N_8950,N_668,N_1473);
or U8951 (N_8951,N_2837,N_3957);
nand U8952 (N_8952,N_662,N_1744);
or U8953 (N_8953,N_2804,N_1676);
nand U8954 (N_8954,N_2096,N_3930);
nor U8955 (N_8955,N_4348,N_767);
nor U8956 (N_8956,N_4671,N_3561);
xor U8957 (N_8957,N_4882,N_4123);
nand U8958 (N_8958,N_3101,N_4117);
nand U8959 (N_8959,N_3894,N_2867);
and U8960 (N_8960,N_614,N_3299);
xor U8961 (N_8961,N_321,N_2559);
or U8962 (N_8962,N_2467,N_1339);
and U8963 (N_8963,N_3455,N_2421);
nor U8964 (N_8964,N_2760,N_2379);
and U8965 (N_8965,N_414,N_3084);
or U8966 (N_8966,N_3023,N_2139);
or U8967 (N_8967,N_908,N_2732);
nand U8968 (N_8968,N_1451,N_4527);
or U8969 (N_8969,N_4226,N_4549);
nor U8970 (N_8970,N_1976,N_396);
and U8971 (N_8971,N_230,N_71);
xnor U8972 (N_8972,N_4398,N_1485);
nor U8973 (N_8973,N_462,N_3616);
xnor U8974 (N_8974,N_1127,N_1509);
nand U8975 (N_8975,N_3603,N_2189);
nand U8976 (N_8976,N_493,N_705);
nor U8977 (N_8977,N_2658,N_3166);
and U8978 (N_8978,N_3769,N_1023);
or U8979 (N_8979,N_2490,N_178);
nand U8980 (N_8980,N_4730,N_2263);
or U8981 (N_8981,N_4328,N_2872);
nor U8982 (N_8982,N_836,N_319);
and U8983 (N_8983,N_4731,N_91);
and U8984 (N_8984,N_279,N_3763);
nor U8985 (N_8985,N_1848,N_3891);
xor U8986 (N_8986,N_376,N_2763);
nor U8987 (N_8987,N_200,N_723);
nor U8988 (N_8988,N_3469,N_72);
xor U8989 (N_8989,N_603,N_1604);
or U8990 (N_8990,N_331,N_4979);
nor U8991 (N_8991,N_4660,N_1664);
nor U8992 (N_8992,N_4538,N_3154);
nand U8993 (N_8993,N_346,N_1174);
nor U8994 (N_8994,N_3281,N_177);
xnor U8995 (N_8995,N_3741,N_2823);
or U8996 (N_8996,N_3987,N_2524);
or U8997 (N_8997,N_1701,N_1892);
nor U8998 (N_8998,N_4361,N_4364);
nand U8999 (N_8999,N_1974,N_2962);
nor U9000 (N_9000,N_416,N_2402);
and U9001 (N_9001,N_2896,N_3220);
nor U9002 (N_9002,N_3207,N_1932);
nand U9003 (N_9003,N_1789,N_4647);
nor U9004 (N_9004,N_2567,N_3128);
xor U9005 (N_9005,N_2289,N_1504);
nor U9006 (N_9006,N_4401,N_3058);
and U9007 (N_9007,N_1540,N_1994);
and U9008 (N_9008,N_3479,N_3749);
nand U9009 (N_9009,N_554,N_4690);
and U9010 (N_9010,N_3465,N_2172);
and U9011 (N_9011,N_1796,N_1387);
nor U9012 (N_9012,N_1696,N_1852);
nand U9013 (N_9013,N_4812,N_4345);
and U9014 (N_9014,N_240,N_2998);
nor U9015 (N_9015,N_2247,N_2752);
nor U9016 (N_9016,N_551,N_1308);
nand U9017 (N_9017,N_424,N_471);
nor U9018 (N_9018,N_4672,N_1580);
and U9019 (N_9019,N_3788,N_1634);
or U9020 (N_9020,N_830,N_3739);
and U9021 (N_9021,N_1329,N_2160);
or U9022 (N_9022,N_2943,N_2237);
nand U9023 (N_9023,N_726,N_89);
and U9024 (N_9024,N_1128,N_1298);
nand U9025 (N_9025,N_4421,N_104);
or U9026 (N_9026,N_1888,N_375);
or U9027 (N_9027,N_3159,N_1528);
nand U9028 (N_9028,N_2060,N_4799);
and U9029 (N_9029,N_1808,N_1921);
xor U9030 (N_9030,N_821,N_1651);
nand U9031 (N_9031,N_4342,N_4107);
or U9032 (N_9032,N_1777,N_3642);
xnor U9033 (N_9033,N_324,N_2304);
or U9034 (N_9034,N_2720,N_2583);
xor U9035 (N_9035,N_3248,N_307);
or U9036 (N_9036,N_904,N_1463);
and U9037 (N_9037,N_4055,N_2825);
or U9038 (N_9038,N_3977,N_2720);
xor U9039 (N_9039,N_626,N_775);
xor U9040 (N_9040,N_2903,N_2467);
nor U9041 (N_9041,N_2828,N_1230);
or U9042 (N_9042,N_4314,N_4910);
and U9043 (N_9043,N_2534,N_3834);
nor U9044 (N_9044,N_4941,N_873);
xor U9045 (N_9045,N_65,N_4292);
xnor U9046 (N_9046,N_1413,N_1900);
nand U9047 (N_9047,N_2368,N_4499);
or U9048 (N_9048,N_4002,N_1282);
nand U9049 (N_9049,N_2842,N_3953);
xnor U9050 (N_9050,N_4003,N_3545);
nor U9051 (N_9051,N_787,N_3647);
xnor U9052 (N_9052,N_1903,N_2198);
or U9053 (N_9053,N_947,N_3496);
xnor U9054 (N_9054,N_3605,N_3479);
xor U9055 (N_9055,N_4423,N_1137);
or U9056 (N_9056,N_730,N_2698);
and U9057 (N_9057,N_4451,N_740);
nor U9058 (N_9058,N_80,N_3223);
or U9059 (N_9059,N_2738,N_1058);
xor U9060 (N_9060,N_83,N_2118);
nand U9061 (N_9061,N_4347,N_4593);
or U9062 (N_9062,N_3495,N_2234);
nor U9063 (N_9063,N_4683,N_2880);
and U9064 (N_9064,N_2722,N_98);
nand U9065 (N_9065,N_3171,N_4404);
or U9066 (N_9066,N_4461,N_687);
nand U9067 (N_9067,N_3104,N_4686);
nand U9068 (N_9068,N_458,N_2568);
nor U9069 (N_9069,N_315,N_4511);
nor U9070 (N_9070,N_4510,N_4291);
or U9071 (N_9071,N_2062,N_4660);
nor U9072 (N_9072,N_873,N_1876);
xnor U9073 (N_9073,N_1816,N_1787);
xor U9074 (N_9074,N_1282,N_3333);
or U9075 (N_9075,N_1430,N_3849);
nand U9076 (N_9076,N_977,N_3989);
xor U9077 (N_9077,N_3129,N_3813);
nand U9078 (N_9078,N_1419,N_4768);
nand U9079 (N_9079,N_1293,N_2911);
or U9080 (N_9080,N_4576,N_3140);
or U9081 (N_9081,N_2042,N_3336);
nor U9082 (N_9082,N_2974,N_1535);
nand U9083 (N_9083,N_2956,N_375);
nand U9084 (N_9084,N_2430,N_1154);
nor U9085 (N_9085,N_1144,N_4617);
nand U9086 (N_9086,N_1868,N_255);
nand U9087 (N_9087,N_1040,N_809);
nor U9088 (N_9088,N_4662,N_4833);
nand U9089 (N_9089,N_3352,N_2049);
or U9090 (N_9090,N_3231,N_603);
nor U9091 (N_9091,N_560,N_4042);
or U9092 (N_9092,N_700,N_2392);
xnor U9093 (N_9093,N_4003,N_4240);
xnor U9094 (N_9094,N_446,N_2844);
and U9095 (N_9095,N_888,N_224);
and U9096 (N_9096,N_746,N_4790);
xnor U9097 (N_9097,N_4568,N_206);
nor U9098 (N_9098,N_1191,N_355);
and U9099 (N_9099,N_1606,N_2590);
and U9100 (N_9100,N_1815,N_4797);
nor U9101 (N_9101,N_3660,N_2928);
and U9102 (N_9102,N_1803,N_1564);
nand U9103 (N_9103,N_3378,N_2194);
xor U9104 (N_9104,N_697,N_4892);
nand U9105 (N_9105,N_1421,N_4996);
nand U9106 (N_9106,N_1179,N_960);
nor U9107 (N_9107,N_1106,N_4239);
nor U9108 (N_9108,N_2762,N_4084);
nand U9109 (N_9109,N_3777,N_2742);
nand U9110 (N_9110,N_1113,N_4963);
xnor U9111 (N_9111,N_2931,N_1723);
or U9112 (N_9112,N_2881,N_4471);
xor U9113 (N_9113,N_2483,N_82);
xnor U9114 (N_9114,N_4015,N_1217);
and U9115 (N_9115,N_4203,N_4);
nand U9116 (N_9116,N_625,N_1312);
or U9117 (N_9117,N_1341,N_2271);
xnor U9118 (N_9118,N_3682,N_3932);
or U9119 (N_9119,N_3756,N_4538);
nand U9120 (N_9120,N_4688,N_1038);
or U9121 (N_9121,N_1036,N_2587);
xor U9122 (N_9122,N_4432,N_4783);
xnor U9123 (N_9123,N_532,N_1272);
nand U9124 (N_9124,N_138,N_1689);
nand U9125 (N_9125,N_3551,N_35);
xor U9126 (N_9126,N_2311,N_1748);
xor U9127 (N_9127,N_2084,N_995);
and U9128 (N_9128,N_674,N_3065);
and U9129 (N_9129,N_4441,N_2700);
xor U9130 (N_9130,N_439,N_422);
xor U9131 (N_9131,N_1690,N_3518);
or U9132 (N_9132,N_4619,N_4525);
nand U9133 (N_9133,N_2632,N_594);
nor U9134 (N_9134,N_1683,N_318);
nor U9135 (N_9135,N_4484,N_1217);
nand U9136 (N_9136,N_1528,N_4408);
nor U9137 (N_9137,N_2307,N_3760);
nand U9138 (N_9138,N_1903,N_1459);
nand U9139 (N_9139,N_656,N_2635);
and U9140 (N_9140,N_2898,N_1897);
nor U9141 (N_9141,N_531,N_2792);
or U9142 (N_9142,N_1811,N_2658);
xnor U9143 (N_9143,N_783,N_609);
nand U9144 (N_9144,N_2974,N_4498);
xnor U9145 (N_9145,N_3087,N_685);
nor U9146 (N_9146,N_3542,N_898);
or U9147 (N_9147,N_3705,N_4370);
nand U9148 (N_9148,N_2460,N_1933);
and U9149 (N_9149,N_4666,N_4703);
and U9150 (N_9150,N_3025,N_4847);
or U9151 (N_9151,N_2783,N_2970);
or U9152 (N_9152,N_1041,N_2908);
and U9153 (N_9153,N_2182,N_2446);
xnor U9154 (N_9154,N_1155,N_3326);
nand U9155 (N_9155,N_2173,N_2302);
nand U9156 (N_9156,N_882,N_2135);
or U9157 (N_9157,N_2641,N_1403);
or U9158 (N_9158,N_2413,N_3853);
nor U9159 (N_9159,N_1321,N_1687);
xnor U9160 (N_9160,N_2353,N_2106);
nor U9161 (N_9161,N_1959,N_4266);
xnor U9162 (N_9162,N_3919,N_3872);
and U9163 (N_9163,N_3700,N_599);
and U9164 (N_9164,N_4357,N_4607);
and U9165 (N_9165,N_2157,N_3957);
nand U9166 (N_9166,N_4201,N_2340);
and U9167 (N_9167,N_4456,N_2950);
or U9168 (N_9168,N_2654,N_6);
nand U9169 (N_9169,N_2760,N_2918);
or U9170 (N_9170,N_2980,N_386);
nor U9171 (N_9171,N_3046,N_3087);
xor U9172 (N_9172,N_3227,N_4188);
nor U9173 (N_9173,N_2076,N_4802);
nor U9174 (N_9174,N_519,N_4491);
and U9175 (N_9175,N_2263,N_4793);
nand U9176 (N_9176,N_4721,N_1528);
nor U9177 (N_9177,N_1761,N_2463);
nand U9178 (N_9178,N_2984,N_3253);
and U9179 (N_9179,N_1820,N_32);
and U9180 (N_9180,N_2821,N_2302);
or U9181 (N_9181,N_1539,N_4911);
or U9182 (N_9182,N_2532,N_4769);
or U9183 (N_9183,N_3542,N_2767);
nand U9184 (N_9184,N_578,N_1628);
and U9185 (N_9185,N_4624,N_1670);
and U9186 (N_9186,N_4270,N_2000);
nand U9187 (N_9187,N_1438,N_2379);
and U9188 (N_9188,N_2031,N_435);
nor U9189 (N_9189,N_3472,N_253);
nor U9190 (N_9190,N_4432,N_2633);
or U9191 (N_9191,N_1924,N_4986);
or U9192 (N_9192,N_556,N_2134);
and U9193 (N_9193,N_2194,N_1763);
nor U9194 (N_9194,N_3247,N_525);
xnor U9195 (N_9195,N_1989,N_907);
xor U9196 (N_9196,N_578,N_4051);
xor U9197 (N_9197,N_3796,N_3281);
or U9198 (N_9198,N_283,N_1207);
nor U9199 (N_9199,N_1746,N_2150);
and U9200 (N_9200,N_2938,N_3792);
and U9201 (N_9201,N_1192,N_420);
or U9202 (N_9202,N_3533,N_4900);
nor U9203 (N_9203,N_3900,N_2203);
xnor U9204 (N_9204,N_4368,N_3961);
nor U9205 (N_9205,N_1638,N_3664);
or U9206 (N_9206,N_3714,N_1890);
or U9207 (N_9207,N_2302,N_3488);
and U9208 (N_9208,N_3151,N_1538);
and U9209 (N_9209,N_2535,N_2399);
xnor U9210 (N_9210,N_1652,N_2965);
or U9211 (N_9211,N_2558,N_4498);
and U9212 (N_9212,N_371,N_1322);
and U9213 (N_9213,N_4161,N_3585);
or U9214 (N_9214,N_3743,N_1596);
nor U9215 (N_9215,N_4784,N_4052);
nand U9216 (N_9216,N_118,N_2793);
or U9217 (N_9217,N_914,N_1727);
nand U9218 (N_9218,N_1315,N_3795);
and U9219 (N_9219,N_4782,N_2591);
xnor U9220 (N_9220,N_2544,N_3557);
and U9221 (N_9221,N_3296,N_4054);
and U9222 (N_9222,N_2651,N_2033);
or U9223 (N_9223,N_1947,N_2774);
or U9224 (N_9224,N_2376,N_1278);
nor U9225 (N_9225,N_602,N_2060);
nand U9226 (N_9226,N_498,N_4451);
nand U9227 (N_9227,N_4713,N_1003);
xnor U9228 (N_9228,N_2657,N_3084);
and U9229 (N_9229,N_3334,N_3569);
nand U9230 (N_9230,N_1116,N_2412);
xnor U9231 (N_9231,N_4680,N_3782);
nor U9232 (N_9232,N_2735,N_3537);
nand U9233 (N_9233,N_4327,N_1174);
nor U9234 (N_9234,N_3616,N_4013);
or U9235 (N_9235,N_572,N_1707);
nand U9236 (N_9236,N_1051,N_2329);
or U9237 (N_9237,N_4030,N_2023);
and U9238 (N_9238,N_4472,N_429);
and U9239 (N_9239,N_1512,N_2714);
nor U9240 (N_9240,N_2261,N_2437);
or U9241 (N_9241,N_2377,N_3071);
nor U9242 (N_9242,N_1620,N_4370);
and U9243 (N_9243,N_2227,N_458);
nor U9244 (N_9244,N_1414,N_154);
or U9245 (N_9245,N_4685,N_3332);
nor U9246 (N_9246,N_530,N_1504);
nand U9247 (N_9247,N_4738,N_2520);
nor U9248 (N_9248,N_4177,N_2643);
nor U9249 (N_9249,N_3273,N_4156);
nand U9250 (N_9250,N_95,N_4508);
xor U9251 (N_9251,N_3040,N_668);
xor U9252 (N_9252,N_3102,N_4277);
nor U9253 (N_9253,N_3656,N_2069);
xnor U9254 (N_9254,N_1676,N_2460);
nand U9255 (N_9255,N_4658,N_2121);
nand U9256 (N_9256,N_4830,N_340);
nor U9257 (N_9257,N_313,N_4757);
and U9258 (N_9258,N_186,N_2661);
xor U9259 (N_9259,N_4851,N_3136);
and U9260 (N_9260,N_1677,N_1114);
and U9261 (N_9261,N_1532,N_3809);
nand U9262 (N_9262,N_418,N_1727);
nor U9263 (N_9263,N_3808,N_1079);
or U9264 (N_9264,N_2972,N_2769);
and U9265 (N_9265,N_167,N_4984);
xor U9266 (N_9266,N_444,N_801);
xnor U9267 (N_9267,N_4082,N_2539);
nand U9268 (N_9268,N_4136,N_1838);
xnor U9269 (N_9269,N_4947,N_1571);
nand U9270 (N_9270,N_3705,N_3304);
and U9271 (N_9271,N_2936,N_4571);
and U9272 (N_9272,N_312,N_4923);
or U9273 (N_9273,N_2805,N_1705);
nand U9274 (N_9274,N_1386,N_2367);
xor U9275 (N_9275,N_4343,N_2447);
or U9276 (N_9276,N_4267,N_311);
xor U9277 (N_9277,N_1528,N_2422);
and U9278 (N_9278,N_73,N_4857);
nor U9279 (N_9279,N_291,N_1950);
nor U9280 (N_9280,N_3825,N_4345);
nand U9281 (N_9281,N_4901,N_4341);
and U9282 (N_9282,N_3685,N_4356);
nand U9283 (N_9283,N_1788,N_4169);
xnor U9284 (N_9284,N_576,N_508);
xnor U9285 (N_9285,N_4311,N_2420);
or U9286 (N_9286,N_179,N_619);
nand U9287 (N_9287,N_3089,N_1247);
xnor U9288 (N_9288,N_1552,N_2307);
nand U9289 (N_9289,N_2026,N_6);
nand U9290 (N_9290,N_1457,N_4424);
nor U9291 (N_9291,N_4069,N_3405);
and U9292 (N_9292,N_1422,N_997);
xnor U9293 (N_9293,N_3232,N_517);
xor U9294 (N_9294,N_1825,N_4553);
nand U9295 (N_9295,N_4862,N_4864);
xor U9296 (N_9296,N_2269,N_3371);
or U9297 (N_9297,N_2136,N_4418);
or U9298 (N_9298,N_1971,N_416);
nand U9299 (N_9299,N_1271,N_437);
nor U9300 (N_9300,N_2927,N_731);
nand U9301 (N_9301,N_206,N_4767);
and U9302 (N_9302,N_4216,N_519);
xor U9303 (N_9303,N_2103,N_1974);
nand U9304 (N_9304,N_4657,N_413);
and U9305 (N_9305,N_4824,N_4034);
xor U9306 (N_9306,N_4869,N_3809);
nor U9307 (N_9307,N_1656,N_3584);
xnor U9308 (N_9308,N_1722,N_4066);
nand U9309 (N_9309,N_3394,N_1532);
nor U9310 (N_9310,N_4628,N_498);
or U9311 (N_9311,N_1165,N_2166);
and U9312 (N_9312,N_1197,N_3798);
nand U9313 (N_9313,N_7,N_582);
nor U9314 (N_9314,N_3608,N_1642);
and U9315 (N_9315,N_3662,N_1515);
and U9316 (N_9316,N_1253,N_4237);
nand U9317 (N_9317,N_176,N_4269);
nor U9318 (N_9318,N_2729,N_536);
nor U9319 (N_9319,N_4633,N_256);
or U9320 (N_9320,N_3177,N_3198);
or U9321 (N_9321,N_61,N_4865);
nand U9322 (N_9322,N_1680,N_2970);
nand U9323 (N_9323,N_3535,N_4425);
nor U9324 (N_9324,N_4939,N_4433);
nor U9325 (N_9325,N_1032,N_4451);
nor U9326 (N_9326,N_2645,N_4584);
nor U9327 (N_9327,N_1697,N_4224);
and U9328 (N_9328,N_3951,N_3788);
xor U9329 (N_9329,N_3580,N_2728);
and U9330 (N_9330,N_2437,N_2410);
xor U9331 (N_9331,N_1468,N_2937);
or U9332 (N_9332,N_3456,N_4833);
nand U9333 (N_9333,N_4228,N_2459);
nand U9334 (N_9334,N_4341,N_3848);
nor U9335 (N_9335,N_732,N_4876);
nor U9336 (N_9336,N_4800,N_4657);
nand U9337 (N_9337,N_2932,N_1740);
nor U9338 (N_9338,N_2899,N_3049);
nor U9339 (N_9339,N_934,N_88);
and U9340 (N_9340,N_3581,N_4135);
and U9341 (N_9341,N_2971,N_3685);
or U9342 (N_9342,N_629,N_1408);
nor U9343 (N_9343,N_1374,N_4221);
or U9344 (N_9344,N_3021,N_3565);
xor U9345 (N_9345,N_2105,N_861);
nand U9346 (N_9346,N_3477,N_4454);
or U9347 (N_9347,N_385,N_4620);
and U9348 (N_9348,N_1585,N_2178);
and U9349 (N_9349,N_858,N_3369);
or U9350 (N_9350,N_3053,N_1166);
nand U9351 (N_9351,N_3762,N_1691);
xnor U9352 (N_9352,N_654,N_844);
and U9353 (N_9353,N_281,N_2758);
or U9354 (N_9354,N_740,N_105);
or U9355 (N_9355,N_3553,N_2251);
nand U9356 (N_9356,N_1699,N_2417);
nand U9357 (N_9357,N_96,N_2017);
nor U9358 (N_9358,N_1106,N_3969);
nor U9359 (N_9359,N_2862,N_1352);
xnor U9360 (N_9360,N_515,N_1266);
and U9361 (N_9361,N_3365,N_470);
and U9362 (N_9362,N_1551,N_3767);
nor U9363 (N_9363,N_2222,N_4496);
and U9364 (N_9364,N_4526,N_2106);
nand U9365 (N_9365,N_1902,N_1514);
nor U9366 (N_9366,N_4567,N_4081);
nand U9367 (N_9367,N_1886,N_3189);
and U9368 (N_9368,N_39,N_4052);
xor U9369 (N_9369,N_3206,N_2183);
xnor U9370 (N_9370,N_627,N_1669);
or U9371 (N_9371,N_1161,N_1831);
or U9372 (N_9372,N_4443,N_908);
or U9373 (N_9373,N_1486,N_1036);
and U9374 (N_9374,N_3988,N_1949);
xnor U9375 (N_9375,N_3907,N_3674);
nor U9376 (N_9376,N_2225,N_3315);
nand U9377 (N_9377,N_491,N_3992);
nor U9378 (N_9378,N_2735,N_3833);
and U9379 (N_9379,N_196,N_2391);
or U9380 (N_9380,N_3020,N_1651);
or U9381 (N_9381,N_2703,N_3905);
or U9382 (N_9382,N_117,N_1905);
or U9383 (N_9383,N_1132,N_4164);
or U9384 (N_9384,N_4181,N_547);
and U9385 (N_9385,N_3679,N_113);
and U9386 (N_9386,N_1846,N_2818);
xor U9387 (N_9387,N_2720,N_4377);
and U9388 (N_9388,N_999,N_1055);
xor U9389 (N_9389,N_4891,N_4174);
xor U9390 (N_9390,N_4228,N_2344);
or U9391 (N_9391,N_2427,N_3588);
nor U9392 (N_9392,N_3744,N_394);
nand U9393 (N_9393,N_1205,N_1727);
nand U9394 (N_9394,N_267,N_987);
nand U9395 (N_9395,N_140,N_662);
or U9396 (N_9396,N_4697,N_410);
or U9397 (N_9397,N_1077,N_2901);
nand U9398 (N_9398,N_2645,N_4636);
nor U9399 (N_9399,N_3007,N_880);
xor U9400 (N_9400,N_63,N_3501);
xnor U9401 (N_9401,N_35,N_314);
xor U9402 (N_9402,N_1253,N_420);
nand U9403 (N_9403,N_1022,N_2313);
or U9404 (N_9404,N_3323,N_2132);
or U9405 (N_9405,N_1537,N_537);
nor U9406 (N_9406,N_235,N_1865);
and U9407 (N_9407,N_4269,N_4339);
nand U9408 (N_9408,N_1973,N_1705);
and U9409 (N_9409,N_3160,N_371);
and U9410 (N_9410,N_4973,N_4942);
xor U9411 (N_9411,N_3122,N_340);
nand U9412 (N_9412,N_410,N_521);
or U9413 (N_9413,N_1840,N_3584);
nor U9414 (N_9414,N_3207,N_1674);
nand U9415 (N_9415,N_1161,N_3359);
nand U9416 (N_9416,N_2551,N_1022);
xor U9417 (N_9417,N_2652,N_317);
xor U9418 (N_9418,N_3086,N_2270);
or U9419 (N_9419,N_3633,N_1085);
nor U9420 (N_9420,N_3099,N_2658);
nor U9421 (N_9421,N_4645,N_3954);
xnor U9422 (N_9422,N_2190,N_1914);
or U9423 (N_9423,N_814,N_2500);
and U9424 (N_9424,N_1179,N_2285);
and U9425 (N_9425,N_2340,N_2231);
or U9426 (N_9426,N_398,N_4514);
or U9427 (N_9427,N_777,N_2753);
and U9428 (N_9428,N_4331,N_772);
nor U9429 (N_9429,N_1509,N_414);
xor U9430 (N_9430,N_3591,N_4388);
nand U9431 (N_9431,N_4737,N_3307);
xor U9432 (N_9432,N_627,N_4142);
nand U9433 (N_9433,N_4532,N_2192);
or U9434 (N_9434,N_4683,N_2911);
xnor U9435 (N_9435,N_2534,N_4538);
nand U9436 (N_9436,N_1418,N_2531);
xnor U9437 (N_9437,N_1603,N_522);
nand U9438 (N_9438,N_3395,N_1423);
and U9439 (N_9439,N_1873,N_2808);
nand U9440 (N_9440,N_744,N_4966);
or U9441 (N_9441,N_4612,N_1588);
xnor U9442 (N_9442,N_4261,N_561);
nor U9443 (N_9443,N_1855,N_3299);
xnor U9444 (N_9444,N_1526,N_1462);
nor U9445 (N_9445,N_4812,N_3182);
or U9446 (N_9446,N_3524,N_4214);
nor U9447 (N_9447,N_2308,N_1625);
and U9448 (N_9448,N_98,N_2550);
nor U9449 (N_9449,N_1724,N_1918);
nor U9450 (N_9450,N_1743,N_84);
nand U9451 (N_9451,N_2675,N_2265);
or U9452 (N_9452,N_1558,N_684);
or U9453 (N_9453,N_716,N_2442);
nand U9454 (N_9454,N_3916,N_4579);
nor U9455 (N_9455,N_2606,N_4481);
or U9456 (N_9456,N_656,N_3623);
xor U9457 (N_9457,N_2991,N_3546);
or U9458 (N_9458,N_1420,N_1490);
or U9459 (N_9459,N_4669,N_2373);
or U9460 (N_9460,N_2977,N_2227);
nand U9461 (N_9461,N_596,N_3924);
and U9462 (N_9462,N_2232,N_4372);
or U9463 (N_9463,N_1652,N_709);
nor U9464 (N_9464,N_1252,N_1065);
nor U9465 (N_9465,N_49,N_1557);
nor U9466 (N_9466,N_1500,N_1171);
xnor U9467 (N_9467,N_1479,N_4873);
or U9468 (N_9468,N_91,N_4976);
or U9469 (N_9469,N_3626,N_2492);
and U9470 (N_9470,N_3557,N_3642);
and U9471 (N_9471,N_1634,N_4862);
nand U9472 (N_9472,N_2164,N_4071);
and U9473 (N_9473,N_2351,N_3576);
and U9474 (N_9474,N_3488,N_2798);
or U9475 (N_9475,N_2900,N_3198);
nand U9476 (N_9476,N_414,N_527);
and U9477 (N_9477,N_3487,N_4598);
and U9478 (N_9478,N_1409,N_2674);
or U9479 (N_9479,N_2346,N_2164);
xor U9480 (N_9480,N_2078,N_975);
and U9481 (N_9481,N_871,N_248);
xor U9482 (N_9482,N_1136,N_4933);
nor U9483 (N_9483,N_3556,N_4886);
and U9484 (N_9484,N_4971,N_1763);
and U9485 (N_9485,N_2972,N_602);
nand U9486 (N_9486,N_3643,N_3325);
nor U9487 (N_9487,N_845,N_4689);
or U9488 (N_9488,N_1287,N_4257);
nand U9489 (N_9489,N_4819,N_890);
and U9490 (N_9490,N_4765,N_1928);
and U9491 (N_9491,N_1832,N_2401);
nor U9492 (N_9492,N_2572,N_185);
nor U9493 (N_9493,N_2355,N_680);
and U9494 (N_9494,N_3492,N_954);
xor U9495 (N_9495,N_43,N_4899);
and U9496 (N_9496,N_4089,N_456);
nand U9497 (N_9497,N_1216,N_1636);
nor U9498 (N_9498,N_1215,N_164);
nor U9499 (N_9499,N_694,N_4591);
nand U9500 (N_9500,N_1476,N_2561);
or U9501 (N_9501,N_4796,N_375);
or U9502 (N_9502,N_2266,N_2470);
nand U9503 (N_9503,N_4392,N_427);
xor U9504 (N_9504,N_2869,N_2709);
nor U9505 (N_9505,N_1056,N_4966);
or U9506 (N_9506,N_595,N_1618);
nor U9507 (N_9507,N_3996,N_4620);
nand U9508 (N_9508,N_3962,N_4673);
nand U9509 (N_9509,N_2764,N_4417);
or U9510 (N_9510,N_2398,N_800);
nor U9511 (N_9511,N_2781,N_1322);
nor U9512 (N_9512,N_3230,N_2222);
or U9513 (N_9513,N_4018,N_132);
or U9514 (N_9514,N_4698,N_1598);
or U9515 (N_9515,N_4268,N_1026);
nor U9516 (N_9516,N_3080,N_3776);
xnor U9517 (N_9517,N_420,N_4017);
or U9518 (N_9518,N_1532,N_3620);
or U9519 (N_9519,N_1591,N_1363);
or U9520 (N_9520,N_40,N_17);
and U9521 (N_9521,N_2905,N_2539);
or U9522 (N_9522,N_1223,N_2717);
and U9523 (N_9523,N_2014,N_3052);
or U9524 (N_9524,N_969,N_1879);
or U9525 (N_9525,N_3915,N_1219);
and U9526 (N_9526,N_391,N_1465);
nand U9527 (N_9527,N_1049,N_813);
nor U9528 (N_9528,N_80,N_1630);
nand U9529 (N_9529,N_2432,N_3003);
or U9530 (N_9530,N_613,N_1903);
or U9531 (N_9531,N_317,N_607);
nor U9532 (N_9532,N_141,N_1060);
xor U9533 (N_9533,N_762,N_4030);
nor U9534 (N_9534,N_2419,N_249);
nor U9535 (N_9535,N_1078,N_1852);
nor U9536 (N_9536,N_2315,N_2446);
xnor U9537 (N_9537,N_1349,N_1878);
nor U9538 (N_9538,N_2583,N_1854);
nor U9539 (N_9539,N_1640,N_2749);
or U9540 (N_9540,N_866,N_4060);
nand U9541 (N_9541,N_2665,N_1675);
xnor U9542 (N_9542,N_3163,N_3942);
xnor U9543 (N_9543,N_3484,N_1548);
and U9544 (N_9544,N_1558,N_1011);
nor U9545 (N_9545,N_3473,N_3069);
nor U9546 (N_9546,N_12,N_1887);
xor U9547 (N_9547,N_1096,N_4918);
nand U9548 (N_9548,N_1731,N_1231);
xor U9549 (N_9549,N_2156,N_2077);
nand U9550 (N_9550,N_3693,N_2680);
or U9551 (N_9551,N_3015,N_2812);
and U9552 (N_9552,N_955,N_337);
or U9553 (N_9553,N_1381,N_4722);
xor U9554 (N_9554,N_153,N_4057);
nor U9555 (N_9555,N_2240,N_3004);
and U9556 (N_9556,N_656,N_4813);
or U9557 (N_9557,N_485,N_2669);
xnor U9558 (N_9558,N_1913,N_828);
xor U9559 (N_9559,N_4495,N_2024);
nand U9560 (N_9560,N_4081,N_4350);
nand U9561 (N_9561,N_1227,N_416);
or U9562 (N_9562,N_2935,N_3698);
nor U9563 (N_9563,N_3265,N_4702);
nor U9564 (N_9564,N_2009,N_1597);
and U9565 (N_9565,N_2102,N_3876);
nor U9566 (N_9566,N_1723,N_3939);
xnor U9567 (N_9567,N_3429,N_1413);
and U9568 (N_9568,N_3075,N_977);
or U9569 (N_9569,N_3783,N_799);
nand U9570 (N_9570,N_4980,N_3713);
xnor U9571 (N_9571,N_4226,N_3070);
and U9572 (N_9572,N_4693,N_1656);
nor U9573 (N_9573,N_792,N_2574);
or U9574 (N_9574,N_4452,N_1696);
nor U9575 (N_9575,N_4359,N_1558);
nand U9576 (N_9576,N_2130,N_3000);
nand U9577 (N_9577,N_824,N_3470);
nor U9578 (N_9578,N_4646,N_152);
nor U9579 (N_9579,N_2394,N_4672);
xnor U9580 (N_9580,N_3566,N_4441);
nor U9581 (N_9581,N_1154,N_800);
or U9582 (N_9582,N_2512,N_3532);
and U9583 (N_9583,N_3731,N_3889);
xnor U9584 (N_9584,N_1864,N_1499);
nand U9585 (N_9585,N_3722,N_2703);
nor U9586 (N_9586,N_2632,N_4863);
nand U9587 (N_9587,N_4439,N_4252);
nor U9588 (N_9588,N_1280,N_3313);
and U9589 (N_9589,N_2358,N_3463);
and U9590 (N_9590,N_77,N_806);
or U9591 (N_9591,N_190,N_1985);
nor U9592 (N_9592,N_428,N_4311);
and U9593 (N_9593,N_1817,N_4242);
and U9594 (N_9594,N_1727,N_2576);
nand U9595 (N_9595,N_4352,N_3374);
or U9596 (N_9596,N_3279,N_1184);
nand U9597 (N_9597,N_2006,N_4714);
xnor U9598 (N_9598,N_2989,N_606);
and U9599 (N_9599,N_649,N_1513);
xnor U9600 (N_9600,N_3535,N_4814);
and U9601 (N_9601,N_1393,N_237);
or U9602 (N_9602,N_2225,N_2233);
or U9603 (N_9603,N_4659,N_4655);
xor U9604 (N_9604,N_3226,N_1099);
xnor U9605 (N_9605,N_3727,N_499);
nor U9606 (N_9606,N_551,N_309);
or U9607 (N_9607,N_4181,N_1229);
nand U9608 (N_9608,N_3808,N_2189);
and U9609 (N_9609,N_4730,N_1574);
or U9610 (N_9610,N_4651,N_2871);
and U9611 (N_9611,N_3963,N_3187);
xnor U9612 (N_9612,N_62,N_725);
nand U9613 (N_9613,N_1558,N_1725);
nand U9614 (N_9614,N_3317,N_2294);
or U9615 (N_9615,N_3675,N_1452);
or U9616 (N_9616,N_4135,N_2459);
nand U9617 (N_9617,N_4653,N_4968);
nor U9618 (N_9618,N_1612,N_2877);
xor U9619 (N_9619,N_2036,N_4623);
nor U9620 (N_9620,N_4254,N_591);
or U9621 (N_9621,N_1090,N_3480);
or U9622 (N_9622,N_4288,N_1182);
nor U9623 (N_9623,N_3060,N_4689);
and U9624 (N_9624,N_1475,N_4957);
nand U9625 (N_9625,N_1503,N_957);
xnor U9626 (N_9626,N_3533,N_131);
nand U9627 (N_9627,N_3686,N_1939);
or U9628 (N_9628,N_4030,N_989);
nor U9629 (N_9629,N_4188,N_2032);
xnor U9630 (N_9630,N_2603,N_4043);
or U9631 (N_9631,N_3605,N_4304);
or U9632 (N_9632,N_4567,N_786);
nor U9633 (N_9633,N_2779,N_329);
or U9634 (N_9634,N_4634,N_3919);
nand U9635 (N_9635,N_2139,N_676);
nand U9636 (N_9636,N_4739,N_3554);
and U9637 (N_9637,N_4320,N_4404);
nand U9638 (N_9638,N_276,N_639);
and U9639 (N_9639,N_3371,N_2998);
nand U9640 (N_9640,N_4439,N_2554);
xnor U9641 (N_9641,N_2079,N_3077);
and U9642 (N_9642,N_4309,N_3525);
and U9643 (N_9643,N_1537,N_4907);
nand U9644 (N_9644,N_4814,N_1671);
nand U9645 (N_9645,N_1230,N_2551);
or U9646 (N_9646,N_2085,N_4498);
and U9647 (N_9647,N_3366,N_4628);
xnor U9648 (N_9648,N_1184,N_4546);
nor U9649 (N_9649,N_2741,N_821);
nand U9650 (N_9650,N_1563,N_1975);
or U9651 (N_9651,N_4652,N_2517);
xnor U9652 (N_9652,N_2598,N_3705);
nand U9653 (N_9653,N_4321,N_4811);
and U9654 (N_9654,N_177,N_977);
nor U9655 (N_9655,N_2159,N_4679);
nor U9656 (N_9656,N_1071,N_953);
and U9657 (N_9657,N_2190,N_4211);
and U9658 (N_9658,N_569,N_2053);
nor U9659 (N_9659,N_2251,N_4544);
and U9660 (N_9660,N_1545,N_174);
nor U9661 (N_9661,N_163,N_2656);
nand U9662 (N_9662,N_2646,N_3569);
nor U9663 (N_9663,N_4677,N_723);
nor U9664 (N_9664,N_3060,N_3137);
nor U9665 (N_9665,N_1278,N_2451);
nor U9666 (N_9666,N_4212,N_4605);
and U9667 (N_9667,N_3914,N_4673);
nor U9668 (N_9668,N_3976,N_4259);
nand U9669 (N_9669,N_268,N_1821);
or U9670 (N_9670,N_1668,N_459);
nand U9671 (N_9671,N_4564,N_4266);
and U9672 (N_9672,N_4241,N_122);
nand U9673 (N_9673,N_2510,N_809);
nand U9674 (N_9674,N_771,N_291);
nand U9675 (N_9675,N_3961,N_1118);
nor U9676 (N_9676,N_187,N_2569);
nand U9677 (N_9677,N_3734,N_508);
xnor U9678 (N_9678,N_2764,N_2070);
xnor U9679 (N_9679,N_3945,N_4439);
or U9680 (N_9680,N_3057,N_3879);
xor U9681 (N_9681,N_4096,N_1536);
nand U9682 (N_9682,N_2371,N_78);
and U9683 (N_9683,N_3017,N_2424);
nor U9684 (N_9684,N_598,N_4915);
or U9685 (N_9685,N_4033,N_4583);
nor U9686 (N_9686,N_1846,N_2328);
nand U9687 (N_9687,N_2822,N_2160);
or U9688 (N_9688,N_1999,N_4008);
or U9689 (N_9689,N_2781,N_459);
nor U9690 (N_9690,N_3096,N_2273);
or U9691 (N_9691,N_1782,N_1221);
or U9692 (N_9692,N_1416,N_792);
xor U9693 (N_9693,N_2476,N_3880);
and U9694 (N_9694,N_335,N_332);
xor U9695 (N_9695,N_2184,N_3444);
xnor U9696 (N_9696,N_4832,N_4736);
nor U9697 (N_9697,N_2771,N_1793);
and U9698 (N_9698,N_3612,N_3926);
or U9699 (N_9699,N_2823,N_1359);
nand U9700 (N_9700,N_1330,N_3842);
or U9701 (N_9701,N_1056,N_533);
or U9702 (N_9702,N_3891,N_2929);
nor U9703 (N_9703,N_4801,N_4532);
nand U9704 (N_9704,N_4820,N_3033);
xnor U9705 (N_9705,N_1231,N_394);
xor U9706 (N_9706,N_2136,N_2372);
or U9707 (N_9707,N_1587,N_331);
xnor U9708 (N_9708,N_2414,N_1430);
and U9709 (N_9709,N_4938,N_2446);
or U9710 (N_9710,N_4880,N_2868);
nand U9711 (N_9711,N_4516,N_2456);
and U9712 (N_9712,N_4380,N_4467);
xnor U9713 (N_9713,N_1058,N_3431);
or U9714 (N_9714,N_4337,N_4104);
nor U9715 (N_9715,N_3889,N_2383);
and U9716 (N_9716,N_1310,N_1432);
nor U9717 (N_9717,N_2794,N_1941);
nor U9718 (N_9718,N_2698,N_358);
or U9719 (N_9719,N_870,N_1777);
xor U9720 (N_9720,N_1449,N_1798);
nor U9721 (N_9721,N_4003,N_3968);
xnor U9722 (N_9722,N_3883,N_3256);
xnor U9723 (N_9723,N_3992,N_1942);
xor U9724 (N_9724,N_4985,N_4573);
or U9725 (N_9725,N_4183,N_2106);
nand U9726 (N_9726,N_3590,N_4335);
or U9727 (N_9727,N_3859,N_2387);
nand U9728 (N_9728,N_3483,N_4276);
xor U9729 (N_9729,N_1260,N_2563);
xor U9730 (N_9730,N_2460,N_1437);
nand U9731 (N_9731,N_3556,N_1583);
nand U9732 (N_9732,N_3525,N_659);
or U9733 (N_9733,N_2621,N_1002);
nand U9734 (N_9734,N_3323,N_1685);
xor U9735 (N_9735,N_3872,N_3350);
nor U9736 (N_9736,N_659,N_129);
nand U9737 (N_9737,N_4792,N_2200);
xnor U9738 (N_9738,N_3490,N_2113);
nor U9739 (N_9739,N_4518,N_3181);
nand U9740 (N_9740,N_4975,N_895);
and U9741 (N_9741,N_111,N_3505);
and U9742 (N_9742,N_3454,N_1117);
nor U9743 (N_9743,N_879,N_1681);
and U9744 (N_9744,N_3998,N_2798);
or U9745 (N_9745,N_4378,N_1362);
nand U9746 (N_9746,N_1161,N_3850);
nor U9747 (N_9747,N_3643,N_1266);
nor U9748 (N_9748,N_1263,N_2552);
and U9749 (N_9749,N_3176,N_1151);
nor U9750 (N_9750,N_1969,N_370);
nand U9751 (N_9751,N_1535,N_2694);
nand U9752 (N_9752,N_3860,N_1535);
xnor U9753 (N_9753,N_1344,N_4334);
and U9754 (N_9754,N_4622,N_1740);
and U9755 (N_9755,N_3717,N_4204);
nor U9756 (N_9756,N_1577,N_811);
and U9757 (N_9757,N_4683,N_174);
or U9758 (N_9758,N_2054,N_664);
nand U9759 (N_9759,N_147,N_3258);
nor U9760 (N_9760,N_182,N_4008);
and U9761 (N_9761,N_1141,N_1194);
and U9762 (N_9762,N_2955,N_4940);
or U9763 (N_9763,N_1211,N_355);
nand U9764 (N_9764,N_35,N_194);
or U9765 (N_9765,N_4181,N_4649);
nand U9766 (N_9766,N_1271,N_2918);
nand U9767 (N_9767,N_3811,N_3031);
nand U9768 (N_9768,N_3379,N_1352);
or U9769 (N_9769,N_4628,N_652);
xnor U9770 (N_9770,N_3828,N_1159);
xnor U9771 (N_9771,N_1384,N_2930);
and U9772 (N_9772,N_2643,N_4353);
xnor U9773 (N_9773,N_1266,N_963);
nand U9774 (N_9774,N_1523,N_3783);
nor U9775 (N_9775,N_3582,N_1966);
nor U9776 (N_9776,N_4717,N_1183);
or U9777 (N_9777,N_2166,N_1717);
or U9778 (N_9778,N_196,N_1439);
or U9779 (N_9779,N_3225,N_2027);
or U9780 (N_9780,N_524,N_4177);
and U9781 (N_9781,N_2077,N_1916);
and U9782 (N_9782,N_2013,N_4425);
nand U9783 (N_9783,N_1097,N_4842);
or U9784 (N_9784,N_2845,N_2477);
or U9785 (N_9785,N_695,N_2383);
and U9786 (N_9786,N_1174,N_4587);
xor U9787 (N_9787,N_3356,N_2784);
xnor U9788 (N_9788,N_3223,N_1105);
xor U9789 (N_9789,N_1465,N_486);
or U9790 (N_9790,N_2055,N_3605);
and U9791 (N_9791,N_3133,N_3553);
and U9792 (N_9792,N_567,N_144);
and U9793 (N_9793,N_2721,N_2298);
or U9794 (N_9794,N_4183,N_3131);
nor U9795 (N_9795,N_305,N_2746);
nand U9796 (N_9796,N_2313,N_2580);
xnor U9797 (N_9797,N_2693,N_1019);
xnor U9798 (N_9798,N_3334,N_4733);
nor U9799 (N_9799,N_4791,N_4582);
and U9800 (N_9800,N_538,N_3081);
or U9801 (N_9801,N_972,N_112);
and U9802 (N_9802,N_1068,N_2151);
nor U9803 (N_9803,N_1137,N_4044);
xnor U9804 (N_9804,N_4622,N_2611);
or U9805 (N_9805,N_3294,N_849);
nand U9806 (N_9806,N_4720,N_2901);
nand U9807 (N_9807,N_1955,N_19);
xnor U9808 (N_9808,N_2012,N_2301);
xnor U9809 (N_9809,N_2204,N_578);
nand U9810 (N_9810,N_1954,N_4210);
or U9811 (N_9811,N_2305,N_1804);
xor U9812 (N_9812,N_1353,N_3931);
nor U9813 (N_9813,N_679,N_2462);
nand U9814 (N_9814,N_1336,N_1661);
and U9815 (N_9815,N_3095,N_915);
and U9816 (N_9816,N_3201,N_486);
xnor U9817 (N_9817,N_4830,N_4418);
xnor U9818 (N_9818,N_4500,N_3268);
nor U9819 (N_9819,N_2457,N_544);
nand U9820 (N_9820,N_205,N_1203);
and U9821 (N_9821,N_4371,N_287);
and U9822 (N_9822,N_3501,N_4183);
nand U9823 (N_9823,N_901,N_4519);
and U9824 (N_9824,N_1320,N_3698);
or U9825 (N_9825,N_3926,N_1369);
or U9826 (N_9826,N_2814,N_2556);
nor U9827 (N_9827,N_1884,N_708);
and U9828 (N_9828,N_1067,N_3501);
and U9829 (N_9829,N_1399,N_4193);
xnor U9830 (N_9830,N_1345,N_2507);
and U9831 (N_9831,N_3150,N_2301);
xnor U9832 (N_9832,N_3930,N_1848);
nor U9833 (N_9833,N_3450,N_1916);
xnor U9834 (N_9834,N_169,N_1682);
and U9835 (N_9835,N_3289,N_3878);
or U9836 (N_9836,N_2190,N_3999);
nand U9837 (N_9837,N_1803,N_2001);
nand U9838 (N_9838,N_4388,N_4918);
nand U9839 (N_9839,N_4582,N_1872);
xor U9840 (N_9840,N_1380,N_3417);
xor U9841 (N_9841,N_3420,N_1925);
nor U9842 (N_9842,N_2718,N_1924);
xnor U9843 (N_9843,N_1486,N_2286);
xor U9844 (N_9844,N_3011,N_1157);
nand U9845 (N_9845,N_3781,N_2369);
and U9846 (N_9846,N_2985,N_504);
nor U9847 (N_9847,N_2553,N_3804);
nor U9848 (N_9848,N_4939,N_1957);
or U9849 (N_9849,N_1887,N_4749);
nor U9850 (N_9850,N_3722,N_4560);
and U9851 (N_9851,N_1829,N_52);
and U9852 (N_9852,N_605,N_2584);
and U9853 (N_9853,N_2935,N_100);
nor U9854 (N_9854,N_1882,N_962);
xor U9855 (N_9855,N_3260,N_2459);
xnor U9856 (N_9856,N_1595,N_2783);
or U9857 (N_9857,N_3481,N_3092);
nor U9858 (N_9858,N_735,N_4220);
or U9859 (N_9859,N_872,N_1033);
nand U9860 (N_9860,N_4925,N_873);
or U9861 (N_9861,N_607,N_3861);
xor U9862 (N_9862,N_63,N_1961);
xor U9863 (N_9863,N_341,N_2052);
nor U9864 (N_9864,N_3916,N_3069);
or U9865 (N_9865,N_1543,N_236);
nor U9866 (N_9866,N_4078,N_4409);
and U9867 (N_9867,N_4670,N_3288);
nor U9868 (N_9868,N_3210,N_2940);
xnor U9869 (N_9869,N_3497,N_0);
or U9870 (N_9870,N_1360,N_3963);
and U9871 (N_9871,N_4466,N_3663);
xor U9872 (N_9872,N_2852,N_2250);
nand U9873 (N_9873,N_4670,N_4682);
xor U9874 (N_9874,N_3263,N_2838);
nand U9875 (N_9875,N_422,N_3313);
nand U9876 (N_9876,N_80,N_4969);
or U9877 (N_9877,N_867,N_1689);
nor U9878 (N_9878,N_838,N_4057);
nand U9879 (N_9879,N_2545,N_3509);
nand U9880 (N_9880,N_581,N_76);
and U9881 (N_9881,N_685,N_3058);
nand U9882 (N_9882,N_592,N_1234);
nand U9883 (N_9883,N_3559,N_2354);
and U9884 (N_9884,N_890,N_4036);
and U9885 (N_9885,N_1093,N_1114);
nor U9886 (N_9886,N_3086,N_3050);
nor U9887 (N_9887,N_3835,N_234);
nand U9888 (N_9888,N_2634,N_1247);
xnor U9889 (N_9889,N_1554,N_4937);
or U9890 (N_9890,N_1038,N_4106);
and U9891 (N_9891,N_1048,N_1722);
nor U9892 (N_9892,N_1667,N_1405);
or U9893 (N_9893,N_3847,N_2972);
nand U9894 (N_9894,N_2085,N_1281);
nand U9895 (N_9895,N_3789,N_933);
and U9896 (N_9896,N_2548,N_3112);
and U9897 (N_9897,N_3780,N_3863);
nand U9898 (N_9898,N_4401,N_1516);
and U9899 (N_9899,N_244,N_4544);
nor U9900 (N_9900,N_889,N_4455);
nor U9901 (N_9901,N_1229,N_63);
nand U9902 (N_9902,N_4666,N_1853);
or U9903 (N_9903,N_2641,N_2958);
nor U9904 (N_9904,N_4969,N_1619);
or U9905 (N_9905,N_870,N_1463);
nand U9906 (N_9906,N_2612,N_3586);
nand U9907 (N_9907,N_2356,N_550);
and U9908 (N_9908,N_1210,N_3964);
nor U9909 (N_9909,N_4047,N_975);
nand U9910 (N_9910,N_263,N_1562);
or U9911 (N_9911,N_3140,N_4329);
and U9912 (N_9912,N_1267,N_4353);
and U9913 (N_9913,N_3643,N_2892);
and U9914 (N_9914,N_4539,N_4309);
xnor U9915 (N_9915,N_3493,N_4535);
nor U9916 (N_9916,N_4583,N_4201);
or U9917 (N_9917,N_3061,N_1753);
or U9918 (N_9918,N_2518,N_1122);
xnor U9919 (N_9919,N_337,N_4816);
xor U9920 (N_9920,N_4068,N_3288);
xnor U9921 (N_9921,N_75,N_2109);
or U9922 (N_9922,N_1863,N_4858);
or U9923 (N_9923,N_3100,N_4905);
and U9924 (N_9924,N_1265,N_255);
nand U9925 (N_9925,N_4573,N_1999);
or U9926 (N_9926,N_376,N_1063);
nand U9927 (N_9927,N_655,N_684);
and U9928 (N_9928,N_708,N_2513);
nor U9929 (N_9929,N_3082,N_3853);
nand U9930 (N_9930,N_1758,N_803);
xnor U9931 (N_9931,N_4916,N_3181);
xor U9932 (N_9932,N_918,N_4601);
nand U9933 (N_9933,N_2813,N_2703);
nor U9934 (N_9934,N_1840,N_1609);
xnor U9935 (N_9935,N_394,N_4325);
nand U9936 (N_9936,N_2273,N_2112);
or U9937 (N_9937,N_1191,N_3198);
and U9938 (N_9938,N_27,N_4318);
nand U9939 (N_9939,N_353,N_296);
nand U9940 (N_9940,N_2705,N_2558);
or U9941 (N_9941,N_4043,N_2468);
or U9942 (N_9942,N_3668,N_4641);
or U9943 (N_9943,N_4055,N_516);
nand U9944 (N_9944,N_4772,N_3852);
or U9945 (N_9945,N_1632,N_2430);
and U9946 (N_9946,N_4393,N_663);
xnor U9947 (N_9947,N_1723,N_338);
and U9948 (N_9948,N_4239,N_4112);
or U9949 (N_9949,N_1070,N_4773);
xnor U9950 (N_9950,N_3742,N_4256);
nand U9951 (N_9951,N_4394,N_3305);
or U9952 (N_9952,N_1816,N_2374);
or U9953 (N_9953,N_2899,N_4540);
and U9954 (N_9954,N_311,N_3087);
xor U9955 (N_9955,N_4431,N_1291);
xnor U9956 (N_9956,N_4434,N_4055);
nand U9957 (N_9957,N_2212,N_1325);
xor U9958 (N_9958,N_2378,N_416);
and U9959 (N_9959,N_2834,N_3369);
or U9960 (N_9960,N_661,N_353);
and U9961 (N_9961,N_3897,N_288);
and U9962 (N_9962,N_2591,N_4787);
and U9963 (N_9963,N_3882,N_4173);
or U9964 (N_9964,N_4590,N_3128);
or U9965 (N_9965,N_2100,N_3450);
and U9966 (N_9966,N_4763,N_2984);
xnor U9967 (N_9967,N_3888,N_3200);
xor U9968 (N_9968,N_3606,N_2174);
xnor U9969 (N_9969,N_1901,N_387);
and U9970 (N_9970,N_3200,N_3341);
nor U9971 (N_9971,N_89,N_46);
and U9972 (N_9972,N_381,N_2240);
xor U9973 (N_9973,N_2157,N_3651);
or U9974 (N_9974,N_1346,N_1135);
xnor U9975 (N_9975,N_1922,N_3739);
or U9976 (N_9976,N_1386,N_1244);
nor U9977 (N_9977,N_1007,N_4088);
and U9978 (N_9978,N_1540,N_3153);
nand U9979 (N_9979,N_610,N_1373);
or U9980 (N_9980,N_3700,N_3178);
and U9981 (N_9981,N_3133,N_2754);
xor U9982 (N_9982,N_4948,N_561);
nand U9983 (N_9983,N_3339,N_151);
and U9984 (N_9984,N_1432,N_3754);
nor U9985 (N_9985,N_2163,N_4101);
and U9986 (N_9986,N_1841,N_1022);
or U9987 (N_9987,N_4821,N_1955);
or U9988 (N_9988,N_2655,N_1456);
xnor U9989 (N_9989,N_4282,N_4587);
nor U9990 (N_9990,N_2463,N_1729);
xnor U9991 (N_9991,N_3690,N_3794);
nand U9992 (N_9992,N_3070,N_3483);
or U9993 (N_9993,N_3544,N_305);
or U9994 (N_9994,N_1648,N_1478);
or U9995 (N_9995,N_758,N_2711);
nor U9996 (N_9996,N_1773,N_1247);
xnor U9997 (N_9997,N_2177,N_2508);
or U9998 (N_9998,N_3390,N_4164);
or U9999 (N_9999,N_1024,N_2202);
xor U10000 (N_10000,N_7504,N_7756);
and U10001 (N_10001,N_7176,N_6659);
nand U10002 (N_10002,N_6707,N_6121);
nand U10003 (N_10003,N_7640,N_7952);
nand U10004 (N_10004,N_9032,N_6559);
and U10005 (N_10005,N_5024,N_8730);
nand U10006 (N_10006,N_9322,N_9903);
nor U10007 (N_10007,N_9979,N_6806);
nor U10008 (N_10008,N_5184,N_8173);
nand U10009 (N_10009,N_7975,N_7413);
nand U10010 (N_10010,N_5653,N_5889);
nor U10011 (N_10011,N_5754,N_6952);
nand U10012 (N_10012,N_5171,N_9277);
or U10013 (N_10013,N_7336,N_8484);
or U10014 (N_10014,N_5051,N_8994);
or U10015 (N_10015,N_8181,N_6704);
nand U10016 (N_10016,N_8851,N_8027);
or U10017 (N_10017,N_6630,N_5652);
and U10018 (N_10018,N_7401,N_8132);
nor U10019 (N_10019,N_5718,N_5032);
nand U10020 (N_10020,N_7350,N_8237);
nor U10021 (N_10021,N_8198,N_5529);
or U10022 (N_10022,N_6266,N_6591);
and U10023 (N_10023,N_9215,N_8899);
and U10024 (N_10024,N_9489,N_9835);
nand U10025 (N_10025,N_9605,N_9775);
xnor U10026 (N_10026,N_6508,N_7390);
nor U10027 (N_10027,N_9448,N_7935);
nand U10028 (N_10028,N_5021,N_5660);
nor U10029 (N_10029,N_5702,N_5404);
nor U10030 (N_10030,N_6299,N_5814);
nor U10031 (N_10031,N_5793,N_5412);
xor U10032 (N_10032,N_8457,N_7383);
nand U10033 (N_10033,N_6723,N_8210);
or U10034 (N_10034,N_8863,N_5855);
xor U10035 (N_10035,N_6878,N_8244);
nor U10036 (N_10036,N_9680,N_7110);
xor U10037 (N_10037,N_7473,N_7137);
or U10038 (N_10038,N_8679,N_9583);
xor U10039 (N_10039,N_8665,N_7923);
nand U10040 (N_10040,N_8180,N_8540);
or U10041 (N_10041,N_6535,N_9989);
nand U10042 (N_10042,N_8068,N_7204);
xor U10043 (N_10043,N_8407,N_6349);
nand U10044 (N_10044,N_5017,N_9899);
and U10045 (N_10045,N_8432,N_6692);
xnor U10046 (N_10046,N_6141,N_6946);
and U10047 (N_10047,N_8718,N_7932);
nor U10048 (N_10048,N_7910,N_8885);
xnor U10049 (N_10049,N_6588,N_5837);
or U10050 (N_10050,N_7684,N_9932);
nor U10051 (N_10051,N_9953,N_8460);
xnor U10052 (N_10052,N_9314,N_8059);
nand U10053 (N_10053,N_9201,N_6291);
nor U10054 (N_10054,N_7856,N_8448);
nor U10055 (N_10055,N_7356,N_8979);
and U10056 (N_10056,N_5294,N_5708);
and U10057 (N_10057,N_8462,N_8552);
nand U10058 (N_10058,N_8169,N_5535);
nor U10059 (N_10059,N_7876,N_5328);
or U10060 (N_10060,N_8263,N_6007);
xnor U10061 (N_10061,N_9531,N_9830);
nand U10062 (N_10062,N_9236,N_7746);
nor U10063 (N_10063,N_8382,N_5756);
or U10064 (N_10064,N_7289,N_5506);
or U10065 (N_10065,N_8528,N_8444);
or U10066 (N_10066,N_9416,N_6875);
nor U10067 (N_10067,N_8592,N_8197);
or U10068 (N_10068,N_8651,N_9450);
and U10069 (N_10069,N_9737,N_6507);
or U10070 (N_10070,N_7001,N_9476);
nand U10071 (N_10071,N_9117,N_6872);
nand U10072 (N_10072,N_9909,N_9611);
and U10073 (N_10073,N_8757,N_6445);
and U10074 (N_10074,N_7596,N_5890);
or U10075 (N_10075,N_8564,N_7706);
nor U10076 (N_10076,N_7308,N_6825);
nand U10077 (N_10077,N_6036,N_7739);
nand U10078 (N_10078,N_8813,N_6877);
and U10079 (N_10079,N_9563,N_9771);
and U10080 (N_10080,N_6844,N_5262);
xnor U10081 (N_10081,N_7243,N_8841);
nand U10082 (N_10082,N_9658,N_5533);
or U10083 (N_10083,N_7084,N_9631);
nor U10084 (N_10084,N_5170,N_9482);
xnor U10085 (N_10085,N_6705,N_8423);
or U10086 (N_10086,N_9804,N_5422);
nor U10087 (N_10087,N_5720,N_9836);
nor U10088 (N_10088,N_7688,N_7995);
xor U10089 (N_10089,N_7482,N_6841);
or U10090 (N_10090,N_8337,N_9037);
nand U10091 (N_10091,N_9128,N_9139);
nand U10092 (N_10092,N_7961,N_7208);
or U10093 (N_10093,N_8005,N_7934);
xnor U10094 (N_10094,N_6370,N_6218);
nand U10095 (N_10095,N_8390,N_6799);
xor U10096 (N_10096,N_8127,N_5210);
xor U10097 (N_10097,N_6197,N_6966);
xnor U10098 (N_10098,N_8419,N_5492);
and U10099 (N_10099,N_7116,N_6736);
xnor U10100 (N_10100,N_5717,N_5540);
nor U10101 (N_10101,N_8040,N_6161);
and U10102 (N_10102,N_7302,N_6363);
nor U10103 (N_10103,N_7380,N_8982);
or U10104 (N_10104,N_7346,N_9831);
nand U10105 (N_10105,N_8375,N_8194);
nor U10106 (N_10106,N_6654,N_6290);
and U10107 (N_10107,N_9475,N_5704);
or U10108 (N_10108,N_8230,N_9012);
or U10109 (N_10109,N_5835,N_5621);
or U10110 (N_10110,N_9387,N_8912);
and U10111 (N_10111,N_8031,N_8305);
xnor U10112 (N_10112,N_7912,N_8856);
nor U10113 (N_10113,N_5330,N_9084);
nand U10114 (N_10114,N_8107,N_9817);
nand U10115 (N_10115,N_6594,N_6770);
nor U10116 (N_10116,N_8538,N_6375);
nor U10117 (N_10117,N_9480,N_5045);
xnor U10118 (N_10118,N_7382,N_9440);
and U10119 (N_10119,N_6400,N_7462);
nor U10120 (N_10120,N_6830,N_9954);
or U10121 (N_10121,N_9855,N_8170);
nor U10122 (N_10122,N_8214,N_6509);
nor U10123 (N_10123,N_9133,N_8357);
nor U10124 (N_10124,N_7916,N_9283);
or U10125 (N_10125,N_9213,N_8531);
nand U10126 (N_10126,N_5074,N_9860);
nand U10127 (N_10127,N_5500,N_8304);
and U10128 (N_10128,N_5972,N_9821);
nand U10129 (N_10129,N_8545,N_9513);
xor U10130 (N_10130,N_6404,N_9261);
xor U10131 (N_10131,N_8036,N_7698);
xor U10132 (N_10132,N_5596,N_8478);
xnor U10133 (N_10133,N_6420,N_8971);
xnor U10134 (N_10134,N_6279,N_6766);
nor U10135 (N_10135,N_7458,N_9842);
or U10136 (N_10136,N_8355,N_9091);
nor U10137 (N_10137,N_8501,N_9704);
or U10138 (N_10138,N_6516,N_7157);
and U10139 (N_10139,N_6193,N_6503);
xnor U10140 (N_10140,N_8111,N_5005);
and U10141 (N_10141,N_5926,N_7284);
or U10142 (N_10142,N_7550,N_9711);
nand U10143 (N_10143,N_9022,N_6146);
or U10144 (N_10144,N_5900,N_5898);
or U10145 (N_10145,N_9303,N_5688);
xnor U10146 (N_10146,N_6683,N_8193);
or U10147 (N_10147,N_5914,N_7148);
or U10148 (N_10148,N_7993,N_8678);
nor U10149 (N_10149,N_8591,N_7446);
nor U10150 (N_10150,N_8482,N_7930);
nand U10151 (N_10151,N_9991,N_9025);
or U10152 (N_10152,N_7141,N_6037);
nand U10153 (N_10153,N_5950,N_8535);
and U10154 (N_10154,N_8314,N_7701);
or U10155 (N_10155,N_6694,N_7854);
nand U10156 (N_10156,N_9594,N_9079);
and U10157 (N_10157,N_9384,N_9529);
nor U10158 (N_10158,N_7601,N_5090);
nor U10159 (N_10159,N_6437,N_6016);
nor U10160 (N_10160,N_9090,N_9871);
nand U10161 (N_10161,N_9030,N_6988);
xor U10162 (N_10162,N_6747,N_8009);
nor U10163 (N_10163,N_5435,N_8511);
nand U10164 (N_10164,N_5558,N_6769);
and U10165 (N_10165,N_9016,N_9595);
and U10166 (N_10166,N_8090,N_5942);
nand U10167 (N_10167,N_8496,N_7655);
nor U10168 (N_10168,N_6274,N_7852);
nand U10169 (N_10169,N_5456,N_7206);
or U10170 (N_10170,N_5602,N_7161);
or U10171 (N_10171,N_9707,N_5482);
nor U10172 (N_10172,N_7341,N_6607);
xor U10173 (N_10173,N_6906,N_8265);
and U10174 (N_10174,N_9397,N_6265);
nand U10175 (N_10175,N_6923,N_6724);
xnor U10176 (N_10176,N_8882,N_7461);
nor U10177 (N_10177,N_9179,N_6213);
and U10178 (N_10178,N_8119,N_8183);
and U10179 (N_10179,N_9069,N_7966);
xnor U10180 (N_10180,N_5515,N_6870);
nand U10181 (N_10181,N_7285,N_5508);
nor U10182 (N_10182,N_7794,N_9156);
nor U10183 (N_10183,N_9327,N_6293);
nand U10184 (N_10184,N_9718,N_9134);
and U10185 (N_10185,N_7659,N_9412);
and U10186 (N_10186,N_9578,N_5548);
or U10187 (N_10187,N_8532,N_7787);
nor U10188 (N_10188,N_5901,N_8354);
nand U10189 (N_10189,N_5925,N_7223);
and U10190 (N_10190,N_6640,N_8056);
and U10191 (N_10191,N_8109,N_8960);
nand U10192 (N_10192,N_7928,N_6795);
nand U10193 (N_10193,N_8363,N_5603);
nor U10194 (N_10194,N_8224,N_8003);
or U10195 (N_10195,N_8365,N_6609);
xor U10196 (N_10196,N_7705,N_9269);
nor U10197 (N_10197,N_7133,N_5661);
nor U10198 (N_10198,N_8200,N_8114);
xnor U10199 (N_10199,N_9459,N_8603);
xor U10200 (N_10200,N_7047,N_5313);
and U10201 (N_10201,N_5745,N_6805);
and U10202 (N_10202,N_5115,N_8820);
xor U10203 (N_10203,N_7730,N_6267);
nor U10204 (N_10204,N_9875,N_8739);
xor U10205 (N_10205,N_8724,N_9323);
nand U10206 (N_10206,N_8586,N_6040);
xnor U10207 (N_10207,N_9306,N_6765);
or U10208 (N_10208,N_6925,N_6709);
nand U10209 (N_10209,N_6316,N_8245);
xnor U10210 (N_10210,N_8459,N_9735);
nor U10211 (N_10211,N_7445,N_7715);
or U10212 (N_10212,N_5218,N_9382);
nor U10213 (N_10213,N_5611,N_5086);
nor U10214 (N_10214,N_9944,N_7272);
and U10215 (N_10215,N_9174,N_5764);
nand U10216 (N_10216,N_7201,N_5546);
xor U10217 (N_10217,N_7604,N_6668);
nor U10218 (N_10218,N_8233,N_5655);
xor U10219 (N_10219,N_7263,N_9422);
xnor U10220 (N_10220,N_6542,N_5189);
or U10221 (N_10221,N_8774,N_5429);
xor U10222 (N_10222,N_7740,N_8389);
nor U10223 (N_10223,N_9806,N_7632);
or U10224 (N_10224,N_9266,N_5577);
or U10225 (N_10225,N_8935,N_9977);
xor U10226 (N_10226,N_5430,N_6170);
nor U10227 (N_10227,N_9437,N_5600);
or U10228 (N_10228,N_6530,N_8218);
nor U10229 (N_10229,N_5928,N_7094);
or U10230 (N_10230,N_9939,N_6350);
and U10231 (N_10231,N_7301,N_7828);
xor U10232 (N_10232,N_6063,N_7873);
nor U10233 (N_10233,N_8674,N_8662);
xor U10234 (N_10234,N_5573,N_6617);
nor U10235 (N_10235,N_9366,N_8034);
or U10236 (N_10236,N_7388,N_7674);
nand U10237 (N_10237,N_5344,N_6545);
nor U10238 (N_10238,N_7503,N_5531);
or U10239 (N_10239,N_9714,N_7191);
and U10240 (N_10240,N_9158,N_6354);
and U10241 (N_10241,N_7188,N_8556);
nand U10242 (N_10242,N_5638,N_5125);
or U10243 (N_10243,N_9495,N_8356);
nor U10244 (N_10244,N_6379,N_6132);
nor U10245 (N_10245,N_9547,N_5428);
or U10246 (N_10246,N_9003,N_7115);
nand U10247 (N_10247,N_6775,N_9007);
nor U10248 (N_10248,N_9941,N_8991);
or U10249 (N_10249,N_5331,N_7754);
nand U10250 (N_10250,N_7597,N_7300);
nand U10251 (N_10251,N_9668,N_6092);
and U10252 (N_10252,N_9031,N_8915);
xnor U10253 (N_10253,N_7216,N_9479);
or U10254 (N_10254,N_8738,N_5303);
and U10255 (N_10255,N_8806,N_9884);
and U10256 (N_10256,N_8252,N_7024);
and U10257 (N_10257,N_8765,N_9191);
xnor U10258 (N_10258,N_9596,N_6169);
nor U10259 (N_10259,N_7868,N_9061);
nor U10260 (N_10260,N_5766,N_7048);
nand U10261 (N_10261,N_7986,N_5700);
nand U10262 (N_10262,N_5671,N_7150);
nor U10263 (N_10263,N_9592,N_6285);
nand U10264 (N_10264,N_8551,N_7907);
or U10265 (N_10265,N_7689,N_5574);
xor U10266 (N_10266,N_5247,N_6103);
nand U10267 (N_10267,N_9978,N_7998);
or U10268 (N_10268,N_8996,N_7066);
xnor U10269 (N_10269,N_5259,N_9181);
and U10270 (N_10270,N_9305,N_5785);
or U10271 (N_10271,N_5453,N_8274);
xnor U10272 (N_10272,N_7325,N_7205);
and U10273 (N_10273,N_9048,N_6105);
nor U10274 (N_10274,N_8828,N_9271);
xnor U10275 (N_10275,N_5378,N_8986);
nor U10276 (N_10276,N_6821,N_6271);
nand U10277 (N_10277,N_7065,N_5784);
nand U10278 (N_10278,N_6432,N_8334);
nand U10279 (N_10279,N_6236,N_6322);
xnor U10280 (N_10280,N_9843,N_5160);
or U10281 (N_10281,N_5368,N_6577);
and U10282 (N_10282,N_6468,N_8761);
nor U10283 (N_10283,N_6690,N_5727);
and U10284 (N_10284,N_6065,N_8782);
xor U10285 (N_10285,N_8387,N_9799);
nor U10286 (N_10286,N_9778,N_9560);
and U10287 (N_10287,N_8393,N_6761);
and U10288 (N_10288,N_7328,N_9644);
and U10289 (N_10289,N_9273,N_6960);
nand U10290 (N_10290,N_8083,N_7421);
xor U10291 (N_10291,N_7843,N_6685);
nor U10292 (N_10292,N_6111,N_8420);
xor U10293 (N_10293,N_7281,N_9197);
xnor U10294 (N_10294,N_6081,N_8957);
nor U10295 (N_10295,N_6819,N_9113);
or U10296 (N_10296,N_7524,N_5758);
xor U10297 (N_10297,N_8211,N_6599);
or U10298 (N_10298,N_6084,N_9601);
nor U10299 (N_10299,N_6373,N_5995);
and U10300 (N_10300,N_8698,N_5128);
xor U10301 (N_10301,N_5141,N_9790);
nor U10302 (N_10302,N_7013,N_9343);
and U10303 (N_10303,N_5178,N_9958);
nor U10304 (N_10304,N_7766,N_8521);
nand U10305 (N_10305,N_9324,N_7927);
nor U10306 (N_10306,N_6651,N_6013);
and U10307 (N_10307,N_7997,N_5085);
nand U10308 (N_10308,N_7290,N_5131);
or U10309 (N_10309,N_8020,N_5214);
or U10310 (N_10310,N_7186,N_7653);
and U10311 (N_10311,N_9603,N_9498);
nand U10312 (N_10312,N_7909,N_7118);
nand U10313 (N_10313,N_5716,N_8923);
nor U10314 (N_10314,N_9756,N_5988);
xnor U10315 (N_10315,N_7112,N_6855);
nand U10316 (N_10316,N_7718,N_8687);
xor U10317 (N_10317,N_5846,N_6751);
or U10318 (N_10318,N_8424,N_9912);
nand U10319 (N_10319,N_5077,N_7077);
or U10320 (N_10320,N_9593,N_8617);
nand U10321 (N_10321,N_5291,N_9086);
and U10322 (N_10322,N_9577,N_9677);
xnor U10323 (N_10323,N_8134,N_8342);
or U10324 (N_10324,N_7123,N_6954);
nand U10325 (N_10325,N_5477,N_5954);
or U10326 (N_10326,N_9268,N_5615);
nor U10327 (N_10327,N_8519,N_5843);
xnor U10328 (N_10328,N_9674,N_5173);
xor U10329 (N_10329,N_9740,N_6076);
or U10330 (N_10330,N_7344,N_5049);
nand U10331 (N_10331,N_8153,N_7100);
xor U10332 (N_10332,N_6777,N_6048);
and U10333 (N_10333,N_6614,N_6242);
and U10334 (N_10334,N_9405,N_7915);
or U10335 (N_10335,N_8092,N_5955);
nand U10336 (N_10336,N_9754,N_5640);
nand U10337 (N_10337,N_8347,N_7512);
xor U10338 (N_10338,N_5795,N_5290);
and U10339 (N_10339,N_9795,N_7732);
and U10340 (N_10340,N_7426,N_9500);
or U10341 (N_10341,N_8486,N_9759);
xor U10342 (N_10342,N_7731,N_7500);
nor U10343 (N_10343,N_5812,N_9962);
xnor U10344 (N_10344,N_5877,N_5683);
or U10345 (N_10345,N_8965,N_5202);
nor U10346 (N_10346,N_6014,N_9969);
nor U10347 (N_10347,N_6713,N_9661);
nor U10348 (N_10348,N_5356,N_6849);
nand U10349 (N_10349,N_6301,N_9539);
nor U10350 (N_10350,N_6125,N_9591);
xnor U10351 (N_10351,N_6674,N_8610);
and U10352 (N_10352,N_6544,N_5695);
xor U10353 (N_10353,N_9921,N_7457);
or U10354 (N_10354,N_9087,N_6377);
or U10355 (N_10355,N_8714,N_5176);
nand U10356 (N_10356,N_9812,N_7145);
xor U10357 (N_10357,N_7054,N_7428);
nand U10358 (N_10358,N_7343,N_9581);
nand U10359 (N_10359,N_7941,N_8789);
nand U10360 (N_10360,N_5466,N_8149);
nand U10361 (N_10361,N_7536,N_9811);
xnor U10362 (N_10362,N_5333,N_7189);
or U10363 (N_10363,N_5188,N_6961);
or U10364 (N_10364,N_8522,N_5132);
xor U10365 (N_10365,N_5973,N_7257);
nor U10366 (N_10366,N_6304,N_5880);
or U10367 (N_10367,N_5617,N_6181);
or U10368 (N_10368,N_9410,N_6309);
and U10369 (N_10369,N_6405,N_9130);
or U10370 (N_10370,N_8825,N_6429);
xor U10371 (N_10371,N_8438,N_7403);
and U10372 (N_10372,N_5627,N_6112);
and U10373 (N_10373,N_6919,N_6001);
xor U10374 (N_10374,N_5732,N_7567);
and U10375 (N_10375,N_5116,N_8992);
or U10376 (N_10376,N_5989,N_6053);
nand U10377 (N_10377,N_7443,N_7763);
nor U10378 (N_10378,N_6323,N_5552);
nor U10379 (N_10379,N_5134,N_9034);
nor U10380 (N_10380,N_6757,N_9217);
and U10381 (N_10381,N_9006,N_8888);
nor U10382 (N_10382,N_7874,N_9454);
xor U10383 (N_10383,N_5020,N_8029);
xor U10384 (N_10384,N_7464,N_6671);
nor U10385 (N_10385,N_6850,N_9700);
and U10386 (N_10386,N_6984,N_6366);
xnor U10387 (N_10387,N_7518,N_5357);
xor U10388 (N_10388,N_7889,N_8947);
nand U10389 (N_10389,N_8756,N_8572);
and U10390 (N_10390,N_5042,N_9575);
xnor U10391 (N_10391,N_5455,N_8931);
xnor U10392 (N_10392,N_9224,N_9634);
nor U10393 (N_10393,N_7082,N_7316);
and U10394 (N_10394,N_6598,N_6527);
or U10395 (N_10395,N_5912,N_8008);
and U10396 (N_10396,N_7075,N_7260);
and U10397 (N_10397,N_8483,N_8509);
and U10398 (N_10398,N_7603,N_6273);
xnor U10399 (N_10399,N_5576,N_9966);
or U10400 (N_10400,N_5868,N_9911);
nor U10401 (N_10401,N_8588,N_9846);
and U10402 (N_10402,N_9227,N_6768);
or U10403 (N_10403,N_6629,N_6655);
and U10404 (N_10404,N_7859,N_8631);
nor U10405 (N_10405,N_7989,N_9237);
xnor U10406 (N_10406,N_6931,N_7072);
or U10407 (N_10407,N_7848,N_7817);
and U10408 (N_10408,N_8001,N_6744);
nand U10409 (N_10409,N_8859,N_6180);
nand U10410 (N_10410,N_6532,N_5951);
xor U10411 (N_10411,N_7644,N_8386);
nand U10412 (N_10412,N_9585,N_7449);
nand U10413 (N_10413,N_5298,N_6525);
xnor U10414 (N_10414,N_5271,N_6257);
and U10415 (N_10415,N_5364,N_7575);
xor U10416 (N_10416,N_6179,N_9630);
or U10417 (N_10417,N_7347,N_7637);
nand U10418 (N_10418,N_8557,N_6427);
or U10419 (N_10419,N_7835,N_8061);
and U10420 (N_10420,N_8704,N_8668);
or U10421 (N_10421,N_9905,N_8425);
xnor U10422 (N_10422,N_8475,N_7359);
xnor U10423 (N_10423,N_8158,N_9663);
and U10424 (N_10424,N_8801,N_6742);
xnor U10425 (N_10425,N_6650,N_5336);
and U10426 (N_10426,N_8434,N_8791);
and U10427 (N_10427,N_5886,N_6077);
and U10428 (N_10428,N_5075,N_8493);
xor U10429 (N_10429,N_9112,N_8070);
nor U10430 (N_10430,N_6455,N_7861);
or U10431 (N_10431,N_9586,N_8209);
or U10432 (N_10432,N_8440,N_9880);
nand U10433 (N_10433,N_5823,N_7781);
or U10434 (N_10434,N_5484,N_7969);
xor U10435 (N_10435,N_6666,N_5036);
or U10436 (N_10436,N_9250,N_5557);
and U10437 (N_10437,N_5337,N_6421);
nor U10438 (N_10438,N_8732,N_6512);
and U10439 (N_10439,N_9436,N_8327);
nor U10440 (N_10440,N_8227,N_5934);
nand U10441 (N_10441,N_6340,N_6985);
and U10442 (N_10442,N_9533,N_7090);
or U10443 (N_10443,N_8161,N_9355);
or U10444 (N_10444,N_5320,N_8293);
xnor U10445 (N_10445,N_7080,N_8400);
nor U10446 (N_10446,N_9329,N_7565);
xnor U10447 (N_10447,N_8156,N_9121);
and U10448 (N_10448,N_9072,N_6277);
xor U10449 (N_10449,N_8388,N_8422);
nand U10450 (N_10450,N_6556,N_7515);
or U10451 (N_10451,N_8843,N_5605);
nor U10452 (N_10452,N_5919,N_5470);
nand U10453 (N_10453,N_8259,N_5885);
or U10454 (N_10454,N_8660,N_9670);
and U10455 (N_10455,N_5816,N_8473);
or U10456 (N_10456,N_8394,N_8666);
or U10457 (N_10457,N_7944,N_5142);
nand U10458 (N_10458,N_9056,N_6246);
nand U10459 (N_10459,N_8467,N_8944);
nand U10460 (N_10460,N_8137,N_7178);
xor U10461 (N_10461,N_7508,N_9379);
xor U10462 (N_10462,N_9528,N_8159);
and U10463 (N_10463,N_9745,N_6163);
nand U10464 (N_10464,N_5146,N_9253);
xor U10465 (N_10465,N_8164,N_6049);
xnor U10466 (N_10466,N_8372,N_6823);
or U10467 (N_10467,N_5097,N_7288);
or U10468 (N_10468,N_6151,N_5003);
or U10469 (N_10469,N_6064,N_9994);
and U10470 (N_10470,N_5866,N_6857);
xor U10471 (N_10471,N_8973,N_6911);
nor U10472 (N_10472,N_7436,N_6465);
and U10473 (N_10473,N_8256,N_5463);
xor U10474 (N_10474,N_8795,N_8812);
nor U10475 (N_10475,N_5102,N_7905);
or U10476 (N_10476,N_7045,N_9627);
nand U10477 (N_10477,N_6886,N_7824);
or U10478 (N_10478,N_5607,N_8690);
nor U10479 (N_10479,N_6470,N_5936);
and U10480 (N_10480,N_6166,N_8103);
nand U10481 (N_10481,N_8606,N_5643);
nor U10482 (N_10482,N_7262,N_6029);
xor U10483 (N_10483,N_6409,N_8968);
xor U10484 (N_10484,N_6456,N_5938);
nand U10485 (N_10485,N_7842,N_7950);
nor U10486 (N_10486,N_9693,N_9936);
nor U10487 (N_10487,N_9484,N_6403);
xnor U10488 (N_10488,N_7822,N_6167);
xor U10489 (N_10489,N_5476,N_6000);
or U10490 (N_10490,N_5117,N_9341);
or U10491 (N_10491,N_9794,N_5489);
or U10492 (N_10492,N_5068,N_6815);
xor U10493 (N_10493,N_5724,N_6862);
xor U10494 (N_10494,N_6968,N_7858);
nor U10495 (N_10495,N_6533,N_9168);
and U10496 (N_10496,N_5873,N_8144);
or U10497 (N_10497,N_6200,N_8299);
and U10498 (N_10498,N_6263,N_8673);
or U10499 (N_10499,N_5610,N_8891);
xor U10500 (N_10500,N_8258,N_8167);
or U10501 (N_10501,N_9111,N_6506);
nand U10502 (N_10502,N_8909,N_5359);
nor U10503 (N_10503,N_8504,N_6009);
nor U10504 (N_10504,N_6871,N_5760);
or U10505 (N_10505,N_7744,N_8913);
and U10506 (N_10506,N_7078,N_6737);
xnor U10507 (N_10507,N_8763,N_6904);
nor U10508 (N_10508,N_5209,N_7267);
or U10509 (N_10509,N_7673,N_5984);
nor U10510 (N_10510,N_9873,N_9572);
nor U10511 (N_10511,N_5355,N_7320);
or U10512 (N_10512,N_9272,N_6555);
nor U10513 (N_10513,N_7179,N_6518);
or U10514 (N_10514,N_5465,N_5385);
or U10515 (N_10515,N_8232,N_8039);
and U10516 (N_10516,N_9774,N_7311);
xor U10517 (N_10517,N_8613,N_6498);
xnor U10518 (N_10518,N_8653,N_6526);
nor U10519 (N_10519,N_9059,N_7389);
or U10520 (N_10520,N_5806,N_6428);
and U10521 (N_10521,N_8614,N_9772);
or U10522 (N_10522,N_9096,N_9851);
and U10523 (N_10523,N_9850,N_8966);
or U10524 (N_10524,N_8582,N_8488);
nor U10525 (N_10525,N_9350,N_6492);
nor U10526 (N_10526,N_7166,N_6884);
and U10527 (N_10527,N_8223,N_7357);
and U10528 (N_10528,N_8974,N_9546);
and U10529 (N_10529,N_5311,N_6239);
xnor U10530 (N_10530,N_7541,N_8562);
xnor U10531 (N_10531,N_9141,N_7782);
xor U10532 (N_10532,N_5139,N_6991);
nor U10533 (N_10533,N_7624,N_8886);
xor U10534 (N_10534,N_6469,N_6973);
nor U10535 (N_10535,N_7943,N_6944);
nand U10536 (N_10536,N_6208,N_6188);
xnor U10537 (N_10537,N_5300,N_9276);
and U10538 (N_10538,N_9400,N_9424);
nor U10539 (N_10539,N_7361,N_8284);
and U10540 (N_10540,N_5730,N_9282);
and U10541 (N_10541,N_8202,N_5585);
xor U10542 (N_10542,N_7299,N_6453);
or U10543 (N_10543,N_8458,N_7460);
and U10544 (N_10544,N_6779,N_7778);
or U10545 (N_10545,N_9984,N_6303);
or U10546 (N_10546,N_6625,N_6441);
nand U10547 (N_10547,N_6873,N_8840);
nor U10548 (N_10548,N_5443,N_6670);
nor U10549 (N_10549,N_5895,N_8560);
xor U10550 (N_10550,N_9166,N_9260);
or U10551 (N_10551,N_7785,N_8905);
nand U10552 (N_10552,N_7083,N_8967);
xor U10553 (N_10553,N_6930,N_5062);
nand U10554 (N_10554,N_8253,N_6572);
nor U10555 (N_10555,N_8712,N_6619);
nor U10556 (N_10556,N_9917,N_9678);
or U10557 (N_10557,N_6926,N_9401);
xnor U10558 (N_10558,N_9981,N_7059);
xor U10559 (N_10559,N_8243,N_7440);
and U10560 (N_10560,N_6646,N_6573);
or U10561 (N_10561,N_8702,N_9615);
and U10562 (N_10562,N_6462,N_7439);
and U10563 (N_10563,N_5436,N_8087);
xor U10564 (N_10564,N_6259,N_6109);
nand U10565 (N_10565,N_9973,N_7154);
or U10566 (N_10566,N_9636,N_7496);
and U10567 (N_10567,N_6051,N_7207);
xor U10568 (N_10568,N_5796,N_6296);
nand U10569 (N_10569,N_9033,N_8946);
nand U10570 (N_10570,N_8866,N_8620);
nand U10571 (N_10571,N_5315,N_7015);
or U10572 (N_10572,N_6156,N_9334);
and U10573 (N_10573,N_7748,N_7904);
and U10574 (N_10574,N_7563,N_5808);
xnor U10575 (N_10575,N_9363,N_6869);
and U10576 (N_10576,N_8696,N_9026);
nand U10577 (N_10577,N_5111,N_7530);
xnor U10578 (N_10578,N_8650,N_6721);
nor U10579 (N_10579,N_8038,N_8634);
or U10580 (N_10580,N_9935,N_9182);
or U10581 (N_10581,N_8685,N_7182);
or U10582 (N_10582,N_5287,N_5567);
nor U10583 (N_10583,N_5402,N_8670);
xnor U10584 (N_10584,N_9751,N_6703);
or U10585 (N_10585,N_8839,N_8953);
xor U10586 (N_10586,N_6412,N_6893);
nand U10587 (N_10587,N_9226,N_5836);
nand U10588 (N_10588,N_9296,N_9151);
xor U10589 (N_10589,N_6514,N_9573);
and U10590 (N_10590,N_6858,N_9598);
nor U10591 (N_10591,N_9619,N_9231);
and U10592 (N_10592,N_8071,N_6853);
xor U10593 (N_10593,N_9750,N_5595);
nand U10594 (N_10594,N_6194,N_7002);
xnor U10595 (N_10595,N_9785,N_7435);
and U10596 (N_10596,N_8077,N_9262);
and U10597 (N_10597,N_5509,N_5274);
xnor U10598 (N_10598,N_5304,N_8833);
nand U10599 (N_10599,N_5152,N_6936);
or U10600 (N_10600,N_6458,N_6397);
nor U10601 (N_10601,N_9175,N_7074);
or U10602 (N_10602,N_9055,N_6511);
xnor U10603 (N_10603,N_8078,N_5821);
xor U10604 (N_10604,N_8465,N_8018);
and U10605 (N_10605,N_6333,N_8404);
or U10606 (N_10606,N_8803,N_7324);
nand U10607 (N_10607,N_9837,N_5064);
xor U10608 (N_10608,N_9402,N_7168);
xnor U10609 (N_10609,N_7830,N_7577);
and U10610 (N_10610,N_6673,N_5159);
nor U10611 (N_10611,N_8207,N_7661);
nor U10612 (N_10612,N_6368,N_6475);
or U10613 (N_10613,N_9946,N_5316);
and U10614 (N_10614,N_8776,N_7716);
or U10615 (N_10615,N_7703,N_5459);
nor U10616 (N_10616,N_9512,N_7619);
xor U10617 (N_10617,N_8536,N_6782);
or U10618 (N_10618,N_8601,N_7035);
nand U10619 (N_10619,N_6901,N_8959);
or U10620 (N_10620,N_9109,N_7404);
nor U10621 (N_10621,N_8045,N_7812);
xor U10622 (N_10622,N_8626,N_5985);
nand U10623 (N_10623,N_8884,N_9612);
nand U10624 (N_10624,N_9834,N_9216);
nand U10625 (N_10625,N_5269,N_6079);
and U10626 (N_10626,N_6028,N_5279);
and U10627 (N_10627,N_5232,N_6434);
nor U10628 (N_10628,N_9847,N_7869);
and U10629 (N_10629,N_5016,N_9990);
nor U10630 (N_10630,N_8442,N_8579);
nor U10631 (N_10631,N_7580,N_8939);
nor U10632 (N_10632,N_9203,N_7921);
and U10633 (N_10633,N_7979,N_7738);
and U10634 (N_10634,N_5767,N_5033);
xor U10635 (N_10635,N_8716,N_9752);
and U10636 (N_10636,N_5738,N_5183);
nor U10637 (N_10637,N_7999,N_7845);
nand U10638 (N_10638,N_7122,N_5952);
nor U10639 (N_10639,N_6648,N_5707);
or U10640 (N_10640,N_6827,N_9725);
and U10641 (N_10641,N_8186,N_6186);
xnor U10642 (N_10642,N_9083,N_6128);
nor U10643 (N_10643,N_8399,N_7773);
xnor U10644 (N_10644,N_6743,N_5687);
or U10645 (N_10645,N_8561,N_5281);
xnor U10646 (N_10646,N_6224,N_7067);
nand U10647 (N_10647,N_7888,N_5961);
xnor U10648 (N_10648,N_7735,N_9617);
nand U10649 (N_10649,N_6365,N_7321);
or U10650 (N_10650,N_8141,N_5186);
nor U10651 (N_10651,N_9439,N_5550);
nand U10652 (N_10652,N_5608,N_5322);
or U10653 (N_10653,N_8846,N_8700);
nand U10654 (N_10654,N_8711,N_9225);
nor U10655 (N_10655,N_7268,N_7903);
xor U10656 (N_10656,N_7723,N_9219);
nor U10657 (N_10657,N_9381,N_9569);
and U10658 (N_10658,N_7937,N_6463);
nand U10659 (N_10659,N_7867,N_8006);
xnor U10660 (N_10660,N_9659,N_5493);
nor U10661 (N_10661,N_8499,N_5306);
nand U10662 (N_10662,N_6593,N_7049);
and U10663 (N_10663,N_9694,N_9009);
or U10664 (N_10664,N_7254,N_6042);
or U10665 (N_10665,N_6287,N_8847);
nand U10666 (N_10666,N_7070,N_8958);
xor U10667 (N_10667,N_6933,N_7222);
xor U10668 (N_10668,N_9274,N_5609);
nor U10669 (N_10669,N_9988,N_7334);
xor U10670 (N_10670,N_6847,N_8283);
and U10671 (N_10671,N_9124,N_9768);
xor U10672 (N_10672,N_5348,N_5968);
nand U10673 (N_10673,N_6826,N_8281);
or U10674 (N_10674,N_5902,N_7545);
xnor U10675 (N_10675,N_7398,N_7764);
xor U10676 (N_10676,N_9165,N_7489);
xor U10677 (N_10677,N_6975,N_7831);
or U10678 (N_10678,N_7906,N_7038);
and U10679 (N_10679,N_8628,N_9690);
and U10680 (N_10680,N_7227,N_5397);
or U10681 (N_10681,N_6226,N_9805);
and U10682 (N_10682,N_8403,N_6772);
nor U10683 (N_10683,N_6927,N_6436);
xnor U10684 (N_10684,N_8580,N_8566);
nor U10685 (N_10685,N_5241,N_8916);
xnor U10686 (N_10686,N_8837,N_6488);
or U10687 (N_10687,N_8770,N_8409);
xor U10688 (N_10688,N_5601,N_8600);
or U10689 (N_10689,N_6863,N_5243);
nand U10690 (N_10690,N_6061,N_5023);
xor U10691 (N_10691,N_6295,N_8546);
or U10692 (N_10692,N_8172,N_8883);
or U10693 (N_10693,N_8858,N_9892);
or U10694 (N_10694,N_6558,N_6330);
xor U10695 (N_10695,N_7276,N_9195);
xnor U10696 (N_10696,N_5310,N_7452);
xnor U10697 (N_10697,N_5309,N_9386);
and U10698 (N_10698,N_7177,N_7450);
or U10699 (N_10699,N_9496,N_8827);
or U10700 (N_10700,N_7419,N_9148);
nand U10701 (N_10701,N_6816,N_7917);
nor U10702 (N_10702,N_9609,N_5460);
and U10703 (N_10703,N_7434,N_7198);
nand U10704 (N_10704,N_9154,N_5648);
xnor U10705 (N_10705,N_7224,N_5445);
and U10706 (N_10706,N_5996,N_6031);
xnor U10707 (N_10707,N_8857,N_6686);
nor U10708 (N_10708,N_7309,N_8832);
nand U10709 (N_10709,N_7612,N_5781);
nor U10710 (N_10710,N_6062,N_7691);
xnor U10711 (N_10711,N_9861,N_9503);
nor U10712 (N_10712,N_9625,N_8849);
nand U10713 (N_10713,N_8615,N_9319);
nor U10714 (N_10714,N_9516,N_7200);
or U10715 (N_10715,N_6140,N_5711);
and U10716 (N_10716,N_8309,N_6536);
nand U10717 (N_10717,N_9106,N_8529);
and U10718 (N_10718,N_5105,N_9776);
nor U10719 (N_10719,N_8513,N_7980);
nand U10720 (N_10720,N_9613,N_8025);
or U10721 (N_10721,N_7555,N_8043);
and U10722 (N_10722,N_6123,N_8758);
or U10723 (N_10723,N_6137,N_7600);
and U10724 (N_10724,N_7893,N_7000);
and U10725 (N_10725,N_9844,N_5370);
or U10726 (N_10726,N_5551,N_7922);
nor U10727 (N_10727,N_8175,N_6615);
or U10728 (N_10728,N_5759,N_6101);
nor U10729 (N_10729,N_6489,N_8861);
or U10730 (N_10730,N_6261,N_7338);
or U10731 (N_10731,N_7850,N_9904);
nor U10732 (N_10732,N_5407,N_7658);
nand U10733 (N_10733,N_9732,N_7033);
xor U10734 (N_10734,N_6962,N_7860);
nor U10735 (N_10735,N_6391,N_5865);
or U10736 (N_10736,N_9542,N_8385);
nand U10737 (N_10737,N_8405,N_5987);
xnor U10738 (N_10738,N_8246,N_9256);
nor U10739 (N_10739,N_8559,N_7479);
and U10740 (N_10740,N_5570,N_9900);
or U10741 (N_10741,N_5983,N_6091);
xnor U10742 (N_10742,N_6367,N_5494);
nor U10743 (N_10743,N_6328,N_6684);
nand U10744 (N_10744,N_9654,N_7396);
nand U10745 (N_10745,N_7467,N_6579);
xnor U10746 (N_10746,N_7983,N_9545);
or U10747 (N_10747,N_7502,N_7441);
xnor U10748 (N_10748,N_9403,N_5314);
and U10749 (N_10749,N_6306,N_8166);
nand U10750 (N_10750,N_5425,N_8629);
xnor U10751 (N_10751,N_6073,N_7402);
nor U10752 (N_10752,N_7772,N_5472);
xnor U10753 (N_10753,N_8768,N_6131);
nor U10754 (N_10754,N_8932,N_5257);
or U10755 (N_10755,N_7152,N_5897);
nand U10756 (N_10756,N_5012,N_8658);
xor U10757 (N_10757,N_6124,N_7582);
nor U10758 (N_10758,N_6129,N_5969);
nand U10759 (N_10759,N_6977,N_6638);
or U10760 (N_10760,N_9640,N_7432);
or U10761 (N_10761,N_6471,N_5478);
nor U10762 (N_10762,N_5437,N_8046);
nor U10763 (N_10763,N_8604,N_6114);
nand U10764 (N_10764,N_5564,N_5216);
nand U10765 (N_10765,N_8085,N_9713);
xor U10766 (N_10766,N_7468,N_6341);
nand U10767 (N_10767,N_8033,N_7671);
nand U10768 (N_10768,N_7322,N_7976);
xnor U10769 (N_10769,N_8506,N_9963);
nand U10770 (N_10770,N_5832,N_6459);
and U10771 (N_10771,N_5915,N_9447);
or U10772 (N_10772,N_5677,N_7506);
xor U10773 (N_10773,N_7849,N_7120);
nor U10774 (N_10774,N_6289,N_9041);
nor U10775 (N_10775,N_5872,N_9075);
and U10776 (N_10776,N_7886,N_8168);
and U10777 (N_10777,N_7591,N_8080);
xnor U10778 (N_10778,N_6788,N_5706);
and U10779 (N_10779,N_8853,N_6814);
xor U10780 (N_10780,N_5169,N_9527);
or U10781 (N_10781,N_7607,N_7345);
and U10782 (N_10782,N_6487,N_7362);
xnor U10783 (N_10783,N_7028,N_6086);
and U10784 (N_10784,N_5668,N_5848);
nand U10785 (N_10785,N_8267,N_6055);
xor U10786 (N_10786,N_9378,N_6351);
nor U10787 (N_10787,N_8809,N_9777);
xor U10788 (N_10788,N_5071,N_6895);
or U10789 (N_10789,N_9064,N_8815);
or U10790 (N_10790,N_9081,N_5670);
or U10791 (N_10791,N_9241,N_5842);
nor U10792 (N_10792,N_9211,N_9832);
nor U10793 (N_10793,N_9122,N_7990);
or U10794 (N_10794,N_8094,N_7693);
or U10795 (N_10795,N_7367,N_9856);
xor U10796 (N_10796,N_8624,N_9819);
and U10797 (N_10797,N_7261,N_5518);
and U10798 (N_10798,N_6138,N_7594);
or U10799 (N_10799,N_5046,N_5312);
and U10800 (N_10800,N_9080,N_5783);
or U10801 (N_10801,N_8491,N_6568);
nor U10802 (N_10802,N_5135,N_5678);
xnor U10803 (N_10803,N_8140,N_5345);
nand U10804 (N_10804,N_6269,N_7081);
or U10805 (N_10805,N_5599,N_7725);
and U10806 (N_10806,N_8220,N_9865);
or U10807 (N_10807,N_7310,N_9252);
nor U10808 (N_10808,N_6406,N_6235);
nand U10809 (N_10809,N_7899,N_6740);
and U10810 (N_10810,N_5826,N_5002);
nand U10811 (N_10811,N_5266,N_5507);
and U10812 (N_10812,N_7621,N_5976);
or U10813 (N_10813,N_8276,N_8241);
nor U10814 (N_10814,N_9894,N_7509);
or U10815 (N_10815,N_7349,N_5031);
nor U10816 (N_10816,N_7660,N_9841);
or U10817 (N_10817,N_7071,N_8630);
nand U10818 (N_10818,N_9645,N_5712);
nor U10819 (N_10819,N_9814,N_9717);
xnor U10820 (N_10820,N_8050,N_8452);
nor U10821 (N_10821,N_6244,N_6089);
or U10822 (N_10822,N_5473,N_5680);
xor U10823 (N_10823,N_6126,N_6249);
nor U10824 (N_10824,N_9029,N_9050);
xor U10825 (N_10825,N_6440,N_6153);
and U10826 (N_10826,N_8799,N_8049);
nor U10827 (N_10827,N_6030,N_8814);
and U10828 (N_10828,N_8249,N_9021);
nand U10829 (N_10829,N_5941,N_8681);
xnor U10830 (N_10830,N_8517,N_7377);
nand U10831 (N_10831,N_8142,N_5674);
nor U10832 (N_10832,N_8428,N_9483);
nor U10833 (N_10833,N_8900,N_8010);
nor U10834 (N_10834,N_9551,N_7030);
and U10835 (N_10835,N_7974,N_9862);
nor U10836 (N_10836,N_5249,N_9541);
or U10837 (N_10837,N_8095,N_7760);
and U10838 (N_10838,N_7096,N_8012);
and U10839 (N_10839,N_7708,N_5561);
xor U10840 (N_10840,N_9689,N_7239);
or U10841 (N_10841,N_7588,N_5238);
and U10842 (N_10842,N_9010,N_8358);
xnor U10843 (N_10843,N_8229,N_6726);
nand U10844 (N_10844,N_5544,N_7587);
nand U10845 (N_10845,N_6172,N_8898);
xor U10846 (N_10846,N_6045,N_5193);
or U10847 (N_10847,N_5924,N_7777);
nor U10848 (N_10848,N_5999,N_6139);
xnor U10849 (N_10849,N_6907,N_7749);
nor U10850 (N_10850,N_5434,N_6955);
and U10851 (N_10851,N_5349,N_7495);
or U10852 (N_10852,N_9968,N_7111);
nor U10853 (N_10853,N_8295,N_8196);
xor U10854 (N_10854,N_8645,N_6564);
nor U10855 (N_10855,N_9235,N_6150);
nand U10856 (N_10856,N_9394,N_5927);
nand U10857 (N_10857,N_5956,N_5497);
nor U10858 (N_10858,N_6822,N_6539);
nor U10859 (N_10859,N_7164,N_8000);
and U10860 (N_10860,N_7385,N_8845);
or U10861 (N_10861,N_6656,N_9367);
nor U10862 (N_10862,N_6896,N_9934);
nor U10863 (N_10863,N_8835,N_7679);
xor U10864 (N_10864,N_8771,N_8583);
or U10865 (N_10865,N_9267,N_8346);
xnor U10866 (N_10866,N_9417,N_7172);
xor U10867 (N_10867,N_8015,N_8451);
nand U10868 (N_10868,N_7933,N_6538);
nor U10869 (N_10869,N_5391,N_9361);
and U10870 (N_10870,N_5859,N_6892);
xor U10871 (N_10871,N_9042,N_5395);
and U10872 (N_10872,N_6361,N_6932);
nand U10873 (N_10873,N_9947,N_7135);
nand U10874 (N_10874,N_9230,N_8602);
nand U10875 (N_10875,N_7631,N_7617);
nand U10876 (N_10876,N_8993,N_8391);
xor U10877 (N_10877,N_8213,N_5844);
or U10878 (N_10878,N_9698,N_6848);
xnor U10879 (N_10879,N_7491,N_9922);
xnor U10880 (N_10880,N_6056,N_9681);
and U10881 (N_10881,N_7378,N_7866);
and U10882 (N_10882,N_6362,N_9443);
nor U10883 (N_10883,N_5761,N_7971);
nor U10884 (N_10884,N_5150,N_8823);
nor U10885 (N_10885,N_6023,N_9399);
and U10886 (N_10886,N_8047,N_8587);
or U10887 (N_10887,N_6940,N_9325);
xnor U10888 (N_10888,N_6552,N_9407);
nand U10889 (N_10889,N_5164,N_9458);
and U10890 (N_10890,N_9952,N_6482);
or U10891 (N_10891,N_9053,N_9210);
or U10892 (N_10892,N_9614,N_8599);
nand U10893 (N_10893,N_5566,N_5631);
nor U10894 (N_10894,N_7752,N_7783);
and U10895 (N_10895,N_8864,N_5854);
nand U10896 (N_10896,N_5966,N_9809);
or U10897 (N_10897,N_7306,N_8359);
nor U10898 (N_10898,N_5606,N_9045);
and U10899 (N_10899,N_7681,N_8904);
and U10900 (N_10900,N_9015,N_9888);
or U10901 (N_10901,N_9800,N_5048);
xnor U10902 (N_10902,N_5426,N_7298);
and U10903 (N_10903,N_5722,N_9425);
xnor U10904 (N_10904,N_5408,N_5423);
nand U10905 (N_10905,N_5786,N_5526);
nor U10906 (N_10906,N_6943,N_9082);
nand U10907 (N_10907,N_9824,N_5251);
nand U10908 (N_10908,N_5339,N_6606);
xnor U10909 (N_10909,N_7884,N_8228);
and U10910 (N_10910,N_6047,N_9132);
nor U10911 (N_10911,N_6217,N_5136);
and U10912 (N_10912,N_9221,N_5180);
nor U10913 (N_10913,N_7142,N_7392);
xor U10914 (N_10914,N_9699,N_7469);
nor U10915 (N_10915,N_7678,N_9797);
nor U10916 (N_10916,N_6329,N_5659);
nand U10917 (N_10917,N_7882,N_9432);
or U10918 (N_10918,N_9576,N_7610);
nor U10919 (N_10919,N_9473,N_6390);
and U10920 (N_10920,N_9118,N_6749);
nand U10921 (N_10921,N_6326,N_6374);
xnor U10922 (N_10922,N_7470,N_7400);
or U10923 (N_10923,N_5639,N_8250);
nand U10924 (N_10924,N_5035,N_7417);
and U10925 (N_10925,N_8477,N_9971);
and U10926 (N_10926,N_9451,N_8989);
nand U10927 (N_10927,N_5041,N_5907);
nor U10928 (N_10928,N_7147,N_9320);
xor U10929 (N_10929,N_7215,N_7803);
nand U10930 (N_10930,N_6719,N_6155);
xnor U10931 (N_10931,N_5204,N_7444);
xnor U10932 (N_10932,N_8412,N_7043);
xnor U10933 (N_10933,N_5616,N_9927);
nor U10934 (N_10934,N_9882,N_7089);
nor U10935 (N_10935,N_5480,N_6416);
or U10936 (N_10936,N_7901,N_6067);
and U10937 (N_10937,N_6637,N_8271);
nand U10938 (N_10938,N_9587,N_8854);
xor U10939 (N_10939,N_8970,N_6937);
nor U10940 (N_10940,N_6384,N_6052);
xor U10941 (N_10941,N_7605,N_7258);
xor U10942 (N_10942,N_7062,N_9561);
and U10943 (N_10943,N_8726,N_7124);
or U10944 (N_10944,N_9682,N_9852);
xor U10945 (N_10945,N_7162,N_8810);
xor U10946 (N_10946,N_8683,N_7516);
nor U10947 (N_10947,N_7699,N_8336);
xnor U10948 (N_10948,N_8990,N_9146);
or U10949 (N_10949,N_7676,N_7836);
nand U10950 (N_10950,N_9504,N_6885);
and U10951 (N_10951,N_7232,N_9147);
nor U10952 (N_10952,N_8524,N_8417);
xor U10953 (N_10953,N_5645,N_9684);
nand U10954 (N_10954,N_6691,N_6813);
or U10955 (N_10955,N_9390,N_9727);
nor U10956 (N_10956,N_5415,N_7657);
or U10957 (N_10957,N_9499,N_5734);
nand U10958 (N_10958,N_8456,N_9955);
nor U10959 (N_10959,N_7963,N_9145);
xor U10960 (N_10960,N_6998,N_9701);
nor U10961 (N_10961,N_6058,N_7581);
and U10962 (N_10962,N_7755,N_7840);
nand U10963 (N_10963,N_9421,N_6439);
nor U10964 (N_10964,N_8692,N_9908);
nor U10965 (N_10965,N_5103,N_9823);
xor U10966 (N_10966,N_7026,N_9308);
and U10967 (N_10967,N_7533,N_7370);
xor U10968 (N_10968,N_6722,N_5361);
nand U10969 (N_10969,N_7663,N_7454);
and U10970 (N_10970,N_8818,N_5469);
or U10971 (N_10971,N_9558,N_9370);
nand U10972 (N_10972,N_7851,N_5481);
or U10973 (N_10973,N_7196,N_6902);
xnor U10974 (N_10974,N_6335,N_8048);
and U10975 (N_10975,N_7429,N_7412);
or U10976 (N_10976,N_5083,N_8288);
or U10977 (N_10977,N_6626,N_9002);
xnor U10978 (N_10978,N_9736,N_6281);
and U10979 (N_10979,N_6935,N_8133);
nor U10980 (N_10980,N_7235,N_6865);
xnor U10981 (N_10981,N_9298,N_5750);
xor U10982 (N_10982,N_7682,N_7230);
and U10983 (N_10983,N_6582,N_7729);
xor U10984 (N_10984,N_9116,N_7525);
or U10985 (N_10985,N_6325,N_6251);
and U10986 (N_10986,N_6553,N_8563);
and U10987 (N_10987,N_5752,N_5056);
or U10988 (N_10988,N_7982,N_8026);
xnor U10989 (N_10989,N_6760,N_9290);
xor U10990 (N_10990,N_8406,N_7471);
xor U10991 (N_10991,N_9919,N_6106);
xnor U10992 (N_10992,N_6921,N_6881);
nor U10993 (N_10993,N_6622,N_5299);
or U10994 (N_10994,N_9105,N_6038);
or U10995 (N_10995,N_5158,N_9095);
and U10996 (N_10996,N_5810,N_7058);
and U10997 (N_10997,N_6143,N_9309);
xor U10998 (N_10998,N_6324,N_7474);
or U10999 (N_10999,N_9442,N_8632);
xnor U11000 (N_11000,N_5076,N_8680);
or U11001 (N_11001,N_5694,N_8684);
nor U11002 (N_11002,N_5225,N_5381);
or U11003 (N_11003,N_6494,N_6478);
and U11004 (N_11004,N_5679,N_6070);
nor U11005 (N_11005,N_5517,N_9463);
xor U11006 (N_11006,N_6754,N_8792);
xor U11007 (N_11007,N_8294,N_5822);
xnor U11008 (N_11008,N_5433,N_5669);
or U11009 (N_11009,N_7034,N_9233);
or U11010 (N_11010,N_5070,N_5651);
nand U11011 (N_11011,N_6423,N_7105);
nor U11012 (N_11012,N_8100,N_8921);
nand U11013 (N_11013,N_5977,N_7391);
xnor U11014 (N_11014,N_6177,N_8659);
nor U11015 (N_11015,N_7337,N_5380);
or U11016 (N_11016,N_7245,N_5211);
nand U11017 (N_11017,N_9734,N_9380);
or U11018 (N_11018,N_8877,N_8266);
and U11019 (N_11019,N_8844,N_5133);
or U11020 (N_11020,N_6612,N_7226);
or U11021 (N_11021,N_5082,N_7542);
xor U11022 (N_11022,N_7633,N_8366);
and U11023 (N_11023,N_8902,N_7480);
or U11024 (N_11024,N_6620,N_6780);
nand U11025 (N_11025,N_9624,N_8383);
and U11026 (N_11026,N_8703,N_9046);
and U11027 (N_11027,N_9067,N_7704);
or U11028 (N_11028,N_9312,N_9588);
nand U11029 (N_11029,N_8222,N_5100);
or U11030 (N_11030,N_5664,N_7642);
or U11031 (N_11031,N_7734,N_5263);
and U11032 (N_11032,N_5122,N_9649);
xnor U11033 (N_11033,N_9285,N_7797);
nand U11034 (N_11034,N_9434,N_5148);
nand U11035 (N_11035,N_5130,N_8999);
nand U11036 (N_11036,N_7877,N_7741);
or U11037 (N_11037,N_9945,N_6088);
xor U11038 (N_11038,N_8231,N_9604);
or U11039 (N_11039,N_8699,N_6807);
nor U11040 (N_11040,N_8199,N_8978);
or U11041 (N_11041,N_8326,N_5301);
nor U11042 (N_11042,N_9199,N_7102);
or U11043 (N_11043,N_7806,N_6981);
nor U11044 (N_11044,N_8800,N_7513);
and U11045 (N_11045,N_6339,N_7751);
xor U11046 (N_11046,N_5019,N_7256);
nor U11047 (N_11047,N_8908,N_6256);
xnor U11048 (N_11048,N_5420,N_8526);
and U11049 (N_11049,N_8367,N_8976);
nor U11050 (N_11050,N_6820,N_8195);
and U11051 (N_11051,N_9982,N_9005);
nor U11052 (N_11052,N_9018,N_7895);
xnor U11053 (N_11053,N_9127,N_8242);
nand U11054 (N_11054,N_9924,N_7839);
and U11055 (N_11055,N_9748,N_9656);
xor U11056 (N_11056,N_7109,N_8798);
nor U11057 (N_11057,N_5475,N_5066);
or U11058 (N_11058,N_9753,N_9877);
nor U11059 (N_11059,N_5015,N_7578);
xnor U11060 (N_11060,N_8066,N_5948);
or U11061 (N_11061,N_5227,N_6702);
or U11062 (N_11062,N_5114,N_5265);
nor U11063 (N_11063,N_6476,N_8598);
or U11064 (N_11064,N_5980,N_8490);
or U11065 (N_11065,N_8596,N_9258);
nor U11066 (N_11066,N_6248,N_6202);
or U11067 (N_11067,N_9950,N_9559);
nor U11068 (N_11068,N_7960,N_7900);
nor U11069 (N_11069,N_6725,N_6311);
and U11070 (N_11070,N_5044,N_7972);
nor U11071 (N_11071,N_7353,N_8790);
nor U11072 (N_11072,N_8163,N_7387);
nor U11073 (N_11073,N_8951,N_9464);
and U11074 (N_11074,N_7046,N_5235);
xnor U11075 (N_11075,N_7837,N_9536);
nor U11076 (N_11076,N_8189,N_9626);
xor U11077 (N_11077,N_8239,N_5782);
xor U11078 (N_11078,N_9910,N_5719);
and U11079 (N_11079,N_9891,N_7862);
and U11080 (N_11080,N_5280,N_7569);
and U11081 (N_11081,N_5773,N_5619);
and U11082 (N_11082,N_6005,N_8722);
nand U11083 (N_11083,N_7136,N_7786);
and U11084 (N_11084,N_8067,N_8481);
nor U11085 (N_11085,N_8101,N_9781);
or U11086 (N_11086,N_9628,N_8362);
nor U11087 (N_11087,N_9263,N_7622);
and U11088 (N_11088,N_6750,N_8942);
nor U11089 (N_11089,N_8429,N_8285);
or U11090 (N_11090,N_8413,N_9408);
xor U11091 (N_11091,N_9567,N_7332);
nand U11092 (N_11092,N_9093,N_5248);
xor U11093 (N_11093,N_7319,N_5656);
nand U11094 (N_11094,N_7964,N_8268);
nor U11095 (N_11095,N_5633,N_5366);
or U11096 (N_11096,N_7568,N_5882);
nor U11097 (N_11097,N_7539,N_8929);
nor U11098 (N_11098,N_9687,N_8638);
nor U11099 (N_11099,N_7634,N_5909);
or U11100 (N_11100,N_6835,N_8235);
nand U11101 (N_11101,N_5403,N_6836);
or U11102 (N_11102,N_8431,N_7376);
nand U11103 (N_11103,N_8190,N_7242);
nand U11104 (N_11104,N_6422,N_5862);
nor U11105 (N_11105,N_8622,N_6554);
or U11106 (N_11106,N_5805,N_5112);
nand U11107 (N_11107,N_7292,N_7061);
xor U11108 (N_11108,N_8819,N_8723);
or U11109 (N_11109,N_7914,N_7282);
and U11110 (N_11110,N_7050,N_6831);
xnor U11111 (N_11111,N_7213,N_7174);
and U11112 (N_11112,N_9943,N_5945);
nand U11113 (N_11113,N_9765,N_5658);
nand U11114 (N_11114,N_6957,N_5905);
nor U11115 (N_11115,N_5091,N_9071);
and U11116 (N_11116,N_8151,N_6164);
xor U11117 (N_11117,N_9119,N_9347);
or U11118 (N_11118,N_5374,N_9967);
or U11119 (N_11119,N_8298,N_5212);
nand U11120 (N_11120,N_7274,N_6590);
nor U11121 (N_11121,N_8280,N_5932);
or U11122 (N_11122,N_7270,N_7553);
or U11123 (N_11123,N_7920,N_5860);
or U11124 (N_11124,N_6087,N_9388);
xor U11125 (N_11125,N_9196,N_9715);
nand U11126 (N_11126,N_8257,N_8741);
xor U11127 (N_11127,N_5072,N_9169);
xor U11128 (N_11128,N_9494,N_8433);
nand U11129 (N_11129,N_7225,N_8278);
xor U11130 (N_11130,N_8411,N_9446);
or U11131 (N_11131,N_5834,N_7865);
nand U11132 (N_11132,N_7700,N_8922);
xor U11133 (N_11133,N_9535,N_5096);
and U11134 (N_11134,N_5462,N_9173);
nor U11135 (N_11135,N_7991,N_7131);
and U11136 (N_11136,N_7776,N_7488);
and U11137 (N_11137,N_9716,N_9089);
or U11138 (N_11138,N_6627,N_6733);
nor U11139 (N_11139,N_9317,N_9249);
nor U11140 (N_11140,N_6513,N_6574);
xnor U11141 (N_11141,N_5205,N_6268);
nor U11142 (N_11142,N_8570,N_8487);
or U11143 (N_11143,N_9784,N_8577);
xor U11144 (N_11144,N_8694,N_5334);
and U11145 (N_11145,N_9764,N_6302);
nor U11146 (N_11146,N_6093,N_9346);
and U11147 (N_11147,N_8497,N_8495);
nor U11148 (N_11148,N_9671,N_6196);
nor U11149 (N_11149,N_8784,N_6837);
and U11150 (N_11150,N_5222,N_5512);
or U11151 (N_11151,N_7472,N_7958);
and U11152 (N_11152,N_6909,N_7278);
nand U11153 (N_11153,N_5733,N_6611);
xor U11154 (N_11154,N_7892,N_5154);
and U11155 (N_11155,N_5884,N_8155);
or U11156 (N_11156,N_6900,N_5811);
nand U11157 (N_11157,N_8147,N_7894);
xor U11158 (N_11158,N_6232,N_9923);
or U11159 (N_11159,N_6210,N_8042);
nor U11160 (N_11160,N_8568,N_8627);
or U11161 (N_11161,N_6158,N_6262);
nor U11162 (N_11162,N_6216,N_5467);
and U11163 (N_11163,N_7890,N_5236);
nor U11164 (N_11164,N_6272,N_5904);
or U11165 (N_11165,N_9423,N_9062);
or U11166 (N_11166,N_6118,N_8876);
or U11167 (N_11167,N_9184,N_7953);
and U11168 (N_11168,N_8555,N_7193);
nor U11169 (N_11169,N_6501,N_6219);
nor U11170 (N_11170,N_5123,N_7586);
and U11171 (N_11171,N_5253,N_9125);
nor U11172 (N_11172,N_7668,N_8955);
nor U11173 (N_11173,N_9730,N_9695);
nand U11174 (N_11174,N_8612,N_8715);
and U11175 (N_11175,N_5689,N_7476);
nor U11176 (N_11176,N_5513,N_9193);
nand U11177 (N_11177,N_5026,N_7598);
nor U11178 (N_11178,N_9639,N_6393);
or U11179 (N_11179,N_8745,N_9461);
nand U11180 (N_11180,N_7408,N_7326);
and U11181 (N_11181,N_9686,N_5807);
or U11182 (N_11182,N_5181,N_9014);
nor U11183 (N_11183,N_7220,N_7720);
nand U11184 (N_11184,N_6108,N_6672);
xnor U11185 (N_11185,N_6120,N_9035);
nand U11186 (N_11186,N_5084,N_6371);
nand U11187 (N_11187,N_6657,N_8084);
xor U11188 (N_11188,N_8530,N_8247);
and U11189 (N_11189,N_6173,N_5254);
and U11190 (N_11190,N_7121,N_8804);
or U11191 (N_11191,N_8105,N_7795);
and U11192 (N_11192,N_8427,N_9339);
or U11193 (N_11193,N_7139,N_9415);
nand U11194 (N_11194,N_5673,N_5802);
xnor U11195 (N_11195,N_7259,N_9518);
nor U11196 (N_11196,N_5833,N_5383);
or U11197 (N_11197,N_7548,N_7294);
nand U11198 (N_11198,N_6145,N_6097);
xor U11199 (N_11199,N_8605,N_5325);
or U11200 (N_11200,N_8122,N_8081);
nor U11201 (N_11201,N_5830,N_7770);
and U11202 (N_11202,N_7173,N_9720);
or U11203 (N_11203,N_6915,N_9709);
or U11204 (N_11204,N_5229,N_9264);
and U11205 (N_11205,N_6965,N_8652);
and U11206 (N_11206,N_8208,N_5034);
nor U11207 (N_11207,N_8130,N_5191);
nor U11208 (N_11208,N_7532,N_8343);
and U11209 (N_11209,N_5779,N_8980);
and U11210 (N_11210,N_9331,N_8755);
nor U11211 (N_11211,N_7846,N_9827);
xor U11212 (N_11212,N_8351,N_9456);
or U11213 (N_11213,N_5365,N_5047);
and U11214 (N_11214,N_7093,N_9300);
and U11215 (N_11215,N_9474,N_8576);
xnor U11216 (N_11216,N_6182,N_6891);
nand U11217 (N_11217,N_5853,N_5398);
xnor U11218 (N_11218,N_6602,N_6889);
or U11219 (N_11219,N_8508,N_7531);
or U11220 (N_11220,N_8075,N_6298);
nor U11221 (N_11221,N_9866,N_6898);
xor U11222 (N_11222,N_6206,N_7792);
and U11223 (N_11223,N_5735,N_8498);
nor U11224 (N_11224,N_7247,N_5957);
nand U11225 (N_11225,N_8079,N_7561);
xnor U11226 (N_11226,N_6122,N_5974);
and U11227 (N_11227,N_8672,N_5618);
or U11228 (N_11228,N_6359,N_6356);
xor U11229 (N_11229,N_6253,N_9543);
xor U11230 (N_11230,N_6083,N_6457);
nand U11231 (N_11231,N_8518,N_7203);
xor U11232 (N_11232,N_6148,N_7181);
nor U11233 (N_11233,N_7014,N_6165);
xnor U11234 (N_11234,N_7085,N_5264);
and U11235 (N_11235,N_9076,N_9705);
and U11236 (N_11236,N_6461,N_7540);
nor U11237 (N_11237,N_8191,N_6288);
nor U11238 (N_11238,N_6992,N_8074);
xnor U11239 (N_11239,N_7608,N_9060);
nand U11240 (N_11240,N_5127,N_9265);
nor U11241 (N_11241,N_8279,N_9247);
or U11242 (N_11242,N_6569,N_5483);
nor U11243 (N_11243,N_5534,N_5982);
or U11244 (N_11244,N_6337,N_7649);
nand U11245 (N_11245,N_7171,N_6398);
nand U11246 (N_11246,N_9633,N_7202);
and U11247 (N_11247,N_8578,N_7623);
or U11248 (N_11248,N_8797,N_5572);
and U11249 (N_11249,N_9728,N_8948);
nand U11250 (N_11250,N_6793,N_8852);
nor U11251 (N_11251,N_8369,N_5376);
or U11252 (N_11252,N_5055,N_7870);
xnor U11253 (N_11253,N_5104,N_8510);
or U11254 (N_11254,N_9311,N_5063);
or U11255 (N_11255,N_9744,N_6433);
xnor U11256 (N_11256,N_5275,N_7219);
nor U11257 (N_11257,N_5118,N_7799);
and U11258 (N_11258,N_8834,N_5501);
xnor U11259 (N_11259,N_7132,N_6969);
xor U11260 (N_11260,N_7052,N_6004);
nand U11261 (N_11261,N_9351,N_8353);
or U11262 (N_11262,N_7437,N_5208);
xor U11263 (N_11263,N_9244,N_5581);
xor U11264 (N_11264,N_9085,N_5997);
xor U11265 (N_11265,N_7044,N_8489);
and U11266 (N_11266,N_9826,N_8512);
xor U11267 (N_11267,N_7427,N_8565);
or U11268 (N_11268,N_9895,N_5379);
nand U11269 (N_11269,N_6313,N_9655);
nand U11270 (N_11270,N_8554,N_8717);
xnor U11271 (N_11271,N_7277,N_9679);
and U11272 (N_11272,N_6773,N_7039);
or U11273 (N_11273,N_7386,N_5014);
or U11274 (N_11274,N_6353,N_5892);
and U11275 (N_11275,N_9501,N_6198);
xor U11276 (N_11276,N_6039,N_6191);
or U11277 (N_11277,N_5891,N_7004);
nand U11278 (N_11278,N_5479,N_7616);
xnor U11279 (N_11279,N_8082,N_9313);
nor U11280 (N_11280,N_9092,N_8919);
and U11281 (N_11281,N_7710,N_6669);
or U11282 (N_11282,N_6949,N_6993);
or U11283 (N_11283,N_9697,N_8426);
or U11284 (N_11284,N_7106,N_8035);
or U11285 (N_11285,N_7522,N_5875);
nor U11286 (N_11286,N_8317,N_7144);
nand U11287 (N_11287,N_7130,N_5946);
xnor U11288 (N_11288,N_5327,N_8523);
nor U11289 (N_11289,N_6861,N_8255);
and U11290 (N_11290,N_8254,N_6549);
or U11291 (N_11291,N_6415,N_7064);
and U11292 (N_11292,N_9020,N_9885);
or U11293 (N_11293,N_5285,N_7595);
nand U11294 (N_11294,N_9364,N_6418);
or U11295 (N_11295,N_7880,N_8926);
xnor U11296 (N_11296,N_8962,N_5728);
or U11297 (N_11297,N_6204,N_9796);
and U11298 (N_11298,N_9326,N_5282);
xor U11299 (N_11299,N_5448,N_7068);
nor U11300 (N_11300,N_6608,N_9365);
and U11301 (N_11301,N_8633,N_5009);
nand U11302 (N_11302,N_7233,N_9926);
xor U11303 (N_11303,N_9066,N_5008);
nor U11304 (N_11304,N_5864,N_9449);
nand U11305 (N_11305,N_6446,N_8930);
or U11306 (N_11306,N_8414,N_6600);
xor U11307 (N_11307,N_9218,N_8185);
nand U11308 (N_11308,N_6708,N_9571);
nor U11309 (N_11309,N_5329,N_6789);
and U11310 (N_11310,N_7790,N_7051);
and U11311 (N_11311,N_6763,N_6616);
or U11312 (N_11312,N_5335,N_8646);
nor U11313 (N_11313,N_7017,N_9925);
nand U11314 (N_11314,N_6801,N_5138);
xor U11315 (N_11315,N_6942,N_5636);
xnor U11316 (N_11316,N_8069,N_8016);
or U11317 (N_11317,N_7675,N_7572);
nor U11318 (N_11318,N_9637,N_6447);
nand U11319 (N_11319,N_6934,N_7291);
nor U11320 (N_11320,N_8480,N_5749);
and U11321 (N_11321,N_9052,N_6922);
nor U11322 (N_11322,N_6460,N_8824);
or U11323 (N_11323,N_8871,N_5373);
or U11324 (N_11324,N_9937,N_7881);
nand U11325 (N_11325,N_9646,N_8215);
xnor U11326 (N_11326,N_5233,N_5078);
and U11327 (N_11327,N_7951,N_5965);
nor U11328 (N_11328,N_8102,N_7101);
xnor U11329 (N_11329,N_7453,N_6385);
nor U11330 (N_11330,N_6066,N_5081);
xnor U11331 (N_11331,N_7360,N_8319);
nand U11332 (N_11332,N_9371,N_9688);
and U11333 (N_11333,N_7218,N_5625);
xor U11334 (N_11334,N_7234,N_8324);
and U11335 (N_11335,N_5237,N_5960);
nor U11336 (N_11336,N_8418,N_7988);
or U11337 (N_11337,N_8030,N_8146);
nor U11338 (N_11338,N_5421,N_5929);
and U11339 (N_11339,N_9931,N_9288);
or U11340 (N_11340,N_8786,N_6950);
xnor U11341 (N_11341,N_9998,N_5815);
nor U11342 (N_11342,N_5396,N_5145);
and U11343 (N_11343,N_9859,N_7696);
nand U11344 (N_11344,N_6964,N_9150);
nor U11345 (N_11345,N_8917,N_5568);
or U11346 (N_11346,N_9185,N_7717);
nor U11347 (N_11347,N_6803,N_9766);
xnor U11348 (N_11348,N_8956,N_6480);
xor U11349 (N_11349,N_9302,N_7965);
nor U11350 (N_11350,N_6728,N_8934);
nand U11351 (N_11351,N_8408,N_7992);
and U11352 (N_11352,N_7743,N_5387);
or U11353 (N_11353,N_5583,N_8410);
or U11354 (N_11354,N_9840,N_7891);
nand U11355 (N_11355,N_9522,N_8262);
or U11356 (N_11356,N_5959,N_5427);
nand U11357 (N_11357,N_6610,N_7304);
or U11358 (N_11358,N_6134,N_5556);
nand U11359 (N_11359,N_8963,N_5743);
and U11360 (N_11360,N_5911,N_6107);
and U11361 (N_11361,N_6095,N_8112);
xnor U11362 (N_11362,N_6451,N_9762);
nand U11363 (N_11363,N_9524,N_9321);
xnor U11364 (N_11364,N_7855,N_6809);
nor U11365 (N_11365,N_8742,N_7762);
or U11366 (N_11366,N_6791,N_8667);
or U11367 (N_11367,N_9810,N_6649);
nor U11368 (N_11368,N_8306,N_6897);
xnor U11369 (N_11369,N_7296,N_8264);
xnor U11370 (N_11370,N_9393,N_5007);
and U11371 (N_11371,N_6002,N_5296);
and U11372 (N_11372,N_9887,N_5937);
or U11373 (N_11373,N_5894,N_8881);
and U11374 (N_11374,N_5059,N_8721);
nor U11375 (N_11375,N_7012,N_7929);
or U11376 (N_11376,N_9470,N_6874);
nand U11377 (N_11377,N_5360,N_6127);
nand U11378 (N_11378,N_7802,N_6430);
nand U11379 (N_11379,N_9246,N_6730);
xnor U11380 (N_11380,N_9719,N_9537);
or U11381 (N_11381,N_6438,N_8816);
or U11382 (N_11382,N_7448,N_8041);
xor U11383 (N_11383,N_8380,N_5753);
or U11384 (N_11384,N_8928,N_9011);
and U11385 (N_11385,N_9724,N_9157);
and U11386 (N_11386,N_5794,N_8933);
or U11387 (N_11387,N_8549,N_5394);
nor U11388 (N_11388,N_7807,N_9552);
or U11389 (N_11389,N_9916,N_7571);
and U11390 (N_11390,N_6980,N_8028);
xor U11391 (N_11391,N_5571,N_5234);
nor U11392 (N_11392,N_5847,N_5721);
or U11393 (N_11393,N_8544,N_8675);
nor U11394 (N_11394,N_5527,N_6832);
xor U11395 (N_11395,N_7269,N_7511);
or U11396 (N_11396,N_6565,N_6982);
or U11397 (N_11397,N_7163,N_9629);
xor U11398 (N_11398,N_5109,N_7559);
xor U11399 (N_11399,N_7639,N_7520);
or U11400 (N_11400,N_6678,N_6410);
or U11401 (N_11401,N_7918,N_7711);
or U11402 (N_11402,N_5705,N_5818);
nand U11403 (N_11403,N_6162,N_9077);
nor U11404 (N_11404,N_8772,N_6017);
nand U11405 (N_11405,N_5006,N_9209);
and U11406 (N_11406,N_5495,N_7628);
or U11407 (N_11407,N_8277,N_7733);
and U11408 (N_11408,N_9280,N_6136);
nor U11409 (N_11409,N_7366,N_5432);
or U11410 (N_11410,N_8936,N_9579);
nand U11411 (N_11411,N_5172,N_6444);
or U11412 (N_11412,N_9574,N_8987);
xor U11413 (N_11413,N_9520,N_5099);
nor U11414 (N_11414,N_8850,N_5414);
nor U11415 (N_11415,N_6414,N_7638);
or U11416 (N_11416,N_6399,N_9746);
and U11417 (N_11417,N_9683,N_9782);
and U11418 (N_11418,N_7924,N_6201);
or U11419 (N_11419,N_7841,N_7365);
nand U11420 (N_11420,N_6027,N_9490);
nor U11421 (N_11421,N_8778,N_9702);
nor U11422 (N_11422,N_5940,N_8807);
and U11423 (N_11423,N_9607,N_7939);
or U11424 (N_11424,N_7498,N_9703);
nand U11425 (N_11425,N_6376,N_6714);
nor U11426 (N_11426,N_7492,N_7447);
or U11427 (N_11427,N_9207,N_5731);
and U11428 (N_11428,N_6802,N_9584);
and U11429 (N_11429,N_6521,N_8575);
nand U11430 (N_11430,N_7092,N_7497);
xnor U11431 (N_11431,N_9238,N_9332);
nor U11432 (N_11432,N_8248,N_8805);
xnor U11433 (N_11433,N_7973,N_8688);
xor U11434 (N_11434,N_7946,N_8641);
xnor U11435 (N_11435,N_5326,N_7962);
and U11436 (N_11436,N_9360,N_6491);
xor U11437 (N_11437,N_7534,N_9825);
nand U11438 (N_11438,N_9153,N_8907);
or U11439 (N_11439,N_8447,N_7420);
nand U11440 (N_11440,N_8316,N_6477);
nand U11441 (N_11441,N_6621,N_5490);
nand U11442 (N_11442,N_6787,N_6187);
nand U11443 (N_11443,N_5852,N_5710);
nor U11444 (N_11444,N_6072,N_5177);
nand U11445 (N_11445,N_7246,N_6976);
or U11446 (N_11446,N_8204,N_8938);
and U11447 (N_11447,N_6534,N_7107);
nor U11448 (N_11448,N_8719,N_9813);
or U11449 (N_11449,N_7665,N_9599);
or U11450 (N_11450,N_8330,N_9335);
nand U11451 (N_11451,N_7543,N_7827);
nor U11452 (N_11452,N_8870,N_9564);
or U11453 (N_11453,N_5119,N_7771);
or U11454 (N_11454,N_7908,N_5080);
xnor U11455 (N_11455,N_9997,N_6225);
nand U11456 (N_11456,N_8454,N_7237);
and U11457 (N_11457,N_5372,N_6560);
or U11458 (N_11458,N_9600,N_8311);
and U11459 (N_11459,N_5692,N_8542);
nand U11460 (N_11460,N_5881,N_6859);
nor U11461 (N_11461,N_9743,N_7652);
nor U11462 (N_11462,N_5992,N_9928);
xor U11463 (N_11463,N_7593,N_8764);
nand U11464 (N_11464,N_5293,N_7606);
or U11465 (N_11465,N_7060,N_5174);
nand U11466 (N_11466,N_6502,N_5273);
xor U11467 (N_11467,N_8340,N_7381);
nand U11468 (N_11468,N_9289,N_5555);
and U11469 (N_11469,N_8401,N_6320);
xor U11470 (N_11470,N_6025,N_9152);
nand U11471 (N_11471,N_7249,N_7007);
nand U11472 (N_11472,N_8752,N_7297);
xor U11473 (N_11473,N_9420,N_5845);
and U11474 (N_11474,N_5377,N_6082);
xor U11475 (N_11475,N_5450,N_5588);
and U11476 (N_11476,N_6011,N_9441);
xor U11477 (N_11477,N_8793,N_9557);
or U11478 (N_11478,N_9187,N_5737);
xnor U11479 (N_11479,N_7303,N_5654);
nand U11480 (N_11480,N_6394,N_9995);
nor U11481 (N_11481,N_7333,N_6810);
and U11482 (N_11482,N_7707,N_7714);
or U11483 (N_11483,N_8106,N_8439);
nand U11484 (N_11484,N_6144,N_5755);
nand U11485 (N_11485,N_6229,N_8437);
nor U11486 (N_11486,N_6338,N_7414);
nand U11487 (N_11487,N_6643,N_6018);
nand U11488 (N_11488,N_5215,N_8088);
or U11489 (N_11489,N_9337,N_5030);
and U11490 (N_11490,N_8338,N_5751);
and U11491 (N_11491,N_7364,N_6207);
or U11492 (N_11492,N_5829,N_6762);
or U11493 (N_11493,N_5772,N_5307);
nor U11494 (N_11494,N_8872,N_5681);
and U11495 (N_11495,N_8014,N_9465);
and U11496 (N_11496,N_8585,N_9027);
and U11497 (N_11497,N_5569,N_6318);
nand U11498 (N_11498,N_6948,N_6843);
nand U11499 (N_11499,N_8379,N_9511);
nand U11500 (N_11500,N_7327,N_7187);
xor U11501 (N_11501,N_5931,N_7073);
or U11502 (N_11502,N_6020,N_9427);
xnor U11503 (N_11503,N_8416,N_9142);
or U11504 (N_11504,N_9507,N_7709);
or U11505 (N_11505,N_8647,N_7801);
and U11506 (N_11506,N_6050,N_7329);
nor U11507 (N_11507,N_9070,N_8619);
xor U11508 (N_11508,N_9202,N_8669);
nor U11509 (N_11509,N_5161,N_6383);
or U11510 (N_11510,N_5828,N_6021);
and U11511 (N_11511,N_5565,N_7523);
nor U11512 (N_11512,N_7759,N_8300);
xnor U11513 (N_11513,N_5471,N_5532);
or U11514 (N_11514,N_9848,N_8720);
or U11515 (N_11515,N_7475,N_8240);
nor U11516 (N_11516,N_7354,N_8867);
xnor U11517 (N_11517,N_6382,N_9126);
nand U11518 (N_11518,N_5871,N_7864);
nor U11519 (N_11519,N_5748,N_8341);
or U11520 (N_11520,N_6715,N_5449);
or U11521 (N_11521,N_8952,N_5763);
nor U11522 (N_11522,N_7956,N_5825);
and U11523 (N_11523,N_9471,N_5918);
nand U11524 (N_11524,N_6613,N_6854);
and U11525 (N_11525,N_7775,N_6307);
xnor U11526 (N_11526,N_7538,N_6756);
nand U11527 (N_11527,N_6358,N_8708);
or U11528 (N_11528,N_6576,N_7104);
xnor U11529 (N_11529,N_7212,N_8838);
nor U11530 (N_11530,N_5182,N_6537);
nand U11531 (N_11531,N_7217,N_7063);
or U11532 (N_11532,N_9000,N_8261);
nor U11533 (N_11533,N_8307,N_7724);
nand U11534 (N_11534,N_6275,N_9097);
or U11535 (N_11535,N_5858,N_7086);
and U11536 (N_11536,N_6426,N_8640);
nand U11537 (N_11537,N_9131,N_5147);
xnor U11538 (N_11538,N_9357,N_6592);
xnor U11539 (N_11539,N_5219,N_5560);
nor U11540 (N_11540,N_8301,N_9426);
nor U11541 (N_11541,N_8750,N_9383);
and U11542 (N_11542,N_7006,N_7769);
nor U11543 (N_11543,N_8430,N_6044);
nand U11544 (N_11544,N_9345,N_6496);
nand U11545 (N_11545,N_6033,N_6652);
and U11546 (N_11546,N_9291,N_6880);
nand U11547 (N_11547,N_5284,N_5226);
and U11548 (N_11548,N_5196,N_8292);
or U11549 (N_11549,N_8450,N_9455);
nand U11550 (N_11550,N_7342,N_7602);
xnor U11551 (N_11551,N_7925,N_5389);
or U11552 (N_11552,N_7236,N_8760);
or U11553 (N_11553,N_8713,N_9101);
or U11554 (N_11554,N_5413,N_5903);
and U11555 (N_11555,N_8590,N_5098);
xnor U11556 (N_11556,N_9063,N_9957);
nor U11557 (N_11557,N_7687,N_5198);
and U11558 (N_11558,N_6633,N_5255);
and U11559 (N_11559,N_8981,N_9304);
and U11560 (N_11560,N_7409,N_5883);
or U11561 (N_11561,N_5637,N_9566);
or U11562 (N_11562,N_5095,N_9530);
xor U11563 (N_11563,N_5559,N_7813);
and U11564 (N_11564,N_6154,N_5073);
nand U11565 (N_11565,N_6276,N_9722);
and U11566 (N_11566,N_9257,N_9889);
xnor U11567 (N_11567,N_8743,N_9243);
xor U11568 (N_11568,N_8443,N_7823);
or U11569 (N_11569,N_7853,N_8328);
nor U11570 (N_11570,N_9466,N_7727);
xnor U11571 (N_11571,N_6310,N_5774);
and U11572 (N_11572,N_8073,N_8251);
nor U11573 (N_11573,N_7719,N_8206);
or U11574 (N_11574,N_6342,N_8007);
nand U11575 (N_11575,N_9519,N_6195);
nor U11576 (N_11576,N_8333,N_5746);
nor U11577 (N_11577,N_9008,N_6282);
or U11578 (N_11578,N_8469,N_9807);
xor U11579 (N_11579,N_6442,N_8830);
xor U11580 (N_11580,N_8855,N_9548);
nand U11581 (N_11581,N_8516,N_8055);
nand U11582 (N_11582,N_9758,N_5634);
nor U11583 (N_11583,N_9239,N_6695);
nand U11584 (N_11584,N_7395,N_6517);
xnor U11585 (N_11585,N_8767,N_8643);
and U11586 (N_11586,N_7919,N_8032);
and U11587 (N_11587,N_6828,N_6584);
xnor U11588 (N_11588,N_7620,N_6133);
xor U11589 (N_11589,N_7318,N_7287);
nor U11590 (N_11590,N_8148,N_6240);
nor U11591 (N_11591,N_5228,N_6696);
xor U11592 (N_11592,N_5324,N_5986);
nand U11593 (N_11593,N_5242,N_9284);
and U11594 (N_11594,N_6589,N_5856);
nand U11595 (N_11595,N_6636,N_9747);
or U11596 (N_11596,N_7863,N_7031);
nand U11597 (N_11597,N_5245,N_9763);
xnor U11598 (N_11598,N_7314,N_7143);
or U11599 (N_11599,N_8920,N_7985);
nand U11600 (N_11600,N_6223,N_7556);
nand U11601 (N_11601,N_6676,N_7127);
and U11602 (N_11602,N_8731,N_9635);
xnor U11603 (N_11603,N_8123,N_8654);
and U11604 (N_11604,N_9525,N_9550);
nand U11605 (N_11605,N_8862,N_6386);
nand U11606 (N_11606,N_8360,N_6524);
or U11607 (N_11607,N_6840,N_5088);
nand U11608 (N_11608,N_5958,N_7008);
xnor U11609 (N_11609,N_6057,N_5575);
nand U11610 (N_11610,N_6867,N_9462);
nor U11611 (N_11611,N_8139,N_5839);
xor U11612 (N_11612,N_8618,N_6175);
nand U11613 (N_11613,N_6541,N_9176);
and U11614 (N_11614,N_9149,N_8961);
xor U11615 (N_11615,N_5849,N_6818);
nor U11616 (N_11616,N_9138,N_9094);
nand U11617 (N_11617,N_8897,N_8361);
xor U11618 (N_11618,N_9354,N_5991);
nand U11619 (N_11619,N_7897,N_6176);
and U11620 (N_11620,N_8120,N_6570);
xnor U11621 (N_11621,N_5054,N_8044);
xor U11622 (N_11622,N_8644,N_6258);
nor U11623 (N_11623,N_7119,N_8943);
xor U11624 (N_11624,N_8453,N_6758);
nor U11625 (N_11625,N_8777,N_7820);
xnor U11626 (N_11626,N_8746,N_6130);
nor U11627 (N_11627,N_5340,N_7369);
or U11628 (N_11628,N_7955,N_5240);
nand U11629 (N_11629,N_5278,N_7153);
xor U11630 (N_11630,N_9359,N_5343);
nor U11631 (N_11631,N_6947,N_9389);
nand U11632 (N_11632,N_5906,N_5124);
nand U11633 (N_11633,N_6531,N_6174);
or U11634 (N_11634,N_8808,N_5768);
nor U11635 (N_11635,N_6008,N_6540);
and U11636 (N_11636,N_6019,N_5604);
or U11637 (N_11637,N_7053,N_9368);
nor U11638 (N_11638,N_7056,N_6490);
or U11639 (N_11639,N_7315,N_9155);
nand U11640 (N_11640,N_7358,N_6075);
and U11641 (N_11641,N_7662,N_6563);
nand U11642 (N_11642,N_6183,N_6221);
xnor U11643 (N_11643,N_9223,N_5120);
nand U11644 (N_11644,N_5168,N_8869);
nand U11645 (N_11645,N_7757,N_5143);
xnor U11646 (N_11646,N_6211,N_5776);
or U11647 (N_11647,N_6999,N_9338);
nor U11648 (N_11648,N_9172,N_8625);
nand U11649 (N_11649,N_8145,N_8051);
nand U11650 (N_11650,N_5028,N_5545);
nand U11651 (N_11651,N_7271,N_7507);
or U11652 (N_11652,N_7431,N_5672);
nor U11653 (N_11653,N_5725,N_5440);
and U11654 (N_11654,N_8236,N_7252);
nor U11655 (N_11655,N_6887,N_7180);
xor U11656 (N_11656,N_5107,N_9457);
or U11657 (N_11657,N_7800,N_6205);
nor U11658 (N_11658,N_5696,N_5065);
or U11659 (N_11659,N_6425,N_8879);
nand U11660 (N_11660,N_9780,N_9980);
xor U11661 (N_11661,N_8187,N_5292);
xnor U11662 (N_11662,N_8021,N_5338);
nand U11663 (N_11663,N_8502,N_9742);
xor U11664 (N_11664,N_9164,N_6970);
nor U11665 (N_11665,N_8023,N_6888);
nor U11666 (N_11666,N_6876,N_6152);
or U11667 (N_11667,N_6192,N_9136);
or U11668 (N_11668,N_7948,N_7517);
nor U11669 (N_11669,N_9878,N_7774);
and U11670 (N_11670,N_7750,N_5563);
xor U11671 (N_11671,N_5401,N_9208);
and U11672 (N_11672,N_9616,N_8312);
or U11673 (N_11673,N_9951,N_7829);
nor U11674 (N_11674,N_9956,N_5231);
xor U11675 (N_11675,N_8152,N_5027);
xor U11676 (N_11676,N_5406,N_6829);
nand U11677 (N_11677,N_6587,N_9414);
nand U11678 (N_11678,N_6252,N_7134);
and U11679 (N_11679,N_8097,N_6209);
nand U11680 (N_11680,N_5431,N_5067);
xor U11681 (N_11681,N_5126,N_7967);
or U11682 (N_11682,N_8217,N_5149);
or U11683 (N_11683,N_7040,N_7613);
xor U11684 (N_11684,N_9180,N_8368);
xor U11685 (N_11685,N_5623,N_9723);
nor U11686 (N_11686,N_8874,N_9706);
or U11687 (N_11687,N_7722,N_8415);
or U11688 (N_11688,N_9532,N_7211);
nand U11689 (N_11689,N_5101,N_8376);
xor U11690 (N_11690,N_6644,N_6711);
and U11691 (N_11691,N_8335,N_9820);
or U11692 (N_11692,N_9770,N_6212);
nand U11693 (N_11693,N_5213,N_8927);
nor U11694 (N_11694,N_9372,N_6929);
or U11695 (N_11695,N_7692,N_9114);
xnor U11696 (N_11696,N_5800,N_7160);
or U11697 (N_11697,N_9167,N_8664);
nor U11698 (N_11698,N_8995,N_9879);
or U11699 (N_11699,N_8344,N_9205);
and U11700 (N_11700,N_8104,N_9281);
nor U11701 (N_11701,N_8058,N_8466);
nor U11702 (N_11702,N_6913,N_7399);
nand U11703 (N_11703,N_7238,N_7758);
nor U11704 (N_11704,N_9692,N_6467);
and U11705 (N_11705,N_5744,N_8325);
nor U11706 (N_11706,N_8736,N_9521);
or U11707 (N_11707,N_9769,N_7609);
nand U11708 (N_11708,N_8574,N_6119);
or U11709 (N_11709,N_5050,N_7241);
nand U11710 (N_11710,N_6631,N_5930);
or U11711 (N_11711,N_9622,N_6522);
xor U11712 (N_11712,N_6308,N_8988);
nand U11713 (N_11713,N_7883,N_7959);
and U11714 (N_11714,N_9342,N_5547);
xnor U11715 (N_11715,N_5690,N_9712);
nand U11716 (N_11716,N_9088,N_7003);
and U11717 (N_11717,N_6347,N_7275);
xor U11718 (N_11718,N_6222,N_8594);
and U11719 (N_11719,N_8053,N_9890);
xnor U11720 (N_11720,N_6718,N_5022);
and U11721 (N_11721,N_5342,N_7406);
nor U11722 (N_11722,N_8129,N_8607);
nor U11723 (N_11723,N_6115,N_8179);
nand U11724 (N_11724,N_7499,N_6015);
nand U11725 (N_11725,N_7815,N_9468);
nand U11726 (N_11726,N_8260,N_7560);
xnor U11727 (N_11727,N_8779,N_7745);
nor U11728 (N_11728,N_8656,N_5939);
nand U11729 (N_11729,N_6003,N_6752);
and U11730 (N_11730,N_6454,N_5878);
or U11731 (N_11731,N_9741,N_8893);
xnor U11732 (N_11732,N_5622,N_5686);
and U11733 (N_11733,N_6452,N_6315);
nand U11734 (N_11734,N_7694,N_5628);
nand U11735 (N_11735,N_9660,N_7529);
or U11736 (N_11736,N_5922,N_5011);
nand U11737 (N_11737,N_6667,N_7016);
nor U11738 (N_11738,N_7685,N_7635);
or U11739 (N_11739,N_5967,N_5510);
and U11740 (N_11740,N_8520,N_6074);
and U11741 (N_11741,N_7630,N_7273);
or U11742 (N_11742,N_6408,N_8472);
nor U11743 (N_11743,N_9413,N_6785);
or U11744 (N_11744,N_8695,N_5578);
nor U11745 (N_11745,N_6586,N_6658);
xor U11746 (N_11746,N_9553,N_5140);
and U11747 (N_11747,N_7670,N_6963);
xnor U11748 (N_11748,N_8945,N_7340);
or U11749 (N_11749,N_6894,N_8616);
xnor U11750 (N_11750,N_8072,N_9100);
or U11751 (N_11751,N_9352,N_5267);
nor U11752 (N_11752,N_7011,N_8671);
nor U11753 (N_11753,N_7885,N_9234);
xnor U11754 (N_11754,N_9857,N_5346);
xor U11755 (N_11755,N_6381,N_5350);
and U11756 (N_11756,N_6774,N_8543);
or U11757 (N_11757,N_8371,N_9676);
and U11758 (N_11758,N_8348,N_6804);
and U11759 (N_11759,N_5121,N_5319);
and U11760 (N_11760,N_9918,N_5069);
xnor U11761 (N_11761,N_7570,N_9445);
or U11762 (N_11762,N_7970,N_7098);
and U11763 (N_11763,N_6505,N_5110);
nand U11764 (N_11764,N_6635,N_5486);
or U11765 (N_11765,N_9369,N_6041);
xor U11766 (N_11766,N_6022,N_7742);
nand U11767 (N_11767,N_5789,N_6852);
xor U11768 (N_11768,N_5410,N_8013);
nor U11769 (N_11769,N_6413,N_9618);
nand U11770 (N_11770,N_6596,N_6472);
xor U11771 (N_11771,N_5000,N_5709);
nand U11772 (N_11772,N_9073,N_6851);
nor U11773 (N_11773,N_7931,N_9760);
and U11774 (N_11774,N_9869,N_6567);
or U11775 (N_11775,N_7099,N_7129);
or U11776 (N_11776,N_8584,N_7117);
nor U11777 (N_11777,N_6543,N_8895);
and U11778 (N_11778,N_8744,N_8270);
xnor U11779 (N_11779,N_5351,N_9259);
xnor U11780 (N_11780,N_8303,N_6746);
xnor U11781 (N_11781,N_9930,N_8753);
xor U11782 (N_11782,N_5318,N_7947);
or U11783 (N_11783,N_9460,N_8910);
nor U11784 (N_11784,N_9589,N_5582);
and U11785 (N_11785,N_7250,N_8364);
nand U11786 (N_11786,N_5155,N_5971);
and U11787 (N_11787,N_7323,N_9487);
nor U11788 (N_11788,N_5224,N_8985);
and U11789 (N_11789,N_6292,N_8635);
xnor U11790 (N_11790,N_9801,N_9538);
xor U11791 (N_11791,N_9171,N_9853);
xor U11792 (N_11792,N_9886,N_7521);
and U11793 (N_11793,N_8234,N_9038);
and U11794 (N_11794,N_8269,N_6378);
and U11795 (N_11795,N_9597,N_6331);
xnor U11796 (N_11796,N_6297,N_5539);
nor U11797 (N_11797,N_7407,N_5038);
or U11798 (N_11798,N_8089,N_5876);
xnor U11799 (N_11799,N_8076,N_8655);
and U11800 (N_11800,N_9523,N_6233);
xor U11801 (N_11801,N_9143,N_8310);
nor U11802 (N_11802,N_8608,N_7646);
xnor U11803 (N_11803,N_5913,N_6284);
or U11804 (N_11804,N_5457,N_5975);
xnor U11805 (N_11805,N_7636,N_9430);
and U11806 (N_11806,N_6283,N_5203);
nand U11807 (N_11807,N_9040,N_5165);
xnor U11808 (N_11808,N_5323,N_8216);
nor U11809 (N_11809,N_5061,N_9307);
or U11810 (N_11810,N_6026,N_8890);
or U11811 (N_11811,N_7415,N_5990);
or U11812 (N_11812,N_6094,N_8115);
nor U11813 (N_11813,N_8595,N_6278);
nor U11814 (N_11814,N_7808,N_6411);
nand U11815 (N_11815,N_8398,N_5382);
or U11816 (N_11816,N_9188,N_5964);
xnor U11817 (N_11817,N_7645,N_7654);
or U11818 (N_11818,N_8573,N_5649);
and U11819 (N_11819,N_7079,N_7753);
or U11820 (N_11820,N_9485,N_6113);
or U11821 (N_11821,N_9186,N_5163);
nand U11822 (N_11822,N_6796,N_8225);
and U11823 (N_11823,N_6312,N_5590);
or U11824 (N_11824,N_7126,N_7355);
nand U11825 (N_11825,N_7184,N_5487);
nor U11826 (N_11826,N_6431,N_7155);
xnor U11827 (N_11827,N_9568,N_8911);
and U11828 (N_11828,N_8290,N_9554);
or U11829 (N_11829,N_8950,N_6228);
and U11830 (N_11830,N_7789,N_6234);
xor U11831 (N_11831,N_5775,N_5920);
nor U11832 (N_11832,N_7728,N_6321);
xor U11833 (N_11833,N_6300,N_9001);
or U11834 (N_11834,N_9104,N_5684);
nor U11835 (N_11835,N_8829,N_9438);
xor U11836 (N_11836,N_7564,N_9318);
nand U11837 (N_11837,N_5375,N_8553);
nor U11838 (N_11838,N_7690,N_9510);
nand U11839 (N_11839,N_7557,N_7158);
and U11840 (N_11840,N_9395,N_9815);
or U11841 (N_11841,N_7018,N_5514);
nand U11842 (N_11842,N_9392,N_7095);
or U11843 (N_11843,N_8868,N_5792);
or U11844 (N_11844,N_6500,N_8135);
nand U11845 (N_11845,N_7528,N_9472);
and U11846 (N_11846,N_8781,N_7466);
nand U11847 (N_11847,N_6110,N_9330);
nand U11848 (N_11848,N_5258,N_7021);
or U11849 (N_11849,N_9867,N_8463);
or U11850 (N_11850,N_8117,N_8402);
or U11851 (N_11851,N_9731,N_7379);
nor U11852 (N_11852,N_5598,N_8773);
or U11853 (N_11853,N_7825,N_6185);
nand U11854 (N_11854,N_8796,N_6784);
or U11855 (N_11855,N_5675,N_5418);
nor U11856 (N_11856,N_5217,N_7037);
or U11857 (N_11857,N_5288,N_8975);
or U11858 (N_11858,N_7579,N_6986);
or U11859 (N_11859,N_5246,N_6928);
nand U11860 (N_11860,N_9914,N_7455);
or U11861 (N_11861,N_8954,N_9240);
or U11862 (N_11862,N_8308,N_5106);
nand U11863 (N_11863,N_9078,N_6214);
nand U11864 (N_11864,N_5579,N_6245);
and U11865 (N_11865,N_9818,N_8637);
nand U11866 (N_11866,N_5850,N_5405);
and U11867 (N_11867,N_8705,N_7228);
and U11868 (N_11868,N_7913,N_5770);
nor U11869 (N_11869,N_6771,N_6348);
and U11870 (N_11870,N_9787,N_9602);
xnor U11871 (N_11871,N_9444,N_7149);
and U11872 (N_11872,N_7796,N_9964);
or U11873 (N_11873,N_8275,N_6355);
xnor U11874 (N_11874,N_9054,N_8725);
and U11875 (N_11875,N_8997,N_6664);
nor U11876 (N_11876,N_7170,N_7424);
nand U11877 (N_11877,N_8550,N_5162);
nor U11878 (N_11878,N_5419,N_6735);
or U11879 (N_11879,N_5635,N_6068);
nand U11880 (N_11880,N_7857,N_6142);
nor U11881 (N_11881,N_9431,N_8727);
nand U11882 (N_11882,N_6951,N_7798);
nor U11883 (N_11883,N_9942,N_8848);
and U11884 (N_11884,N_5392,N_7397);
and U11885 (N_11885,N_5179,N_8178);
and U11886 (N_11886,N_5840,N_6149);
or U11887 (N_11887,N_9652,N_9486);
xor U11888 (N_11888,N_9514,N_7902);
or U11889 (N_11889,N_8507,N_9491);
and U11890 (N_11890,N_7984,N_5629);
nand U11891 (N_11891,N_9212,N_9358);
xnor U11892 (N_11892,N_8766,N_5703);
nor U11893 (N_11893,N_5297,N_5039);
and U11894 (N_11894,N_7199,N_9992);
or U11895 (N_11895,N_6520,N_5813);
or U11896 (N_11896,N_5592,N_6231);
nand U11897 (N_11897,N_7585,N_8160);
nand U11898 (N_11898,N_6528,N_9163);
nand U11899 (N_11899,N_8381,N_8157);
or U11900 (N_11900,N_5270,N_7683);
nor U11901 (N_11901,N_9452,N_6634);
or U11902 (N_11902,N_8091,N_7510);
or U11903 (N_11903,N_6866,N_5393);
or U11904 (N_11904,N_9985,N_5474);
or U11905 (N_11905,N_8541,N_9540);
nor U11906 (N_11906,N_8836,N_6781);
xnor U11907 (N_11907,N_8794,N_8446);
and U11908 (N_11908,N_5762,N_8345);
nor U11909 (N_11909,N_7108,N_5851);
nor U11910 (N_11910,N_6317,N_7584);
nand U11911 (N_11911,N_6641,N_9621);
nor U11912 (N_11912,N_9883,N_5321);
xor U11913 (N_11913,N_8273,N_8065);
xor U11914 (N_11914,N_6168,N_5058);
nor U11915 (N_11915,N_7027,N_9198);
nor U11916 (N_11916,N_7747,N_5630);
nor U11917 (N_11917,N_9299,N_8441);
nor U11918 (N_11918,N_6994,N_5685);
and U11919 (N_11919,N_5624,N_8527);
nand U11920 (N_11920,N_5390,N_9293);
xor U11921 (N_11921,N_8709,N_7057);
xnor U11922 (N_11922,N_9065,N_7210);
or U11923 (N_11923,N_6566,N_9375);
and U11924 (N_11924,N_7438,N_9788);
xor U11925 (N_11925,N_9691,N_5714);
nand U11926 (N_11926,N_8589,N_6716);
nor U11927 (N_11927,N_6956,N_5879);
nor U11928 (N_11928,N_9726,N_9242);
or U11929 (N_11929,N_7195,N_6388);
nor U11930 (N_11930,N_8811,N_5522);
and U11931 (N_11931,N_6682,N_9279);
or U11932 (N_11932,N_7266,N_6485);
xor U11933 (N_11933,N_5642,N_7375);
or U11934 (N_11934,N_9348,N_6903);
nand U11935 (N_11935,N_8751,N_9398);
or U11936 (N_11936,N_6220,N_5347);
xor U11937 (N_11937,N_8286,N_8395);
or U11938 (N_11938,N_8729,N_8099);
or U11939 (N_11939,N_5769,N_5144);
nor U11940 (N_11940,N_5447,N_7411);
or U11941 (N_11941,N_5614,N_9643);
and U11942 (N_11942,N_9534,N_8623);
and U11943 (N_11943,N_5200,N_8547);
and U11944 (N_11944,N_6845,N_8880);
xor U11945 (N_11945,N_6618,N_6953);
nand U11946 (N_11946,N_6732,N_8377);
or U11947 (N_11947,N_7936,N_7280);
nor U11948 (N_11948,N_7629,N_6910);
nand U11949 (N_11949,N_5589,N_6294);
and U11950 (N_11950,N_8949,N_9749);
or U11951 (N_11951,N_5185,N_9685);
or U11952 (N_11952,N_5831,N_6706);
nor U11953 (N_11953,N_7113,N_5013);
or U11954 (N_11954,N_9200,N_5194);
nand U11955 (N_11955,N_9665,N_9610);
nor U11956 (N_11956,N_8329,N_7373);
or U11957 (N_11957,N_8098,N_6035);
and U11958 (N_11958,N_9120,N_7020);
or U11959 (N_11959,N_8128,N_5998);
or U11960 (N_11960,N_7151,N_7667);
or U11961 (N_11961,N_5451,N_9517);
nand U11962 (N_11962,N_9789,N_8205);
or U11963 (N_11963,N_6959,N_9893);
nor U11964 (N_11964,N_6102,N_6941);
nand U11965 (N_11965,N_7552,N_6717);
and U11966 (N_11966,N_7055,N_9232);
nor U11967 (N_11967,N_8136,N_8392);
nor U11968 (N_11968,N_9786,N_6069);
nor U11969 (N_11969,N_7478,N_5893);
xor U11970 (N_11970,N_5799,N_5698);
nor U11971 (N_11971,N_9428,N_9294);
or U11972 (N_11972,N_9876,N_6135);
nand U11973 (N_11973,N_9493,N_6581);
and U11974 (N_11974,N_6755,N_7240);
or U11975 (N_11975,N_7167,N_5530);
and U11976 (N_11976,N_7194,N_5949);
nand U11977 (N_11977,N_5736,N_5667);
nand U11978 (N_11978,N_9385,N_8374);
xnor U11979 (N_11979,N_8086,N_6995);
and U11980 (N_11980,N_5741,N_9965);
xor U11981 (N_11981,N_6059,N_9972);
nand U11982 (N_11982,N_6745,N_7898);
or U11983 (N_11983,N_8378,N_6184);
or U11984 (N_11984,N_6006,N_5887);
nand U11985 (N_11985,N_7394,N_6401);
or U11986 (N_11986,N_9254,N_7551);
xnor U11987 (N_11987,N_8188,N_8639);
and U11988 (N_11988,N_9783,N_9110);
nor U11989 (N_11989,N_7029,N_8017);
xnor U11990 (N_11990,N_5543,N_8710);
nor U11991 (N_11991,N_7726,N_9641);
and U11992 (N_11992,N_7650,N_5521);
nor U11993 (N_11993,N_5332,N_8282);
and U11994 (N_11994,N_5819,N_6407);
xor U11995 (N_11995,N_5283,N_5092);
and U11996 (N_11996,N_8468,N_8313);
xor U11997 (N_11997,N_5439,N_6918);
or U11998 (N_11998,N_5693,N_5803);
or U11999 (N_11999,N_8525,N_8479);
nand U12000 (N_12000,N_5765,N_8054);
and U12001 (N_12001,N_7159,N_8184);
xor U12002 (N_12002,N_8697,N_6838);
and U12003 (N_12003,N_9502,N_6833);
nor U12004 (N_12004,N_5896,N_8455);
or U12005 (N_12005,N_8977,N_8002);
or U12006 (N_12006,N_9453,N_9481);
nor U12007 (N_12007,N_6764,N_6473);
xnor U12008 (N_12008,N_9194,N_9648);
nand U12009 (N_12009,N_7527,N_7265);
nand U12010 (N_12010,N_8780,N_5525);
nand U12011 (N_12011,N_6842,N_6967);
nor U12012 (N_12012,N_6595,N_9739);
nand U12013 (N_12013,N_6495,N_5797);
and U12014 (N_12014,N_7547,N_7363);
nand U12015 (N_12015,N_6741,N_7165);
or U12016 (N_12016,N_8875,N_8972);
nor U12017 (N_12017,N_5944,N_7010);
nor U12018 (N_12018,N_6883,N_9975);
or U12019 (N_12019,N_6585,N_5620);
nand U12020 (N_12020,N_9043,N_9023);
and U12021 (N_12021,N_6043,N_8691);
or U12022 (N_12022,N_6753,N_7872);
nand U12023 (N_12023,N_5820,N_9868);
nand U12024 (N_12024,N_5244,N_5276);
and U12025 (N_12025,N_9286,N_9344);
or U12026 (N_12026,N_6090,N_6419);
xnor U12027 (N_12027,N_5499,N_7994);
nand U12028 (N_12028,N_7317,N_9773);
or U12029 (N_12029,N_6899,N_8063);
and U12030 (N_12030,N_5817,N_9429);
or U12031 (N_12031,N_9833,N_9647);
or U12032 (N_12032,N_8332,N_5220);
nand U12033 (N_12033,N_6504,N_6449);
nor U12034 (N_12034,N_6519,N_9803);
or U12035 (N_12035,N_8162,N_8318);
and U12036 (N_12036,N_7614,N_5018);
xnor U12037 (N_12037,N_8350,N_8182);
and U12038 (N_12038,N_9477,N_8505);
and U12039 (N_12039,N_6679,N_7535);
nor U12040 (N_12040,N_6551,N_8821);
or U12041 (N_12041,N_5874,N_5260);
or U12042 (N_12042,N_8116,N_9509);
xor U12043 (N_12043,N_9666,N_6474);
nor U12044 (N_12044,N_8315,N_9673);
and U12045 (N_12045,N_6790,N_5153);
or U12046 (N_12046,N_7549,N_7330);
nand U12047 (N_12047,N_8219,N_5358);
and U12048 (N_12048,N_5562,N_9099);
and U12049 (N_12049,N_8609,N_8873);
and U12050 (N_12050,N_7023,N_8192);
and U12051 (N_12051,N_8110,N_8889);
and U12052 (N_12052,N_7248,N_8062);
xor U12053 (N_12053,N_9638,N_7793);
nor U12054 (N_12054,N_7456,N_7847);
xor U12055 (N_12055,N_6215,N_7283);
nand U12056 (N_12056,N_7146,N_5867);
nor U12057 (N_12057,N_7372,N_5129);
nor U12058 (N_12058,N_5863,N_5699);
nand U12059 (N_12059,N_8500,N_6905);
nor U12060 (N_12060,N_8492,N_8302);
xnor U12061 (N_12061,N_8052,N_8373);
xor U12062 (N_12062,N_9580,N_9374);
nand U12063 (N_12063,N_9488,N_7809);
nor U12064 (N_12064,N_7721,N_6571);
and U12065 (N_12065,N_9409,N_7611);
and U12066 (N_12066,N_9976,N_5094);
and U12067 (N_12067,N_6997,N_8203);
and U12068 (N_12068,N_9757,N_8485);
or U12069 (N_12069,N_8177,N_6817);
nand U12070 (N_12070,N_9102,N_8896);
nand U12071 (N_12071,N_6515,N_9623);
and U12072 (N_12072,N_6920,N_6402);
and U12073 (N_12073,N_5641,N_8533);
and U12074 (N_12074,N_9292,N_6392);
and U12075 (N_12075,N_6147,N_5354);
xnor U12076 (N_12076,N_8636,N_5632);
nand U12077 (N_12077,N_9028,N_9565);
and U12078 (N_12078,N_7264,N_5626);
nand U12079 (N_12079,N_8642,N_8064);
nor U12080 (N_12080,N_7810,N_7526);
and U12081 (N_12081,N_8754,N_7821);
xnor U12082 (N_12082,N_9822,N_7583);
nand U12083 (N_12083,N_6116,N_5108);
nand U12084 (N_12084,N_5468,N_7544);
nor U12085 (N_12085,N_8597,N_6677);
nor U12086 (N_12086,N_6623,N_9902);
and U12087 (N_12087,N_8941,N_7712);
nand U12088 (N_12088,N_6479,N_6178);
xnor U12089 (N_12089,N_6681,N_9373);
or U12090 (N_12090,N_5962,N_7589);
or U12091 (N_12091,N_7626,N_9255);
xor U12092 (N_12092,N_5978,N_5221);
nor U12093 (N_12093,N_5697,N_6241);
or U12094 (N_12094,N_5305,N_7295);
or U12095 (N_12095,N_5029,N_9733);
xor U12096 (N_12096,N_8940,N_5916);
and U12097 (N_12097,N_5923,N_5650);
or U12098 (N_12098,N_6798,N_9287);
or U12099 (N_12099,N_7425,N_6435);
or U12100 (N_12100,N_7680,N_8121);
and U12101 (N_12101,N_7651,N_6839);
nor U12102 (N_12102,N_6698,N_9544);
nor U12103 (N_12103,N_8435,N_8748);
xor U12104 (N_12104,N_9160,N_8011);
nor U12105 (N_12105,N_6280,N_9137);
nor U12106 (N_12106,N_6605,N_7834);
and U12107 (N_12107,N_8165,N_9036);
xnor U12108 (N_12108,N_6493,N_7244);
xnor U12109 (N_12109,N_7041,N_6661);
and U12110 (N_12110,N_5953,N_6237);
nand U12111 (N_12111,N_9907,N_9245);
and U12112 (N_12112,N_7279,N_9183);
and U12113 (N_12113,N_5268,N_6792);
or U12114 (N_12114,N_7451,N_6104);
or U12115 (N_12115,N_5591,N_7832);
nor U12116 (N_12116,N_9906,N_6914);
xor U12117 (N_12117,N_8474,N_5646);
nand U12118 (N_12118,N_8901,N_9970);
xor U12119 (N_12119,N_8494,N_6247);
nand U12120 (N_12120,N_7430,N_5053);
and U12121 (N_12121,N_6778,N_9107);
and U12122 (N_12122,N_8914,N_7761);
nand U12123 (N_12123,N_5994,N_5190);
nor U12124 (N_12124,N_7175,N_9159);
nand U12125 (N_12125,N_6336,N_9024);
nor U12126 (N_12126,N_7957,N_8174);
nor U12127 (N_12127,N_5461,N_7005);
nand U12128 (N_12128,N_7339,N_8176);
and U12129 (N_12129,N_8842,N_9898);
or U12130 (N_12130,N_6012,N_6450);
xnor U12131 (N_12131,N_7255,N_5715);
and U12132 (N_12132,N_8037,N_7968);
or U12133 (N_12133,N_6958,N_5726);
or U12134 (N_12134,N_9590,N_8649);
or U12135 (N_12135,N_8621,N_9651);
nand U12136 (N_12136,N_9019,N_7558);
nor U12137 (N_12137,N_5870,N_9961);
and U12138 (N_12138,N_7221,N_6230);
and U12139 (N_12139,N_7253,N_5536);
xor U12140 (N_12140,N_5454,N_6700);
or U12141 (N_12141,N_9872,N_7335);
xor U12142 (N_12142,N_5528,N_5308);
or U12143 (N_12143,N_7926,N_5040);
xor U12144 (N_12144,N_7546,N_9549);
xor U12145 (N_12145,N_7209,N_5777);
and U12146 (N_12146,N_7574,N_5542);
nor U12147 (N_12147,N_5594,N_9816);
nor U12148 (N_12148,N_9650,N_8701);
nor U12149 (N_12149,N_5025,N_8611);
and U12150 (N_12150,N_6739,N_8096);
nor U12151 (N_12151,N_5613,N_6912);
xor U12152 (N_12152,N_7805,N_5052);
or U12153 (N_12153,N_9642,N_8323);
xnor U12154 (N_12154,N_5771,N_6360);
xor U12155 (N_12155,N_5933,N_9562);
xnor U12156 (N_12156,N_5485,N_6117);
xor U12157 (N_12157,N_6908,N_8539);
nand U12158 (N_12158,N_9874,N_5662);
or U12159 (N_12159,N_6034,N_8998);
nand U12160 (N_12160,N_6550,N_8822);
and U12161 (N_12161,N_9515,N_5888);
and U12162 (N_12162,N_6578,N_6254);
and U12163 (N_12163,N_9933,N_5277);
and U12164 (N_12164,N_6380,N_8802);
and U12165 (N_12165,N_8352,N_5498);
xor U12166 (N_12166,N_7103,N_9506);
or U12167 (N_12167,N_6628,N_8937);
nor U12168 (N_12168,N_8515,N_7767);
or U12169 (N_12169,N_7648,N_5935);
or U12170 (N_12170,N_5917,N_5252);
or U12171 (N_12171,N_9632,N_7459);
nor U12172 (N_12172,N_6972,N_5060);
nand U12173 (N_12173,N_9391,N_6546);
nor U12174 (N_12174,N_5442,N_9275);
xor U12175 (N_12175,N_5549,N_9418);
nor U12176 (N_12176,N_5827,N_7695);
and U12177 (N_12177,N_7505,N_9708);
xnor U12178 (N_12178,N_6783,N_6484);
nor U12179 (N_12179,N_6601,N_5861);
or U12180 (N_12180,N_6660,N_6808);
xor U12181 (N_12181,N_9297,N_7736);
nor U12182 (N_12182,N_7087,N_6080);
and U12183 (N_12183,N_7091,N_5644);
nand U12184 (N_12184,N_6270,N_8817);
xnor U12185 (N_12185,N_7185,N_7592);
or U12186 (N_12186,N_9098,N_5742);
nor U12187 (N_12187,N_6486,N_6917);
or U12188 (N_12188,N_9478,N_5341);
nor U12189 (N_12189,N_5156,N_6448);
and U12190 (N_12190,N_6264,N_8289);
and U12191 (N_12191,N_8663,N_7190);
xnor U12192 (N_12192,N_5943,N_7554);
nor U12193 (N_12193,N_8860,N_8887);
nand U12194 (N_12194,N_8906,N_6890);
nor U12195 (N_12195,N_5388,N_6748);
and U12196 (N_12196,N_8126,N_6687);
and U12197 (N_12197,N_9845,N_8131);
xnor U12198 (N_12198,N_7463,N_8238);
nor U12199 (N_12199,N_7618,N_6983);
and U12200 (N_12200,N_9017,N_9135);
or U12201 (N_12201,N_6054,N_7487);
xor U12202 (N_12202,N_6575,N_7214);
and U12203 (N_12203,N_8370,N_5580);
xnor U12204 (N_12204,N_6160,N_9929);
or U12205 (N_12205,N_5166,N_9190);
nor U12206 (N_12206,N_9582,N_9870);
xor U12207 (N_12207,N_5757,N_5286);
xor U12208 (N_12208,N_9996,N_9058);
or U12209 (N_12209,N_6561,N_9049);
nand U12210 (N_12210,N_8272,N_8686);
or U12211 (N_12211,N_8661,N_5261);
or U12212 (N_12212,N_5438,N_9662);
and U12213 (N_12213,N_5809,N_5411);
nor U12214 (N_12214,N_6693,N_6868);
nor U12215 (N_12215,N_9664,N_6238);
or U12216 (N_12216,N_7371,N_7494);
and U12217 (N_12217,N_8537,N_7814);
nand U12218 (N_12218,N_8775,N_7348);
and U12219 (N_12219,N_7625,N_7666);
or U12220 (N_12220,N_7422,N_9356);
xor U12221 (N_12221,N_7019,N_5584);
xor U12222 (N_12222,N_6243,N_8397);
and U12223 (N_12223,N_5363,N_7978);
or U12224 (N_12224,N_6856,N_9074);
nor U12225 (N_12225,N_5452,N_6096);
or U12226 (N_12226,N_6971,N_7128);
nor U12227 (N_12227,N_7875,N_9222);
nor U12228 (N_12228,N_9310,N_9896);
nand U12229 (N_12229,N_6938,N_6305);
or U12230 (N_12230,N_7954,N_6060);
or U12231 (N_12231,N_6483,N_5093);
or U12232 (N_12232,N_5838,N_5057);
nand U12233 (N_12233,N_9404,N_7231);
xor U12234 (N_12234,N_6583,N_8648);
nand U12235 (N_12235,N_9170,N_9328);
nor U12236 (N_12236,N_9940,N_5175);
nor U12237 (N_12237,N_9949,N_7977);
xnor U12238 (N_12238,N_9838,N_6688);
nor U12239 (N_12239,N_9411,N_9419);
nand U12240 (N_12240,N_5553,N_8735);
nand U12241 (N_12241,N_9901,N_6010);
nand U12242 (N_12242,N_7784,N_8749);
nor U12243 (N_12243,N_5089,N_5496);
or U12244 (N_12244,N_7713,N_6647);
and U12245 (N_12245,N_7069,N_9798);
nor U12246 (N_12246,N_8783,N_8331);
xor U12247 (N_12247,N_8878,N_5201);
nand U12248 (N_12248,N_9938,N_7702);
xnor U12249 (N_12249,N_9987,N_9913);
nand U12250 (N_12250,N_5239,N_8212);
nand U12251 (N_12251,N_8436,N_9672);
nand U12252 (N_12252,N_5043,N_7833);
xor U12253 (N_12253,N_8964,N_5739);
nor U12254 (N_12254,N_6603,N_8740);
xor U12255 (N_12255,N_5302,N_6710);
and U12256 (N_12256,N_8567,N_5824);
nand U12257 (N_12257,N_7818,N_5537);
nor U12258 (N_12258,N_9974,N_5593);
and U12259 (N_12259,N_5491,N_8396);
nand U12260 (N_12260,N_7981,N_5386);
nand U12261 (N_12261,N_6343,N_5223);
xor U12262 (N_12262,N_7987,N_8476);
or U12263 (N_12263,N_9828,N_5538);
and U12264 (N_12264,N_6078,N_8384);
and U12265 (N_12265,N_7305,N_8657);
or U12266 (N_12266,N_8296,N_6882);
or U12267 (N_12267,N_8291,N_5113);
nand U12268 (N_12268,N_5663,N_7656);
xnor U12269 (N_12269,N_9396,N_7838);
nor U12270 (N_12270,N_7940,N_6987);
nand U12271 (N_12271,N_8024,N_6689);
xnor U12272 (N_12272,N_5666,N_7819);
or U12273 (N_12273,N_8449,N_6864);
or U12274 (N_12274,N_5399,N_7811);
or U12275 (N_12275,N_7352,N_5713);
or U12276 (N_12276,N_7293,N_9336);
xnor U12277 (N_12277,N_8124,N_9270);
xnor U12278 (N_12278,N_9620,N_6767);
or U12279 (N_12279,N_5541,N_9608);
nor U12280 (N_12280,N_9204,N_9433);
nor U12281 (N_12281,N_6642,N_5187);
or U12282 (N_12282,N_8226,N_8320);
nand U12283 (N_12283,N_6396,N_6286);
nand U12284 (N_12284,N_8593,N_6389);
xor U12285 (N_12285,N_5516,N_8534);
and U12286 (N_12286,N_9248,N_5921);
or U12287 (N_12287,N_7140,N_9767);
or U12288 (N_12288,N_9948,N_5289);
xnor U12289 (N_12289,N_5801,N_6699);
xor U12290 (N_12290,N_9729,N_6978);
or U12291 (N_12291,N_6372,N_8421);
nor U12292 (N_12292,N_5441,N_6260);
and U12293 (N_12293,N_8143,N_5446);
or U12294 (N_12294,N_6731,N_8548);
and U12295 (N_12295,N_6653,N_9406);
xor U12296 (N_12296,N_5197,N_5362);
and U12297 (N_12297,N_5665,N_7737);
xnor U12298 (N_12298,N_6227,N_8826);
and U12299 (N_12299,N_9999,N_8925);
xor U12300 (N_12300,N_6974,N_8569);
nor U12301 (N_12301,N_8682,N_6786);
nand U12302 (N_12302,N_9435,N_6604);
nor U12303 (N_12303,N_5857,N_7384);
xnor U12304 (N_12304,N_7896,N_9129);
xor U12305 (N_12305,N_7076,N_8171);
nor U12306 (N_12306,N_9047,N_6776);
and U12307 (N_12307,N_7615,N_6171);
xor U12308 (N_12308,N_6529,N_5295);
and U12309 (N_12309,N_7911,N_7949);
or U12310 (N_12310,N_9108,N_7844);
and U12311 (N_12311,N_7938,N_9377);
and U12312 (N_12312,N_6417,N_5691);
xor U12313 (N_12313,N_9959,N_9854);
nand U12314 (N_12314,N_6794,N_8108);
or U12315 (N_12315,N_5910,N_6797);
nand U12316 (N_12316,N_7433,N_5503);
or U12317 (N_12317,N_8558,N_9278);
xnor U12318 (N_12318,N_6557,N_6523);
nand U12319 (N_12319,N_8322,N_6424);
nand U12320 (N_12320,N_8154,N_5367);
nor U12321 (N_12321,N_5788,N_7286);
and U12322 (N_12322,N_8581,N_9497);
nand U12323 (N_12323,N_5424,N_5151);
nand U12324 (N_12324,N_5317,N_7576);
xor U12325 (N_12325,N_7477,N_6675);
and U12326 (N_12326,N_6046,N_8060);
nor U12327 (N_12327,N_5010,N_6024);
nand U12328 (N_12328,N_5250,N_5869);
nand U12329 (N_12329,N_6255,N_6662);
nor U12330 (N_12330,N_7697,N_9669);
nand U12331 (N_12331,N_9802,N_8689);
nand U12332 (N_12332,N_9555,N_8118);
xnor U12333 (N_12333,N_7307,N_8019);
nor U12334 (N_12334,N_9340,N_5256);
xnor U12335 (N_12335,N_9505,N_7519);
and U12336 (N_12336,N_8093,N_7627);
xnor U12337 (N_12337,N_6562,N_6364);
or U12338 (N_12338,N_7493,N_5087);
nand U12339 (N_12339,N_5787,N_5657);
and U12340 (N_12340,N_5037,N_9192);
nand U12341 (N_12341,N_6846,N_6834);
nand U12342 (N_12342,N_6334,N_7483);
nand U12343 (N_12343,N_5676,N_5458);
nor U12344 (N_12344,N_8571,N_6811);
nand U12345 (N_12345,N_6499,N_8894);
nor U12346 (N_12346,N_5230,N_7788);
nor U12347 (N_12347,N_6387,N_7878);
or U12348 (N_12348,N_5369,N_7484);
xnor U12349 (N_12349,N_7156,N_8503);
nand U12350 (N_12350,N_5554,N_8728);
nor U12351 (N_12351,N_7088,N_7879);
nand U12352 (N_12352,N_6548,N_9881);
or U12353 (N_12353,N_7169,N_6580);
xor U12354 (N_12354,N_7566,N_7036);
nor U12355 (N_12355,N_9177,N_9214);
nand U12356 (N_12356,N_7197,N_9162);
or U12357 (N_12357,N_6395,N_7945);
or U12358 (N_12358,N_6879,N_5740);
and U12359 (N_12359,N_8514,N_5597);
nor U12360 (N_12360,N_6800,N_8706);
and U12361 (N_12361,N_9057,N_7192);
and U12362 (N_12362,N_5384,N_5079);
nor U12363 (N_12363,N_7942,N_5798);
xor U12364 (N_12364,N_6250,N_7229);
xor U12365 (N_12365,N_7647,N_7686);
or U12366 (N_12366,N_5524,N_5353);
and U12367 (N_12367,N_6860,N_8004);
nor U12368 (N_12368,N_7410,N_9829);
nand U12369 (N_12369,N_9993,N_9526);
and U12370 (N_12370,N_8734,N_8113);
or U12371 (N_12371,N_7826,N_5979);
nand U12372 (N_12372,N_7418,N_6443);
nand U12373 (N_12373,N_6759,N_5701);
nor U12374 (N_12374,N_9051,N_6812);
or U12375 (N_12375,N_5899,N_9606);
and U12376 (N_12376,N_5488,N_9920);
nand U12377 (N_12377,N_9492,N_9863);
and U12378 (N_12378,N_7022,N_7804);
or U12379 (N_12379,N_6203,N_9657);
and U12380 (N_12380,N_6099,N_5993);
nor U12381 (N_12381,N_6547,N_5004);
or U12382 (N_12382,N_8865,N_9189);
xor U12383 (N_12383,N_8924,N_6624);
nand U12384 (N_12384,N_5947,N_7643);
and U12385 (N_12385,N_7042,N_5804);
and U12386 (N_12386,N_9295,N_8984);
nand U12387 (N_12387,N_6510,N_6738);
nand U12388 (N_12388,N_8464,N_5519);
and U12389 (N_12389,N_7025,N_7677);
xnor U12390 (N_12390,N_7465,N_6680);
and U12391 (N_12391,N_5586,N_9376);
and U12392 (N_12392,N_9362,N_9206);
xnor U12393 (N_12393,N_8918,N_5791);
nor U12394 (N_12394,N_5723,N_7768);
or U12395 (N_12395,N_7490,N_6727);
nor U12396 (N_12396,N_7138,N_5371);
nand U12397 (N_12397,N_6464,N_7183);
xor U12398 (N_12398,N_9068,N_7537);
or U12399 (N_12399,N_5167,N_6632);
or U12400 (N_12400,N_5504,N_9103);
or U12401 (N_12401,N_7312,N_6729);
or U12402 (N_12402,N_8445,N_7816);
or U12403 (N_12403,N_6332,N_7009);
and U12404 (N_12404,N_7331,N_5520);
nor U12405 (N_12405,N_8969,N_9353);
or U12406 (N_12406,N_5272,N_9983);
or U12407 (N_12407,N_7486,N_9469);
nor U12408 (N_12408,N_9220,N_9858);
and U12409 (N_12409,N_5729,N_6344);
xor U12410 (N_12410,N_9710,N_7442);
or U12411 (N_12411,N_6319,N_7672);
nand U12412 (N_12412,N_7573,N_8057);
xnor U12413 (N_12413,N_8297,N_5790);
or U12414 (N_12414,N_5511,N_6327);
or U12415 (N_12415,N_8461,N_9140);
or U12416 (N_12416,N_6314,N_9251);
and U12417 (N_12417,N_5841,N_5001);
and U12418 (N_12418,N_8201,N_9144);
and U12419 (N_12419,N_7791,N_6071);
or U12420 (N_12420,N_7405,N_7032);
xnor U12421 (N_12421,N_5206,N_7501);
nand U12422 (N_12422,N_6100,N_5400);
nand U12423 (N_12423,N_9793,N_6345);
nand U12424 (N_12424,N_6352,N_9115);
xnor U12425 (N_12425,N_8287,N_5502);
or U12426 (N_12426,N_6697,N_9228);
or U12427 (N_12427,N_9653,N_7313);
and U12428 (N_12428,N_6824,N_6663);
xnor U12429 (N_12429,N_6989,N_6466);
or U12430 (N_12430,N_5417,N_9349);
and U12431 (N_12431,N_9808,N_9864);
nor U12432 (N_12432,N_7114,N_5464);
xor U12433 (N_12433,N_7669,N_9667);
nor U12434 (N_12434,N_8892,N_6346);
xnor U12435 (N_12435,N_7351,N_8470);
or U12436 (N_12436,N_6098,N_9721);
and U12437 (N_12437,N_8138,N_8759);
and U12438 (N_12438,N_9849,N_5199);
nand U12439 (N_12439,N_8693,N_9960);
xnor U12440 (N_12440,N_7481,N_8769);
and U12441 (N_12441,N_6945,N_5587);
and U12442 (N_12442,N_6665,N_6916);
nand U12443 (N_12443,N_8339,N_5747);
nand U12444 (N_12444,N_5682,N_9696);
or U12445 (N_12445,N_7996,N_5195);
nand U12446 (N_12446,N_5352,N_7779);
and U12447 (N_12447,N_7590,N_9839);
and U12448 (N_12448,N_9508,N_7780);
xor U12449 (N_12449,N_8022,N_5970);
and U12450 (N_12450,N_7251,N_6190);
nor U12451 (N_12451,N_9039,N_6085);
nand U12452 (N_12452,N_9161,N_7368);
xor U12453 (N_12453,N_5409,N_6996);
xnor U12454 (N_12454,N_6924,N_9755);
or U12455 (N_12455,N_5505,N_7765);
nor U12456 (N_12456,N_5778,N_7599);
and U12457 (N_12457,N_7641,N_8471);
xnor U12458 (N_12458,N_7514,N_9013);
nor U12459 (N_12459,N_8150,N_9675);
and U12460 (N_12460,N_6990,N_9915);
nor U12461 (N_12461,N_5416,N_9467);
xnor U12462 (N_12462,N_6712,N_9761);
xnor U12463 (N_12463,N_6199,N_7374);
nand U12464 (N_12464,N_6357,N_8762);
nor U12465 (N_12465,N_5207,N_6979);
or U12466 (N_12466,N_6645,N_8787);
nor U12467 (N_12467,N_9004,N_6157);
nor U12468 (N_12468,N_6720,N_9315);
or U12469 (N_12469,N_8733,N_8785);
or U12470 (N_12470,N_7097,N_7485);
and U12471 (N_12471,N_5908,N_7562);
or U12472 (N_12472,N_8737,N_5444);
or U12473 (N_12473,N_8321,N_9738);
nand U12474 (N_12474,N_6497,N_9570);
and U12475 (N_12475,N_8349,N_7664);
and U12476 (N_12476,N_5780,N_5963);
and U12477 (N_12477,N_5157,N_5192);
and U12478 (N_12478,N_8676,N_9556);
and U12479 (N_12479,N_6032,N_7871);
xnor U12480 (N_12480,N_6734,N_8831);
and U12481 (N_12481,N_9316,N_9229);
nand U12482 (N_12482,N_6481,N_6701);
nor U12483 (N_12483,N_9779,N_9123);
nor U12484 (N_12484,N_9986,N_8221);
nor U12485 (N_12485,N_7393,N_6159);
nand U12486 (N_12486,N_7887,N_5523);
nor U12487 (N_12487,N_8747,N_7423);
nand U12488 (N_12488,N_9792,N_5137);
xor U12489 (N_12489,N_8788,N_8677);
nor U12490 (N_12490,N_6189,N_8125);
or U12491 (N_12491,N_5981,N_6369);
nor U12492 (N_12492,N_9791,N_8903);
xnor U12493 (N_12493,N_6597,N_9301);
nor U12494 (N_12494,N_7125,N_6939);
and U12495 (N_12495,N_5612,N_9333);
nor U12496 (N_12496,N_6639,N_9897);
nand U12497 (N_12497,N_9044,N_5647);
nor U12498 (N_12498,N_9178,N_7416);
or U12499 (N_12499,N_8983,N_8707);
and U12500 (N_12500,N_6489,N_5497);
or U12501 (N_12501,N_5888,N_8827);
nand U12502 (N_12502,N_7731,N_7072);
nor U12503 (N_12503,N_5553,N_5521);
and U12504 (N_12504,N_8426,N_6680);
nand U12505 (N_12505,N_9193,N_9148);
nand U12506 (N_12506,N_6590,N_8360);
nand U12507 (N_12507,N_7063,N_6526);
or U12508 (N_12508,N_8098,N_7258);
nand U12509 (N_12509,N_6274,N_6022);
or U12510 (N_12510,N_9311,N_8873);
xor U12511 (N_12511,N_7902,N_6761);
xor U12512 (N_12512,N_5694,N_7976);
nand U12513 (N_12513,N_6246,N_5777);
xnor U12514 (N_12514,N_6815,N_5579);
nand U12515 (N_12515,N_7217,N_7487);
and U12516 (N_12516,N_8512,N_6494);
or U12517 (N_12517,N_6237,N_8567);
and U12518 (N_12518,N_8797,N_9861);
and U12519 (N_12519,N_5151,N_6071);
nor U12520 (N_12520,N_7828,N_6984);
xor U12521 (N_12521,N_6907,N_9114);
and U12522 (N_12522,N_7335,N_7500);
or U12523 (N_12523,N_6363,N_8672);
xnor U12524 (N_12524,N_8438,N_9742);
xnor U12525 (N_12525,N_6405,N_6810);
xor U12526 (N_12526,N_7207,N_8911);
nor U12527 (N_12527,N_7245,N_9816);
and U12528 (N_12528,N_7823,N_7245);
and U12529 (N_12529,N_5234,N_6310);
nor U12530 (N_12530,N_8363,N_9508);
xor U12531 (N_12531,N_6670,N_8699);
and U12532 (N_12532,N_5523,N_7270);
nor U12533 (N_12533,N_9404,N_6235);
xor U12534 (N_12534,N_5869,N_7857);
and U12535 (N_12535,N_7657,N_6600);
nor U12536 (N_12536,N_9472,N_9614);
nor U12537 (N_12537,N_5505,N_5449);
nand U12538 (N_12538,N_6074,N_7596);
or U12539 (N_12539,N_6408,N_9085);
or U12540 (N_12540,N_5016,N_7585);
or U12541 (N_12541,N_5866,N_6098);
nor U12542 (N_12542,N_9132,N_7154);
nor U12543 (N_12543,N_8617,N_7988);
nor U12544 (N_12544,N_7797,N_7785);
and U12545 (N_12545,N_9067,N_8573);
xnor U12546 (N_12546,N_8500,N_6954);
xnor U12547 (N_12547,N_8769,N_9189);
xor U12548 (N_12548,N_6979,N_9947);
or U12549 (N_12549,N_8824,N_6572);
and U12550 (N_12550,N_5966,N_8905);
and U12551 (N_12551,N_9982,N_7209);
and U12552 (N_12552,N_5889,N_9780);
or U12553 (N_12553,N_8185,N_6791);
xnor U12554 (N_12554,N_7372,N_8910);
nor U12555 (N_12555,N_8590,N_5857);
nor U12556 (N_12556,N_7896,N_9282);
nor U12557 (N_12557,N_9652,N_9211);
nor U12558 (N_12558,N_8478,N_9764);
nand U12559 (N_12559,N_7572,N_9704);
nor U12560 (N_12560,N_7052,N_8250);
nor U12561 (N_12561,N_7083,N_8456);
or U12562 (N_12562,N_9295,N_6468);
xor U12563 (N_12563,N_6755,N_7121);
or U12564 (N_12564,N_6170,N_9725);
or U12565 (N_12565,N_6461,N_6569);
or U12566 (N_12566,N_7971,N_8032);
xor U12567 (N_12567,N_7043,N_9296);
nand U12568 (N_12568,N_9212,N_5144);
nand U12569 (N_12569,N_7023,N_8601);
xnor U12570 (N_12570,N_9421,N_6234);
nor U12571 (N_12571,N_5543,N_6995);
nand U12572 (N_12572,N_5541,N_9947);
nand U12573 (N_12573,N_6713,N_9787);
or U12574 (N_12574,N_8161,N_6685);
nand U12575 (N_12575,N_7589,N_5315);
nor U12576 (N_12576,N_9356,N_6570);
and U12577 (N_12577,N_8481,N_5091);
nand U12578 (N_12578,N_5775,N_7254);
nor U12579 (N_12579,N_7841,N_8573);
xnor U12580 (N_12580,N_9302,N_6156);
nor U12581 (N_12581,N_6157,N_8372);
nor U12582 (N_12582,N_8923,N_9433);
or U12583 (N_12583,N_6747,N_6298);
or U12584 (N_12584,N_6010,N_9397);
nor U12585 (N_12585,N_9908,N_6763);
and U12586 (N_12586,N_5951,N_8209);
or U12587 (N_12587,N_9893,N_8836);
or U12588 (N_12588,N_6721,N_9965);
xnor U12589 (N_12589,N_5960,N_7801);
or U12590 (N_12590,N_7103,N_5556);
nand U12591 (N_12591,N_6999,N_5381);
nor U12592 (N_12592,N_5335,N_9923);
xor U12593 (N_12593,N_9819,N_8084);
and U12594 (N_12594,N_7307,N_7197);
and U12595 (N_12595,N_5134,N_8231);
nand U12596 (N_12596,N_6582,N_5527);
or U12597 (N_12597,N_5984,N_7495);
or U12598 (N_12598,N_9092,N_8014);
or U12599 (N_12599,N_5275,N_8591);
nor U12600 (N_12600,N_8071,N_7430);
or U12601 (N_12601,N_6847,N_7802);
nor U12602 (N_12602,N_5954,N_5511);
or U12603 (N_12603,N_8817,N_7540);
nand U12604 (N_12604,N_6271,N_9945);
xor U12605 (N_12605,N_8845,N_9924);
or U12606 (N_12606,N_9377,N_9235);
nor U12607 (N_12607,N_6524,N_7723);
nor U12608 (N_12608,N_7383,N_5449);
nor U12609 (N_12609,N_7530,N_5446);
nor U12610 (N_12610,N_7061,N_6043);
xor U12611 (N_12611,N_5307,N_5830);
and U12612 (N_12612,N_5730,N_9311);
xor U12613 (N_12613,N_6230,N_7379);
nand U12614 (N_12614,N_9329,N_6961);
nor U12615 (N_12615,N_5490,N_8244);
or U12616 (N_12616,N_6677,N_9099);
or U12617 (N_12617,N_8480,N_7543);
or U12618 (N_12618,N_9036,N_6467);
or U12619 (N_12619,N_8990,N_9912);
xor U12620 (N_12620,N_7511,N_8222);
xor U12621 (N_12621,N_6273,N_6570);
nand U12622 (N_12622,N_6252,N_8532);
and U12623 (N_12623,N_7131,N_5492);
xnor U12624 (N_12624,N_9274,N_9521);
or U12625 (N_12625,N_5302,N_5591);
xor U12626 (N_12626,N_7944,N_8143);
nor U12627 (N_12627,N_5866,N_6515);
nor U12628 (N_12628,N_6157,N_9965);
and U12629 (N_12629,N_7534,N_5440);
nand U12630 (N_12630,N_6220,N_6837);
and U12631 (N_12631,N_5952,N_6805);
nand U12632 (N_12632,N_9625,N_6904);
nand U12633 (N_12633,N_5624,N_5676);
or U12634 (N_12634,N_9517,N_7479);
nand U12635 (N_12635,N_8688,N_5694);
and U12636 (N_12636,N_7461,N_6629);
nand U12637 (N_12637,N_5687,N_9114);
nand U12638 (N_12638,N_6135,N_5014);
nand U12639 (N_12639,N_5115,N_9396);
or U12640 (N_12640,N_8121,N_7246);
or U12641 (N_12641,N_9886,N_9607);
nand U12642 (N_12642,N_7011,N_9398);
or U12643 (N_12643,N_9899,N_7900);
or U12644 (N_12644,N_9876,N_8613);
xnor U12645 (N_12645,N_5679,N_9541);
nor U12646 (N_12646,N_7826,N_5910);
and U12647 (N_12647,N_7997,N_9162);
nand U12648 (N_12648,N_7019,N_6282);
nand U12649 (N_12649,N_9499,N_5383);
nand U12650 (N_12650,N_6817,N_6021);
nand U12651 (N_12651,N_5504,N_9848);
and U12652 (N_12652,N_5221,N_8242);
nand U12653 (N_12653,N_8279,N_6440);
and U12654 (N_12654,N_8408,N_8344);
nand U12655 (N_12655,N_9934,N_7682);
and U12656 (N_12656,N_8395,N_6454);
nor U12657 (N_12657,N_7486,N_8723);
and U12658 (N_12658,N_9790,N_9947);
and U12659 (N_12659,N_7728,N_6453);
and U12660 (N_12660,N_7254,N_6870);
and U12661 (N_12661,N_8592,N_8751);
or U12662 (N_12662,N_8903,N_5191);
and U12663 (N_12663,N_7463,N_9168);
and U12664 (N_12664,N_5458,N_6007);
and U12665 (N_12665,N_5633,N_9742);
nand U12666 (N_12666,N_7382,N_9723);
or U12667 (N_12667,N_9450,N_9224);
nor U12668 (N_12668,N_6063,N_6022);
xnor U12669 (N_12669,N_6686,N_8015);
or U12670 (N_12670,N_5816,N_9799);
and U12671 (N_12671,N_5046,N_7389);
nand U12672 (N_12672,N_7767,N_7239);
nor U12673 (N_12673,N_9267,N_6753);
nor U12674 (N_12674,N_9883,N_8201);
nand U12675 (N_12675,N_7905,N_7762);
xnor U12676 (N_12676,N_7177,N_8605);
nor U12677 (N_12677,N_7419,N_5516);
nor U12678 (N_12678,N_7439,N_7021);
xnor U12679 (N_12679,N_5678,N_6633);
nand U12680 (N_12680,N_5411,N_8216);
nor U12681 (N_12681,N_8394,N_7636);
xnor U12682 (N_12682,N_7409,N_9521);
or U12683 (N_12683,N_5879,N_6285);
nor U12684 (N_12684,N_7144,N_6933);
and U12685 (N_12685,N_7562,N_9761);
nor U12686 (N_12686,N_7649,N_6402);
xor U12687 (N_12687,N_5002,N_7169);
nor U12688 (N_12688,N_6017,N_7741);
nor U12689 (N_12689,N_8890,N_7286);
or U12690 (N_12690,N_5853,N_7337);
and U12691 (N_12691,N_8464,N_7311);
xor U12692 (N_12692,N_7474,N_8115);
xnor U12693 (N_12693,N_8748,N_9713);
nand U12694 (N_12694,N_5595,N_9463);
xnor U12695 (N_12695,N_7968,N_9077);
or U12696 (N_12696,N_7015,N_5915);
nor U12697 (N_12697,N_9048,N_7975);
nand U12698 (N_12698,N_7510,N_8321);
xnor U12699 (N_12699,N_5380,N_5036);
or U12700 (N_12700,N_5755,N_6764);
nor U12701 (N_12701,N_9627,N_6751);
or U12702 (N_12702,N_7688,N_5546);
and U12703 (N_12703,N_8378,N_7912);
nor U12704 (N_12704,N_7622,N_5614);
nand U12705 (N_12705,N_6554,N_8425);
or U12706 (N_12706,N_7434,N_8744);
xnor U12707 (N_12707,N_8539,N_8479);
nor U12708 (N_12708,N_9296,N_8715);
or U12709 (N_12709,N_8975,N_8429);
nor U12710 (N_12710,N_6752,N_8999);
xnor U12711 (N_12711,N_8764,N_6838);
nor U12712 (N_12712,N_9146,N_9086);
or U12713 (N_12713,N_7767,N_6671);
xnor U12714 (N_12714,N_9833,N_8402);
and U12715 (N_12715,N_6211,N_7542);
xor U12716 (N_12716,N_9427,N_6759);
nand U12717 (N_12717,N_5568,N_6146);
or U12718 (N_12718,N_9549,N_5442);
xor U12719 (N_12719,N_6190,N_8122);
nand U12720 (N_12720,N_8507,N_6760);
or U12721 (N_12721,N_9182,N_8419);
or U12722 (N_12722,N_6695,N_6709);
and U12723 (N_12723,N_6194,N_7092);
and U12724 (N_12724,N_9387,N_8060);
xor U12725 (N_12725,N_8893,N_5151);
and U12726 (N_12726,N_6813,N_6495);
nor U12727 (N_12727,N_8048,N_5993);
xnor U12728 (N_12728,N_6223,N_7680);
nor U12729 (N_12729,N_5314,N_7123);
xnor U12730 (N_12730,N_8666,N_7256);
nand U12731 (N_12731,N_9177,N_5414);
or U12732 (N_12732,N_5151,N_9955);
or U12733 (N_12733,N_9154,N_7877);
and U12734 (N_12734,N_8543,N_5380);
nand U12735 (N_12735,N_9923,N_7148);
and U12736 (N_12736,N_9891,N_9485);
nor U12737 (N_12737,N_7059,N_7300);
or U12738 (N_12738,N_7381,N_6997);
nand U12739 (N_12739,N_8619,N_9937);
or U12740 (N_12740,N_7736,N_8284);
nand U12741 (N_12741,N_8039,N_7250);
or U12742 (N_12742,N_8824,N_9112);
xor U12743 (N_12743,N_7413,N_8917);
nor U12744 (N_12744,N_8892,N_8532);
nor U12745 (N_12745,N_6540,N_9826);
and U12746 (N_12746,N_6570,N_7056);
or U12747 (N_12747,N_5055,N_5307);
nor U12748 (N_12748,N_8030,N_5643);
nand U12749 (N_12749,N_6793,N_6498);
or U12750 (N_12750,N_5232,N_5029);
or U12751 (N_12751,N_5306,N_6264);
nor U12752 (N_12752,N_6979,N_7630);
nand U12753 (N_12753,N_7279,N_9463);
and U12754 (N_12754,N_7049,N_7640);
or U12755 (N_12755,N_5496,N_8279);
or U12756 (N_12756,N_5884,N_7843);
xor U12757 (N_12757,N_9102,N_9952);
nor U12758 (N_12758,N_9169,N_9413);
and U12759 (N_12759,N_6112,N_5085);
or U12760 (N_12760,N_7006,N_5703);
nand U12761 (N_12761,N_7150,N_5418);
or U12762 (N_12762,N_6898,N_5398);
nand U12763 (N_12763,N_8595,N_8598);
or U12764 (N_12764,N_7295,N_7748);
nand U12765 (N_12765,N_7439,N_5883);
nor U12766 (N_12766,N_9024,N_8351);
or U12767 (N_12767,N_7426,N_5852);
and U12768 (N_12768,N_8457,N_8482);
and U12769 (N_12769,N_6915,N_5570);
nand U12770 (N_12770,N_9495,N_7411);
nor U12771 (N_12771,N_9834,N_9455);
or U12772 (N_12772,N_6794,N_9265);
and U12773 (N_12773,N_5309,N_5947);
and U12774 (N_12774,N_6506,N_7967);
nand U12775 (N_12775,N_6360,N_9318);
nand U12776 (N_12776,N_8634,N_6816);
xnor U12777 (N_12777,N_5054,N_8582);
xnor U12778 (N_12778,N_5483,N_5784);
or U12779 (N_12779,N_5394,N_7062);
or U12780 (N_12780,N_5566,N_6043);
or U12781 (N_12781,N_8236,N_6771);
nand U12782 (N_12782,N_7696,N_5157);
nand U12783 (N_12783,N_6824,N_7953);
and U12784 (N_12784,N_7037,N_8350);
or U12785 (N_12785,N_6106,N_8762);
xor U12786 (N_12786,N_5167,N_8647);
nand U12787 (N_12787,N_8731,N_7386);
or U12788 (N_12788,N_9057,N_7059);
nand U12789 (N_12789,N_7927,N_6553);
xnor U12790 (N_12790,N_6857,N_7957);
and U12791 (N_12791,N_9135,N_7772);
nor U12792 (N_12792,N_8486,N_9501);
nor U12793 (N_12793,N_5485,N_7691);
nor U12794 (N_12794,N_8307,N_8455);
and U12795 (N_12795,N_6923,N_9251);
nand U12796 (N_12796,N_5098,N_5814);
nor U12797 (N_12797,N_9223,N_8101);
or U12798 (N_12798,N_9178,N_8626);
nand U12799 (N_12799,N_6911,N_6761);
xor U12800 (N_12800,N_8372,N_6386);
or U12801 (N_12801,N_6249,N_5084);
and U12802 (N_12802,N_9107,N_5322);
or U12803 (N_12803,N_7514,N_6197);
nand U12804 (N_12804,N_9246,N_9913);
and U12805 (N_12805,N_9380,N_6761);
nor U12806 (N_12806,N_5776,N_5901);
xor U12807 (N_12807,N_5038,N_8249);
xnor U12808 (N_12808,N_9610,N_5667);
nand U12809 (N_12809,N_9664,N_7566);
and U12810 (N_12810,N_6689,N_7420);
or U12811 (N_12811,N_5823,N_6280);
nand U12812 (N_12812,N_8923,N_6726);
or U12813 (N_12813,N_7799,N_8114);
or U12814 (N_12814,N_9831,N_5857);
nor U12815 (N_12815,N_8885,N_8484);
or U12816 (N_12816,N_8796,N_5137);
xnor U12817 (N_12817,N_9880,N_6098);
nand U12818 (N_12818,N_9595,N_5338);
nand U12819 (N_12819,N_8044,N_7053);
nor U12820 (N_12820,N_6361,N_5251);
nor U12821 (N_12821,N_8745,N_8518);
or U12822 (N_12822,N_6675,N_8208);
xor U12823 (N_12823,N_6279,N_5300);
and U12824 (N_12824,N_7386,N_5096);
nand U12825 (N_12825,N_5971,N_5745);
and U12826 (N_12826,N_7010,N_8972);
nor U12827 (N_12827,N_5858,N_6926);
xor U12828 (N_12828,N_8562,N_7527);
nor U12829 (N_12829,N_9353,N_7161);
nor U12830 (N_12830,N_7493,N_8998);
nand U12831 (N_12831,N_6102,N_7721);
or U12832 (N_12832,N_7631,N_9846);
or U12833 (N_12833,N_9550,N_6434);
xnor U12834 (N_12834,N_9457,N_6158);
nand U12835 (N_12835,N_8290,N_8636);
and U12836 (N_12836,N_8166,N_7695);
nor U12837 (N_12837,N_7882,N_8424);
xor U12838 (N_12838,N_9023,N_5139);
or U12839 (N_12839,N_9676,N_9079);
and U12840 (N_12840,N_5600,N_6079);
xnor U12841 (N_12841,N_9590,N_6847);
and U12842 (N_12842,N_8768,N_6025);
nor U12843 (N_12843,N_5820,N_8533);
or U12844 (N_12844,N_8495,N_9491);
nand U12845 (N_12845,N_5880,N_7731);
or U12846 (N_12846,N_7222,N_6266);
xor U12847 (N_12847,N_8536,N_9953);
or U12848 (N_12848,N_6185,N_6935);
and U12849 (N_12849,N_9417,N_5807);
nand U12850 (N_12850,N_6105,N_9002);
nor U12851 (N_12851,N_5129,N_9210);
and U12852 (N_12852,N_6476,N_7550);
xor U12853 (N_12853,N_6142,N_6370);
and U12854 (N_12854,N_8171,N_8559);
xnor U12855 (N_12855,N_5099,N_9363);
xnor U12856 (N_12856,N_7170,N_7777);
xor U12857 (N_12857,N_9500,N_8698);
xnor U12858 (N_12858,N_8540,N_5849);
and U12859 (N_12859,N_6595,N_9447);
and U12860 (N_12860,N_5512,N_6013);
xor U12861 (N_12861,N_5169,N_6981);
nand U12862 (N_12862,N_7184,N_9081);
and U12863 (N_12863,N_5041,N_9124);
nor U12864 (N_12864,N_6755,N_6790);
nor U12865 (N_12865,N_6509,N_5778);
or U12866 (N_12866,N_8227,N_6997);
or U12867 (N_12867,N_9123,N_8798);
nand U12868 (N_12868,N_7749,N_8419);
nand U12869 (N_12869,N_9288,N_6192);
and U12870 (N_12870,N_9684,N_9530);
nand U12871 (N_12871,N_6679,N_8307);
xnor U12872 (N_12872,N_5841,N_8439);
and U12873 (N_12873,N_6345,N_7852);
nor U12874 (N_12874,N_5624,N_9111);
and U12875 (N_12875,N_5461,N_7332);
and U12876 (N_12876,N_8664,N_8135);
xnor U12877 (N_12877,N_6220,N_6461);
or U12878 (N_12878,N_6355,N_5214);
or U12879 (N_12879,N_7460,N_6584);
or U12880 (N_12880,N_5558,N_9551);
and U12881 (N_12881,N_8826,N_6799);
or U12882 (N_12882,N_8104,N_8944);
nand U12883 (N_12883,N_5953,N_6299);
xor U12884 (N_12884,N_5795,N_5405);
and U12885 (N_12885,N_8954,N_8585);
and U12886 (N_12886,N_9336,N_6447);
nand U12887 (N_12887,N_6210,N_6177);
or U12888 (N_12888,N_8121,N_5513);
or U12889 (N_12889,N_6523,N_6574);
nand U12890 (N_12890,N_9859,N_8068);
nor U12891 (N_12891,N_5263,N_6709);
and U12892 (N_12892,N_9182,N_8664);
xnor U12893 (N_12893,N_5906,N_8221);
or U12894 (N_12894,N_9403,N_9706);
nor U12895 (N_12895,N_7952,N_8359);
and U12896 (N_12896,N_6244,N_6239);
or U12897 (N_12897,N_8081,N_9706);
or U12898 (N_12898,N_8375,N_9690);
nor U12899 (N_12899,N_8804,N_9738);
and U12900 (N_12900,N_5667,N_6712);
and U12901 (N_12901,N_5269,N_5080);
or U12902 (N_12902,N_9660,N_5240);
nor U12903 (N_12903,N_8671,N_7244);
xnor U12904 (N_12904,N_9796,N_8486);
and U12905 (N_12905,N_6962,N_8277);
and U12906 (N_12906,N_7302,N_9743);
and U12907 (N_12907,N_9448,N_7008);
xor U12908 (N_12908,N_6971,N_5456);
xor U12909 (N_12909,N_8440,N_8941);
nor U12910 (N_12910,N_5292,N_8378);
xnor U12911 (N_12911,N_6062,N_8479);
or U12912 (N_12912,N_7578,N_6888);
nand U12913 (N_12913,N_5929,N_9846);
or U12914 (N_12914,N_6993,N_8491);
nor U12915 (N_12915,N_9548,N_5175);
or U12916 (N_12916,N_9811,N_8012);
or U12917 (N_12917,N_8088,N_7820);
nand U12918 (N_12918,N_7964,N_8757);
and U12919 (N_12919,N_6626,N_6528);
nand U12920 (N_12920,N_9696,N_8675);
and U12921 (N_12921,N_5280,N_9299);
and U12922 (N_12922,N_9516,N_9572);
or U12923 (N_12923,N_8832,N_8188);
nand U12924 (N_12924,N_6962,N_8812);
and U12925 (N_12925,N_8810,N_9120);
nor U12926 (N_12926,N_9239,N_7482);
or U12927 (N_12927,N_8441,N_5360);
nand U12928 (N_12928,N_6213,N_9584);
nand U12929 (N_12929,N_7557,N_8985);
and U12930 (N_12930,N_7345,N_8426);
nand U12931 (N_12931,N_9081,N_8829);
xnor U12932 (N_12932,N_5962,N_6679);
or U12933 (N_12933,N_9952,N_6733);
nand U12934 (N_12934,N_7578,N_6772);
or U12935 (N_12935,N_9596,N_9434);
nand U12936 (N_12936,N_7671,N_9619);
and U12937 (N_12937,N_7638,N_6920);
or U12938 (N_12938,N_6697,N_5805);
or U12939 (N_12939,N_6117,N_7845);
or U12940 (N_12940,N_5332,N_7839);
nor U12941 (N_12941,N_7637,N_8958);
and U12942 (N_12942,N_8105,N_7903);
nand U12943 (N_12943,N_6533,N_5526);
nor U12944 (N_12944,N_6313,N_9143);
nor U12945 (N_12945,N_9501,N_5646);
xor U12946 (N_12946,N_8637,N_6830);
or U12947 (N_12947,N_5419,N_6712);
and U12948 (N_12948,N_8147,N_9998);
xor U12949 (N_12949,N_6034,N_6486);
nand U12950 (N_12950,N_5228,N_6716);
or U12951 (N_12951,N_9937,N_8219);
and U12952 (N_12952,N_8430,N_9464);
nand U12953 (N_12953,N_9964,N_7727);
or U12954 (N_12954,N_6571,N_7004);
xor U12955 (N_12955,N_7999,N_8152);
xnor U12956 (N_12956,N_5695,N_6134);
or U12957 (N_12957,N_8883,N_5583);
nor U12958 (N_12958,N_8373,N_6060);
nand U12959 (N_12959,N_9969,N_7931);
or U12960 (N_12960,N_5084,N_6921);
xnor U12961 (N_12961,N_6385,N_7307);
nand U12962 (N_12962,N_8019,N_7879);
nor U12963 (N_12963,N_6322,N_5135);
and U12964 (N_12964,N_6203,N_6123);
xor U12965 (N_12965,N_6622,N_8379);
nor U12966 (N_12966,N_5624,N_6216);
nor U12967 (N_12967,N_5854,N_5271);
nor U12968 (N_12968,N_6002,N_8119);
or U12969 (N_12969,N_5527,N_7448);
nand U12970 (N_12970,N_7311,N_6920);
xnor U12971 (N_12971,N_7382,N_6452);
nor U12972 (N_12972,N_9792,N_8097);
nor U12973 (N_12973,N_9531,N_9566);
or U12974 (N_12974,N_9006,N_6858);
xnor U12975 (N_12975,N_7881,N_5880);
and U12976 (N_12976,N_6902,N_5957);
nor U12977 (N_12977,N_8549,N_9650);
nor U12978 (N_12978,N_8690,N_6732);
nor U12979 (N_12979,N_8172,N_9710);
nor U12980 (N_12980,N_7392,N_6070);
xor U12981 (N_12981,N_9352,N_5740);
or U12982 (N_12982,N_8796,N_9562);
xnor U12983 (N_12983,N_7253,N_9458);
nand U12984 (N_12984,N_5656,N_8349);
nand U12985 (N_12985,N_8967,N_7597);
nand U12986 (N_12986,N_8220,N_9296);
nand U12987 (N_12987,N_7417,N_7361);
and U12988 (N_12988,N_7917,N_5004);
and U12989 (N_12989,N_6978,N_5799);
xnor U12990 (N_12990,N_6334,N_5409);
xnor U12991 (N_12991,N_8722,N_9507);
nand U12992 (N_12992,N_6485,N_6376);
nand U12993 (N_12993,N_8836,N_6388);
nor U12994 (N_12994,N_8961,N_8013);
nand U12995 (N_12995,N_9210,N_8398);
nand U12996 (N_12996,N_8022,N_9088);
nor U12997 (N_12997,N_6996,N_7328);
nand U12998 (N_12998,N_8110,N_7721);
and U12999 (N_12999,N_9543,N_8250);
xor U13000 (N_13000,N_5113,N_8111);
or U13001 (N_13001,N_9267,N_6881);
and U13002 (N_13002,N_5815,N_5210);
nand U13003 (N_13003,N_6159,N_8157);
nor U13004 (N_13004,N_5924,N_8501);
nand U13005 (N_13005,N_5688,N_5192);
or U13006 (N_13006,N_6121,N_6378);
nand U13007 (N_13007,N_8649,N_7103);
and U13008 (N_13008,N_5177,N_5348);
xnor U13009 (N_13009,N_6561,N_7227);
xnor U13010 (N_13010,N_9196,N_8999);
and U13011 (N_13011,N_8657,N_6915);
nand U13012 (N_13012,N_9598,N_7023);
nand U13013 (N_13013,N_6902,N_9952);
nand U13014 (N_13014,N_6033,N_6105);
nor U13015 (N_13015,N_7359,N_6397);
nand U13016 (N_13016,N_8047,N_6238);
nor U13017 (N_13017,N_8507,N_5226);
xnor U13018 (N_13018,N_5109,N_7121);
xor U13019 (N_13019,N_7619,N_7145);
nor U13020 (N_13020,N_5256,N_9022);
or U13021 (N_13021,N_8249,N_9923);
xor U13022 (N_13022,N_9567,N_6899);
xnor U13023 (N_13023,N_8881,N_9077);
or U13024 (N_13024,N_7042,N_5517);
nand U13025 (N_13025,N_8560,N_8202);
nand U13026 (N_13026,N_9798,N_5815);
nor U13027 (N_13027,N_9166,N_9362);
nand U13028 (N_13028,N_8235,N_7616);
and U13029 (N_13029,N_5944,N_9512);
or U13030 (N_13030,N_7484,N_5653);
or U13031 (N_13031,N_6695,N_8945);
and U13032 (N_13032,N_9688,N_6422);
and U13033 (N_13033,N_8649,N_5537);
xor U13034 (N_13034,N_5208,N_8349);
nor U13035 (N_13035,N_9096,N_6963);
and U13036 (N_13036,N_6149,N_8187);
xor U13037 (N_13037,N_6421,N_9205);
and U13038 (N_13038,N_8639,N_7204);
nand U13039 (N_13039,N_9554,N_6641);
or U13040 (N_13040,N_7394,N_7928);
nand U13041 (N_13041,N_6995,N_8285);
nor U13042 (N_13042,N_9396,N_5231);
xnor U13043 (N_13043,N_9698,N_6439);
xor U13044 (N_13044,N_9916,N_6160);
and U13045 (N_13045,N_9533,N_5556);
nand U13046 (N_13046,N_6083,N_7736);
and U13047 (N_13047,N_8039,N_6777);
and U13048 (N_13048,N_7301,N_9299);
xor U13049 (N_13049,N_7648,N_6074);
and U13050 (N_13050,N_5352,N_6028);
and U13051 (N_13051,N_5522,N_8215);
nand U13052 (N_13052,N_7749,N_8048);
and U13053 (N_13053,N_5690,N_8014);
nor U13054 (N_13054,N_7261,N_6245);
or U13055 (N_13055,N_6007,N_9594);
and U13056 (N_13056,N_8539,N_5399);
or U13057 (N_13057,N_7366,N_9828);
or U13058 (N_13058,N_6586,N_5449);
xor U13059 (N_13059,N_5824,N_9029);
nor U13060 (N_13060,N_6703,N_6383);
nor U13061 (N_13061,N_9223,N_9977);
or U13062 (N_13062,N_6388,N_7016);
nand U13063 (N_13063,N_7738,N_9974);
and U13064 (N_13064,N_7628,N_6728);
nand U13065 (N_13065,N_9197,N_8697);
or U13066 (N_13066,N_6492,N_7308);
or U13067 (N_13067,N_9950,N_5066);
or U13068 (N_13068,N_6257,N_9116);
nor U13069 (N_13069,N_8977,N_6316);
nor U13070 (N_13070,N_6668,N_9077);
nor U13071 (N_13071,N_7702,N_6266);
and U13072 (N_13072,N_6180,N_7149);
xor U13073 (N_13073,N_5651,N_8407);
nand U13074 (N_13074,N_9729,N_8058);
or U13075 (N_13075,N_8645,N_9699);
and U13076 (N_13076,N_8607,N_8688);
nor U13077 (N_13077,N_8304,N_7976);
xnor U13078 (N_13078,N_7518,N_9202);
nand U13079 (N_13079,N_6857,N_7088);
nor U13080 (N_13080,N_5320,N_5326);
or U13081 (N_13081,N_7713,N_7282);
or U13082 (N_13082,N_6787,N_8559);
xnor U13083 (N_13083,N_7366,N_8153);
nand U13084 (N_13084,N_9566,N_5093);
or U13085 (N_13085,N_9051,N_5107);
xor U13086 (N_13086,N_7600,N_9830);
nand U13087 (N_13087,N_9517,N_9170);
and U13088 (N_13088,N_7443,N_8647);
nor U13089 (N_13089,N_8557,N_9114);
xnor U13090 (N_13090,N_6817,N_9370);
xor U13091 (N_13091,N_7523,N_8914);
nor U13092 (N_13092,N_6211,N_9789);
xnor U13093 (N_13093,N_6969,N_7824);
xor U13094 (N_13094,N_9408,N_9286);
xnor U13095 (N_13095,N_9594,N_8050);
or U13096 (N_13096,N_9356,N_8403);
nor U13097 (N_13097,N_9276,N_6154);
or U13098 (N_13098,N_6651,N_8952);
nor U13099 (N_13099,N_7535,N_6222);
xor U13100 (N_13100,N_5825,N_6238);
xor U13101 (N_13101,N_9371,N_8849);
nor U13102 (N_13102,N_8809,N_6154);
nand U13103 (N_13103,N_7782,N_6323);
or U13104 (N_13104,N_9906,N_6334);
or U13105 (N_13105,N_8737,N_9025);
nor U13106 (N_13106,N_9609,N_6038);
or U13107 (N_13107,N_7114,N_5907);
nand U13108 (N_13108,N_9266,N_6879);
xor U13109 (N_13109,N_5899,N_9958);
and U13110 (N_13110,N_5119,N_6030);
nand U13111 (N_13111,N_7095,N_5210);
nand U13112 (N_13112,N_9025,N_8909);
and U13113 (N_13113,N_5545,N_7561);
nor U13114 (N_13114,N_5696,N_6572);
xor U13115 (N_13115,N_9291,N_8654);
nor U13116 (N_13116,N_7411,N_7936);
xor U13117 (N_13117,N_8629,N_7107);
nand U13118 (N_13118,N_5899,N_5756);
and U13119 (N_13119,N_8737,N_9919);
xnor U13120 (N_13120,N_5074,N_6630);
or U13121 (N_13121,N_8656,N_6144);
xnor U13122 (N_13122,N_8250,N_9442);
nor U13123 (N_13123,N_9584,N_9365);
nor U13124 (N_13124,N_9208,N_9376);
or U13125 (N_13125,N_7629,N_9627);
xor U13126 (N_13126,N_6001,N_8457);
nor U13127 (N_13127,N_5785,N_7227);
nand U13128 (N_13128,N_8481,N_8066);
and U13129 (N_13129,N_8960,N_6424);
xor U13130 (N_13130,N_6905,N_9053);
xnor U13131 (N_13131,N_6022,N_7516);
nor U13132 (N_13132,N_6424,N_9748);
and U13133 (N_13133,N_5731,N_7401);
nand U13134 (N_13134,N_9249,N_5793);
nor U13135 (N_13135,N_9881,N_6860);
xor U13136 (N_13136,N_5749,N_5364);
and U13137 (N_13137,N_7577,N_6393);
and U13138 (N_13138,N_7578,N_5469);
or U13139 (N_13139,N_8983,N_7313);
xor U13140 (N_13140,N_5901,N_6971);
and U13141 (N_13141,N_8896,N_9611);
or U13142 (N_13142,N_7452,N_8489);
or U13143 (N_13143,N_6175,N_7546);
or U13144 (N_13144,N_9140,N_9287);
nand U13145 (N_13145,N_5494,N_6535);
and U13146 (N_13146,N_8047,N_6439);
nor U13147 (N_13147,N_7111,N_9918);
nand U13148 (N_13148,N_8026,N_7593);
and U13149 (N_13149,N_5607,N_7757);
nand U13150 (N_13150,N_6313,N_9202);
nand U13151 (N_13151,N_6699,N_5432);
or U13152 (N_13152,N_9024,N_9456);
or U13153 (N_13153,N_7106,N_9448);
xor U13154 (N_13154,N_8452,N_8206);
xnor U13155 (N_13155,N_7189,N_5671);
xor U13156 (N_13156,N_5786,N_9947);
nand U13157 (N_13157,N_6727,N_9849);
and U13158 (N_13158,N_6332,N_8448);
and U13159 (N_13159,N_9632,N_5459);
nand U13160 (N_13160,N_7261,N_8500);
nand U13161 (N_13161,N_7897,N_8907);
or U13162 (N_13162,N_6083,N_8611);
and U13163 (N_13163,N_5849,N_8665);
xnor U13164 (N_13164,N_7293,N_7049);
and U13165 (N_13165,N_8610,N_6095);
or U13166 (N_13166,N_7318,N_7193);
nor U13167 (N_13167,N_5461,N_6047);
nor U13168 (N_13168,N_8895,N_7256);
and U13169 (N_13169,N_5341,N_6924);
xor U13170 (N_13170,N_7347,N_5343);
or U13171 (N_13171,N_9512,N_6961);
or U13172 (N_13172,N_7116,N_7876);
nor U13173 (N_13173,N_5077,N_7305);
and U13174 (N_13174,N_9747,N_6427);
or U13175 (N_13175,N_7207,N_7435);
and U13176 (N_13176,N_9763,N_9141);
or U13177 (N_13177,N_9226,N_6943);
nand U13178 (N_13178,N_8171,N_5401);
and U13179 (N_13179,N_6391,N_9590);
xnor U13180 (N_13180,N_8878,N_6687);
xnor U13181 (N_13181,N_7602,N_9694);
xnor U13182 (N_13182,N_9038,N_6547);
nand U13183 (N_13183,N_6351,N_8115);
or U13184 (N_13184,N_8030,N_5124);
xor U13185 (N_13185,N_7503,N_9505);
nor U13186 (N_13186,N_8726,N_8340);
xnor U13187 (N_13187,N_6145,N_5835);
xor U13188 (N_13188,N_8561,N_5915);
xor U13189 (N_13189,N_9973,N_5718);
xnor U13190 (N_13190,N_7585,N_8707);
nand U13191 (N_13191,N_7474,N_9807);
nor U13192 (N_13192,N_7906,N_7095);
nor U13193 (N_13193,N_6879,N_7702);
xnor U13194 (N_13194,N_6191,N_9372);
nand U13195 (N_13195,N_8462,N_6852);
and U13196 (N_13196,N_8965,N_7279);
or U13197 (N_13197,N_6210,N_7655);
nor U13198 (N_13198,N_6901,N_5743);
and U13199 (N_13199,N_7098,N_7348);
nand U13200 (N_13200,N_9427,N_6894);
and U13201 (N_13201,N_6847,N_6336);
nand U13202 (N_13202,N_5177,N_7289);
nor U13203 (N_13203,N_8063,N_7260);
nor U13204 (N_13204,N_5475,N_6907);
nand U13205 (N_13205,N_6765,N_6537);
nand U13206 (N_13206,N_6425,N_7955);
and U13207 (N_13207,N_6936,N_5783);
and U13208 (N_13208,N_5233,N_7867);
xnor U13209 (N_13209,N_9791,N_9417);
or U13210 (N_13210,N_7865,N_5695);
xor U13211 (N_13211,N_7846,N_7301);
nor U13212 (N_13212,N_5598,N_7773);
nand U13213 (N_13213,N_8231,N_9545);
xnor U13214 (N_13214,N_7260,N_7042);
xnor U13215 (N_13215,N_5369,N_7487);
nand U13216 (N_13216,N_5047,N_8795);
xnor U13217 (N_13217,N_5981,N_7176);
nor U13218 (N_13218,N_8485,N_5023);
xor U13219 (N_13219,N_9302,N_7860);
or U13220 (N_13220,N_6794,N_6464);
xor U13221 (N_13221,N_9632,N_8867);
nor U13222 (N_13222,N_7052,N_5439);
and U13223 (N_13223,N_7696,N_6636);
or U13224 (N_13224,N_5660,N_5070);
and U13225 (N_13225,N_7024,N_7655);
and U13226 (N_13226,N_6815,N_9255);
or U13227 (N_13227,N_7022,N_9078);
nor U13228 (N_13228,N_7738,N_7515);
or U13229 (N_13229,N_6178,N_7237);
and U13230 (N_13230,N_6099,N_8092);
nand U13231 (N_13231,N_5610,N_8080);
nor U13232 (N_13232,N_7598,N_8603);
nor U13233 (N_13233,N_9227,N_8188);
and U13234 (N_13234,N_5356,N_8084);
and U13235 (N_13235,N_8975,N_9915);
or U13236 (N_13236,N_9372,N_7278);
or U13237 (N_13237,N_9465,N_8136);
or U13238 (N_13238,N_8736,N_9250);
xnor U13239 (N_13239,N_6243,N_6853);
or U13240 (N_13240,N_9202,N_7159);
or U13241 (N_13241,N_6624,N_6051);
nand U13242 (N_13242,N_5574,N_9035);
xnor U13243 (N_13243,N_9342,N_5247);
nor U13244 (N_13244,N_7379,N_9562);
xnor U13245 (N_13245,N_9573,N_6309);
or U13246 (N_13246,N_6056,N_7844);
nand U13247 (N_13247,N_7216,N_9809);
nand U13248 (N_13248,N_9274,N_6304);
nor U13249 (N_13249,N_5140,N_8172);
or U13250 (N_13250,N_5828,N_9526);
xor U13251 (N_13251,N_5845,N_8598);
nor U13252 (N_13252,N_7008,N_5745);
and U13253 (N_13253,N_6816,N_9321);
or U13254 (N_13254,N_9372,N_9846);
xnor U13255 (N_13255,N_7486,N_8745);
xor U13256 (N_13256,N_9375,N_7120);
nand U13257 (N_13257,N_8947,N_5416);
and U13258 (N_13258,N_8697,N_7152);
nand U13259 (N_13259,N_6416,N_6927);
nor U13260 (N_13260,N_6988,N_6172);
xor U13261 (N_13261,N_8235,N_5831);
nor U13262 (N_13262,N_7595,N_7239);
nand U13263 (N_13263,N_8883,N_7978);
xnor U13264 (N_13264,N_7935,N_6977);
xor U13265 (N_13265,N_8911,N_6298);
and U13266 (N_13266,N_8524,N_9894);
and U13267 (N_13267,N_7181,N_8886);
xnor U13268 (N_13268,N_6830,N_5428);
nor U13269 (N_13269,N_5408,N_6303);
xnor U13270 (N_13270,N_9132,N_7175);
and U13271 (N_13271,N_5072,N_7071);
xnor U13272 (N_13272,N_7774,N_8309);
or U13273 (N_13273,N_7774,N_5071);
nand U13274 (N_13274,N_5024,N_6542);
xor U13275 (N_13275,N_8506,N_8499);
nand U13276 (N_13276,N_9369,N_5630);
and U13277 (N_13277,N_6586,N_9528);
nor U13278 (N_13278,N_5219,N_5889);
nor U13279 (N_13279,N_9894,N_8171);
xnor U13280 (N_13280,N_6042,N_6626);
or U13281 (N_13281,N_9485,N_6437);
or U13282 (N_13282,N_9723,N_9267);
xnor U13283 (N_13283,N_6912,N_6446);
nand U13284 (N_13284,N_6274,N_8576);
xor U13285 (N_13285,N_7310,N_8595);
nand U13286 (N_13286,N_5807,N_6136);
nand U13287 (N_13287,N_9090,N_6843);
nand U13288 (N_13288,N_8343,N_7193);
or U13289 (N_13289,N_5144,N_6602);
nand U13290 (N_13290,N_6382,N_9025);
or U13291 (N_13291,N_6329,N_7118);
xnor U13292 (N_13292,N_9188,N_6427);
and U13293 (N_13293,N_9075,N_8457);
nand U13294 (N_13294,N_8743,N_5132);
nand U13295 (N_13295,N_8552,N_9517);
or U13296 (N_13296,N_5451,N_9293);
xor U13297 (N_13297,N_9727,N_5723);
nor U13298 (N_13298,N_6799,N_5612);
xor U13299 (N_13299,N_7399,N_7515);
xnor U13300 (N_13300,N_9774,N_6454);
and U13301 (N_13301,N_7280,N_6628);
xor U13302 (N_13302,N_5197,N_5678);
and U13303 (N_13303,N_8287,N_5610);
nand U13304 (N_13304,N_6355,N_5930);
nor U13305 (N_13305,N_6138,N_5673);
or U13306 (N_13306,N_7847,N_8021);
or U13307 (N_13307,N_8808,N_9002);
and U13308 (N_13308,N_8465,N_7383);
and U13309 (N_13309,N_9526,N_5506);
and U13310 (N_13310,N_9285,N_6883);
or U13311 (N_13311,N_9758,N_6873);
xor U13312 (N_13312,N_9888,N_7542);
nand U13313 (N_13313,N_9937,N_8171);
and U13314 (N_13314,N_6882,N_6098);
and U13315 (N_13315,N_7756,N_6590);
nor U13316 (N_13316,N_7639,N_8423);
or U13317 (N_13317,N_5646,N_6155);
xor U13318 (N_13318,N_6098,N_6401);
and U13319 (N_13319,N_5653,N_8117);
xnor U13320 (N_13320,N_9633,N_6722);
and U13321 (N_13321,N_5133,N_5220);
and U13322 (N_13322,N_7944,N_8177);
nand U13323 (N_13323,N_8834,N_5429);
or U13324 (N_13324,N_8965,N_9058);
and U13325 (N_13325,N_5137,N_6929);
xnor U13326 (N_13326,N_5612,N_7417);
nand U13327 (N_13327,N_6875,N_6119);
and U13328 (N_13328,N_6627,N_6223);
or U13329 (N_13329,N_7243,N_6103);
nand U13330 (N_13330,N_8245,N_6297);
nor U13331 (N_13331,N_9931,N_7624);
nand U13332 (N_13332,N_6143,N_9766);
xnor U13333 (N_13333,N_9507,N_6913);
nor U13334 (N_13334,N_7794,N_7315);
and U13335 (N_13335,N_5718,N_9036);
and U13336 (N_13336,N_6987,N_5650);
xor U13337 (N_13337,N_8674,N_7725);
xor U13338 (N_13338,N_6746,N_5445);
xnor U13339 (N_13339,N_7147,N_7486);
or U13340 (N_13340,N_7043,N_8409);
and U13341 (N_13341,N_6869,N_8284);
xnor U13342 (N_13342,N_8241,N_7923);
nor U13343 (N_13343,N_5356,N_6033);
nor U13344 (N_13344,N_6707,N_8952);
or U13345 (N_13345,N_9752,N_8260);
and U13346 (N_13346,N_9545,N_6249);
or U13347 (N_13347,N_9692,N_8396);
or U13348 (N_13348,N_8768,N_8172);
or U13349 (N_13349,N_9713,N_7022);
and U13350 (N_13350,N_9284,N_9930);
xnor U13351 (N_13351,N_9774,N_7402);
and U13352 (N_13352,N_8988,N_9107);
or U13353 (N_13353,N_5546,N_7885);
and U13354 (N_13354,N_8075,N_6236);
nor U13355 (N_13355,N_5789,N_6861);
or U13356 (N_13356,N_7253,N_8165);
nand U13357 (N_13357,N_8279,N_5986);
xnor U13358 (N_13358,N_7101,N_9251);
or U13359 (N_13359,N_5820,N_7339);
and U13360 (N_13360,N_7152,N_8587);
or U13361 (N_13361,N_9500,N_5592);
and U13362 (N_13362,N_6544,N_8359);
and U13363 (N_13363,N_7048,N_6492);
nor U13364 (N_13364,N_6203,N_9310);
nand U13365 (N_13365,N_7382,N_6227);
nand U13366 (N_13366,N_9366,N_8028);
or U13367 (N_13367,N_9960,N_7103);
nand U13368 (N_13368,N_5862,N_6479);
and U13369 (N_13369,N_6272,N_9852);
nand U13370 (N_13370,N_9218,N_7720);
xor U13371 (N_13371,N_8134,N_9813);
xor U13372 (N_13372,N_9275,N_9031);
and U13373 (N_13373,N_9426,N_9847);
or U13374 (N_13374,N_6558,N_8685);
and U13375 (N_13375,N_9321,N_9225);
xnor U13376 (N_13376,N_7501,N_7955);
nand U13377 (N_13377,N_5517,N_7129);
or U13378 (N_13378,N_8337,N_6630);
nand U13379 (N_13379,N_8725,N_8684);
and U13380 (N_13380,N_7086,N_8340);
or U13381 (N_13381,N_9534,N_9421);
nand U13382 (N_13382,N_5973,N_7394);
or U13383 (N_13383,N_5516,N_6734);
and U13384 (N_13384,N_5418,N_6415);
nand U13385 (N_13385,N_6587,N_8881);
xnor U13386 (N_13386,N_8890,N_8174);
and U13387 (N_13387,N_6475,N_7460);
nand U13388 (N_13388,N_9528,N_8025);
or U13389 (N_13389,N_6595,N_6323);
or U13390 (N_13390,N_7644,N_7384);
or U13391 (N_13391,N_7508,N_9254);
or U13392 (N_13392,N_7020,N_9367);
xnor U13393 (N_13393,N_8088,N_5506);
xor U13394 (N_13394,N_9779,N_8374);
nand U13395 (N_13395,N_6991,N_6474);
nand U13396 (N_13396,N_7317,N_8324);
xor U13397 (N_13397,N_9026,N_7856);
nor U13398 (N_13398,N_5470,N_5946);
nand U13399 (N_13399,N_5015,N_9107);
nand U13400 (N_13400,N_8036,N_7734);
or U13401 (N_13401,N_9187,N_6588);
or U13402 (N_13402,N_7133,N_5379);
nor U13403 (N_13403,N_7552,N_8921);
nor U13404 (N_13404,N_8667,N_8317);
and U13405 (N_13405,N_8784,N_7290);
nand U13406 (N_13406,N_5807,N_8864);
or U13407 (N_13407,N_5927,N_8064);
nand U13408 (N_13408,N_9331,N_9429);
or U13409 (N_13409,N_5540,N_7645);
nor U13410 (N_13410,N_6465,N_5385);
and U13411 (N_13411,N_8370,N_8218);
nor U13412 (N_13412,N_5872,N_5566);
nand U13413 (N_13413,N_6974,N_7712);
and U13414 (N_13414,N_9045,N_9387);
or U13415 (N_13415,N_7931,N_5627);
nand U13416 (N_13416,N_5187,N_7942);
nor U13417 (N_13417,N_9342,N_6332);
and U13418 (N_13418,N_9029,N_8382);
nand U13419 (N_13419,N_9006,N_9338);
or U13420 (N_13420,N_7162,N_5565);
nor U13421 (N_13421,N_5812,N_6590);
nand U13422 (N_13422,N_6842,N_9584);
xnor U13423 (N_13423,N_5671,N_9496);
nor U13424 (N_13424,N_5178,N_7588);
or U13425 (N_13425,N_5323,N_8085);
nor U13426 (N_13426,N_8879,N_9995);
nand U13427 (N_13427,N_7191,N_7958);
nor U13428 (N_13428,N_9086,N_7500);
nor U13429 (N_13429,N_5979,N_9172);
or U13430 (N_13430,N_6471,N_6067);
nor U13431 (N_13431,N_5437,N_7500);
nor U13432 (N_13432,N_6985,N_8359);
nand U13433 (N_13433,N_8692,N_6486);
nor U13434 (N_13434,N_9762,N_5585);
or U13435 (N_13435,N_8108,N_9410);
or U13436 (N_13436,N_8943,N_9755);
nand U13437 (N_13437,N_8797,N_7314);
xnor U13438 (N_13438,N_9716,N_7868);
nand U13439 (N_13439,N_8185,N_7928);
nand U13440 (N_13440,N_7729,N_7578);
or U13441 (N_13441,N_8921,N_9892);
xnor U13442 (N_13442,N_5506,N_9935);
and U13443 (N_13443,N_7197,N_8179);
xnor U13444 (N_13444,N_9867,N_9427);
and U13445 (N_13445,N_5845,N_9323);
nand U13446 (N_13446,N_7611,N_5985);
nor U13447 (N_13447,N_6601,N_7162);
nand U13448 (N_13448,N_8026,N_9987);
and U13449 (N_13449,N_7723,N_7043);
nor U13450 (N_13450,N_5651,N_9253);
nand U13451 (N_13451,N_5346,N_9697);
nand U13452 (N_13452,N_5680,N_8110);
xnor U13453 (N_13453,N_6924,N_6978);
and U13454 (N_13454,N_7952,N_7161);
nand U13455 (N_13455,N_7087,N_7109);
or U13456 (N_13456,N_7060,N_6181);
nand U13457 (N_13457,N_9993,N_6105);
or U13458 (N_13458,N_9952,N_5951);
or U13459 (N_13459,N_6991,N_9554);
or U13460 (N_13460,N_9982,N_8969);
and U13461 (N_13461,N_7653,N_8585);
or U13462 (N_13462,N_8204,N_7032);
or U13463 (N_13463,N_5485,N_6918);
nor U13464 (N_13464,N_9564,N_5809);
nand U13465 (N_13465,N_8169,N_6744);
or U13466 (N_13466,N_6034,N_8776);
nand U13467 (N_13467,N_9593,N_5036);
nor U13468 (N_13468,N_6821,N_7653);
or U13469 (N_13469,N_5333,N_5891);
nor U13470 (N_13470,N_5379,N_9949);
xor U13471 (N_13471,N_6119,N_8721);
or U13472 (N_13472,N_7229,N_6656);
and U13473 (N_13473,N_8744,N_8958);
or U13474 (N_13474,N_6764,N_5001);
or U13475 (N_13475,N_9506,N_8802);
nor U13476 (N_13476,N_8465,N_7862);
nor U13477 (N_13477,N_8833,N_6175);
nor U13478 (N_13478,N_6645,N_9190);
nor U13479 (N_13479,N_7034,N_7889);
nor U13480 (N_13480,N_9403,N_5477);
xnor U13481 (N_13481,N_6344,N_9244);
nand U13482 (N_13482,N_5061,N_8382);
and U13483 (N_13483,N_9476,N_8695);
and U13484 (N_13484,N_7230,N_8077);
nor U13485 (N_13485,N_7813,N_8713);
xnor U13486 (N_13486,N_9069,N_8751);
xor U13487 (N_13487,N_8237,N_7346);
and U13488 (N_13488,N_7847,N_5479);
and U13489 (N_13489,N_7621,N_5542);
or U13490 (N_13490,N_7225,N_8544);
and U13491 (N_13491,N_5182,N_8120);
and U13492 (N_13492,N_7320,N_5853);
nand U13493 (N_13493,N_8300,N_7195);
and U13494 (N_13494,N_6085,N_8570);
nand U13495 (N_13495,N_6193,N_6933);
nand U13496 (N_13496,N_7184,N_8784);
and U13497 (N_13497,N_9983,N_8139);
or U13498 (N_13498,N_6581,N_5300);
or U13499 (N_13499,N_7658,N_9403);
xnor U13500 (N_13500,N_8341,N_9415);
nand U13501 (N_13501,N_8525,N_5839);
or U13502 (N_13502,N_9357,N_5717);
xnor U13503 (N_13503,N_8645,N_5590);
nor U13504 (N_13504,N_9289,N_7817);
nand U13505 (N_13505,N_5683,N_9636);
and U13506 (N_13506,N_6038,N_9062);
xnor U13507 (N_13507,N_7358,N_5736);
nor U13508 (N_13508,N_6897,N_5735);
and U13509 (N_13509,N_6520,N_7417);
nor U13510 (N_13510,N_6051,N_8791);
or U13511 (N_13511,N_7527,N_7410);
nor U13512 (N_13512,N_9427,N_6547);
and U13513 (N_13513,N_5891,N_6053);
and U13514 (N_13514,N_7764,N_7174);
xor U13515 (N_13515,N_8162,N_8325);
nand U13516 (N_13516,N_5321,N_5032);
nand U13517 (N_13517,N_6465,N_7528);
xor U13518 (N_13518,N_7910,N_9566);
or U13519 (N_13519,N_9829,N_7686);
and U13520 (N_13520,N_5416,N_9840);
nand U13521 (N_13521,N_5905,N_9715);
or U13522 (N_13522,N_7744,N_6834);
and U13523 (N_13523,N_8163,N_8207);
nand U13524 (N_13524,N_6173,N_7062);
nand U13525 (N_13525,N_8471,N_8735);
xnor U13526 (N_13526,N_5702,N_5720);
xor U13527 (N_13527,N_7098,N_6320);
or U13528 (N_13528,N_6215,N_5154);
xnor U13529 (N_13529,N_5671,N_7422);
xor U13530 (N_13530,N_7264,N_6532);
and U13531 (N_13531,N_8103,N_5217);
xnor U13532 (N_13532,N_9757,N_8441);
nor U13533 (N_13533,N_5676,N_6192);
nand U13534 (N_13534,N_9841,N_8961);
and U13535 (N_13535,N_5967,N_7051);
nor U13536 (N_13536,N_6304,N_9822);
and U13537 (N_13537,N_8010,N_7960);
and U13538 (N_13538,N_9565,N_8441);
and U13539 (N_13539,N_9180,N_8159);
nor U13540 (N_13540,N_9680,N_9316);
xor U13541 (N_13541,N_9288,N_8899);
nor U13542 (N_13542,N_9220,N_9180);
nand U13543 (N_13543,N_6775,N_7730);
and U13544 (N_13544,N_5654,N_9482);
or U13545 (N_13545,N_5813,N_9691);
and U13546 (N_13546,N_9116,N_8505);
or U13547 (N_13547,N_8405,N_7631);
or U13548 (N_13548,N_9246,N_7337);
nand U13549 (N_13549,N_8185,N_6638);
nand U13550 (N_13550,N_7092,N_9339);
or U13551 (N_13551,N_6556,N_7811);
or U13552 (N_13552,N_9286,N_5496);
or U13553 (N_13553,N_5763,N_7181);
nand U13554 (N_13554,N_8339,N_5245);
and U13555 (N_13555,N_5511,N_8634);
xor U13556 (N_13556,N_7911,N_6551);
xor U13557 (N_13557,N_6387,N_6944);
nor U13558 (N_13558,N_9105,N_9691);
or U13559 (N_13559,N_6226,N_9534);
or U13560 (N_13560,N_8921,N_5190);
nand U13561 (N_13561,N_6906,N_5419);
nor U13562 (N_13562,N_7703,N_9986);
or U13563 (N_13563,N_5031,N_5507);
and U13564 (N_13564,N_5315,N_5372);
and U13565 (N_13565,N_7859,N_6851);
and U13566 (N_13566,N_7527,N_6111);
and U13567 (N_13567,N_7735,N_7757);
nand U13568 (N_13568,N_7416,N_7194);
or U13569 (N_13569,N_9682,N_9504);
and U13570 (N_13570,N_6729,N_5398);
and U13571 (N_13571,N_8963,N_5387);
nor U13572 (N_13572,N_5907,N_8302);
nor U13573 (N_13573,N_9009,N_9320);
or U13574 (N_13574,N_7291,N_8493);
nor U13575 (N_13575,N_5225,N_7538);
nand U13576 (N_13576,N_7920,N_7760);
and U13577 (N_13577,N_7915,N_8283);
or U13578 (N_13578,N_6168,N_5206);
or U13579 (N_13579,N_7648,N_6757);
xor U13580 (N_13580,N_6910,N_9838);
xor U13581 (N_13581,N_5486,N_5076);
or U13582 (N_13582,N_7677,N_8918);
nor U13583 (N_13583,N_5582,N_9884);
nand U13584 (N_13584,N_5974,N_7777);
nor U13585 (N_13585,N_6359,N_6478);
nand U13586 (N_13586,N_5037,N_7874);
xnor U13587 (N_13587,N_5054,N_9768);
and U13588 (N_13588,N_6343,N_6455);
nor U13589 (N_13589,N_8968,N_8294);
nor U13590 (N_13590,N_7001,N_8426);
xor U13591 (N_13591,N_9903,N_8150);
or U13592 (N_13592,N_9079,N_9852);
nor U13593 (N_13593,N_5089,N_5090);
and U13594 (N_13594,N_9846,N_5583);
nand U13595 (N_13595,N_5445,N_5390);
xnor U13596 (N_13596,N_7809,N_7583);
nand U13597 (N_13597,N_9838,N_9062);
and U13598 (N_13598,N_5442,N_5570);
or U13599 (N_13599,N_9044,N_8825);
and U13600 (N_13600,N_6162,N_5804);
or U13601 (N_13601,N_8048,N_8075);
or U13602 (N_13602,N_9728,N_5963);
and U13603 (N_13603,N_9417,N_7641);
nand U13604 (N_13604,N_9506,N_5504);
xnor U13605 (N_13605,N_9933,N_5459);
xor U13606 (N_13606,N_7164,N_8225);
or U13607 (N_13607,N_6502,N_7967);
or U13608 (N_13608,N_8588,N_9351);
xor U13609 (N_13609,N_7190,N_7779);
and U13610 (N_13610,N_7475,N_5684);
nor U13611 (N_13611,N_5522,N_5861);
xnor U13612 (N_13612,N_6226,N_7348);
nand U13613 (N_13613,N_9066,N_6443);
and U13614 (N_13614,N_5097,N_8659);
and U13615 (N_13615,N_9600,N_8112);
xor U13616 (N_13616,N_9298,N_5076);
or U13617 (N_13617,N_8428,N_7882);
nor U13618 (N_13618,N_8762,N_8226);
nor U13619 (N_13619,N_6650,N_5407);
nand U13620 (N_13620,N_7213,N_9564);
xnor U13621 (N_13621,N_8086,N_6958);
and U13622 (N_13622,N_6251,N_5913);
nand U13623 (N_13623,N_8563,N_7675);
or U13624 (N_13624,N_7680,N_7856);
nand U13625 (N_13625,N_7690,N_6855);
nor U13626 (N_13626,N_8863,N_5997);
or U13627 (N_13627,N_8247,N_5232);
or U13628 (N_13628,N_6560,N_6873);
nand U13629 (N_13629,N_9623,N_6563);
or U13630 (N_13630,N_5339,N_7317);
nor U13631 (N_13631,N_8967,N_7136);
nor U13632 (N_13632,N_8810,N_7209);
xor U13633 (N_13633,N_9540,N_8952);
and U13634 (N_13634,N_5502,N_8937);
nand U13635 (N_13635,N_7740,N_7547);
nand U13636 (N_13636,N_8723,N_8399);
xor U13637 (N_13637,N_9232,N_7514);
or U13638 (N_13638,N_7996,N_6368);
nand U13639 (N_13639,N_7410,N_5198);
and U13640 (N_13640,N_6257,N_6988);
nand U13641 (N_13641,N_9899,N_5062);
nand U13642 (N_13642,N_6897,N_6650);
nand U13643 (N_13643,N_8977,N_7579);
or U13644 (N_13644,N_6876,N_5490);
nand U13645 (N_13645,N_5955,N_8774);
xor U13646 (N_13646,N_5251,N_5898);
nand U13647 (N_13647,N_8127,N_5229);
xnor U13648 (N_13648,N_7364,N_8450);
nor U13649 (N_13649,N_8668,N_9364);
nor U13650 (N_13650,N_6762,N_7537);
xor U13651 (N_13651,N_9196,N_9033);
and U13652 (N_13652,N_7477,N_8899);
nand U13653 (N_13653,N_6606,N_7943);
or U13654 (N_13654,N_6995,N_5700);
and U13655 (N_13655,N_8532,N_7300);
nor U13656 (N_13656,N_5771,N_9967);
nor U13657 (N_13657,N_6243,N_8608);
xor U13658 (N_13658,N_7757,N_7762);
nand U13659 (N_13659,N_6466,N_5221);
and U13660 (N_13660,N_6052,N_9945);
nor U13661 (N_13661,N_9766,N_5780);
or U13662 (N_13662,N_8655,N_8125);
nand U13663 (N_13663,N_5486,N_9034);
nand U13664 (N_13664,N_7357,N_8307);
nand U13665 (N_13665,N_9321,N_5191);
nor U13666 (N_13666,N_6544,N_5279);
or U13667 (N_13667,N_5095,N_6981);
xnor U13668 (N_13668,N_6508,N_6266);
and U13669 (N_13669,N_6876,N_7380);
nor U13670 (N_13670,N_7539,N_9926);
xnor U13671 (N_13671,N_5494,N_9805);
xnor U13672 (N_13672,N_9559,N_8255);
xor U13673 (N_13673,N_5992,N_9840);
xor U13674 (N_13674,N_9693,N_8889);
or U13675 (N_13675,N_9668,N_9889);
xor U13676 (N_13676,N_6679,N_5875);
nand U13677 (N_13677,N_6564,N_8438);
xnor U13678 (N_13678,N_6906,N_9353);
or U13679 (N_13679,N_5996,N_6113);
or U13680 (N_13680,N_5646,N_7138);
xor U13681 (N_13681,N_9855,N_6917);
nor U13682 (N_13682,N_8173,N_6624);
nand U13683 (N_13683,N_6131,N_5048);
or U13684 (N_13684,N_8802,N_9586);
xnor U13685 (N_13685,N_5774,N_9943);
or U13686 (N_13686,N_8885,N_8614);
xnor U13687 (N_13687,N_7716,N_7034);
nand U13688 (N_13688,N_9040,N_7272);
nor U13689 (N_13689,N_5704,N_9240);
xor U13690 (N_13690,N_5318,N_6040);
or U13691 (N_13691,N_7720,N_7547);
and U13692 (N_13692,N_6895,N_9781);
or U13693 (N_13693,N_6055,N_7396);
and U13694 (N_13694,N_9677,N_7786);
xnor U13695 (N_13695,N_6806,N_6533);
xor U13696 (N_13696,N_9866,N_7094);
and U13697 (N_13697,N_7632,N_7908);
xor U13698 (N_13698,N_5760,N_7732);
nor U13699 (N_13699,N_5067,N_7823);
xnor U13700 (N_13700,N_8342,N_7398);
nand U13701 (N_13701,N_6943,N_8031);
xnor U13702 (N_13702,N_5597,N_9501);
xnor U13703 (N_13703,N_8498,N_9369);
xor U13704 (N_13704,N_7691,N_9502);
or U13705 (N_13705,N_6971,N_5276);
nand U13706 (N_13706,N_6300,N_6626);
nor U13707 (N_13707,N_6727,N_5857);
and U13708 (N_13708,N_8054,N_5445);
xor U13709 (N_13709,N_8212,N_6466);
or U13710 (N_13710,N_7631,N_8994);
nor U13711 (N_13711,N_6887,N_9975);
nor U13712 (N_13712,N_7763,N_7881);
nor U13713 (N_13713,N_9371,N_5885);
nor U13714 (N_13714,N_6540,N_9824);
nand U13715 (N_13715,N_8004,N_5497);
or U13716 (N_13716,N_5197,N_8465);
and U13717 (N_13717,N_5317,N_9798);
nand U13718 (N_13718,N_9889,N_8593);
or U13719 (N_13719,N_5817,N_5799);
or U13720 (N_13720,N_6618,N_9815);
nor U13721 (N_13721,N_7461,N_6346);
nor U13722 (N_13722,N_5296,N_7028);
xnor U13723 (N_13723,N_5881,N_6799);
and U13724 (N_13724,N_8954,N_9846);
or U13725 (N_13725,N_7172,N_5020);
and U13726 (N_13726,N_7737,N_9869);
xnor U13727 (N_13727,N_8555,N_5995);
or U13728 (N_13728,N_9113,N_5476);
nand U13729 (N_13729,N_6013,N_6102);
or U13730 (N_13730,N_7028,N_8177);
xor U13731 (N_13731,N_7010,N_9922);
nand U13732 (N_13732,N_9207,N_5651);
and U13733 (N_13733,N_8318,N_8618);
xnor U13734 (N_13734,N_5198,N_8597);
nor U13735 (N_13735,N_5057,N_9856);
nand U13736 (N_13736,N_8575,N_9639);
or U13737 (N_13737,N_8489,N_9543);
nand U13738 (N_13738,N_6164,N_6388);
nand U13739 (N_13739,N_6546,N_7755);
nand U13740 (N_13740,N_7424,N_8062);
xnor U13741 (N_13741,N_8485,N_6574);
or U13742 (N_13742,N_9062,N_7910);
or U13743 (N_13743,N_7830,N_9351);
nand U13744 (N_13744,N_8886,N_6023);
nor U13745 (N_13745,N_6986,N_8836);
xor U13746 (N_13746,N_8863,N_5865);
nor U13747 (N_13747,N_8688,N_9397);
and U13748 (N_13748,N_6524,N_6876);
xor U13749 (N_13749,N_8692,N_7760);
or U13750 (N_13750,N_6376,N_8900);
nand U13751 (N_13751,N_6842,N_5858);
xnor U13752 (N_13752,N_5790,N_8180);
xor U13753 (N_13753,N_5655,N_6289);
xnor U13754 (N_13754,N_6326,N_6492);
nand U13755 (N_13755,N_8523,N_9179);
nand U13756 (N_13756,N_6804,N_9046);
or U13757 (N_13757,N_6378,N_8403);
nand U13758 (N_13758,N_5075,N_8122);
or U13759 (N_13759,N_7608,N_8011);
xnor U13760 (N_13760,N_7286,N_6423);
or U13761 (N_13761,N_8339,N_6559);
nand U13762 (N_13762,N_8281,N_8709);
nand U13763 (N_13763,N_5174,N_7712);
and U13764 (N_13764,N_9950,N_9939);
nor U13765 (N_13765,N_9880,N_9795);
or U13766 (N_13766,N_5746,N_8053);
nand U13767 (N_13767,N_7979,N_6502);
xnor U13768 (N_13768,N_9500,N_7264);
nor U13769 (N_13769,N_7666,N_7961);
and U13770 (N_13770,N_7058,N_5687);
nand U13771 (N_13771,N_5798,N_5157);
nor U13772 (N_13772,N_5206,N_5653);
and U13773 (N_13773,N_7333,N_8413);
xnor U13774 (N_13774,N_6536,N_6823);
nand U13775 (N_13775,N_5802,N_7315);
and U13776 (N_13776,N_7405,N_5475);
nor U13777 (N_13777,N_8581,N_6819);
xor U13778 (N_13778,N_5752,N_5202);
or U13779 (N_13779,N_8897,N_5223);
nor U13780 (N_13780,N_9235,N_6865);
and U13781 (N_13781,N_8132,N_8497);
nand U13782 (N_13782,N_6702,N_7994);
or U13783 (N_13783,N_6382,N_5269);
nand U13784 (N_13784,N_6676,N_9590);
nand U13785 (N_13785,N_6707,N_9970);
nor U13786 (N_13786,N_6848,N_7449);
xor U13787 (N_13787,N_5874,N_6514);
or U13788 (N_13788,N_9748,N_8953);
xor U13789 (N_13789,N_5134,N_6151);
xor U13790 (N_13790,N_8365,N_9857);
nand U13791 (N_13791,N_5696,N_5034);
nor U13792 (N_13792,N_9673,N_6670);
or U13793 (N_13793,N_8306,N_7963);
nand U13794 (N_13794,N_6468,N_8517);
and U13795 (N_13795,N_7795,N_5459);
nand U13796 (N_13796,N_8966,N_9251);
nand U13797 (N_13797,N_6815,N_5703);
nor U13798 (N_13798,N_8472,N_7509);
and U13799 (N_13799,N_8399,N_6407);
nor U13800 (N_13800,N_5429,N_9792);
or U13801 (N_13801,N_7458,N_9614);
xnor U13802 (N_13802,N_7295,N_7352);
or U13803 (N_13803,N_6918,N_9905);
xnor U13804 (N_13804,N_6275,N_8959);
or U13805 (N_13805,N_9636,N_6810);
xnor U13806 (N_13806,N_5198,N_9145);
nand U13807 (N_13807,N_8718,N_5971);
nor U13808 (N_13808,N_7378,N_8875);
nand U13809 (N_13809,N_8876,N_6576);
xnor U13810 (N_13810,N_5590,N_9783);
or U13811 (N_13811,N_7810,N_9161);
xor U13812 (N_13812,N_6754,N_5514);
nor U13813 (N_13813,N_9145,N_7870);
and U13814 (N_13814,N_8471,N_5565);
xor U13815 (N_13815,N_8580,N_9428);
or U13816 (N_13816,N_9951,N_7162);
or U13817 (N_13817,N_6984,N_5916);
and U13818 (N_13818,N_8308,N_8783);
or U13819 (N_13819,N_8796,N_5216);
or U13820 (N_13820,N_6855,N_5976);
nor U13821 (N_13821,N_7813,N_5737);
nor U13822 (N_13822,N_8644,N_5955);
or U13823 (N_13823,N_6199,N_9507);
nor U13824 (N_13824,N_7283,N_7458);
xnor U13825 (N_13825,N_8905,N_6003);
or U13826 (N_13826,N_9973,N_8101);
or U13827 (N_13827,N_9888,N_8345);
nand U13828 (N_13828,N_8756,N_6122);
or U13829 (N_13829,N_6203,N_7035);
xnor U13830 (N_13830,N_8930,N_5185);
or U13831 (N_13831,N_6409,N_8848);
nor U13832 (N_13832,N_5637,N_6659);
and U13833 (N_13833,N_6308,N_7865);
and U13834 (N_13834,N_5264,N_7172);
nor U13835 (N_13835,N_5795,N_8036);
nor U13836 (N_13836,N_9374,N_6374);
nand U13837 (N_13837,N_9920,N_6046);
or U13838 (N_13838,N_5968,N_8278);
nand U13839 (N_13839,N_6480,N_9262);
nor U13840 (N_13840,N_6979,N_7247);
nand U13841 (N_13841,N_8462,N_8134);
nand U13842 (N_13842,N_5697,N_9395);
and U13843 (N_13843,N_7135,N_8147);
nand U13844 (N_13844,N_7649,N_8895);
or U13845 (N_13845,N_8392,N_8913);
or U13846 (N_13846,N_6397,N_5931);
xor U13847 (N_13847,N_5559,N_9753);
nand U13848 (N_13848,N_6027,N_6411);
nor U13849 (N_13849,N_9723,N_8024);
or U13850 (N_13850,N_7310,N_5824);
or U13851 (N_13851,N_5893,N_5680);
nor U13852 (N_13852,N_9840,N_7622);
or U13853 (N_13853,N_6843,N_7333);
nand U13854 (N_13854,N_7762,N_6928);
and U13855 (N_13855,N_8035,N_5271);
nor U13856 (N_13856,N_6935,N_5176);
nor U13857 (N_13857,N_5243,N_7887);
xnor U13858 (N_13858,N_5896,N_5073);
and U13859 (N_13859,N_8294,N_7528);
and U13860 (N_13860,N_5975,N_9610);
and U13861 (N_13861,N_5632,N_6137);
and U13862 (N_13862,N_7267,N_5039);
xor U13863 (N_13863,N_9655,N_9738);
and U13864 (N_13864,N_5743,N_7231);
nand U13865 (N_13865,N_8981,N_6436);
nor U13866 (N_13866,N_6163,N_5391);
or U13867 (N_13867,N_9978,N_7234);
nand U13868 (N_13868,N_6027,N_8104);
and U13869 (N_13869,N_6014,N_6769);
xor U13870 (N_13870,N_5457,N_8904);
nor U13871 (N_13871,N_8181,N_9410);
nor U13872 (N_13872,N_9187,N_9718);
or U13873 (N_13873,N_7893,N_5000);
and U13874 (N_13874,N_7652,N_6255);
xor U13875 (N_13875,N_5009,N_5581);
xnor U13876 (N_13876,N_9779,N_8227);
nand U13877 (N_13877,N_8891,N_5192);
or U13878 (N_13878,N_8625,N_6011);
and U13879 (N_13879,N_7386,N_8765);
nor U13880 (N_13880,N_9311,N_7652);
or U13881 (N_13881,N_7394,N_5138);
or U13882 (N_13882,N_9567,N_6607);
nor U13883 (N_13883,N_9222,N_8378);
and U13884 (N_13884,N_7582,N_6083);
xnor U13885 (N_13885,N_5233,N_8404);
or U13886 (N_13886,N_9955,N_9978);
xnor U13887 (N_13887,N_9974,N_7338);
and U13888 (N_13888,N_9592,N_8431);
nor U13889 (N_13889,N_5571,N_6673);
or U13890 (N_13890,N_7937,N_9539);
xor U13891 (N_13891,N_5453,N_6521);
nand U13892 (N_13892,N_8025,N_6742);
and U13893 (N_13893,N_9030,N_7045);
xnor U13894 (N_13894,N_8226,N_9989);
xor U13895 (N_13895,N_6457,N_7426);
nor U13896 (N_13896,N_5440,N_7309);
or U13897 (N_13897,N_8788,N_6467);
and U13898 (N_13898,N_6285,N_6156);
nand U13899 (N_13899,N_6373,N_5833);
nor U13900 (N_13900,N_8840,N_5018);
or U13901 (N_13901,N_6223,N_9907);
and U13902 (N_13902,N_6497,N_7874);
or U13903 (N_13903,N_5065,N_9483);
or U13904 (N_13904,N_8735,N_5507);
nand U13905 (N_13905,N_7573,N_8137);
nand U13906 (N_13906,N_7460,N_7968);
nand U13907 (N_13907,N_6598,N_9306);
nand U13908 (N_13908,N_7276,N_8499);
nor U13909 (N_13909,N_8319,N_8114);
or U13910 (N_13910,N_8124,N_5819);
xor U13911 (N_13911,N_5393,N_5564);
nand U13912 (N_13912,N_5571,N_8994);
and U13913 (N_13913,N_6281,N_6735);
and U13914 (N_13914,N_7366,N_9628);
nand U13915 (N_13915,N_8315,N_8697);
or U13916 (N_13916,N_8703,N_6454);
and U13917 (N_13917,N_8158,N_8816);
and U13918 (N_13918,N_5111,N_7116);
nor U13919 (N_13919,N_9927,N_6943);
nor U13920 (N_13920,N_6098,N_7851);
and U13921 (N_13921,N_5378,N_8532);
nor U13922 (N_13922,N_5989,N_6835);
and U13923 (N_13923,N_9631,N_9952);
nand U13924 (N_13924,N_6473,N_6854);
nand U13925 (N_13925,N_7786,N_6029);
or U13926 (N_13926,N_8648,N_7220);
and U13927 (N_13927,N_7193,N_6799);
or U13928 (N_13928,N_8494,N_7034);
and U13929 (N_13929,N_8350,N_7044);
or U13930 (N_13930,N_6018,N_5041);
and U13931 (N_13931,N_7757,N_6483);
nor U13932 (N_13932,N_8084,N_8591);
nand U13933 (N_13933,N_5983,N_7129);
or U13934 (N_13934,N_5425,N_8831);
nor U13935 (N_13935,N_6862,N_7638);
or U13936 (N_13936,N_5798,N_7344);
xor U13937 (N_13937,N_8259,N_6108);
nor U13938 (N_13938,N_8915,N_8379);
or U13939 (N_13939,N_5654,N_8429);
nand U13940 (N_13940,N_8736,N_7158);
nand U13941 (N_13941,N_8082,N_5983);
or U13942 (N_13942,N_5523,N_6380);
nor U13943 (N_13943,N_6181,N_8846);
and U13944 (N_13944,N_8714,N_7176);
nor U13945 (N_13945,N_5738,N_8783);
or U13946 (N_13946,N_7868,N_8220);
nor U13947 (N_13947,N_7712,N_6961);
and U13948 (N_13948,N_8282,N_9748);
nor U13949 (N_13949,N_5789,N_9854);
or U13950 (N_13950,N_9110,N_7855);
and U13951 (N_13951,N_5974,N_8095);
nor U13952 (N_13952,N_5162,N_7534);
or U13953 (N_13953,N_9067,N_9729);
nor U13954 (N_13954,N_9161,N_8836);
or U13955 (N_13955,N_6220,N_7258);
nor U13956 (N_13956,N_9660,N_7312);
nand U13957 (N_13957,N_7346,N_8761);
or U13958 (N_13958,N_5166,N_5456);
or U13959 (N_13959,N_5523,N_5153);
xnor U13960 (N_13960,N_8836,N_8554);
nand U13961 (N_13961,N_8711,N_8094);
nor U13962 (N_13962,N_9334,N_7762);
nand U13963 (N_13963,N_9876,N_5382);
nor U13964 (N_13964,N_5821,N_8419);
xnor U13965 (N_13965,N_8533,N_8334);
or U13966 (N_13966,N_7597,N_5492);
xor U13967 (N_13967,N_9569,N_7273);
or U13968 (N_13968,N_7878,N_5574);
and U13969 (N_13969,N_6085,N_8750);
or U13970 (N_13970,N_5239,N_7879);
or U13971 (N_13971,N_8878,N_7013);
nand U13972 (N_13972,N_5063,N_7675);
and U13973 (N_13973,N_7789,N_7081);
or U13974 (N_13974,N_8087,N_5194);
nor U13975 (N_13975,N_6484,N_7428);
and U13976 (N_13976,N_9413,N_8788);
nor U13977 (N_13977,N_5677,N_9323);
nor U13978 (N_13978,N_6444,N_8643);
nand U13979 (N_13979,N_5849,N_7946);
nor U13980 (N_13980,N_6987,N_5569);
and U13981 (N_13981,N_8170,N_9712);
and U13982 (N_13982,N_8759,N_7053);
xor U13983 (N_13983,N_5097,N_6991);
and U13984 (N_13984,N_7238,N_6765);
and U13985 (N_13985,N_9113,N_8856);
nor U13986 (N_13986,N_5063,N_9579);
or U13987 (N_13987,N_6739,N_8024);
or U13988 (N_13988,N_7469,N_8452);
or U13989 (N_13989,N_8553,N_5098);
and U13990 (N_13990,N_5552,N_6324);
and U13991 (N_13991,N_7538,N_5365);
xnor U13992 (N_13992,N_6891,N_9739);
or U13993 (N_13993,N_7019,N_5136);
nand U13994 (N_13994,N_5426,N_6579);
nor U13995 (N_13995,N_9992,N_8252);
xnor U13996 (N_13996,N_8788,N_6150);
nand U13997 (N_13997,N_6207,N_6338);
nor U13998 (N_13998,N_7782,N_6960);
and U13999 (N_13999,N_8763,N_9175);
nand U14000 (N_14000,N_5510,N_6851);
nand U14001 (N_14001,N_8911,N_9637);
xnor U14002 (N_14002,N_5952,N_6491);
or U14003 (N_14003,N_5332,N_7205);
or U14004 (N_14004,N_8884,N_7832);
and U14005 (N_14005,N_6217,N_6597);
nand U14006 (N_14006,N_5573,N_5630);
xnor U14007 (N_14007,N_5618,N_7678);
or U14008 (N_14008,N_6162,N_7461);
xor U14009 (N_14009,N_9230,N_5394);
or U14010 (N_14010,N_9469,N_5112);
xor U14011 (N_14011,N_9830,N_9842);
or U14012 (N_14012,N_9333,N_9160);
or U14013 (N_14013,N_7815,N_6012);
or U14014 (N_14014,N_7061,N_8387);
xor U14015 (N_14015,N_8000,N_8525);
and U14016 (N_14016,N_5740,N_5965);
or U14017 (N_14017,N_9089,N_7622);
or U14018 (N_14018,N_9435,N_9691);
and U14019 (N_14019,N_7242,N_7140);
or U14020 (N_14020,N_7665,N_6970);
nor U14021 (N_14021,N_9872,N_7963);
nor U14022 (N_14022,N_5114,N_7658);
or U14023 (N_14023,N_5206,N_9918);
xor U14024 (N_14024,N_5032,N_9025);
or U14025 (N_14025,N_7598,N_8217);
nand U14026 (N_14026,N_5927,N_9081);
and U14027 (N_14027,N_9777,N_9526);
nor U14028 (N_14028,N_6018,N_6152);
or U14029 (N_14029,N_6923,N_7295);
nand U14030 (N_14030,N_6569,N_9189);
xnor U14031 (N_14031,N_7522,N_8459);
xor U14032 (N_14032,N_9532,N_7746);
xor U14033 (N_14033,N_6078,N_5980);
nand U14034 (N_14034,N_9262,N_6338);
nor U14035 (N_14035,N_9682,N_6204);
and U14036 (N_14036,N_7994,N_8757);
nand U14037 (N_14037,N_5858,N_8001);
or U14038 (N_14038,N_8660,N_8212);
xnor U14039 (N_14039,N_6538,N_8605);
nand U14040 (N_14040,N_7143,N_8521);
nor U14041 (N_14041,N_5025,N_9494);
and U14042 (N_14042,N_5546,N_5462);
nor U14043 (N_14043,N_8240,N_9750);
and U14044 (N_14044,N_7711,N_8388);
or U14045 (N_14045,N_6625,N_7767);
or U14046 (N_14046,N_9522,N_8257);
nor U14047 (N_14047,N_6885,N_7430);
and U14048 (N_14048,N_8323,N_8221);
or U14049 (N_14049,N_5916,N_7105);
nor U14050 (N_14050,N_7015,N_5451);
nand U14051 (N_14051,N_6331,N_9534);
xnor U14052 (N_14052,N_7454,N_5854);
and U14053 (N_14053,N_8513,N_7548);
xnor U14054 (N_14054,N_5201,N_8079);
and U14055 (N_14055,N_8616,N_9441);
or U14056 (N_14056,N_5867,N_7084);
or U14057 (N_14057,N_9382,N_6647);
or U14058 (N_14058,N_7663,N_8342);
xor U14059 (N_14059,N_9191,N_6744);
and U14060 (N_14060,N_6339,N_9986);
nor U14061 (N_14061,N_6994,N_7019);
nand U14062 (N_14062,N_9086,N_8706);
nor U14063 (N_14063,N_5386,N_5214);
or U14064 (N_14064,N_6777,N_9482);
nand U14065 (N_14065,N_9999,N_9391);
and U14066 (N_14066,N_8902,N_9023);
and U14067 (N_14067,N_5015,N_9910);
and U14068 (N_14068,N_8118,N_5912);
nor U14069 (N_14069,N_8510,N_8757);
nand U14070 (N_14070,N_8920,N_7719);
nand U14071 (N_14071,N_5653,N_7452);
nand U14072 (N_14072,N_7889,N_6805);
or U14073 (N_14073,N_8658,N_8463);
nand U14074 (N_14074,N_7199,N_6341);
nand U14075 (N_14075,N_6316,N_5016);
or U14076 (N_14076,N_6597,N_9786);
or U14077 (N_14077,N_9272,N_9706);
and U14078 (N_14078,N_7632,N_5572);
nor U14079 (N_14079,N_5168,N_5917);
nand U14080 (N_14080,N_5066,N_6868);
xor U14081 (N_14081,N_6221,N_5029);
nor U14082 (N_14082,N_9525,N_6814);
and U14083 (N_14083,N_5241,N_6563);
and U14084 (N_14084,N_8606,N_8945);
nor U14085 (N_14085,N_7703,N_6337);
or U14086 (N_14086,N_9616,N_9309);
or U14087 (N_14087,N_6985,N_7100);
or U14088 (N_14088,N_7458,N_6187);
nor U14089 (N_14089,N_9778,N_8238);
nand U14090 (N_14090,N_7877,N_5147);
nor U14091 (N_14091,N_8737,N_6873);
nand U14092 (N_14092,N_9860,N_9092);
xnor U14093 (N_14093,N_8112,N_8076);
xnor U14094 (N_14094,N_9754,N_5399);
or U14095 (N_14095,N_5193,N_7063);
nand U14096 (N_14096,N_5402,N_6776);
and U14097 (N_14097,N_6055,N_5899);
and U14098 (N_14098,N_8743,N_7813);
and U14099 (N_14099,N_9381,N_9157);
nor U14100 (N_14100,N_7597,N_9732);
nand U14101 (N_14101,N_8863,N_8571);
or U14102 (N_14102,N_6542,N_5280);
nor U14103 (N_14103,N_5701,N_7164);
nand U14104 (N_14104,N_9137,N_5853);
nand U14105 (N_14105,N_9361,N_7846);
and U14106 (N_14106,N_9271,N_9965);
or U14107 (N_14107,N_8146,N_9813);
xor U14108 (N_14108,N_8106,N_6207);
nor U14109 (N_14109,N_7307,N_6554);
and U14110 (N_14110,N_8055,N_9524);
and U14111 (N_14111,N_8126,N_9624);
or U14112 (N_14112,N_8564,N_9775);
nor U14113 (N_14113,N_6362,N_9078);
nand U14114 (N_14114,N_9307,N_9992);
or U14115 (N_14115,N_9338,N_7601);
nand U14116 (N_14116,N_9198,N_5487);
nor U14117 (N_14117,N_5012,N_9033);
xnor U14118 (N_14118,N_9826,N_5239);
nand U14119 (N_14119,N_9235,N_9547);
or U14120 (N_14120,N_9719,N_9045);
nand U14121 (N_14121,N_6163,N_7831);
nor U14122 (N_14122,N_7846,N_7797);
xor U14123 (N_14123,N_6365,N_8433);
or U14124 (N_14124,N_6890,N_6134);
xnor U14125 (N_14125,N_6326,N_5806);
xnor U14126 (N_14126,N_8487,N_7535);
and U14127 (N_14127,N_7844,N_8102);
and U14128 (N_14128,N_7914,N_7091);
xnor U14129 (N_14129,N_5393,N_8036);
nand U14130 (N_14130,N_6581,N_5600);
nor U14131 (N_14131,N_7013,N_5540);
nor U14132 (N_14132,N_7039,N_8227);
nand U14133 (N_14133,N_6373,N_5617);
nand U14134 (N_14134,N_8811,N_9401);
and U14135 (N_14135,N_7398,N_9654);
nor U14136 (N_14136,N_9731,N_7570);
and U14137 (N_14137,N_5084,N_7962);
xnor U14138 (N_14138,N_5458,N_6585);
or U14139 (N_14139,N_6803,N_6235);
nand U14140 (N_14140,N_5108,N_5113);
xor U14141 (N_14141,N_9986,N_5737);
or U14142 (N_14142,N_9295,N_8324);
xor U14143 (N_14143,N_8610,N_7538);
and U14144 (N_14144,N_6004,N_5313);
nand U14145 (N_14145,N_6416,N_8951);
xnor U14146 (N_14146,N_7160,N_7862);
nand U14147 (N_14147,N_8467,N_6017);
nor U14148 (N_14148,N_8258,N_7535);
nand U14149 (N_14149,N_7086,N_6420);
and U14150 (N_14150,N_5286,N_9425);
nor U14151 (N_14151,N_8511,N_9564);
xor U14152 (N_14152,N_7191,N_7425);
and U14153 (N_14153,N_9588,N_9520);
or U14154 (N_14154,N_6613,N_6820);
nor U14155 (N_14155,N_9107,N_5264);
xnor U14156 (N_14156,N_8275,N_6631);
and U14157 (N_14157,N_8073,N_6308);
nor U14158 (N_14158,N_8421,N_7491);
nor U14159 (N_14159,N_7591,N_9278);
nor U14160 (N_14160,N_6619,N_9442);
or U14161 (N_14161,N_7221,N_8276);
and U14162 (N_14162,N_9705,N_9758);
and U14163 (N_14163,N_6582,N_8997);
or U14164 (N_14164,N_8749,N_8353);
and U14165 (N_14165,N_8998,N_6392);
and U14166 (N_14166,N_5627,N_7311);
nand U14167 (N_14167,N_5491,N_8015);
and U14168 (N_14168,N_6487,N_8114);
nand U14169 (N_14169,N_8341,N_7944);
and U14170 (N_14170,N_8227,N_9002);
nor U14171 (N_14171,N_6519,N_5464);
xor U14172 (N_14172,N_5497,N_9343);
nor U14173 (N_14173,N_8279,N_9084);
or U14174 (N_14174,N_8419,N_7847);
nor U14175 (N_14175,N_7373,N_9251);
xor U14176 (N_14176,N_7533,N_5220);
or U14177 (N_14177,N_7905,N_9837);
or U14178 (N_14178,N_7422,N_5845);
xnor U14179 (N_14179,N_7872,N_9035);
nor U14180 (N_14180,N_6039,N_7170);
or U14181 (N_14181,N_7236,N_5323);
or U14182 (N_14182,N_9566,N_7478);
or U14183 (N_14183,N_6848,N_6413);
or U14184 (N_14184,N_7027,N_9651);
nand U14185 (N_14185,N_8652,N_8859);
and U14186 (N_14186,N_7910,N_8768);
nand U14187 (N_14187,N_5870,N_6681);
nor U14188 (N_14188,N_8969,N_9509);
and U14189 (N_14189,N_9514,N_9383);
and U14190 (N_14190,N_6695,N_6491);
and U14191 (N_14191,N_6300,N_6768);
xor U14192 (N_14192,N_5232,N_6117);
nor U14193 (N_14193,N_8348,N_9945);
or U14194 (N_14194,N_8833,N_7756);
and U14195 (N_14195,N_7015,N_8737);
nand U14196 (N_14196,N_5932,N_6771);
and U14197 (N_14197,N_6921,N_9349);
nor U14198 (N_14198,N_9773,N_8610);
and U14199 (N_14199,N_6488,N_5411);
and U14200 (N_14200,N_6167,N_5340);
nor U14201 (N_14201,N_8046,N_7131);
or U14202 (N_14202,N_9225,N_8792);
nand U14203 (N_14203,N_8436,N_6851);
or U14204 (N_14204,N_8375,N_9338);
nand U14205 (N_14205,N_5137,N_6592);
and U14206 (N_14206,N_9462,N_7247);
and U14207 (N_14207,N_5177,N_5819);
xnor U14208 (N_14208,N_5162,N_5326);
nor U14209 (N_14209,N_6621,N_5272);
and U14210 (N_14210,N_7099,N_8791);
xnor U14211 (N_14211,N_7950,N_8424);
and U14212 (N_14212,N_9161,N_9184);
nand U14213 (N_14213,N_8864,N_9847);
nand U14214 (N_14214,N_7459,N_8902);
or U14215 (N_14215,N_5181,N_8630);
or U14216 (N_14216,N_5138,N_8893);
or U14217 (N_14217,N_9190,N_6430);
and U14218 (N_14218,N_5677,N_6121);
nand U14219 (N_14219,N_6739,N_8614);
and U14220 (N_14220,N_8873,N_6696);
nand U14221 (N_14221,N_9042,N_9843);
or U14222 (N_14222,N_5193,N_7957);
nand U14223 (N_14223,N_9238,N_5586);
nand U14224 (N_14224,N_9379,N_7978);
and U14225 (N_14225,N_5473,N_9845);
or U14226 (N_14226,N_6299,N_9625);
or U14227 (N_14227,N_9729,N_6666);
nor U14228 (N_14228,N_6264,N_8070);
and U14229 (N_14229,N_6528,N_8726);
xor U14230 (N_14230,N_7437,N_8266);
nand U14231 (N_14231,N_5440,N_9692);
nand U14232 (N_14232,N_9912,N_8021);
xor U14233 (N_14233,N_6291,N_5758);
or U14234 (N_14234,N_8599,N_8084);
or U14235 (N_14235,N_5694,N_8924);
or U14236 (N_14236,N_8525,N_9280);
and U14237 (N_14237,N_9387,N_5366);
nand U14238 (N_14238,N_6870,N_9215);
and U14239 (N_14239,N_6745,N_6446);
and U14240 (N_14240,N_8656,N_9322);
or U14241 (N_14241,N_7555,N_6706);
or U14242 (N_14242,N_6001,N_9411);
xor U14243 (N_14243,N_5966,N_5238);
or U14244 (N_14244,N_6451,N_6268);
or U14245 (N_14245,N_8814,N_8120);
or U14246 (N_14246,N_5973,N_5116);
nor U14247 (N_14247,N_8581,N_8419);
or U14248 (N_14248,N_5438,N_5171);
nand U14249 (N_14249,N_5585,N_8575);
nand U14250 (N_14250,N_5452,N_8971);
xor U14251 (N_14251,N_6184,N_6532);
or U14252 (N_14252,N_7917,N_5324);
xnor U14253 (N_14253,N_6448,N_6590);
or U14254 (N_14254,N_5445,N_8550);
or U14255 (N_14255,N_9804,N_9440);
xor U14256 (N_14256,N_8021,N_5621);
nor U14257 (N_14257,N_7401,N_7076);
nor U14258 (N_14258,N_5674,N_8984);
and U14259 (N_14259,N_6682,N_8836);
nor U14260 (N_14260,N_8100,N_5734);
nand U14261 (N_14261,N_8010,N_9501);
xnor U14262 (N_14262,N_6161,N_5859);
or U14263 (N_14263,N_7037,N_9380);
xor U14264 (N_14264,N_8476,N_8157);
xor U14265 (N_14265,N_9848,N_6399);
xor U14266 (N_14266,N_5036,N_7804);
xor U14267 (N_14267,N_8492,N_5322);
and U14268 (N_14268,N_6149,N_7208);
and U14269 (N_14269,N_8117,N_5403);
xnor U14270 (N_14270,N_5665,N_9753);
nor U14271 (N_14271,N_7628,N_7877);
nand U14272 (N_14272,N_5446,N_6914);
xnor U14273 (N_14273,N_8653,N_8306);
nand U14274 (N_14274,N_8910,N_9560);
and U14275 (N_14275,N_5390,N_5254);
and U14276 (N_14276,N_7445,N_7220);
or U14277 (N_14277,N_8099,N_9108);
xor U14278 (N_14278,N_9271,N_8231);
nor U14279 (N_14279,N_5094,N_9846);
nand U14280 (N_14280,N_9588,N_7614);
nand U14281 (N_14281,N_8925,N_6973);
nand U14282 (N_14282,N_8734,N_6692);
or U14283 (N_14283,N_8387,N_6137);
xnor U14284 (N_14284,N_7233,N_9495);
nand U14285 (N_14285,N_8738,N_6495);
xor U14286 (N_14286,N_7147,N_9607);
or U14287 (N_14287,N_7897,N_6185);
nand U14288 (N_14288,N_6740,N_7929);
and U14289 (N_14289,N_5044,N_8238);
nor U14290 (N_14290,N_9564,N_5294);
xnor U14291 (N_14291,N_5411,N_7840);
and U14292 (N_14292,N_9364,N_7538);
and U14293 (N_14293,N_9811,N_9039);
nand U14294 (N_14294,N_6596,N_6181);
nand U14295 (N_14295,N_6774,N_9394);
xnor U14296 (N_14296,N_7525,N_5696);
or U14297 (N_14297,N_9362,N_6076);
nor U14298 (N_14298,N_8932,N_6414);
nor U14299 (N_14299,N_6341,N_7686);
nor U14300 (N_14300,N_9413,N_6087);
or U14301 (N_14301,N_5181,N_6776);
xnor U14302 (N_14302,N_9196,N_9732);
and U14303 (N_14303,N_6220,N_7103);
and U14304 (N_14304,N_7238,N_9183);
or U14305 (N_14305,N_9034,N_5898);
xor U14306 (N_14306,N_8861,N_6800);
or U14307 (N_14307,N_6824,N_8566);
nor U14308 (N_14308,N_7221,N_8598);
and U14309 (N_14309,N_7154,N_7419);
nor U14310 (N_14310,N_8592,N_7423);
nor U14311 (N_14311,N_7280,N_6629);
nand U14312 (N_14312,N_5809,N_7307);
or U14313 (N_14313,N_7954,N_8073);
or U14314 (N_14314,N_7637,N_7845);
nor U14315 (N_14315,N_5597,N_6764);
and U14316 (N_14316,N_9964,N_6575);
nor U14317 (N_14317,N_9987,N_7411);
xor U14318 (N_14318,N_8927,N_5866);
nor U14319 (N_14319,N_6489,N_5541);
or U14320 (N_14320,N_7823,N_9979);
xor U14321 (N_14321,N_5850,N_7208);
or U14322 (N_14322,N_7544,N_8665);
xor U14323 (N_14323,N_9896,N_8525);
or U14324 (N_14324,N_7521,N_5014);
and U14325 (N_14325,N_5925,N_5918);
or U14326 (N_14326,N_8119,N_7558);
nor U14327 (N_14327,N_9673,N_7993);
nand U14328 (N_14328,N_6973,N_6430);
nor U14329 (N_14329,N_9173,N_5803);
nand U14330 (N_14330,N_6931,N_8108);
xnor U14331 (N_14331,N_8477,N_8190);
xor U14332 (N_14332,N_8701,N_7270);
or U14333 (N_14333,N_7722,N_9230);
or U14334 (N_14334,N_9494,N_8573);
xor U14335 (N_14335,N_5019,N_7273);
xnor U14336 (N_14336,N_8356,N_7228);
nand U14337 (N_14337,N_8958,N_7986);
nand U14338 (N_14338,N_9253,N_9639);
nand U14339 (N_14339,N_8962,N_8795);
nand U14340 (N_14340,N_8648,N_8127);
nor U14341 (N_14341,N_5230,N_9215);
or U14342 (N_14342,N_5017,N_5950);
nor U14343 (N_14343,N_5638,N_7178);
or U14344 (N_14344,N_6972,N_6600);
nand U14345 (N_14345,N_7416,N_8796);
and U14346 (N_14346,N_6749,N_7346);
xnor U14347 (N_14347,N_6322,N_9241);
nand U14348 (N_14348,N_7575,N_8968);
and U14349 (N_14349,N_9739,N_7071);
or U14350 (N_14350,N_7415,N_6272);
or U14351 (N_14351,N_9965,N_9993);
or U14352 (N_14352,N_8064,N_5110);
and U14353 (N_14353,N_6339,N_7670);
or U14354 (N_14354,N_8475,N_8005);
xor U14355 (N_14355,N_7727,N_5665);
and U14356 (N_14356,N_9186,N_7629);
xor U14357 (N_14357,N_7565,N_5813);
nor U14358 (N_14358,N_5062,N_7953);
nor U14359 (N_14359,N_6351,N_7416);
or U14360 (N_14360,N_9374,N_6013);
and U14361 (N_14361,N_8837,N_5025);
and U14362 (N_14362,N_8869,N_7695);
nand U14363 (N_14363,N_5921,N_6991);
or U14364 (N_14364,N_6827,N_6407);
xnor U14365 (N_14365,N_9374,N_5678);
or U14366 (N_14366,N_9287,N_9596);
and U14367 (N_14367,N_5369,N_7536);
nor U14368 (N_14368,N_5996,N_9531);
or U14369 (N_14369,N_6554,N_9852);
nor U14370 (N_14370,N_6439,N_5379);
and U14371 (N_14371,N_8230,N_6883);
and U14372 (N_14372,N_5429,N_9173);
or U14373 (N_14373,N_5420,N_6387);
nand U14374 (N_14374,N_5436,N_7516);
or U14375 (N_14375,N_9578,N_7965);
xor U14376 (N_14376,N_8159,N_9565);
nor U14377 (N_14377,N_5987,N_8930);
and U14378 (N_14378,N_6041,N_7199);
nor U14379 (N_14379,N_8728,N_8995);
nor U14380 (N_14380,N_5691,N_9902);
or U14381 (N_14381,N_6485,N_9473);
or U14382 (N_14382,N_9809,N_5570);
or U14383 (N_14383,N_9711,N_8807);
nand U14384 (N_14384,N_8486,N_6786);
xor U14385 (N_14385,N_6519,N_7373);
or U14386 (N_14386,N_6959,N_6037);
and U14387 (N_14387,N_7837,N_5612);
nor U14388 (N_14388,N_5168,N_8398);
or U14389 (N_14389,N_5481,N_8600);
xor U14390 (N_14390,N_6822,N_8542);
nor U14391 (N_14391,N_5276,N_8108);
or U14392 (N_14392,N_6789,N_7975);
xnor U14393 (N_14393,N_7256,N_8281);
xnor U14394 (N_14394,N_9974,N_9283);
or U14395 (N_14395,N_7505,N_6827);
or U14396 (N_14396,N_9376,N_5945);
nand U14397 (N_14397,N_5400,N_8366);
or U14398 (N_14398,N_8891,N_7675);
nor U14399 (N_14399,N_5869,N_5409);
nand U14400 (N_14400,N_6744,N_8078);
xnor U14401 (N_14401,N_9776,N_8767);
or U14402 (N_14402,N_5782,N_5906);
xnor U14403 (N_14403,N_8787,N_7828);
xor U14404 (N_14404,N_8749,N_5218);
xor U14405 (N_14405,N_6402,N_5466);
nor U14406 (N_14406,N_5095,N_9394);
and U14407 (N_14407,N_8840,N_7029);
and U14408 (N_14408,N_9198,N_9625);
or U14409 (N_14409,N_6101,N_8039);
or U14410 (N_14410,N_5890,N_7167);
and U14411 (N_14411,N_6128,N_8991);
or U14412 (N_14412,N_8681,N_6193);
nor U14413 (N_14413,N_8844,N_6845);
or U14414 (N_14414,N_5038,N_6421);
xor U14415 (N_14415,N_5973,N_7369);
or U14416 (N_14416,N_6948,N_8799);
nor U14417 (N_14417,N_9649,N_5873);
xor U14418 (N_14418,N_8266,N_9085);
or U14419 (N_14419,N_6840,N_9085);
nand U14420 (N_14420,N_9349,N_8947);
xor U14421 (N_14421,N_5817,N_9497);
xor U14422 (N_14422,N_5286,N_6282);
nor U14423 (N_14423,N_9400,N_5086);
nand U14424 (N_14424,N_8450,N_5001);
and U14425 (N_14425,N_7783,N_5403);
xnor U14426 (N_14426,N_6512,N_7975);
or U14427 (N_14427,N_5398,N_5094);
or U14428 (N_14428,N_9736,N_6096);
nor U14429 (N_14429,N_6667,N_6581);
nor U14430 (N_14430,N_8520,N_7993);
nor U14431 (N_14431,N_5945,N_5372);
and U14432 (N_14432,N_9846,N_5486);
or U14433 (N_14433,N_7436,N_9880);
nor U14434 (N_14434,N_6632,N_9264);
and U14435 (N_14435,N_5952,N_5372);
and U14436 (N_14436,N_6317,N_7156);
and U14437 (N_14437,N_6780,N_9959);
or U14438 (N_14438,N_5553,N_9015);
or U14439 (N_14439,N_9013,N_9611);
nor U14440 (N_14440,N_6016,N_8444);
and U14441 (N_14441,N_5787,N_5296);
or U14442 (N_14442,N_9330,N_8091);
xnor U14443 (N_14443,N_5681,N_9504);
and U14444 (N_14444,N_9055,N_5659);
xor U14445 (N_14445,N_5162,N_9517);
xnor U14446 (N_14446,N_7168,N_7254);
nor U14447 (N_14447,N_7585,N_8019);
xor U14448 (N_14448,N_6957,N_6894);
nor U14449 (N_14449,N_7292,N_9704);
xor U14450 (N_14450,N_7480,N_6055);
xor U14451 (N_14451,N_9113,N_6048);
nor U14452 (N_14452,N_6117,N_8076);
nand U14453 (N_14453,N_7486,N_6219);
nor U14454 (N_14454,N_9878,N_6653);
nor U14455 (N_14455,N_8692,N_9510);
nand U14456 (N_14456,N_7037,N_9625);
nor U14457 (N_14457,N_7938,N_5602);
nor U14458 (N_14458,N_9935,N_7731);
or U14459 (N_14459,N_8847,N_5230);
or U14460 (N_14460,N_6664,N_7577);
nand U14461 (N_14461,N_8843,N_6912);
nor U14462 (N_14462,N_9771,N_7010);
and U14463 (N_14463,N_6106,N_6978);
nor U14464 (N_14464,N_9260,N_7869);
or U14465 (N_14465,N_7733,N_6969);
nand U14466 (N_14466,N_8557,N_9756);
nor U14467 (N_14467,N_5211,N_9322);
and U14468 (N_14468,N_5909,N_7430);
xor U14469 (N_14469,N_8893,N_5644);
and U14470 (N_14470,N_7935,N_6546);
nand U14471 (N_14471,N_5238,N_5343);
and U14472 (N_14472,N_9538,N_6688);
xnor U14473 (N_14473,N_8411,N_7035);
xnor U14474 (N_14474,N_9479,N_9402);
nor U14475 (N_14475,N_7148,N_9524);
nor U14476 (N_14476,N_6647,N_6207);
or U14477 (N_14477,N_6997,N_5972);
and U14478 (N_14478,N_7574,N_5044);
xor U14479 (N_14479,N_6831,N_9618);
and U14480 (N_14480,N_5039,N_5070);
nand U14481 (N_14481,N_9246,N_6970);
xor U14482 (N_14482,N_7934,N_7080);
nor U14483 (N_14483,N_5838,N_8664);
xor U14484 (N_14484,N_8020,N_9317);
xnor U14485 (N_14485,N_7759,N_6655);
or U14486 (N_14486,N_5708,N_6049);
and U14487 (N_14487,N_6890,N_8466);
nor U14488 (N_14488,N_9080,N_9801);
xor U14489 (N_14489,N_8848,N_8891);
nand U14490 (N_14490,N_8327,N_9842);
xnor U14491 (N_14491,N_7970,N_8610);
or U14492 (N_14492,N_6938,N_9643);
xor U14493 (N_14493,N_6645,N_8155);
xor U14494 (N_14494,N_5225,N_6564);
nand U14495 (N_14495,N_6942,N_8812);
xor U14496 (N_14496,N_6695,N_5837);
nand U14497 (N_14497,N_8519,N_7633);
nand U14498 (N_14498,N_5841,N_6277);
and U14499 (N_14499,N_5900,N_7363);
nor U14500 (N_14500,N_9407,N_6328);
or U14501 (N_14501,N_5737,N_9185);
nand U14502 (N_14502,N_5530,N_8185);
nor U14503 (N_14503,N_9365,N_6844);
or U14504 (N_14504,N_9297,N_6903);
xnor U14505 (N_14505,N_8318,N_6549);
xor U14506 (N_14506,N_9038,N_5574);
or U14507 (N_14507,N_9368,N_5611);
and U14508 (N_14508,N_8943,N_6108);
xnor U14509 (N_14509,N_7834,N_5423);
xor U14510 (N_14510,N_7729,N_5461);
nor U14511 (N_14511,N_9173,N_7373);
nand U14512 (N_14512,N_7464,N_7968);
nand U14513 (N_14513,N_7951,N_6822);
or U14514 (N_14514,N_7558,N_6766);
and U14515 (N_14515,N_6970,N_8566);
and U14516 (N_14516,N_5130,N_6062);
xor U14517 (N_14517,N_7745,N_5066);
or U14518 (N_14518,N_6080,N_8724);
xnor U14519 (N_14519,N_5270,N_7900);
or U14520 (N_14520,N_6376,N_7743);
or U14521 (N_14521,N_9387,N_9137);
and U14522 (N_14522,N_5574,N_7424);
nor U14523 (N_14523,N_6790,N_7832);
nor U14524 (N_14524,N_6051,N_5125);
nand U14525 (N_14525,N_9278,N_9109);
and U14526 (N_14526,N_5057,N_6140);
or U14527 (N_14527,N_6362,N_7929);
and U14528 (N_14528,N_6745,N_6148);
nor U14529 (N_14529,N_6178,N_6916);
or U14530 (N_14530,N_8830,N_8805);
and U14531 (N_14531,N_7940,N_9933);
xor U14532 (N_14532,N_5201,N_9082);
or U14533 (N_14533,N_7937,N_6684);
and U14534 (N_14534,N_5180,N_8109);
nor U14535 (N_14535,N_8644,N_8992);
and U14536 (N_14536,N_7790,N_8196);
and U14537 (N_14537,N_9612,N_5688);
and U14538 (N_14538,N_9059,N_9246);
nand U14539 (N_14539,N_9397,N_9126);
nor U14540 (N_14540,N_7912,N_9578);
or U14541 (N_14541,N_6074,N_9197);
nand U14542 (N_14542,N_9769,N_8768);
and U14543 (N_14543,N_6716,N_5941);
or U14544 (N_14544,N_9887,N_6870);
xnor U14545 (N_14545,N_6361,N_5852);
and U14546 (N_14546,N_5649,N_9174);
or U14547 (N_14547,N_7762,N_5674);
xnor U14548 (N_14548,N_5477,N_5704);
nand U14549 (N_14549,N_5186,N_9568);
xor U14550 (N_14550,N_8266,N_7071);
or U14551 (N_14551,N_9503,N_7550);
nor U14552 (N_14552,N_9110,N_9767);
nor U14553 (N_14553,N_9895,N_7845);
xor U14554 (N_14554,N_6975,N_5752);
nand U14555 (N_14555,N_7657,N_9320);
or U14556 (N_14556,N_8832,N_8361);
or U14557 (N_14557,N_9012,N_8164);
and U14558 (N_14558,N_7844,N_8113);
or U14559 (N_14559,N_6397,N_5720);
and U14560 (N_14560,N_9168,N_5570);
or U14561 (N_14561,N_5970,N_9883);
xor U14562 (N_14562,N_5512,N_7466);
or U14563 (N_14563,N_8082,N_6395);
nor U14564 (N_14564,N_9188,N_6409);
nor U14565 (N_14565,N_9107,N_9308);
xnor U14566 (N_14566,N_8508,N_8182);
or U14567 (N_14567,N_8522,N_7833);
nand U14568 (N_14568,N_9543,N_7176);
nand U14569 (N_14569,N_5613,N_8040);
or U14570 (N_14570,N_9690,N_8675);
xnor U14571 (N_14571,N_5107,N_8310);
and U14572 (N_14572,N_5947,N_7510);
or U14573 (N_14573,N_8107,N_8386);
nor U14574 (N_14574,N_8848,N_6380);
and U14575 (N_14575,N_6303,N_5911);
nor U14576 (N_14576,N_8166,N_8220);
nor U14577 (N_14577,N_5045,N_7354);
nand U14578 (N_14578,N_6437,N_9578);
nand U14579 (N_14579,N_7685,N_8652);
or U14580 (N_14580,N_9073,N_6264);
xnor U14581 (N_14581,N_9137,N_9360);
or U14582 (N_14582,N_9760,N_7582);
xor U14583 (N_14583,N_5916,N_5972);
nor U14584 (N_14584,N_7050,N_5419);
xor U14585 (N_14585,N_6451,N_7809);
and U14586 (N_14586,N_8949,N_9253);
nand U14587 (N_14587,N_6684,N_8235);
xnor U14588 (N_14588,N_8421,N_8238);
nor U14589 (N_14589,N_5876,N_6322);
xnor U14590 (N_14590,N_9758,N_8525);
and U14591 (N_14591,N_8283,N_9189);
nor U14592 (N_14592,N_8479,N_5247);
nor U14593 (N_14593,N_5003,N_8468);
xnor U14594 (N_14594,N_6085,N_8508);
xor U14595 (N_14595,N_5673,N_7072);
and U14596 (N_14596,N_9358,N_9527);
nand U14597 (N_14597,N_6375,N_7330);
and U14598 (N_14598,N_5792,N_9609);
nor U14599 (N_14599,N_6853,N_5292);
or U14600 (N_14600,N_8735,N_7772);
xor U14601 (N_14601,N_9067,N_8658);
and U14602 (N_14602,N_8980,N_7125);
nand U14603 (N_14603,N_6793,N_9464);
or U14604 (N_14604,N_5333,N_8792);
or U14605 (N_14605,N_7647,N_8691);
and U14606 (N_14606,N_9957,N_7187);
nand U14607 (N_14607,N_8487,N_6349);
nor U14608 (N_14608,N_7222,N_7988);
nor U14609 (N_14609,N_9862,N_9938);
and U14610 (N_14610,N_8055,N_5445);
nor U14611 (N_14611,N_6605,N_7961);
nor U14612 (N_14612,N_7193,N_7584);
or U14613 (N_14613,N_5379,N_5430);
nand U14614 (N_14614,N_6213,N_6817);
nand U14615 (N_14615,N_6465,N_7748);
and U14616 (N_14616,N_9665,N_6695);
nand U14617 (N_14617,N_7597,N_7621);
nor U14618 (N_14618,N_6111,N_5111);
xnor U14619 (N_14619,N_6058,N_9972);
nor U14620 (N_14620,N_7091,N_9669);
nand U14621 (N_14621,N_5990,N_7746);
or U14622 (N_14622,N_8235,N_9435);
or U14623 (N_14623,N_8149,N_6032);
or U14624 (N_14624,N_8769,N_5846);
xor U14625 (N_14625,N_5129,N_5687);
nor U14626 (N_14626,N_8272,N_5121);
nor U14627 (N_14627,N_9337,N_8775);
xnor U14628 (N_14628,N_5024,N_7257);
and U14629 (N_14629,N_7133,N_7729);
or U14630 (N_14630,N_5043,N_8293);
and U14631 (N_14631,N_8848,N_8372);
nand U14632 (N_14632,N_7833,N_5976);
or U14633 (N_14633,N_5626,N_5314);
or U14634 (N_14634,N_5036,N_7841);
nand U14635 (N_14635,N_6050,N_6511);
nand U14636 (N_14636,N_8466,N_5151);
and U14637 (N_14637,N_5813,N_9546);
nor U14638 (N_14638,N_7760,N_8592);
nor U14639 (N_14639,N_9211,N_8822);
or U14640 (N_14640,N_6883,N_5366);
and U14641 (N_14641,N_9062,N_7150);
or U14642 (N_14642,N_7070,N_5195);
nand U14643 (N_14643,N_5377,N_9086);
nand U14644 (N_14644,N_5108,N_6394);
nand U14645 (N_14645,N_5230,N_9841);
or U14646 (N_14646,N_5678,N_8822);
or U14647 (N_14647,N_7176,N_9790);
or U14648 (N_14648,N_5525,N_8204);
and U14649 (N_14649,N_6391,N_8738);
nand U14650 (N_14650,N_8844,N_6804);
nor U14651 (N_14651,N_6735,N_6675);
xnor U14652 (N_14652,N_8627,N_9992);
xnor U14653 (N_14653,N_6258,N_9625);
nand U14654 (N_14654,N_9544,N_8640);
and U14655 (N_14655,N_8593,N_7569);
and U14656 (N_14656,N_7424,N_5120);
nor U14657 (N_14657,N_8065,N_5409);
xor U14658 (N_14658,N_6964,N_8968);
nand U14659 (N_14659,N_9340,N_7957);
xor U14660 (N_14660,N_7666,N_6809);
nand U14661 (N_14661,N_9345,N_7071);
xnor U14662 (N_14662,N_5064,N_8721);
nand U14663 (N_14663,N_7256,N_8258);
or U14664 (N_14664,N_7547,N_8273);
or U14665 (N_14665,N_9770,N_5198);
nand U14666 (N_14666,N_5822,N_5374);
and U14667 (N_14667,N_6050,N_5617);
xnor U14668 (N_14668,N_5593,N_7476);
nand U14669 (N_14669,N_5048,N_7268);
nor U14670 (N_14670,N_6142,N_5430);
or U14671 (N_14671,N_9768,N_5827);
xnor U14672 (N_14672,N_8905,N_6730);
nand U14673 (N_14673,N_9692,N_8513);
and U14674 (N_14674,N_9692,N_9716);
or U14675 (N_14675,N_9804,N_7503);
nor U14676 (N_14676,N_7281,N_9971);
and U14677 (N_14677,N_8442,N_6609);
or U14678 (N_14678,N_5371,N_9289);
or U14679 (N_14679,N_9453,N_5729);
nor U14680 (N_14680,N_8932,N_6675);
xor U14681 (N_14681,N_9679,N_8227);
and U14682 (N_14682,N_9556,N_5023);
and U14683 (N_14683,N_8272,N_5312);
or U14684 (N_14684,N_6471,N_5676);
or U14685 (N_14685,N_7219,N_8721);
nand U14686 (N_14686,N_5381,N_7993);
or U14687 (N_14687,N_8269,N_7411);
nor U14688 (N_14688,N_7666,N_7397);
nor U14689 (N_14689,N_7853,N_5764);
nor U14690 (N_14690,N_8131,N_8537);
or U14691 (N_14691,N_6835,N_9818);
nor U14692 (N_14692,N_9257,N_6909);
xor U14693 (N_14693,N_7113,N_7465);
xnor U14694 (N_14694,N_5146,N_5514);
and U14695 (N_14695,N_9796,N_7662);
xor U14696 (N_14696,N_5493,N_8273);
nor U14697 (N_14697,N_8525,N_7733);
nor U14698 (N_14698,N_5922,N_8230);
nand U14699 (N_14699,N_5051,N_9986);
or U14700 (N_14700,N_8499,N_6603);
or U14701 (N_14701,N_5342,N_6053);
and U14702 (N_14702,N_5336,N_6164);
and U14703 (N_14703,N_6352,N_6152);
xor U14704 (N_14704,N_6903,N_5481);
or U14705 (N_14705,N_9028,N_7749);
and U14706 (N_14706,N_8154,N_8557);
nand U14707 (N_14707,N_5709,N_7927);
nor U14708 (N_14708,N_9597,N_8319);
and U14709 (N_14709,N_7219,N_7928);
and U14710 (N_14710,N_7464,N_5673);
xor U14711 (N_14711,N_8655,N_9845);
xor U14712 (N_14712,N_9667,N_9578);
or U14713 (N_14713,N_7741,N_8427);
or U14714 (N_14714,N_6954,N_6442);
and U14715 (N_14715,N_8007,N_7276);
nand U14716 (N_14716,N_7347,N_7146);
nand U14717 (N_14717,N_5907,N_5391);
and U14718 (N_14718,N_7752,N_7056);
and U14719 (N_14719,N_8699,N_9654);
nand U14720 (N_14720,N_8073,N_7919);
xor U14721 (N_14721,N_7438,N_9021);
xnor U14722 (N_14722,N_6904,N_6696);
nor U14723 (N_14723,N_8319,N_8778);
nor U14724 (N_14724,N_6288,N_5552);
nor U14725 (N_14725,N_5300,N_8107);
nor U14726 (N_14726,N_9406,N_5732);
or U14727 (N_14727,N_8711,N_8932);
nor U14728 (N_14728,N_9612,N_9692);
nor U14729 (N_14729,N_8665,N_5293);
or U14730 (N_14730,N_9942,N_7668);
nor U14731 (N_14731,N_7998,N_7878);
nor U14732 (N_14732,N_6777,N_8605);
nand U14733 (N_14733,N_5327,N_8150);
nor U14734 (N_14734,N_7765,N_5465);
and U14735 (N_14735,N_5784,N_5204);
nand U14736 (N_14736,N_5711,N_7939);
nand U14737 (N_14737,N_6735,N_5973);
nor U14738 (N_14738,N_8613,N_7612);
nand U14739 (N_14739,N_6882,N_9583);
xor U14740 (N_14740,N_5733,N_7002);
and U14741 (N_14741,N_5295,N_6379);
xnor U14742 (N_14742,N_7526,N_8630);
and U14743 (N_14743,N_5351,N_8224);
and U14744 (N_14744,N_5819,N_8569);
or U14745 (N_14745,N_9100,N_6280);
nand U14746 (N_14746,N_9248,N_5281);
nand U14747 (N_14747,N_9047,N_9724);
nor U14748 (N_14748,N_6977,N_8856);
nand U14749 (N_14749,N_9522,N_6676);
nand U14750 (N_14750,N_7337,N_9846);
xnor U14751 (N_14751,N_8564,N_6458);
or U14752 (N_14752,N_9736,N_8619);
or U14753 (N_14753,N_8419,N_7788);
nor U14754 (N_14754,N_8810,N_6604);
nand U14755 (N_14755,N_9709,N_7904);
xnor U14756 (N_14756,N_8202,N_7906);
and U14757 (N_14757,N_7887,N_8595);
xnor U14758 (N_14758,N_6869,N_5533);
nand U14759 (N_14759,N_5407,N_6825);
nand U14760 (N_14760,N_5142,N_7887);
nor U14761 (N_14761,N_6908,N_7865);
nand U14762 (N_14762,N_7508,N_9829);
nand U14763 (N_14763,N_8817,N_5412);
or U14764 (N_14764,N_9065,N_8830);
nor U14765 (N_14765,N_6467,N_5547);
xor U14766 (N_14766,N_5226,N_5975);
nor U14767 (N_14767,N_8872,N_7110);
nor U14768 (N_14768,N_9815,N_9182);
xnor U14769 (N_14769,N_5026,N_6318);
and U14770 (N_14770,N_7571,N_7472);
or U14771 (N_14771,N_6312,N_5234);
nor U14772 (N_14772,N_6658,N_6115);
nor U14773 (N_14773,N_7171,N_6144);
or U14774 (N_14774,N_6328,N_5725);
nand U14775 (N_14775,N_5861,N_6557);
nand U14776 (N_14776,N_6591,N_8672);
nand U14777 (N_14777,N_7195,N_5504);
nand U14778 (N_14778,N_6431,N_7866);
and U14779 (N_14779,N_5817,N_5922);
xnor U14780 (N_14780,N_7321,N_5475);
or U14781 (N_14781,N_6560,N_8708);
and U14782 (N_14782,N_7638,N_9151);
nand U14783 (N_14783,N_6522,N_9618);
xnor U14784 (N_14784,N_7119,N_7178);
nand U14785 (N_14785,N_5972,N_8465);
and U14786 (N_14786,N_9295,N_7762);
xor U14787 (N_14787,N_7448,N_6625);
xor U14788 (N_14788,N_8099,N_5633);
nand U14789 (N_14789,N_7327,N_9050);
nor U14790 (N_14790,N_9830,N_7380);
nand U14791 (N_14791,N_9879,N_6365);
nor U14792 (N_14792,N_5234,N_5986);
nor U14793 (N_14793,N_6549,N_6596);
xor U14794 (N_14794,N_6271,N_5583);
nor U14795 (N_14795,N_8799,N_8922);
and U14796 (N_14796,N_5081,N_6793);
and U14797 (N_14797,N_7473,N_8593);
and U14798 (N_14798,N_9541,N_6590);
and U14799 (N_14799,N_8547,N_8988);
and U14800 (N_14800,N_5682,N_8428);
or U14801 (N_14801,N_6765,N_9582);
nand U14802 (N_14802,N_9598,N_6630);
xnor U14803 (N_14803,N_6445,N_7919);
or U14804 (N_14804,N_8491,N_5497);
nand U14805 (N_14805,N_9091,N_5712);
xor U14806 (N_14806,N_8215,N_7999);
and U14807 (N_14807,N_5715,N_7704);
or U14808 (N_14808,N_5795,N_7337);
or U14809 (N_14809,N_5089,N_9817);
and U14810 (N_14810,N_5003,N_8819);
nand U14811 (N_14811,N_5822,N_8000);
nand U14812 (N_14812,N_5349,N_6227);
xnor U14813 (N_14813,N_5594,N_7468);
xor U14814 (N_14814,N_9069,N_6141);
and U14815 (N_14815,N_9539,N_9267);
xnor U14816 (N_14816,N_9857,N_9867);
or U14817 (N_14817,N_9107,N_9055);
xor U14818 (N_14818,N_8035,N_8303);
nand U14819 (N_14819,N_6936,N_7819);
or U14820 (N_14820,N_5268,N_6474);
nor U14821 (N_14821,N_5629,N_6094);
and U14822 (N_14822,N_9378,N_6935);
nor U14823 (N_14823,N_9166,N_8922);
or U14824 (N_14824,N_5037,N_7176);
or U14825 (N_14825,N_5859,N_9355);
and U14826 (N_14826,N_7791,N_5896);
nor U14827 (N_14827,N_5616,N_5559);
xor U14828 (N_14828,N_6906,N_6059);
nor U14829 (N_14829,N_5031,N_8553);
nand U14830 (N_14830,N_9849,N_9419);
xnor U14831 (N_14831,N_7494,N_7718);
or U14832 (N_14832,N_6078,N_6278);
nor U14833 (N_14833,N_5436,N_9241);
or U14834 (N_14834,N_9481,N_6424);
xor U14835 (N_14835,N_8280,N_8290);
or U14836 (N_14836,N_8968,N_9613);
and U14837 (N_14837,N_7435,N_6215);
and U14838 (N_14838,N_6241,N_6685);
nor U14839 (N_14839,N_5264,N_9378);
nor U14840 (N_14840,N_9069,N_7232);
or U14841 (N_14841,N_8372,N_6180);
nand U14842 (N_14842,N_8706,N_8406);
nor U14843 (N_14843,N_9249,N_8575);
and U14844 (N_14844,N_8923,N_8556);
and U14845 (N_14845,N_6626,N_5844);
nand U14846 (N_14846,N_7721,N_6828);
or U14847 (N_14847,N_8136,N_5768);
nor U14848 (N_14848,N_9650,N_5510);
nand U14849 (N_14849,N_7246,N_9230);
xor U14850 (N_14850,N_8617,N_9574);
xor U14851 (N_14851,N_9124,N_6675);
xor U14852 (N_14852,N_8090,N_9913);
xnor U14853 (N_14853,N_7860,N_6023);
nand U14854 (N_14854,N_5028,N_7121);
xnor U14855 (N_14855,N_9356,N_8928);
or U14856 (N_14856,N_7742,N_5859);
nand U14857 (N_14857,N_6873,N_6999);
nor U14858 (N_14858,N_6839,N_9951);
nand U14859 (N_14859,N_9979,N_6207);
nor U14860 (N_14860,N_5459,N_5874);
nand U14861 (N_14861,N_6318,N_8139);
nand U14862 (N_14862,N_7191,N_8225);
nand U14863 (N_14863,N_5079,N_8891);
nand U14864 (N_14864,N_6741,N_7036);
nand U14865 (N_14865,N_7256,N_7224);
nor U14866 (N_14866,N_6278,N_9524);
or U14867 (N_14867,N_8392,N_5091);
nand U14868 (N_14868,N_9525,N_9283);
or U14869 (N_14869,N_9420,N_5918);
or U14870 (N_14870,N_9519,N_9343);
xnor U14871 (N_14871,N_6808,N_5146);
and U14872 (N_14872,N_8083,N_6918);
and U14873 (N_14873,N_7577,N_8702);
or U14874 (N_14874,N_9443,N_7410);
nand U14875 (N_14875,N_9770,N_9044);
nor U14876 (N_14876,N_6558,N_8445);
nand U14877 (N_14877,N_8752,N_5406);
xnor U14878 (N_14878,N_8603,N_7134);
or U14879 (N_14879,N_7058,N_8021);
and U14880 (N_14880,N_6658,N_6241);
nor U14881 (N_14881,N_6815,N_5726);
xor U14882 (N_14882,N_7841,N_7882);
nand U14883 (N_14883,N_9122,N_9848);
or U14884 (N_14884,N_6936,N_6516);
xor U14885 (N_14885,N_5916,N_5713);
nor U14886 (N_14886,N_9801,N_8191);
and U14887 (N_14887,N_7798,N_9652);
and U14888 (N_14888,N_5288,N_8197);
nand U14889 (N_14889,N_9215,N_5196);
xnor U14890 (N_14890,N_8099,N_6803);
xnor U14891 (N_14891,N_9554,N_9228);
nor U14892 (N_14892,N_6321,N_7638);
xnor U14893 (N_14893,N_7588,N_8179);
nand U14894 (N_14894,N_7431,N_9102);
and U14895 (N_14895,N_8084,N_8064);
xnor U14896 (N_14896,N_6827,N_8006);
nor U14897 (N_14897,N_6436,N_8633);
nand U14898 (N_14898,N_6769,N_6179);
or U14899 (N_14899,N_6002,N_7386);
or U14900 (N_14900,N_9846,N_6110);
and U14901 (N_14901,N_6352,N_9192);
or U14902 (N_14902,N_5554,N_6853);
nor U14903 (N_14903,N_9481,N_8593);
nor U14904 (N_14904,N_6894,N_9537);
xnor U14905 (N_14905,N_6516,N_5448);
and U14906 (N_14906,N_8295,N_5262);
nand U14907 (N_14907,N_6163,N_5338);
or U14908 (N_14908,N_5429,N_9073);
nor U14909 (N_14909,N_9764,N_6107);
and U14910 (N_14910,N_8865,N_8885);
and U14911 (N_14911,N_8726,N_8500);
or U14912 (N_14912,N_5906,N_6752);
nand U14913 (N_14913,N_8759,N_7279);
or U14914 (N_14914,N_5122,N_5884);
and U14915 (N_14915,N_8049,N_5105);
and U14916 (N_14916,N_9949,N_7304);
and U14917 (N_14917,N_7728,N_6470);
xor U14918 (N_14918,N_5098,N_8930);
nand U14919 (N_14919,N_7659,N_8955);
xor U14920 (N_14920,N_7967,N_8032);
nor U14921 (N_14921,N_5049,N_6900);
nand U14922 (N_14922,N_9761,N_6678);
xnor U14923 (N_14923,N_8978,N_5260);
xnor U14924 (N_14924,N_8428,N_5806);
xnor U14925 (N_14925,N_9145,N_8315);
nor U14926 (N_14926,N_7893,N_5196);
nor U14927 (N_14927,N_5723,N_7969);
nand U14928 (N_14928,N_6242,N_7973);
nand U14929 (N_14929,N_8758,N_5778);
and U14930 (N_14930,N_7661,N_9553);
or U14931 (N_14931,N_7370,N_9628);
xnor U14932 (N_14932,N_8980,N_6674);
nor U14933 (N_14933,N_5080,N_5306);
and U14934 (N_14934,N_8387,N_5782);
nor U14935 (N_14935,N_7982,N_9001);
nand U14936 (N_14936,N_7177,N_9046);
nand U14937 (N_14937,N_8612,N_6306);
and U14938 (N_14938,N_8051,N_7701);
or U14939 (N_14939,N_6787,N_7011);
xnor U14940 (N_14940,N_8288,N_7391);
nand U14941 (N_14941,N_7077,N_5037);
and U14942 (N_14942,N_5625,N_5183);
nor U14943 (N_14943,N_7942,N_5332);
xnor U14944 (N_14944,N_5887,N_7192);
xnor U14945 (N_14945,N_6255,N_5412);
xnor U14946 (N_14946,N_5852,N_6170);
and U14947 (N_14947,N_7771,N_6704);
or U14948 (N_14948,N_9899,N_8495);
or U14949 (N_14949,N_7429,N_5583);
or U14950 (N_14950,N_7290,N_6132);
nand U14951 (N_14951,N_7439,N_6203);
xor U14952 (N_14952,N_9689,N_7834);
nor U14953 (N_14953,N_9692,N_8832);
or U14954 (N_14954,N_9699,N_9534);
xor U14955 (N_14955,N_6491,N_6834);
xor U14956 (N_14956,N_7160,N_8728);
or U14957 (N_14957,N_5115,N_8770);
nor U14958 (N_14958,N_8098,N_6613);
or U14959 (N_14959,N_8531,N_5386);
or U14960 (N_14960,N_5801,N_7855);
nand U14961 (N_14961,N_6522,N_5566);
and U14962 (N_14962,N_8490,N_5379);
nand U14963 (N_14963,N_6733,N_5622);
and U14964 (N_14964,N_7054,N_5318);
nand U14965 (N_14965,N_9396,N_9196);
nor U14966 (N_14966,N_8887,N_8817);
nor U14967 (N_14967,N_5450,N_8262);
nor U14968 (N_14968,N_8138,N_7306);
nand U14969 (N_14969,N_9215,N_8597);
nor U14970 (N_14970,N_6141,N_9672);
nand U14971 (N_14971,N_9623,N_6035);
or U14972 (N_14972,N_5048,N_6366);
or U14973 (N_14973,N_5833,N_7469);
nand U14974 (N_14974,N_6355,N_8988);
or U14975 (N_14975,N_5195,N_5579);
xnor U14976 (N_14976,N_5877,N_7386);
nor U14977 (N_14977,N_6610,N_5851);
nor U14978 (N_14978,N_9268,N_7271);
nor U14979 (N_14979,N_8639,N_5365);
nor U14980 (N_14980,N_9086,N_8041);
nor U14981 (N_14981,N_7500,N_6672);
nand U14982 (N_14982,N_9532,N_9500);
and U14983 (N_14983,N_6915,N_9438);
or U14984 (N_14984,N_9641,N_6642);
and U14985 (N_14985,N_5001,N_8775);
xnor U14986 (N_14986,N_6307,N_9436);
xnor U14987 (N_14987,N_6656,N_7160);
nand U14988 (N_14988,N_7453,N_5507);
or U14989 (N_14989,N_9284,N_9865);
or U14990 (N_14990,N_8365,N_5248);
xor U14991 (N_14991,N_7227,N_5065);
and U14992 (N_14992,N_8207,N_7306);
nand U14993 (N_14993,N_7371,N_5599);
or U14994 (N_14994,N_5988,N_8172);
nor U14995 (N_14995,N_9978,N_9871);
or U14996 (N_14996,N_8932,N_5396);
and U14997 (N_14997,N_7582,N_9464);
and U14998 (N_14998,N_9922,N_6970);
or U14999 (N_14999,N_6991,N_5973);
nor U15000 (N_15000,N_13212,N_11792);
and U15001 (N_15001,N_11888,N_13063);
xor U15002 (N_15002,N_13537,N_14198);
nand U15003 (N_15003,N_14875,N_12937);
and U15004 (N_15004,N_14432,N_12965);
xnor U15005 (N_15005,N_14487,N_14442);
nand U15006 (N_15006,N_14829,N_11018);
nor U15007 (N_15007,N_13164,N_10260);
or U15008 (N_15008,N_10598,N_14932);
or U15009 (N_15009,N_12992,N_12847);
nand U15010 (N_15010,N_13036,N_14837);
or U15011 (N_15011,N_12207,N_10132);
or U15012 (N_15012,N_10753,N_13917);
nand U15013 (N_15013,N_12396,N_14688);
xor U15014 (N_15014,N_11641,N_10606);
nor U15015 (N_15015,N_13493,N_13231);
or U15016 (N_15016,N_12841,N_11775);
or U15017 (N_15017,N_13184,N_14209);
or U15018 (N_15018,N_14518,N_11412);
xnor U15019 (N_15019,N_10049,N_13546);
or U15020 (N_15020,N_12318,N_12949);
or U15021 (N_15021,N_14325,N_11349);
nor U15022 (N_15022,N_13750,N_12539);
xor U15023 (N_15023,N_13309,N_11194);
and U15024 (N_15024,N_14006,N_11042);
xnor U15025 (N_15025,N_11920,N_12805);
or U15026 (N_15026,N_11827,N_12900);
nor U15027 (N_15027,N_12511,N_10698);
or U15028 (N_15028,N_13176,N_12080);
and U15029 (N_15029,N_12060,N_11504);
nor U15030 (N_15030,N_14587,N_12178);
xnor U15031 (N_15031,N_10831,N_13699);
xnor U15032 (N_15032,N_14755,N_12001);
or U15033 (N_15033,N_10937,N_10109);
and U15034 (N_15034,N_11308,N_13382);
nor U15035 (N_15035,N_10202,N_10729);
xor U15036 (N_15036,N_10788,N_10657);
nor U15037 (N_15037,N_12485,N_13619);
nand U15038 (N_15038,N_13716,N_13811);
and U15039 (N_15039,N_13919,N_11969);
nand U15040 (N_15040,N_10140,N_12740);
nor U15041 (N_15041,N_13028,N_12295);
xor U15042 (N_15042,N_11232,N_10934);
xnor U15043 (N_15043,N_10785,N_10977);
nand U15044 (N_15044,N_14020,N_10527);
and U15045 (N_15045,N_10866,N_14307);
nor U15046 (N_15046,N_11752,N_13427);
nor U15047 (N_15047,N_14638,N_12758);
and U15048 (N_15048,N_14502,N_13075);
nor U15049 (N_15049,N_12825,N_10387);
or U15050 (N_15050,N_14352,N_10391);
and U15051 (N_15051,N_14053,N_14713);
or U15052 (N_15052,N_13524,N_13383);
nor U15053 (N_15053,N_13853,N_14014);
nand U15054 (N_15054,N_14483,N_14706);
xor U15055 (N_15055,N_13973,N_12643);
or U15056 (N_15056,N_12716,N_12421);
xnor U15057 (N_15057,N_11333,N_12098);
or U15058 (N_15058,N_12623,N_13479);
or U15059 (N_15059,N_10272,N_13453);
nor U15060 (N_15060,N_10286,N_14665);
and U15061 (N_15061,N_14627,N_12192);
nand U15062 (N_15062,N_10065,N_12704);
nor U15063 (N_15063,N_12425,N_10442);
nand U15064 (N_15064,N_13431,N_12345);
nor U15065 (N_15065,N_11320,N_12116);
nand U15066 (N_15066,N_14165,N_14052);
nand U15067 (N_15067,N_11411,N_10943);
and U15068 (N_15068,N_13281,N_13369);
nand U15069 (N_15069,N_12124,N_11521);
nand U15070 (N_15070,N_12050,N_13447);
nand U15071 (N_15071,N_11957,N_12674);
and U15072 (N_15072,N_11597,N_13214);
and U15073 (N_15073,N_12311,N_12607);
nand U15074 (N_15074,N_12392,N_12887);
and U15075 (N_15075,N_13152,N_12486);
xnor U15076 (N_15076,N_12397,N_11904);
nand U15077 (N_15077,N_14366,N_12997);
and U15078 (N_15078,N_14090,N_13577);
or U15079 (N_15079,N_13528,N_13828);
nor U15080 (N_15080,N_10223,N_13580);
nor U15081 (N_15081,N_10329,N_12198);
and U15082 (N_15082,N_11754,N_11576);
nand U15083 (N_15083,N_13804,N_11730);
or U15084 (N_15084,N_11363,N_12430);
or U15085 (N_15085,N_11756,N_10616);
or U15086 (N_15086,N_11898,N_11219);
or U15087 (N_15087,N_13790,N_13554);
and U15088 (N_15088,N_11012,N_11699);
or U15089 (N_15089,N_11686,N_11666);
and U15090 (N_15090,N_10297,N_10972);
and U15091 (N_15091,N_13288,N_14142);
or U15092 (N_15092,N_10405,N_13450);
nand U15093 (N_15093,N_11225,N_11931);
nor U15094 (N_15094,N_10360,N_12833);
and U15095 (N_15095,N_14602,N_14903);
nand U15096 (N_15096,N_10821,N_12102);
nand U15097 (N_15097,N_12559,N_13781);
or U15098 (N_15098,N_11782,N_13882);
and U15099 (N_15099,N_13023,N_10144);
and U15100 (N_15100,N_10030,N_14745);
or U15101 (N_15101,N_14280,N_13012);
nor U15102 (N_15102,N_12380,N_10544);
or U15103 (N_15103,N_10294,N_14027);
xnor U15104 (N_15104,N_10669,N_10740);
xor U15105 (N_15105,N_10678,N_11436);
or U15106 (N_15106,N_13482,N_12158);
and U15107 (N_15107,N_11577,N_12524);
and U15108 (N_15108,N_10760,N_12020);
and U15109 (N_15109,N_14421,N_14469);
nand U15110 (N_15110,N_11068,N_14630);
nand U15111 (N_15111,N_13714,N_13242);
nor U15112 (N_15112,N_11622,N_11335);
or U15113 (N_15113,N_11369,N_14095);
and U15114 (N_15114,N_13838,N_13348);
or U15115 (N_15115,N_12072,N_11184);
nand U15116 (N_15116,N_11464,N_10230);
xor U15117 (N_15117,N_12796,N_10509);
xor U15118 (N_15118,N_11065,N_14309);
xor U15119 (N_15119,N_10855,N_12747);
or U15120 (N_15120,N_12662,N_10533);
nor U15121 (N_15121,N_10692,N_14120);
nand U15122 (N_15122,N_11738,N_14567);
or U15123 (N_15123,N_12016,N_12991);
nand U15124 (N_15124,N_12558,N_11679);
nand U15125 (N_15125,N_13355,N_14299);
nor U15126 (N_15126,N_12159,N_14793);
and U15127 (N_15127,N_10700,N_13994);
nand U15128 (N_15128,N_12071,N_13414);
and U15129 (N_15129,N_12280,N_10026);
xnor U15130 (N_15130,N_14091,N_12096);
and U15131 (N_15131,N_10989,N_13864);
nor U15132 (N_15132,N_11723,N_10474);
or U15133 (N_15133,N_10991,N_12584);
xor U15134 (N_15134,N_10852,N_12544);
and U15135 (N_15135,N_14546,N_13261);
xnor U15136 (N_15136,N_12270,N_11372);
nor U15137 (N_15137,N_11395,N_11088);
xnor U15138 (N_15138,N_14237,N_10809);
nor U15139 (N_15139,N_12785,N_13208);
xor U15140 (N_15140,N_14576,N_12748);
and U15141 (N_15141,N_14653,N_14029);
and U15142 (N_15142,N_13850,N_10521);
or U15143 (N_15143,N_11536,N_11378);
and U15144 (N_15144,N_13048,N_10248);
or U15145 (N_15145,N_14058,N_14075);
nor U15146 (N_15146,N_12580,N_14396);
and U15147 (N_15147,N_13228,N_12382);
nand U15148 (N_15148,N_13576,N_11217);
nand U15149 (N_15149,N_10818,N_13755);
nand U15150 (N_15150,N_10677,N_10167);
and U15151 (N_15151,N_11751,N_14485);
or U15152 (N_15152,N_13454,N_13262);
xor U15153 (N_15153,N_10377,N_14661);
xnor U15154 (N_15154,N_12468,N_13485);
xnor U15155 (N_15155,N_11262,N_12929);
xnor U15156 (N_15156,N_12032,N_14113);
xnor U15157 (N_15157,N_10439,N_10850);
xor U15158 (N_15158,N_12973,N_10104);
or U15159 (N_15159,N_10602,N_14216);
nand U15160 (N_15160,N_11570,N_12540);
nand U15161 (N_15161,N_13291,N_14998);
and U15162 (N_15162,N_11535,N_11853);
xnor U15163 (N_15163,N_12701,N_12051);
nand U15164 (N_15164,N_12187,N_11627);
nor U15165 (N_15165,N_10331,N_13601);
xnor U15166 (N_15166,N_13832,N_13535);
or U15167 (N_15167,N_14874,N_14315);
or U15168 (N_15168,N_10306,N_10607);
nand U15169 (N_15169,N_11505,N_12868);
nand U15170 (N_15170,N_12946,N_13950);
or U15171 (N_15171,N_11470,N_11719);
and U15172 (N_15172,N_14345,N_12452);
and U15173 (N_15173,N_12147,N_12465);
nor U15174 (N_15174,N_14581,N_11935);
nand U15175 (N_15175,N_14966,N_14488);
xor U15176 (N_15176,N_11709,N_10658);
or U15177 (N_15177,N_12971,N_10550);
nand U15178 (N_15178,N_11102,N_11544);
xnor U15179 (N_15179,N_12789,N_11787);
nand U15180 (N_15180,N_13924,N_10252);
and U15181 (N_15181,N_13774,N_11462);
and U15182 (N_15182,N_14431,N_10898);
nor U15183 (N_15183,N_10871,N_12444);
nand U15184 (N_15184,N_12319,N_11506);
and U15185 (N_15185,N_10125,N_10681);
or U15186 (N_15186,N_11166,N_14428);
and U15187 (N_15187,N_13407,N_14583);
and U15188 (N_15188,N_12369,N_12117);
nor U15189 (N_15189,N_14036,N_12707);
nand U15190 (N_15190,N_10895,N_11650);
and U15191 (N_15191,N_11866,N_11024);
nor U15192 (N_15192,N_13923,N_11342);
and U15193 (N_15193,N_13229,N_11909);
or U15194 (N_15194,N_10367,N_11701);
and U15195 (N_15195,N_13791,N_14646);
or U15196 (N_15196,N_14070,N_12669);
nand U15197 (N_15197,N_10584,N_10565);
xnor U15198 (N_15198,N_10307,N_11553);
and U15199 (N_15199,N_12440,N_14687);
and U15200 (N_15200,N_13278,N_14395);
nand U15201 (N_15201,N_10471,N_12548);
and U15202 (N_15202,N_10660,N_14691);
nor U15203 (N_15203,N_11906,N_11094);
nand U15204 (N_15204,N_11207,N_10917);
and U15205 (N_15205,N_12283,N_14462);
or U15206 (N_15206,N_10534,N_10081);
or U15207 (N_15207,N_14704,N_14715);
nor U15208 (N_15208,N_10824,N_10158);
xor U15209 (N_15209,N_10015,N_13929);
nand U15210 (N_15210,N_12981,N_11408);
xnor U15211 (N_15211,N_14479,N_12492);
and U15212 (N_15212,N_11264,N_12732);
nand U15213 (N_15213,N_10668,N_13326);
or U15214 (N_15214,N_14484,N_12671);
and U15215 (N_15215,N_10718,N_14802);
nand U15216 (N_15216,N_14886,N_10772);
or U15217 (N_15217,N_10285,N_10108);
or U15218 (N_15218,N_11446,N_10139);
and U15219 (N_15219,N_11221,N_11864);
nor U15220 (N_15220,N_10756,N_10489);
or U15221 (N_15221,N_10549,N_11240);
xnor U15222 (N_15222,N_13602,N_10399);
and U15223 (N_15223,N_12362,N_10043);
or U15224 (N_15224,N_10354,N_13178);
nand U15225 (N_15225,N_11347,N_10627);
and U15226 (N_15226,N_12140,N_12594);
or U15227 (N_15227,N_12474,N_11897);
xor U15228 (N_15228,N_12568,N_12359);
nor U15229 (N_15229,N_11048,N_13044);
nor U15230 (N_15230,N_14580,N_10919);
or U15231 (N_15231,N_14818,N_13729);
nor U15232 (N_15232,N_13595,N_14424);
nor U15233 (N_15233,N_11238,N_11846);
xor U15234 (N_15234,N_12400,N_13316);
and U15235 (N_15235,N_14520,N_10333);
xnor U15236 (N_15236,N_12509,N_11035);
nand U15237 (N_15237,N_12145,N_12402);
nor U15238 (N_15238,N_13213,N_12363);
nand U15239 (N_15239,N_12749,N_10169);
xor U15240 (N_15240,N_11290,N_10473);
nand U15241 (N_15241,N_10136,N_12448);
and U15242 (N_15242,N_10918,N_14304);
or U15243 (N_15243,N_10336,N_10455);
or U15244 (N_15244,N_10872,N_12123);
nor U15245 (N_15245,N_14413,N_10930);
xor U15246 (N_15246,N_14757,N_14868);
nor U15247 (N_15247,N_11814,N_14898);
and U15248 (N_15248,N_13233,N_11821);
nand U15249 (N_15249,N_13701,N_12293);
xor U15250 (N_15250,N_11800,N_12910);
and U15251 (N_15251,N_10281,N_13342);
or U15252 (N_15252,N_13782,N_12620);
nand U15253 (N_15253,N_12304,N_11081);
nand U15254 (N_15254,N_13905,N_10292);
xnor U15255 (N_15255,N_14012,N_10430);
nand U15256 (N_15256,N_13553,N_14429);
or U15257 (N_15257,N_13708,N_12944);
and U15258 (N_15258,N_11836,N_12995);
xnor U15259 (N_15259,N_14124,N_10123);
or U15260 (N_15260,N_12821,N_10902);
nor U15261 (N_15261,N_10840,N_10596);
xor U15262 (N_15262,N_12472,N_10613);
and U15263 (N_15263,N_10142,N_13557);
nor U15264 (N_15264,N_13312,N_12848);
and U15265 (N_15265,N_10379,N_10813);
or U15266 (N_15266,N_10558,N_14418);
or U15267 (N_15267,N_13787,N_13978);
or U15268 (N_15268,N_10308,N_10433);
xor U15269 (N_15269,N_10887,N_11947);
nor U15270 (N_15270,N_10319,N_14777);
xnor U15271 (N_15271,N_13732,N_14972);
and U15272 (N_15272,N_12510,N_14496);
or U15273 (N_15273,N_14132,N_14221);
xor U15274 (N_15274,N_11959,N_14635);
or U15275 (N_15275,N_12719,N_14823);
and U15276 (N_15276,N_12196,N_10274);
xor U15277 (N_15277,N_11932,N_12697);
and U15278 (N_15278,N_11859,N_10422);
xor U15279 (N_15279,N_14302,N_14836);
nand U15280 (N_15280,N_11565,N_14261);
nor U15281 (N_15281,N_12069,N_10827);
nand U15282 (N_15282,N_10579,N_12600);
or U15283 (N_15283,N_11162,N_13142);
nand U15284 (N_15284,N_10680,N_10176);
or U15285 (N_15285,N_11438,N_14674);
nand U15286 (N_15286,N_12317,N_10854);
nand U15287 (N_15287,N_11244,N_10012);
and U15288 (N_15288,N_14681,N_14541);
xnor U15289 (N_15289,N_11343,N_13368);
and U15290 (N_15290,N_11900,N_10040);
or U15291 (N_15291,N_12156,N_14782);
and U15292 (N_15292,N_11818,N_13592);
and U15293 (N_15293,N_14181,N_13220);
or U15294 (N_15294,N_10996,N_13131);
nor U15295 (N_15295,N_11925,N_11720);
nor U15296 (N_15296,N_12136,N_13661);
xor U15297 (N_15297,N_12921,N_12387);
nor U15298 (N_15298,N_14913,N_13547);
nand U15299 (N_15299,N_12375,N_10894);
and U15300 (N_15300,N_12213,N_13207);
nor U15301 (N_15301,N_13013,N_12045);
and U15302 (N_15302,N_12576,N_11523);
or U15303 (N_15303,N_13377,N_14391);
nor U15304 (N_15304,N_12461,N_14323);
nand U15305 (N_15305,N_14609,N_12893);
or U15306 (N_15306,N_11428,N_14867);
nand U15307 (N_15307,N_12146,N_13252);
or U15308 (N_15308,N_14781,N_11033);
or U15309 (N_15309,N_10041,N_14506);
nand U15310 (N_15310,N_11987,N_12313);
nand U15311 (N_15311,N_10909,N_11868);
nand U15312 (N_15312,N_11386,N_13797);
and U15313 (N_15313,N_10174,N_12763);
or U15314 (N_15314,N_12658,N_11645);
and U15315 (N_15315,N_14059,N_10135);
nor U15316 (N_15316,N_12664,N_10914);
xnor U15317 (N_15317,N_11421,N_12011);
xor U15318 (N_15318,N_13523,N_12347);
and U15319 (N_15319,N_12681,N_14298);
nand U15320 (N_15320,N_11455,N_13789);
nor U15321 (N_15321,N_12809,N_10315);
and U15322 (N_15322,N_12204,N_11041);
nand U15323 (N_15323,N_11360,N_12459);
and U15324 (N_15324,N_12393,N_12226);
nand U15325 (N_15325,N_10611,N_13802);
xnor U15326 (N_15326,N_13632,N_12108);
or U15327 (N_15327,N_13465,N_10722);
xnor U15328 (N_15328,N_12309,N_10774);
and U15329 (N_15329,N_11625,N_13459);
and U15330 (N_15330,N_12592,N_11979);
nor U15331 (N_15331,N_13809,N_12224);
and U15332 (N_15332,N_11885,N_11556);
or U15333 (N_15333,N_13788,N_14288);
or U15334 (N_15334,N_11181,N_13122);
and U15335 (N_15335,N_11668,N_12751);
and U15336 (N_15336,N_10559,N_12877);
nand U15337 (N_15337,N_13135,N_11450);
xor U15338 (N_15338,N_14148,N_10359);
nor U15339 (N_15339,N_10983,N_12711);
nand U15340 (N_15340,N_11953,N_11763);
nor U15341 (N_15341,N_14362,N_14102);
nor U15342 (N_15342,N_10157,N_11522);
nor U15343 (N_15343,N_14416,N_12598);
xor U15344 (N_15344,N_11095,N_10153);
nor U15345 (N_15345,N_13404,N_12673);
and U15346 (N_15346,N_12884,N_10023);
nor U15347 (N_15347,N_13140,N_11323);
or U15348 (N_15348,N_11541,N_13772);
nor U15349 (N_15349,N_13860,N_10290);
nand U15350 (N_15350,N_10148,N_12804);
nor U15351 (N_15351,N_13413,N_10232);
or U15352 (N_15352,N_14814,N_13689);
xnor U15353 (N_15353,N_14458,N_11036);
xor U15354 (N_15354,N_13157,N_11891);
or U15355 (N_15355,N_11591,N_13498);
or U15356 (N_15356,N_13959,N_14785);
and U15357 (N_15357,N_10708,N_14351);
xor U15358 (N_15358,N_10007,N_10776);
nor U15359 (N_15359,N_11237,N_12070);
nor U15360 (N_15360,N_14146,N_13756);
xnor U15361 (N_15361,N_12261,N_14220);
nand U15362 (N_15362,N_13256,N_12322);
xor U15363 (N_15363,N_13292,N_13680);
or U15364 (N_15364,N_12754,N_10221);
nor U15365 (N_15365,N_12963,N_12812);
nor U15366 (N_15366,N_13445,N_14766);
xnor U15367 (N_15367,N_12954,N_12626);
nand U15368 (N_15368,N_12231,N_10721);
or U15369 (N_15369,N_13741,N_14446);
nand U15370 (N_15370,N_12630,N_14608);
or U15371 (N_15371,N_11816,N_10084);
or U15372 (N_15372,N_14667,N_14000);
or U15373 (N_15373,N_10035,N_12634);
nand U15374 (N_15374,N_14791,N_11064);
nor U15375 (N_15375,N_14816,N_10314);
nand U15376 (N_15376,N_14531,N_10633);
nand U15377 (N_15377,N_11881,N_13055);
nor U15378 (N_15378,N_14222,N_12976);
xor U15379 (N_15379,N_14414,N_11243);
and U15380 (N_15380,N_12776,N_14986);
and U15381 (N_15381,N_12989,N_10266);
nor U15382 (N_15382,N_10154,N_11642);
nor U15383 (N_15383,N_11675,N_12341);
or U15384 (N_15384,N_13362,N_13011);
nor U15385 (N_15385,N_10006,N_12481);
xnor U15386 (N_15386,N_14450,N_13399);
or U15387 (N_15387,N_11200,N_13746);
and U15388 (N_15388,N_10392,N_12260);
nand U15389 (N_15389,N_10434,N_13467);
nor U15390 (N_15390,N_12337,N_11587);
nor U15391 (N_15391,N_11497,N_10563);
nand U15392 (N_15392,N_13378,N_14805);
nor U15393 (N_15393,N_10486,N_12277);
nor U15394 (N_15394,N_12238,N_10293);
nor U15395 (N_15395,N_14597,N_13235);
xnor U15396 (N_15396,N_11322,N_10862);
or U15397 (N_15397,N_11129,N_12053);
nand U15398 (N_15398,N_11128,N_14730);
nor U15399 (N_15399,N_13126,N_14285);
nor U15400 (N_15400,N_10141,N_12619);
and U15401 (N_15401,N_10045,N_10039);
nand U15402 (N_15402,N_12281,N_13470);
and U15403 (N_15403,N_13159,N_13080);
or U15404 (N_15404,N_12455,N_13390);
and U15405 (N_15405,N_12890,N_11525);
xnor U15406 (N_15406,N_11390,N_12646);
xnor U15407 (N_15407,N_14154,N_12177);
xor U15408 (N_15408,N_10580,N_11174);
or U15409 (N_15409,N_13848,N_10724);
xor U15410 (N_15410,N_13438,N_14572);
nor U15411 (N_15411,N_14420,N_10402);
and U15412 (N_15412,N_12727,N_14474);
xor U15413 (N_15413,N_12036,N_10755);
nor U15414 (N_15414,N_10072,N_12494);
or U15415 (N_15415,N_10177,N_12487);
or U15416 (N_15416,N_10966,N_12659);
nor U15417 (N_15417,N_10363,N_12314);
or U15418 (N_15418,N_14639,N_10632);
nand U15419 (N_15419,N_12935,N_14566);
xnor U15420 (N_15420,N_14069,N_13452);
or U15421 (N_15421,N_11602,N_14009);
nor U15422 (N_15422,N_11107,N_13678);
and U15423 (N_15423,N_11735,N_10566);
nor U15424 (N_15424,N_12451,N_11008);
nand U15425 (N_15425,N_13890,N_13700);
xnor U15426 (N_15426,N_12133,N_13975);
and U15427 (N_15427,N_12699,N_12447);
nand U15428 (N_15428,N_11314,N_12818);
nor U15429 (N_15429,N_14697,N_11739);
nor U15430 (N_15430,N_14379,N_13628);
xor U15431 (N_15431,N_11996,N_12018);
nor U15432 (N_15432,N_12964,N_13918);
and U15433 (N_15433,N_13087,N_14369);
and U15434 (N_15434,N_14314,N_11119);
and U15435 (N_15435,N_14025,N_11146);
or U15436 (N_15436,N_11376,N_14270);
or U15437 (N_15437,N_10372,N_14321);
nand U15438 (N_15438,N_13515,N_11940);
nand U15439 (N_15439,N_10107,N_11116);
xnor U15440 (N_15440,N_12581,N_13329);
xor U15441 (N_15441,N_13143,N_13879);
nor U15442 (N_15442,N_10665,N_11605);
and U15443 (N_15443,N_14563,N_14437);
xor U15444 (N_15444,N_12729,N_10131);
and U15445 (N_15445,N_13422,N_11942);
nor U15446 (N_15446,N_13107,N_12957);
or U15447 (N_15447,N_12235,N_12230);
or U15448 (N_15448,N_13589,N_13673);
nand U15449 (N_15449,N_14940,N_10697);
and U15450 (N_15450,N_11952,N_14929);
nand U15451 (N_15451,N_13793,N_14751);
nand U15452 (N_15452,N_11626,N_11669);
xor U15453 (N_15453,N_10408,N_12253);
or U15454 (N_15454,N_11430,N_13394);
xnor U15455 (N_15455,N_11911,N_14210);
or U15456 (N_15456,N_11230,N_13743);
or U15457 (N_15457,N_13636,N_12650);
and U15458 (N_15458,N_10370,N_11972);
and U15459 (N_15459,N_11729,N_11380);
nand U15460 (N_15460,N_14834,N_13433);
nand U15461 (N_15461,N_13725,N_10688);
xor U15462 (N_15462,N_11632,N_11362);
nor U15463 (N_15463,N_10373,N_13806);
xnor U15464 (N_15464,N_13110,N_13927);
xor U15465 (N_15465,N_13093,N_10487);
and U15466 (N_15466,N_14460,N_12292);
nand U15467 (N_15467,N_10931,N_12705);
nor U15468 (N_15468,N_11691,N_12516);
and U15469 (N_15469,N_14544,N_14204);
nand U15470 (N_15470,N_11755,N_11848);
nor U15471 (N_15471,N_10126,N_11545);
or U15472 (N_15472,N_11677,N_12582);
xnor U15473 (N_15473,N_14939,N_11757);
nand U15474 (N_15474,N_13150,N_13600);
nand U15475 (N_15475,N_10089,N_12913);
and U15476 (N_15476,N_14441,N_11603);
and U15477 (N_15477,N_14605,N_11265);
or U15478 (N_15478,N_10526,N_12039);
nor U15479 (N_15479,N_13408,N_11580);
nand U15480 (N_15480,N_10949,N_14480);
nand U15481 (N_15481,N_10053,N_11191);
nand U15482 (N_15482,N_12644,N_10298);
xnor U15483 (N_15483,N_11399,N_12786);
nand U15484 (N_15484,N_14253,N_12118);
nand U15485 (N_15485,N_14558,N_12175);
or U15486 (N_15486,N_13133,N_12386);
nand U15487 (N_15487,N_11899,N_14131);
nand U15488 (N_15488,N_10517,N_11798);
and U15489 (N_15489,N_12065,N_13308);
xor U15490 (N_15490,N_13430,N_13519);
nand U15491 (N_15491,N_10767,N_14086);
and U15492 (N_15492,N_13166,N_14108);
xor U15493 (N_15493,N_14650,N_13983);
and U15494 (N_15494,N_13499,N_14974);
nand U15495 (N_15495,N_14957,N_13249);
and U15496 (N_15496,N_10667,N_13129);
nand U15497 (N_15497,N_10215,N_14843);
nand U15498 (N_15498,N_10686,N_14213);
and U15499 (N_15499,N_12885,N_10865);
and U15500 (N_15500,N_14728,N_11053);
nor U15501 (N_15501,N_10102,N_12506);
xnor U15502 (N_15502,N_12267,N_12022);
xnor U15503 (N_15503,N_10552,N_14515);
nand U15504 (N_15504,N_13112,N_10162);
and U15505 (N_15505,N_11070,N_12041);
nor U15506 (N_15506,N_14466,N_11211);
and U15507 (N_15507,N_11529,N_11027);
xnor U15508 (N_15508,N_13964,N_10021);
xnor U15509 (N_15509,N_10357,N_12907);
xnor U15510 (N_15510,N_14177,N_10807);
nor U15511 (N_15511,N_14208,N_12284);
nand U15512 (N_15512,N_12120,N_10743);
nor U15513 (N_15513,N_14349,N_10973);
and U15514 (N_15514,N_11831,N_11612);
nand U15515 (N_15515,N_11158,N_13040);
nor U15516 (N_15516,N_14811,N_11938);
nand U15517 (N_15517,N_10256,N_10537);
nor U15518 (N_15518,N_12325,N_12826);
xor U15519 (N_15519,N_14168,N_11640);
and U15520 (N_15520,N_12040,N_13397);
nor U15521 (N_15521,N_11703,N_14801);
nand U15522 (N_15522,N_13736,N_10725);
nand U15523 (N_15523,N_12859,N_14410);
nand U15524 (N_15524,N_12398,N_10085);
nand U15525 (N_15525,N_10245,N_13079);
nor U15526 (N_15526,N_13984,N_11569);
and U15527 (N_15527,N_12614,N_14409);
nor U15528 (N_15528,N_13359,N_14186);
nor U15529 (N_15529,N_12176,N_14382);
nand U15530 (N_15530,N_12107,N_11133);
nor U15531 (N_15531,N_12531,N_12374);
and U15532 (N_15532,N_12585,N_12256);
xor U15533 (N_15533,N_11209,N_10192);
nand U15534 (N_15534,N_14692,N_13282);
and U15535 (N_15535,N_14953,N_13317);
nor U15536 (N_15536,N_14968,N_13704);
nor U15537 (N_15537,N_13552,N_14830);
and U15538 (N_15538,N_10710,N_14188);
xnor U15539 (N_15539,N_11021,N_13720);
or U15540 (N_15540,N_13775,N_14579);
and U15541 (N_15541,N_11246,N_13718);
nor U15542 (N_15542,N_11708,N_13175);
nand U15543 (N_15543,N_12167,N_14007);
or U15544 (N_15544,N_14087,N_11637);
nor U15545 (N_15545,N_12952,N_12460);
or U15546 (N_15546,N_10662,N_14083);
or U15547 (N_15547,N_11796,N_11748);
nor U15548 (N_15548,N_13878,N_12403);
nor U15549 (N_15549,N_10569,N_14862);
and U15550 (N_15550,N_10720,N_12218);
xor U15551 (N_15551,N_12490,N_12399);
and U15552 (N_15552,N_13768,N_12377);
or U15553 (N_15553,N_12038,N_11649);
nand U15554 (N_15554,N_11279,N_14890);
and U15555 (N_15555,N_13873,N_10560);
nand U15556 (N_15556,N_14195,N_13227);
or U15557 (N_15557,N_12712,N_12932);
xor U15558 (N_15558,N_12810,N_14127);
or U15559 (N_15559,N_12024,N_14164);
nor U15560 (N_15560,N_10418,N_13981);
xnor U15561 (N_15561,N_13551,N_12523);
nor U15562 (N_15562,N_13202,N_13922);
xor U15563 (N_15563,N_11283,N_10656);
xor U15564 (N_15564,N_13588,N_12476);
or U15565 (N_15565,N_11052,N_14130);
nor U15566 (N_15566,N_10382,N_10113);
or U15567 (N_15567,N_13590,N_10097);
xor U15568 (N_15568,N_14332,N_12596);
and U15569 (N_15569,N_14622,N_13200);
or U15570 (N_15570,N_14916,N_11198);
and U15571 (N_15571,N_11375,N_10540);
nor U15572 (N_15572,N_14753,N_14921);
xor U15573 (N_15573,N_11977,N_11773);
xor U15574 (N_15574,N_12252,N_13779);
nor U15575 (N_15575,N_10670,N_13398);
nand U15576 (N_15576,N_11471,N_12526);
nor U15577 (N_15577,N_12811,N_10034);
and U15578 (N_15578,N_10013,N_12410);
nor U15579 (N_15579,N_11031,N_12654);
and U15580 (N_15580,N_10539,N_12379);
xnor U15581 (N_15581,N_10068,N_11539);
or U15582 (N_15582,N_13962,N_12415);
nand U15583 (N_15583,N_11352,N_14386);
xor U15584 (N_15584,N_10477,N_10062);
xnor U15585 (N_15585,N_14350,N_11934);
nand U15586 (N_15586,N_14535,N_14557);
xor U15587 (N_15587,N_10376,N_12099);
nand U15588 (N_15588,N_10150,N_13258);
xnor U15589 (N_15589,N_12349,N_14554);
and U15590 (N_15590,N_13353,N_11946);
or U15591 (N_15591,N_10591,N_14870);
or U15592 (N_15592,N_12285,N_12229);
xnor U15593 (N_15593,N_14367,N_11673);
nand U15594 (N_15594,N_13183,N_14550);
or U15595 (N_15595,N_11617,N_14673);
nand U15596 (N_15596,N_10186,N_12219);
xor U15597 (N_15597,N_11657,N_12622);
nand U15598 (N_15598,N_10096,N_11753);
nand U15599 (N_15599,N_13961,N_11955);
and U15600 (N_15600,N_10646,N_11770);
xnor U15601 (N_15601,N_11875,N_14909);
and U15602 (N_15602,N_11113,N_14822);
or U15603 (N_15603,N_10317,N_12358);
and U15604 (N_15604,N_11171,N_12263);
or U15605 (N_15605,N_10318,N_14804);
xnor U15606 (N_15606,N_10603,N_14902);
xnor U15607 (N_15607,N_10398,N_11419);
nor U15608 (N_15608,N_14928,N_11298);
and U15609 (N_15609,N_10586,N_11377);
xnor U15610 (N_15610,N_11533,N_14227);
xor U15611 (N_15611,N_12835,N_12625);
xor U15612 (N_15612,N_14423,N_12212);
or U15613 (N_15613,N_11253,N_10181);
or U15614 (N_15614,N_10019,N_13645);
nor U15615 (N_15615,N_13480,N_12518);
or U15616 (N_15616,N_11604,N_12499);
nand U15617 (N_15617,N_14085,N_12898);
or U15618 (N_15618,N_11801,N_13409);
xor U15619 (N_15619,N_11697,N_13443);
nor U15620 (N_15620,N_12383,N_10339);
and U15621 (N_15621,N_13786,N_14258);
nand U15622 (N_15622,N_12653,N_10815);
or U15623 (N_15623,N_14039,N_13197);
and U15624 (N_15624,N_11100,N_12908);
xnor U15625 (N_15625,N_13696,N_11954);
xnor U15626 (N_15626,N_13302,N_11862);
xnor U15627 (N_15627,N_13295,N_10371);
nor U15628 (N_15628,N_12865,N_12766);
and U15629 (N_15629,N_10661,N_13198);
nand U15630 (N_15630,N_14894,N_12409);
nand U15631 (N_15631,N_11272,N_13582);
nor U15632 (N_15632,N_11744,N_14670);
or U15633 (N_15633,N_10998,N_13761);
nor U15634 (N_15634,N_11137,N_13889);
xor U15635 (N_15635,N_10780,N_11877);
and U15636 (N_15636,N_12205,N_13260);
and U15637 (N_15637,N_13655,N_13211);
xor U15638 (N_15638,N_12453,N_10829);
or U15639 (N_15639,N_10648,N_13163);
nor U15640 (N_15640,N_13125,N_13286);
nor U15641 (N_15641,N_13475,N_10819);
xnor U15642 (N_15642,N_11694,N_11160);
nand U15643 (N_15643,N_13405,N_14530);
nand U15644 (N_15644,N_10938,N_13403);
xor U15645 (N_15645,N_13340,N_14992);
or U15646 (N_15646,N_10853,N_11620);
nand U15647 (N_15647,N_11676,N_11267);
and U15648 (N_15648,N_13682,N_13649);
xor U15649 (N_15649,N_14675,N_14788);
nor U15650 (N_15650,N_13104,N_13710);
xnor U15651 (N_15651,N_14881,N_10737);
xor U15652 (N_15652,N_14708,N_11190);
nand U15653 (N_15653,N_14393,N_11944);
nand U15654 (N_15654,N_12597,N_13357);
or U15655 (N_15655,N_12591,N_14809);
nand U15656 (N_15656,N_14399,N_14311);
and U15657 (N_15657,N_12160,N_13062);
nand U15658 (N_15658,N_13560,N_13097);
xor U15659 (N_15659,N_13224,N_14246);
xnor U15660 (N_15660,N_10403,N_10445);
or U15661 (N_15661,N_10170,N_13418);
xnor U15662 (N_15662,N_12424,N_12756);
and U15663 (N_15663,N_13641,N_11549);
or U15664 (N_15664,N_12203,N_14319);
and U15665 (N_15665,N_11828,N_10773);
or U15666 (N_15666,N_13834,N_10927);
xnor U15667 (N_15667,N_10312,N_13637);
and U15668 (N_15668,N_11289,N_14604);
nand U15669 (N_15669,N_10243,N_13222);
nand U15670 (N_15670,N_12004,N_11985);
nor U15671 (N_15671,N_13966,N_11495);
nor U15672 (N_15672,N_14370,N_14093);
and U15673 (N_15673,N_10683,N_14243);
xor U15674 (N_15674,N_12228,N_10783);
nor U15675 (N_15675,N_13766,N_12463);
and U15676 (N_15676,N_10187,N_14997);
or U15677 (N_15677,N_14570,N_12477);
nand U15678 (N_15678,N_12560,N_14762);
xor U15679 (N_15679,N_11051,N_10110);
nor U15680 (N_15680,N_11582,N_11874);
nand U15681 (N_15681,N_14754,N_14385);
nor U15682 (N_15682,N_11614,N_11305);
xnor U15683 (N_15683,N_12849,N_13821);
and U15684 (N_15684,N_12894,N_14774);
or U15685 (N_15685,N_11341,N_14672);
xor U15686 (N_15686,N_14628,N_11030);
nor U15687 (N_15687,N_12575,N_11771);
xnor U15688 (N_15688,N_10190,N_12791);
or U15689 (N_15689,N_11537,N_14092);
xnor U15690 (N_15690,N_10707,N_12923);
xor U15691 (N_15691,N_14397,N_12063);
xor U15692 (N_15692,N_11418,N_13870);
xnor U15693 (N_15693,N_11379,N_11026);
nor U15694 (N_15694,N_12469,N_12864);
nor U15695 (N_15695,N_13313,N_14585);
nand U15696 (N_15696,N_12645,N_12479);
xnor U15697 (N_15697,N_10067,N_12371);
xnor U15698 (N_15698,N_11750,N_10806);
nor U15699 (N_15699,N_11254,N_13046);
nor U15700 (N_15700,N_12174,N_14676);
nor U15701 (N_15701,N_12950,N_11354);
xnor U15702 (N_15702,N_13541,N_12850);
nor U15703 (N_15703,N_14153,N_10063);
nor U15704 (N_15704,N_12009,N_14945);
or U15705 (N_15705,N_13172,N_13501);
nor U15706 (N_15706,N_12866,N_12296);
nor U15707 (N_15707,N_12744,N_10936);
nor U15708 (N_15708,N_14456,N_12344);
or U15709 (N_15709,N_13009,N_12982);
nand U15710 (N_15710,N_14252,N_13384);
and U15711 (N_15711,N_12361,N_12760);
or U15712 (N_15712,N_14912,N_14983);
nor U15713 (N_15713,N_10410,N_11177);
and U15714 (N_15714,N_11894,N_14357);
and U15715 (N_15715,N_12642,N_14218);
or U15716 (N_15716,N_11725,N_14738);
or U15717 (N_15717,N_12470,N_10327);
or U15718 (N_15718,N_12953,N_13734);
and U15719 (N_15719,N_12975,N_13026);
nor U15720 (N_15720,N_12794,N_14833);
nor U15721 (N_15721,N_14812,N_11079);
nand U15722 (N_15722,N_13029,N_12886);
nand U15723 (N_15723,N_14101,N_10017);
or U15724 (N_15724,N_14269,N_10615);
and U15725 (N_15725,N_13339,N_12924);
or U15726 (N_15726,N_11109,N_10269);
or U15727 (N_15727,N_14850,N_14401);
or U15728 (N_15728,N_12892,N_13280);
xor U15729 (N_15729,N_13669,N_13204);
nand U15730 (N_15730,N_10846,N_13000);
xor U15731 (N_15731,N_11004,N_11971);
nand U15732 (N_15732,N_11867,N_11213);
and U15733 (N_15733,N_14908,N_12093);
and U15734 (N_15734,N_14135,N_11766);
and U15735 (N_15735,N_14247,N_12148);
xor U15736 (N_15736,N_13245,N_10556);
and U15737 (N_15737,N_10567,N_11978);
xor U15738 (N_15738,N_12273,N_13194);
or U15739 (N_15739,N_10500,N_13325);
nand U15740 (N_15740,N_13380,N_11091);
or U15741 (N_15741,N_11108,N_14118);
xor U15742 (N_15742,N_12179,N_10283);
or U15743 (N_15743,N_10674,N_11639);
xor U15744 (N_15744,N_10165,N_14359);
xnor U15745 (N_15745,N_14888,N_10682);
xnor U15746 (N_15746,N_10739,N_13455);
nand U15747 (N_15747,N_14555,N_14248);
xnor U15748 (N_15748,N_13489,N_12968);
and U15749 (N_15749,N_13957,N_13456);
and U15750 (N_15750,N_11890,N_13875);
nand U15751 (N_15751,N_13154,N_10194);
nand U15752 (N_15752,N_11023,N_12801);
nand U15753 (N_15753,N_11361,N_10207);
nand U15754 (N_15754,N_13921,N_14336);
nand U15755 (N_15755,N_10000,N_14292);
xor U15756 (N_15756,N_13728,N_10758);
nand U15757 (N_15757,N_14950,N_14062);
and U15758 (N_15758,N_13310,N_10672);
nor U15759 (N_15759,N_13440,N_12407);
nand U15760 (N_15760,N_10826,N_12570);
or U15761 (N_15761,N_14098,N_13817);
xnor U15762 (N_15762,N_13694,N_10195);
or U15763 (N_15763,N_10993,N_12528);
nand U15764 (N_15764,N_14229,N_14404);
nand U15765 (N_15765,N_10465,N_12339);
or U15766 (N_15766,N_13967,N_14866);
xnor U15767 (N_15767,N_10304,N_11315);
and U15768 (N_15768,N_12276,N_12134);
nand U15769 (N_15769,N_11963,N_12122);
or U15770 (N_15770,N_13221,N_12110);
xnor U15771 (N_15771,N_10145,N_10590);
xor U15772 (N_15772,N_13945,N_14591);
nor U15773 (N_15773,N_12652,N_10959);
nand U15774 (N_15774,N_11278,N_14990);
nand U15775 (N_15775,N_13928,N_13393);
nand U15776 (N_15776,N_14795,N_10859);
nor U15777 (N_15777,N_14573,N_11226);
and U15778 (N_15778,N_12332,N_14517);
or U15779 (N_15779,N_12142,N_13345);
and U15780 (N_15780,N_11742,N_14961);
nand U15781 (N_15781,N_11255,N_13531);
or U15782 (N_15782,N_10709,N_12665);
xor U15783 (N_15783,N_12227,N_14952);
or U15784 (N_15784,N_11835,N_13130);
nor U15785 (N_15785,N_11772,N_14123);
and U15786 (N_15786,N_14662,N_14582);
and U15787 (N_15787,N_11276,N_10795);
nor U15788 (N_15788,N_12587,N_14882);
or U15789 (N_15789,N_10056,N_12507);
nand U15790 (N_15790,N_13615,N_12942);
nand U15791 (N_15791,N_13311,N_10644);
xnor U15792 (N_15792,N_10870,N_14536);
nand U15793 (N_15793,N_14877,N_13463);
nand U15794 (N_15794,N_14491,N_14071);
and U15795 (N_15795,N_13266,N_14899);
or U15796 (N_15796,N_10099,N_10515);
and U15797 (N_15797,N_12824,N_14141);
xor U15798 (N_15798,N_12702,N_14895);
or U15799 (N_15799,N_11706,N_14434);
nand U15800 (N_15800,N_13674,N_12125);
xnor U15801 (N_15801,N_13021,N_13690);
nand U15802 (N_15802,N_13257,N_14726);
xnor U15803 (N_15803,N_11032,N_13758);
or U15804 (N_15804,N_12977,N_12779);
nor U15805 (N_15805,N_12840,N_14334);
and U15806 (N_15806,N_10801,N_11072);
nor U15807 (N_15807,N_10699,N_10825);
or U15808 (N_15808,N_12217,N_14272);
nand U15809 (N_15809,N_10246,N_13558);
or U15810 (N_15810,N_10001,N_14171);
and U15811 (N_15811,N_11059,N_13293);
nor U15812 (N_15812,N_11989,N_11011);
xnor U15813 (N_15813,N_13795,N_12753);
nor U15814 (N_15814,N_13512,N_14329);
xnor U15815 (N_15815,N_10542,N_12168);
nor U15816 (N_15816,N_13953,N_11945);
or U15817 (N_15817,N_12986,N_11204);
nand U15818 (N_15818,N_13174,N_13191);
and U15819 (N_15819,N_12761,N_12013);
nor U15820 (N_15820,N_14347,N_11385);
and U15821 (N_15821,N_14064,N_11517);
nor U15822 (N_15822,N_13085,N_13045);
and U15823 (N_15823,N_13711,N_10886);
and U15824 (N_15824,N_13672,N_14492);
and U15825 (N_15825,N_10264,N_11664);
and U15826 (N_15826,N_12200,N_14024);
or U15827 (N_15827,N_12917,N_11743);
nor U15828 (N_15828,N_12757,N_14846);
or U15829 (N_15829,N_14575,N_14119);
or U15830 (N_15830,N_13218,N_13992);
or U15831 (N_15831,N_10218,N_12493);
or U15832 (N_15832,N_13705,N_11366);
and U15833 (N_15833,N_11929,N_12289);
or U15834 (N_15834,N_13726,N_14296);
nor U15835 (N_15835,N_10419,N_12074);
and U15836 (N_15836,N_12305,N_13603);
and U15837 (N_15837,N_10845,N_12553);
or U15838 (N_15838,N_11615,N_14937);
or U15839 (N_15839,N_10349,N_10470);
xor U15840 (N_15840,N_12549,N_10171);
or U15841 (N_15841,N_13759,N_12827);
and U15842 (N_15842,N_12366,N_14778);
nor U15843 (N_15843,N_11879,N_11496);
or U15844 (N_15844,N_12948,N_12395);
and U15845 (N_15845,N_12771,N_12373);
or U15846 (N_15846,N_14402,N_12017);
nor U15847 (N_15847,N_11601,N_13607);
nor U15848 (N_15848,N_10935,N_10951);
and U15849 (N_15849,N_11817,N_11991);
nor U15850 (N_15850,N_14324,N_13939);
or U15851 (N_15851,N_13494,N_14649);
nand U15852 (N_15852,N_10146,N_12693);
nand U15853 (N_15853,N_11114,N_14611);
nand U15854 (N_15854,N_14417,N_10957);
or U15855 (N_15855,N_12936,N_13662);
and U15856 (N_15856,N_11058,N_12909);
and U15857 (N_15857,N_10467,N_12101);
and U15858 (N_15858,N_14477,N_10112);
nor U15859 (N_15859,N_12726,N_12666);
nor U15860 (N_15860,N_13757,N_13544);
and U15861 (N_15861,N_11208,N_11045);
nand U15862 (N_15862,N_13439,N_14151);
or U15863 (N_15863,N_12922,N_12299);
nand U15864 (N_15864,N_14962,N_12321);
or U15865 (N_15865,N_14949,N_12483);
xor U15866 (N_15866,N_11075,N_11169);
xor U15867 (N_15867,N_11778,N_11662);
xnor U15868 (N_15868,N_10261,N_13617);
and U15869 (N_15869,N_12286,N_10463);
xnor U15870 (N_15870,N_12037,N_13173);
xnor U15871 (N_15871,N_14403,N_13778);
xnor U15872 (N_15872,N_12564,N_14275);
nor U15873 (N_15873,N_11936,N_12330);
nor U15874 (N_15874,N_14200,N_14637);
nand U15875 (N_15875,N_10415,N_10421);
xnor U15876 (N_15876,N_11937,N_13388);
nand U15877 (N_15877,N_12489,N_14022);
and U15878 (N_15878,N_10982,N_12491);
nor U15879 (N_15879,N_14150,N_14499);
and U15880 (N_15880,N_14040,N_12554);
and U15881 (N_15881,N_10504,N_12327);
nor U15882 (N_15882,N_10625,N_12852);
xor U15883 (N_15883,N_13457,N_13579);
nor U15884 (N_15884,N_12143,N_11077);
nor U15885 (N_15885,N_12298,N_10003);
or U15886 (N_15886,N_13514,N_10198);
nand U15887 (N_15887,N_12272,N_12307);
or U15888 (N_15888,N_10129,N_12355);
nor U15889 (N_15889,N_13321,N_14941);
or U15890 (N_15890,N_12408,N_13199);
nor U15891 (N_15891,N_13849,N_14273);
nand U15892 (N_15892,N_13561,N_11122);
or U15893 (N_15893,N_12955,N_14509);
or U15894 (N_15894,N_14454,N_11690);
or U15895 (N_15895,N_12457,N_11422);
nand U15896 (N_15896,N_14435,N_12682);
xor U15897 (N_15897,N_14079,N_10727);
or U15898 (N_15898,N_14503,N_10480);
xor U15899 (N_15899,N_13098,N_13979);
and U15900 (N_15900,N_10321,N_10652);
nor U15901 (N_15901,N_13290,N_10322);
xor U15902 (N_15902,N_14425,N_11002);
xnor U15903 (N_15903,N_13988,N_12221);
nor U15904 (N_15904,N_12933,N_14300);
xor U15905 (N_15905,N_11749,N_10091);
and U15906 (N_15906,N_12367,N_14107);
or U15907 (N_15907,N_12445,N_10713);
xor U15908 (N_15908,N_11090,N_10388);
nor U15909 (N_15909,N_12816,N_13134);
or U15910 (N_15910,N_13540,N_11003);
or U15911 (N_15911,N_14551,N_14813);
nor U15912 (N_15912,N_11140,N_13091);
xor U15913 (N_15913,N_13925,N_11665);
and U15914 (N_15914,N_14632,N_11988);
xnor U15915 (N_15915,N_11202,N_11608);
nor U15916 (N_15916,N_14657,N_12822);
xor U15917 (N_15917,N_10278,N_14982);
xor U15918 (N_15918,N_14498,N_12996);
and U15919 (N_15919,N_10033,N_10704);
xor U15920 (N_15920,N_11381,N_10302);
xor U15921 (N_15921,N_14242,N_11811);
and U15922 (N_15922,N_12220,N_13372);
nor U15923 (N_15923,N_10952,N_11651);
and U15924 (N_15924,N_13373,N_14008);
xnor U15925 (N_15925,N_11970,N_13338);
and U15926 (N_15926,N_12081,N_10628);
nor U15927 (N_15927,N_14259,N_14931);
or U15928 (N_15928,N_10044,N_10609);
xor U15929 (N_15929,N_10703,N_12775);
or U15930 (N_15930,N_10877,N_10385);
or U15931 (N_15931,N_12773,N_12062);
nand U15932 (N_15932,N_10744,N_12638);
and U15933 (N_15933,N_12047,N_13078);
or U15934 (N_15934,N_13586,N_13958);
xor U15935 (N_15935,N_11758,N_13337);
or U15936 (N_15936,N_13722,N_11224);
or U15937 (N_15937,N_13423,N_14374);
or U15938 (N_15938,N_10134,N_13253);
and U15939 (N_15939,N_11687,N_13076);
nor U15940 (N_15940,N_11528,N_10691);
or U15941 (N_15941,N_14159,N_11882);
and U15942 (N_15942,N_12006,N_10124);
or U15943 (N_15943,N_12052,N_14612);
nor U15944 (N_15944,N_12525,N_11216);
and U15945 (N_15945,N_12030,N_14959);
and U15946 (N_15946,N_11321,N_14106);
xnor U15947 (N_15947,N_11435,N_10375);
xnor U15948 (N_15948,N_10587,N_11078);
xnor U15949 (N_15949,N_12418,N_12488);
or U15950 (N_15950,N_10889,N_10472);
or U15951 (N_15951,N_12201,N_11762);
nor U15952 (N_15952,N_11807,N_10042);
xor U15953 (N_15953,N_12166,N_11813);
xor U15954 (N_15954,N_12684,N_12044);
and U15955 (N_15955,N_14668,N_14838);
or U15956 (N_15956,N_13549,N_11330);
nand U15957 (N_15957,N_14468,N_12715);
xnor U15958 (N_15958,N_14933,N_11300);
or U15959 (N_15959,N_14685,N_10541);
and U15960 (N_15960,N_10457,N_13273);
nand U15961 (N_15961,N_10127,N_10847);
xnor U15962 (N_15962,N_13141,N_14482);
xor U15963 (N_15963,N_10064,N_10994);
xor U15964 (N_15964,N_10926,N_13651);
xnor U15965 (N_15965,N_10835,N_14995);
or U15966 (N_15966,N_11869,N_11905);
and U15967 (N_15967,N_10695,N_10276);
xnor U15968 (N_15968,N_12139,N_11019);
nor U15969 (N_15969,N_11842,N_12423);
xor U15970 (N_15970,N_10495,N_14139);
nand U15971 (N_15971,N_11593,N_10857);
nor U15972 (N_15972,N_12012,N_13247);
nor U15973 (N_15973,N_12519,N_10736);
xor U15974 (N_15974,N_11466,N_11992);
nand U15975 (N_15975,N_14690,N_12294);
nor U15976 (N_15976,N_14647,N_14180);
and U15977 (N_15977,N_13241,N_12714);
nor U15978 (N_15978,N_13017,N_10093);
nand U15979 (N_15979,N_13474,N_13375);
nor U15980 (N_15980,N_13015,N_14748);
xnor U15981 (N_15981,N_14547,N_11006);
xor U15982 (N_15982,N_12417,N_10075);
nor U15983 (N_15983,N_10478,N_13381);
xor U15984 (N_15984,N_12853,N_14018);
and U15985 (N_15985,N_11980,N_12640);
nand U15986 (N_15986,N_10332,N_13283);
and U15987 (N_15987,N_10608,N_11628);
nand U15988 (N_15988,N_11520,N_13301);
or U15989 (N_15989,N_11789,N_11334);
or U15990 (N_15990,N_14043,N_11039);
nand U15991 (N_15991,N_12875,N_13344);
nor U15992 (N_15992,N_13693,N_14849);
and U15993 (N_15993,N_10766,N_14245);
or U15994 (N_15994,N_12741,N_12082);
or U15995 (N_15995,N_10595,N_13647);
and U15996 (N_15996,N_11829,N_11389);
nor U15997 (N_15997,N_12058,N_11722);
or U15998 (N_15998,N_11721,N_13562);
xor U15999 (N_15999,N_10047,N_10689);
or U16000 (N_16000,N_10990,N_14654);
or U16001 (N_16001,N_12164,N_12601);
nand U16002 (N_16002,N_12830,N_14718);
nand U16003 (N_16003,N_10346,N_14731);
nor U16004 (N_16004,N_13751,N_11475);
and U16005 (N_16005,N_11832,N_13449);
nand U16006 (N_16006,N_12326,N_11268);
or U16007 (N_16007,N_10511,N_10953);
nand U16008 (N_16008,N_14694,N_11524);
or U16009 (N_16009,N_14763,N_11968);
and U16010 (N_16010,N_10582,N_12959);
xor U16011 (N_16011,N_11883,N_13862);
or U16012 (N_16012,N_11554,N_14179);
nand U16013 (N_16013,N_12413,N_13416);
and U16014 (N_16014,N_13676,N_13594);
nand U16015 (N_16015,N_10732,N_13304);
and U16016 (N_16016,N_14225,N_11038);
nor U16017 (N_16017,N_11022,N_11926);
nand U16018 (N_16018,N_12974,N_14004);
nand U16019 (N_16019,N_10428,N_11530);
or U16020 (N_16020,N_14308,N_11588);
xnor U16021 (N_16021,N_10962,N_14011);
xnor U16022 (N_16022,N_12338,N_11429);
or U16023 (N_16023,N_13814,N_12302);
and U16024 (N_16024,N_14268,N_13777);
nor U16025 (N_16025,N_12881,N_12828);
xor U16026 (N_16026,N_13920,N_14680);
and U16027 (N_16027,N_14055,N_14219);
nand U16028 (N_16028,N_11515,N_10183);
or U16029 (N_16029,N_14969,N_12500);
nand U16030 (N_16030,N_13251,N_14290);
or U16031 (N_16031,N_14919,N_11239);
nand U16032 (N_16032,N_12232,N_10746);
or U16033 (N_16033,N_14383,N_13611);
xor U16034 (N_16034,N_11355,N_11844);
xor U16035 (N_16035,N_11803,N_11598);
nand U16036 (N_16036,N_12774,N_10975);
xnor U16037 (N_16037,N_14677,N_14089);
or U16038 (N_16038,N_10235,N_13567);
and U16039 (N_16039,N_13037,N_10792);
or U16040 (N_16040,N_12482,N_14338);
and U16041 (N_16041,N_10400,N_13210);
nand U16042 (N_16042,N_14907,N_14175);
nand U16043 (N_16043,N_12103,N_13490);
and U16044 (N_16044,N_14739,N_10771);
and U16045 (N_16045,N_11653,N_14457);
nand U16046 (N_16046,N_14826,N_14408);
or U16047 (N_16047,N_10676,N_13618);
nor U16048 (N_16048,N_14161,N_12246);
or U16049 (N_16049,N_11297,N_14832);
and U16050 (N_16050,N_12381,N_12556);
or U16051 (N_16051,N_12190,N_12687);
nand U16052 (N_16052,N_11852,N_12613);
or U16053 (N_16053,N_11550,N_14987);
xnor U16054 (N_16054,N_14527,N_12042);
or U16055 (N_16055,N_13497,N_13102);
nand U16056 (N_16056,N_11500,N_14516);
nand U16057 (N_16057,N_14109,N_13346);
nor U16058 (N_16058,N_13088,N_13639);
and U16059 (N_16059,N_11313,N_14493);
nand U16060 (N_16060,N_11461,N_11447);
nor U16061 (N_16061,N_10640,N_13970);
or U16062 (N_16062,N_11984,N_10046);
nand U16063 (N_16063,N_12919,N_14624);
or U16064 (N_16064,N_11115,N_12208);
xnor U16065 (N_16065,N_12956,N_14360);
xor U16066 (N_16066,N_14267,N_12475);
and U16067 (N_16067,N_12275,N_11788);
xnor U16068 (N_16068,N_13041,N_10119);
or U16069 (N_16069,N_11359,N_12782);
xor U16070 (N_16070,N_12562,N_11445);
nor U16071 (N_16071,N_12414,N_12767);
or U16072 (N_16072,N_10484,N_11884);
xnor U16073 (N_16073,N_14400,N_11600);
xor U16074 (N_16074,N_14856,N_13819);
nand U16075 (N_16075,N_13525,N_10066);
nand U16076 (N_16076,N_13323,N_14030);
or U16077 (N_16077,N_14746,N_12920);
nand U16078 (N_16078,N_11986,N_11930);
nor U16079 (N_16079,N_10288,N_12765);
and U16080 (N_16080,N_13305,N_14790);
nand U16081 (N_16081,N_10090,N_11696);
nand U16082 (N_16082,N_13509,N_13995);
or U16083 (N_16083,N_13747,N_10522);
or U16084 (N_16084,N_12348,N_11437);
or U16085 (N_16085,N_11976,N_10525);
nand U16086 (N_16086,N_13121,N_13089);
nand U16087 (N_16087,N_12308,N_10447);
or U16088 (N_16088,N_10778,N_14584);
and U16089 (N_16089,N_14543,N_13314);
xnor U16090 (N_16090,N_13675,N_10986);
xor U16091 (N_16091,N_13706,N_14241);
nand U16092 (N_16092,N_12428,N_13030);
nor U16093 (N_16093,N_14702,N_13203);
xnor U16094 (N_16094,N_11148,N_14236);
and U16095 (N_16095,N_11850,N_10137);
or U16096 (N_16096,N_11409,N_10779);
and U16097 (N_16097,N_14254,N_12802);
and U16098 (N_16098,N_13807,N_10967);
xnor U16099 (N_16099,N_12170,N_13350);
nand U16100 (N_16100,N_14946,N_14305);
nand U16101 (N_16101,N_12278,N_11234);
nor U16102 (N_16102,N_14002,N_11768);
nand U16103 (N_16103,N_13370,N_11281);
nor U16104 (N_16104,N_14228,N_11257);
nor U16105 (N_16105,N_12683,N_10249);
nand U16106 (N_16106,N_14914,N_14901);
or U16107 (N_16107,N_10432,N_10641);
xor U16108 (N_16108,N_14771,N_14031);
or U16109 (N_16109,N_12089,N_13366);
and U16110 (N_16110,N_10313,N_12154);
xnor U16111 (N_16111,N_14977,N_10915);
and U16112 (N_16112,N_14244,N_13998);
or U16113 (N_16113,N_10594,N_11621);
and U16114 (N_16114,N_10963,N_14266);
nand U16115 (N_16115,N_14537,N_11712);
or U16116 (N_16116,N_12426,N_10876);
or U16117 (N_16117,N_14750,N_12742);
nand U16118 (N_16118,N_12984,N_11962);
xnor U16119 (N_16119,N_14184,N_13956);
xor U16120 (N_16120,N_13671,N_14684);
nand U16121 (N_16121,N_11420,N_14312);
and U16122 (N_16122,N_14388,N_13216);
and U16123 (N_16123,N_12029,N_13926);
and U16124 (N_16124,N_13158,N_11196);
nor U16125 (N_16125,N_10671,N_13568);
xnor U16126 (N_16126,N_13906,N_14976);
or U16127 (N_16127,N_14355,N_14475);
or U16128 (N_16128,N_13625,N_10921);
and U16129 (N_16129,N_14951,N_10365);
or U16130 (N_16130,N_12401,N_13116);
nand U16131 (N_16131,N_13006,N_10413);
nand U16132 (N_16132,N_13571,N_14038);
xor U16133 (N_16133,N_12194,N_14666);
xor U16134 (N_16134,N_10130,N_14501);
or U16135 (N_16135,N_14775,N_10649);
xor U16136 (N_16136,N_14958,N_10573);
or U16137 (N_16137,N_11981,N_10839);
and U16138 (N_16138,N_10752,N_12151);
and U16139 (N_16139,N_12566,N_14857);
nor U16140 (N_16140,N_10790,N_13481);
and U16141 (N_16141,N_11374,N_10160);
xnor U16142 (N_16142,N_11502,N_13127);
nor U16143 (N_16143,N_11123,N_14965);
or U16144 (N_16144,N_11155,N_11999);
xor U16145 (N_16145,N_10856,N_11302);
and U16146 (N_16146,N_11558,N_10435);
xnor U16147 (N_16147,N_12617,N_13954);
nand U16148 (N_16148,N_11205,N_12723);
and U16149 (N_16149,N_12780,N_13703);
xnor U16150 (N_16150,N_10462,N_14779);
xor U16151 (N_16151,N_12328,N_14807);
nand U16152 (N_16152,N_12484,N_11066);
nand U16153 (N_16153,N_12257,N_13240);
nand U16154 (N_16154,N_14798,N_11050);
and U16155 (N_16155,N_11370,N_14452);
nand U16156 (N_16156,N_12857,N_13715);
xnor U16157 (N_16157,N_14876,N_10701);
nor U16158 (N_16158,N_11425,N_11599);
nor U16159 (N_16159,N_10863,N_14096);
nand U16160 (N_16160,N_13004,N_11804);
and U16161 (N_16161,N_13335,N_10161);
and U16162 (N_16162,N_14686,N_10694);
nand U16163 (N_16163,N_13867,N_13942);
or U16164 (N_16164,N_14523,N_11410);
xnor U16165 (N_16165,N_10599,N_11618);
xnor U16166 (N_16166,N_12404,N_11093);
or U16167 (N_16167,N_13008,N_10969);
or U16168 (N_16168,N_12571,N_14806);
nand U16169 (N_16169,N_13001,N_10719);
nand U16170 (N_16170,N_10369,N_12236);
or U16171 (N_16171,N_11403,N_14556);
and U16172 (N_16172,N_13688,N_13332);
and U16173 (N_16173,N_11201,N_11784);
xor U16174 (N_16174,N_12188,N_12184);
xnor U16175 (N_16175,N_12025,N_13884);
nor U16176 (N_16176,N_14533,N_14615);
or U16177 (N_16177,N_13685,N_12839);
xnor U16178 (N_16178,N_14599,N_11085);
and U16179 (N_16179,N_11413,N_13487);
xor U16180 (N_16180,N_14117,N_14390);
nor U16181 (N_16181,N_11726,N_11901);
xnor U16182 (N_16182,N_11183,N_13681);
nor U16183 (N_16183,N_13533,N_12439);
and U16184 (N_16184,N_11555,N_10121);
nand U16185 (N_16185,N_11020,N_12441);
and U16186 (N_16186,N_13391,N_10992);
nor U16187 (N_16187,N_14542,N_13188);
and U16188 (N_16188,N_10213,N_14652);
and U16189 (N_16189,N_13094,N_11105);
nand U16190 (N_16190,N_14026,N_10437);
or U16191 (N_16191,N_12237,N_12590);
or U16192 (N_16192,N_14787,N_10978);
nor U16193 (N_16193,N_14651,N_11473);
nor U16194 (N_16194,N_11044,N_13599);
nor U16195 (N_16195,N_14863,N_11142);
and U16196 (N_16196,N_10833,N_10745);
xor U16197 (N_16197,N_14289,N_12787);
or U16198 (N_16198,N_11266,N_11112);
and U16199 (N_16199,N_11250,N_14619);
nand U16200 (N_16200,N_11426,N_11433);
nand U16201 (N_16201,N_10118,N_14295);
xor U16202 (N_16202,N_11159,N_14565);
or U16203 (N_16203,N_13949,N_14614);
nor U16204 (N_16204,N_13358,N_12357);
or U16205 (N_16205,N_12906,N_10193);
or U16206 (N_16206,N_10009,N_14893);
nand U16207 (N_16207,N_10955,N_10458);
nand U16208 (N_16208,N_11132,N_14720);
and U16209 (N_16209,N_10896,N_11291);
and U16210 (N_16210,N_13148,N_10182);
and U16211 (N_16211,N_14406,N_13624);
or U16212 (N_16212,N_11073,N_11711);
and U16213 (N_16213,N_11918,N_12878);
or U16214 (N_16214,N_11228,N_12130);
nand U16215 (N_16215,N_10614,N_14964);
nand U16216 (N_16216,N_12605,N_11069);
nand U16217 (N_16217,N_12602,N_11472);
nand U16218 (N_16218,N_13656,N_12739);
nand U16219 (N_16219,N_10414,N_11659);
or U16220 (N_16220,N_12615,N_10100);
xor U16221 (N_16221,N_14384,N_13289);
xnor U16222 (N_16222,N_14224,N_14601);
or U16223 (N_16223,N_13018,N_11825);
nor U16224 (N_16224,N_10932,N_14112);
nor U16225 (N_16225,N_14301,N_14892);
nand U16226 (N_16226,N_13065,N_11414);
nand U16227 (N_16227,N_13887,N_10650);
or U16228 (N_16228,N_12059,N_13486);
or U16229 (N_16229,N_14239,N_11319);
xor U16230 (N_16230,N_11793,N_11655);
and U16231 (N_16231,N_11192,N_11270);
nor U16232 (N_16232,N_12251,N_12735);
nor U16233 (N_16233,N_11913,N_10685);
nor U16234 (N_16234,N_13695,N_11157);
nor U16235 (N_16235,N_13851,N_14330);
or U16236 (N_16236,N_14831,N_13830);
nand U16237 (N_16237,N_13542,N_14915);
xor U16238 (N_16238,N_14589,N_10054);
or U16239 (N_16239,N_13518,N_14606);
and U16240 (N_16240,N_11469,N_11492);
xnor U16241 (N_16241,N_10201,N_13016);
xnor U16242 (N_16242,N_11294,N_10659);
nand U16243 (N_16243,N_13161,N_13351);
or U16244 (N_16244,N_13986,N_13105);
or U16245 (N_16245,N_14828,N_11481);
and U16246 (N_16246,N_14197,N_11172);
or U16247 (N_16247,N_14703,N_14935);
nor U16248 (N_16248,N_12462,N_11973);
nand U16249 (N_16249,N_10092,N_11532);
nor U16250 (N_16250,N_11951,N_12320);
xnor U16251 (N_16251,N_10617,N_14773);
nand U16252 (N_16252,N_12639,N_12248);
xor U16253 (N_16253,N_10851,N_12966);
nor U16254 (N_16254,N_10505,N_10416);
or U16255 (N_16255,N_14810,N_12137);
nor U16256 (N_16256,N_12661,N_10798);
nor U16257 (N_16257,N_14076,N_14897);
xor U16258 (N_16258,N_12034,N_10789);
and U16259 (N_16259,N_11327,N_10468);
xor U16260 (N_16260,N_13111,N_10106);
xor U16261 (N_16261,N_10417,N_12254);
nor U16262 (N_16262,N_10735,N_11141);
or U16263 (N_16263,N_10491,N_12250);
nor U16264 (N_16264,N_11325,N_14411);
xor U16265 (N_16265,N_11824,N_12969);
nand U16266 (N_16266,N_11028,N_12870);
xor U16267 (N_16267,N_10696,N_10328);
nand U16268 (N_16268,N_10891,N_14176);
or U16269 (N_16269,N_11786,N_13763);
nor U16270 (N_16270,N_13049,N_12799);
nor U16271 (N_16271,N_14240,N_11067);
nor U16272 (N_16272,N_12434,N_14532);
and U16273 (N_16273,N_10420,N_10323);
nand U16274 (N_16274,N_14339,N_10816);
nor U16275 (N_16275,N_12331,N_10920);
or U16276 (N_16276,N_10384,N_11110);
nand U16277 (N_16277,N_12225,N_14238);
xor U16278 (N_16278,N_10945,N_11633);
or U16279 (N_16279,N_14235,N_10310);
nor U16280 (N_16280,N_12202,N_12005);
nand U16281 (N_16281,N_14971,N_11304);
nand U16282 (N_16282,N_13068,N_14911);
or U16283 (N_16283,N_12306,N_14160);
xor U16284 (N_16284,N_10159,N_14571);
xor U16285 (N_16285,N_12543,N_14310);
nand U16286 (N_16286,N_14724,N_12067);
xnor U16287 (N_16287,N_14449,N_12817);
or U16288 (N_16288,N_11017,N_11303);
and U16289 (N_16289,N_11040,N_12112);
xnor U16290 (N_16290,N_14065,N_13620);
xor U16291 (N_16291,N_11671,N_12717);
xnor U16292 (N_16292,N_10309,N_10626);
xnor U16293 (N_16293,N_13230,N_11241);
or U16294 (N_16294,N_10247,N_12721);
and U16295 (N_16295,N_10241,N_12947);
and U16296 (N_16296,N_10885,N_14991);
and U16297 (N_16297,N_10551,N_10705);
xnor U16298 (N_16298,N_10987,N_13177);
nor U16299 (N_16299,N_14128,N_13668);
nor U16300 (N_16300,N_10353,N_13002);
nand U16301 (N_16301,N_11329,N_12094);
or U16302 (N_16302,N_12473,N_11493);
or U16303 (N_16303,N_14640,N_11404);
nor U16304 (N_16304,N_10508,N_14344);
and U16305 (N_16305,N_12728,N_14500);
and U16306 (N_16306,N_11165,N_12068);
nand U16307 (N_16307,N_13473,N_14734);
nor U16308 (N_16308,N_10250,N_14398);
and U16309 (N_16309,N_12427,N_10277);
nor U16310 (N_16310,N_10808,N_11474);
and U16311 (N_16311,N_13982,N_11542);
nand U16312 (N_16312,N_14037,N_12513);
or U16313 (N_16313,N_14189,N_11761);
nand U16314 (N_16314,N_11009,N_13460);
xnor U16315 (N_16315,N_13539,N_12315);
or U16316 (N_16316,N_14603,N_13990);
and U16317 (N_16317,N_14072,N_11457);
nand U16318 (N_16318,N_11358,N_14143);
xnor U16319 (N_16319,N_14115,N_10728);
nand U16320 (N_16320,N_12350,N_14287);
nand U16321 (N_16321,N_10948,N_10025);
xor U16322 (N_16322,N_14710,N_11047);
nor U16323 (N_16323,N_10639,N_13762);
xor U16324 (N_16324,N_10184,N_13697);
nand U16325 (N_16325,N_14659,N_12557);
and U16326 (N_16326,N_12028,N_14041);
and U16327 (N_16327,N_11759,N_11218);
or U16328 (N_16328,N_12621,N_11566);
nor U16329 (N_16329,N_12391,N_10675);
or U16330 (N_16330,N_14887,N_12980);
nand U16331 (N_16331,N_10844,N_14461);
xor U16332 (N_16332,N_11995,N_11097);
or U16333 (N_16333,N_10631,N_12000);
and U16334 (N_16334,N_12837,N_13401);
xnor U16335 (N_16335,N_11498,N_11328);
nand U16336 (N_16336,N_14994,N_11387);
xnor U16337 (N_16337,N_13702,N_14752);
nand U16338 (N_16338,N_11927,N_10666);
nor U16339 (N_16339,N_14910,N_13101);
or U16340 (N_16340,N_13320,N_10425);
nand U16341 (N_16341,N_13859,N_13234);
nand U16342 (N_16342,N_14858,N_14440);
or U16343 (N_16343,N_13232,N_12109);
nor U16344 (N_16344,N_12583,N_14507);
xor U16345 (N_16345,N_10828,N_10103);
and U16346 (N_16346,N_12858,N_11485);
or U16347 (N_16347,N_12895,N_11993);
and U16348 (N_16348,N_13885,N_14626);
nor U16349 (N_16349,N_14465,N_10911);
and U16350 (N_16350,N_10837,N_13803);
or U16351 (N_16351,N_14904,N_11175);
xor U16352 (N_16352,N_11456,N_12104);
xor U16353 (N_16353,N_14644,N_13136);
nor U16354 (N_16354,N_11568,N_13083);
and U16355 (N_16355,N_12663,N_11480);
xnor U16356 (N_16356,N_14051,N_13985);
nand U16357 (N_16357,N_10060,N_10228);
or U16358 (N_16358,N_12820,N_13740);
xnor U16359 (N_16359,N_13748,N_12790);
and U16360 (N_16360,N_13527,N_12316);
xnor U16361 (N_16361,N_13660,N_13863);
xnor U16362 (N_16362,N_10149,N_12083);
or U16363 (N_16363,N_13903,N_11714);
and U16364 (N_16364,N_11306,N_14984);
nand U16365 (N_16365,N_14331,N_13491);
or U16366 (N_16366,N_11733,N_11779);
or U16367 (N_16367,N_11685,N_12862);
and U16368 (N_16368,N_13096,N_14817);
nand U16369 (N_16369,N_10343,N_10262);
nor U16370 (N_16370,N_11182,N_11487);
xor U16371 (N_16371,N_11149,N_13846);
nand U16372 (N_16372,N_14157,N_11956);
and U16373 (N_16373,N_14848,N_11540);
nor U16374 (N_16374,N_11299,N_10965);
and U16375 (N_16375,N_14136,N_11716);
xnor U16376 (N_16376,N_11233,N_14825);
or U16377 (N_16377,N_10679,N_14013);
nand U16378 (N_16378,N_12985,N_12003);
nand U16379 (N_16379,N_10200,N_11982);
and U16380 (N_16380,N_10884,N_11919);
or U16381 (N_16381,N_10548,N_12209);
xor U16382 (N_16382,N_13865,N_10014);
or U16383 (N_16383,N_10687,N_10492);
xnor U16384 (N_16384,N_11700,N_13654);
nand U16385 (N_16385,N_13003,N_14861);
and U16386 (N_16386,N_13367,N_11317);
nor U16387 (N_16387,N_10240,N_10929);
and U16388 (N_16388,N_10553,N_13898);
or U16389 (N_16389,N_10796,N_13563);
nor U16390 (N_16390,N_12431,N_13108);
xnor U16391 (N_16391,N_13931,N_12836);
or U16392 (N_16392,N_14740,N_11746);
and U16393 (N_16393,N_12416,N_10204);
xnor U16394 (N_16394,N_12508,N_14819);
and U16395 (N_16395,N_14955,N_10481);
xor U16396 (N_16396,N_10386,N_10337);
or U16397 (N_16397,N_14481,N_13056);
xor U16398 (N_16398,N_11427,N_14707);
or U16399 (N_16399,N_10574,N_13425);
nand U16400 (N_16400,N_10940,N_10812);
nor U16401 (N_16401,N_10910,N_13279);
nor U16402 (N_16402,N_14104,N_10513);
and U16403 (N_16403,N_13155,N_14552);
nor U16404 (N_16404,N_14205,N_13318);
nand U16405 (N_16405,N_13269,N_14464);
nand U16406 (N_16406,N_10185,N_13471);
nor U16407 (N_16407,N_12245,N_13912);
and U16408 (N_16408,N_10562,N_13997);
nand U16409 (N_16409,N_11406,N_12677);
nand U16410 (N_16410,N_12435,N_14044);
and U16411 (N_16411,N_11449,N_14074);
and U16412 (N_16412,N_10601,N_11441);
nand U16413 (N_16413,N_12565,N_10004);
xor U16414 (N_16414,N_14540,N_12266);
nand U16415 (N_16415,N_14616,N_14306);
nand U16416 (N_16416,N_11309,N_10820);
or U16417 (N_16417,N_10922,N_14017);
nor U16418 (N_16418,N_13277,N_10404);
and U16419 (N_16419,N_13845,N_13386);
or U16420 (N_16420,N_11231,N_14010);
nand U16421 (N_16421,N_11702,N_13472);
or U16422 (N_16422,N_12939,N_11046);
xnor U16423 (N_16423,N_14066,N_10485);
or U16424 (N_16424,N_13225,N_10459);
xor U16425 (N_16425,N_12931,N_10155);
or U16426 (N_16426,N_12255,N_11135);
or U16427 (N_16427,N_14820,N_14664);
nand U16428 (N_16428,N_12872,N_13770);
nand U16429 (N_16429,N_12999,N_11259);
and U16430 (N_16430,N_12856,N_13005);
and U16431 (N_16431,N_13185,N_12914);
xor U16432 (N_16432,N_14578,N_14821);
nor U16433 (N_16433,N_11967,N_13483);
or U16434 (N_16434,N_14815,N_10079);
nand U16435 (N_16435,N_13365,N_14427);
and U16436 (N_16436,N_11124,N_13419);
and U16437 (N_16437,N_12647,N_10623);
or U16438 (N_16438,N_14494,N_14765);
xnor U16439 (N_16439,N_14620,N_12144);
xnor U16440 (N_16440,N_13106,N_10168);
or U16441 (N_16441,N_13145,N_10037);
or U16442 (N_16442,N_14764,N_12819);
or U16443 (N_16443,N_10254,N_12342);
and U16444 (N_16444,N_12046,N_13243);
and U16445 (N_16445,N_13417,N_13168);
xor U16446 (N_16446,N_10770,N_10867);
or U16447 (N_16447,N_11834,N_12725);
nand U16448 (N_16448,N_10226,N_13503);
xor U16449 (N_16449,N_10503,N_12368);
xor U16450 (N_16450,N_10520,N_11658);
nor U16451 (N_16451,N_13570,N_10585);
nor U16452 (N_16452,N_10059,N_13564);
nor U16453 (N_16453,N_13007,N_11356);
and U16454 (N_16454,N_12100,N_12737);
xnor U16455 (N_16455,N_10830,N_11477);
and U16456 (N_16456,N_12023,N_11096);
or U16457 (N_16457,N_10878,N_13857);
nand U16458 (N_16458,N_14376,N_14525);
and U16459 (N_16459,N_10268,N_14942);
or U16460 (N_16460,N_13842,N_12569);
and U16461 (N_16461,N_12941,N_14453);
nand U16462 (N_16462,N_14747,N_13698);
xnor U16463 (N_16463,N_11383,N_14346);
or U16464 (N_16464,N_10988,N_11074);
xor U16465 (N_16465,N_12918,N_12514);
xor U16466 (N_16466,N_14459,N_13575);
nor U16467 (N_16467,N_10637,N_12132);
and U16468 (N_16468,N_12686,N_13371);
nor U16469 (N_16469,N_11760,N_12290);
nor U16470 (N_16470,N_11434,N_11667);
or U16471 (N_16471,N_14956,N_14769);
nor U16472 (N_16472,N_13488,N_12031);
nor U16473 (N_16473,N_13767,N_13626);
nor U16474 (N_16474,N_11223,N_13916);
and U16475 (N_16475,N_13032,N_10469);
or U16476 (N_16476,N_13412,N_11514);
xnor U16477 (N_16477,N_14166,N_12106);
nand U16478 (N_16478,N_13987,N_14938);
or U16479 (N_16479,N_11179,N_12346);
or U16480 (N_16480,N_10076,N_14262);
xor U16481 (N_16481,N_13999,N_11654);
nand U16482 (N_16482,N_11368,N_11453);
xor U16483 (N_16483,N_10706,N_13502);
nand U16484 (N_16484,N_12987,N_14736);
and U16485 (N_16485,N_10210,N_13665);
or U16486 (N_16486,N_14046,N_14759);
and U16487 (N_16487,N_10757,N_13014);
or U16488 (N_16488,N_11567,N_13356);
nor U16489 (N_16489,N_11282,N_13123);
and U16490 (N_16490,N_10114,N_14936);
nor U16491 (N_16491,N_12152,N_12648);
or U16492 (N_16492,N_12019,N_14320);
nor U16493 (N_16493,N_14019,N_11252);
nand U16494 (N_16494,N_11161,N_11764);
or U16495 (N_16495,N_13458,N_11054);
and U16496 (N_16496,N_13760,N_10341);
nor U16497 (N_16497,N_12731,N_10979);
nand U16498 (N_16498,N_13156,N_14081);
or U16499 (N_16499,N_12781,N_13349);
nor U16500 (N_16500,N_10188,N_12061);
or U16501 (N_16501,N_14593,N_10303);
xor U16502 (N_16502,N_14100,N_14521);
nand U16503 (N_16503,N_14415,N_14281);
xor U16504 (N_16504,N_10916,N_14979);
xnor U16505 (N_16505,N_12720,N_14975);
nor U16506 (N_16506,N_13429,N_10381);
nand U16507 (N_16507,N_10754,N_10087);
or U16508 (N_16508,N_12343,N_13352);
and U16509 (N_16509,N_13679,N_10189);
nor U16510 (N_16510,N_12249,N_10624);
or U16511 (N_16511,N_14033,N_10747);
nor U16512 (N_16512,N_11010,N_11187);
nor U16513 (N_16513,N_12743,N_12667);
nand U16514 (N_16514,N_14342,N_13205);
and U16515 (N_16515,N_10693,N_13963);
xnor U16516 (N_16516,N_10954,N_10280);
nand U16517 (N_16517,N_10265,N_13952);
nor U16518 (N_16518,N_13960,N_11103);
xor U16519 (N_16519,N_11840,N_12879);
or U16520 (N_16520,N_13861,N_13573);
and U16521 (N_16521,N_13808,N_11367);
and U16522 (N_16522,N_12777,N_13437);
nand U16523 (N_16523,N_12405,N_11512);
or U16524 (N_16524,N_12970,N_14121);
xor U16525 (N_16525,N_12049,N_13608);
nand U16526 (N_16526,N_13652,N_14438);
or U16527 (N_16527,N_13930,N_11892);
nand U16528 (N_16528,N_11519,N_12629);
nand U16529 (N_16529,N_12301,N_13376);
xor U16530 (N_16530,N_10436,N_14564);
nand U16531 (N_16531,N_12279,N_13910);
nand U16532 (N_16532,N_14278,N_11168);
nand U16533 (N_16533,N_11180,N_13100);
nor U16534 (N_16534,N_14028,N_14922);
nor U16535 (N_16535,N_10761,N_12573);
or U16536 (N_16536,N_14196,N_11907);
nand U16537 (N_16537,N_13856,N_10105);
and U16538 (N_16538,N_10380,N_10642);
nor U16539 (N_16539,N_13057,N_12738);
or U16540 (N_16540,N_12692,N_14265);
and U16541 (N_16541,N_13103,N_12419);
or U16542 (N_16542,N_13400,N_13657);
nor U16543 (N_16543,N_14548,N_14199);
nand U16544 (N_16544,N_12464,N_14356);
and U16545 (N_16545,N_12438,N_13117);
xor U16546 (N_16546,N_10345,N_12688);
or U16547 (N_16547,N_13114,N_14042);
xor U16548 (N_16548,N_11397,N_13385);
nor U16549 (N_16549,N_10348,N_14185);
or U16550 (N_16550,N_14284,N_12241);
or U16551 (N_16551,N_13943,N_12378);
nand U16552 (N_16552,N_14803,N_13189);
xor U16553 (N_16553,N_12165,N_13263);
xnor U16554 (N_16554,N_13420,N_13735);
nand U16555 (N_16555,N_13500,N_14061);
nand U16556 (N_16556,N_12938,N_13132);
and U16557 (N_16557,N_11101,N_11393);
nand U16558 (N_16558,N_11371,N_12027);
nand U16559 (N_16559,N_10787,N_10016);
nand U16560 (N_16560,N_12706,N_10424);
and U16561 (N_16561,N_12636,N_12928);
nor U16562 (N_16562,N_10823,N_13971);
or U16563 (N_16563,N_10684,N_11806);
xnor U16564 (N_16564,N_10078,N_10257);
nand U16565 (N_16565,N_10638,N_13996);
and U16566 (N_16566,N_10655,N_10731);
nor U16567 (N_16567,N_13663,N_11644);
nor U16568 (N_16568,N_10214,N_12606);
and U16569 (N_16569,N_13713,N_10716);
and U16570 (N_16570,N_10206,N_14327);
or U16571 (N_16571,N_13874,N_11388);
and U16572 (N_16572,N_11923,N_14430);
nor U16573 (N_16573,N_12624,N_13035);
or U16574 (N_16574,N_14445,N_13276);
or U16575 (N_16575,N_10253,N_14126);
nor U16576 (N_16576,N_11718,N_11136);
and U16577 (N_16577,N_14905,N_11491);
nand U16578 (N_16578,N_11854,N_12983);
and U16579 (N_16579,N_13259,N_10450);
xor U16580 (N_16580,N_12538,N_10397);
and U16581 (N_16581,N_14925,N_14203);
or U16582 (N_16582,N_11964,N_10645);
nand U16583 (N_16583,N_12180,N_11364);
xor U16584 (N_16584,N_10838,N_10446);
nand U16585 (N_16585,N_14077,N_11924);
xnor U16586 (N_16586,N_10912,N_10897);
xnor U16587 (N_16587,N_13820,N_12173);
and U16588 (N_16588,N_10848,N_12271);
xor U16589 (N_16589,N_12578,N_14512);
nor U16590 (N_16590,N_11548,N_10802);
nor U16591 (N_16591,N_13073,N_14631);
and U16592 (N_16592,N_12542,N_14182);
or U16593 (N_16593,N_11483,N_11463);
nand U16594 (N_16594,N_10163,N_14944);
and U16595 (N_16595,N_14088,N_10401);
xor U16596 (N_16596,N_14553,N_13801);
nor U16597 (N_16597,N_11199,N_11301);
and U16598 (N_16598,N_11326,N_10610);
or U16599 (N_16599,N_11156,N_10636);
xnor U16600 (N_16600,N_10229,N_13090);
xor U16601 (N_16601,N_14711,N_14960);
and U16602 (N_16602,N_11482,N_12635);
xnor U16603 (N_16603,N_14559,N_10765);
and U16604 (N_16604,N_11499,N_12353);
and U16605 (N_16605,N_13196,N_13387);
or U16606 (N_16606,N_10605,N_10342);
or U16607 (N_16607,N_14405,N_12703);
nand U16608 (N_16608,N_12831,N_13167);
nor U16609 (N_16609,N_14282,N_12532);
or U16610 (N_16610,N_10443,N_10374);
nor U16611 (N_16611,N_10817,N_12891);
xnor U16612 (N_16612,N_11106,N_12784);
nor U16613 (N_16613,N_10501,N_12572);
nor U16614 (N_16614,N_11423,N_12268);
or U16615 (N_16615,N_14381,N_12541);
xor U16616 (N_16616,N_13614,N_10024);
and U16617 (N_16617,N_12360,N_14629);
xor U16618 (N_16618,N_14015,N_10575);
nor U16619 (N_16619,N_12269,N_12815);
xnor U16620 (N_16620,N_10849,N_14590);
and U16621 (N_16621,N_13691,N_14049);
xor U16622 (N_16622,N_13907,N_14125);
and U16623 (N_16623,N_14663,N_14495);
and U16624 (N_16624,N_12458,N_11501);
nand U16625 (N_16625,N_13683,N_13591);
and U16626 (N_16626,N_10208,N_12537);
nor U16627 (N_16627,N_11284,N_11916);
nand U16628 (N_16628,N_11606,N_14097);
and U16629 (N_16629,N_11791,N_13530);
xor U16630 (N_16630,N_10543,N_10101);
nand U16631 (N_16631,N_13237,N_10389);
and U16632 (N_16632,N_14303,N_12994);
or U16633 (N_16633,N_13517,N_11574);
and U16634 (N_16634,N_11849,N_10205);
or U16635 (N_16635,N_14906,N_10111);
or U16636 (N_16636,N_11949,N_10804);
or U16637 (N_16637,N_10523,N_11802);
nand U16638 (N_16638,N_12432,N_10255);
nand U16639 (N_16639,N_10038,N_14361);
and U16640 (N_16640,N_12829,N_11439);
or U16641 (N_16641,N_10320,N_12354);
and U16642 (N_16642,N_13644,N_12618);
and U16643 (N_16643,N_13099,N_11440);
nor U16644 (N_16644,N_13534,N_13627);
or U16645 (N_16645,N_14879,N_14852);
or U16646 (N_16646,N_12657,N_10083);
nor U16647 (N_16647,N_12223,N_12105);
xor U16648 (N_16648,N_10199,N_13938);
or U16649 (N_16649,N_10456,N_11958);
nand U16650 (N_16650,N_14884,N_12085);
nand U16651 (N_16651,N_11611,N_12577);
or U16652 (N_16652,N_13162,N_12079);
or U16653 (N_16653,N_14883,N_10588);
and U16654 (N_16654,N_11061,N_13991);
nor U16655 (N_16655,N_14116,N_13840);
and U16656 (N_16656,N_14855,N_13052);
xor U16657 (N_16657,N_12517,N_13461);
or U16658 (N_16658,N_13464,N_10519);
xor U16659 (N_16659,N_10273,N_14756);
or U16660 (N_16660,N_14152,N_11071);
and U16661 (N_16661,N_13354,N_11872);
xor U16662 (N_16662,N_10441,N_13937);
nand U16663 (N_16663,N_13334,N_11258);
nor U16664 (N_16664,N_14808,N_11543);
or U16665 (N_16665,N_14035,N_12904);
nor U16666 (N_16666,N_12586,N_13226);
nor U16667 (N_16667,N_14264,N_12871);
and U16668 (N_16668,N_10554,N_12798);
xor U16669 (N_16669,N_14679,N_10612);
and U16670 (N_16670,N_11914,N_11643);
xor U16671 (N_16671,N_10564,N_10098);
xnor U16672 (N_16672,N_13974,N_12214);
nand U16673 (N_16673,N_10448,N_11736);
or U16674 (N_16674,N_10690,N_14032);
and U16675 (N_16675,N_11705,N_13687);
or U16676 (N_16676,N_14574,N_13451);
nand U16677 (N_16677,N_13513,N_12800);
nand U16678 (N_16678,N_11573,N_12433);
nand U16679 (N_16679,N_13737,N_14231);
nor U16680 (N_16680,N_11865,N_13972);
and U16681 (N_16681,N_14155,N_13604);
or U16682 (N_16682,N_13616,N_13192);
or U16683 (N_16683,N_12054,N_12384);
nand U16684 (N_16684,N_14023,N_13206);
nor U16685 (N_16685,N_10242,N_12672);
xor U16686 (N_16686,N_10561,N_11431);
xor U16687 (N_16687,N_14749,N_10390);
or U16688 (N_16688,N_11812,N_10899);
nand U16689 (N_16689,N_13623,N_10908);
xor U16690 (N_16690,N_11741,N_11592);
or U16691 (N_16691,N_10466,N_11346);
nor U16692 (N_16692,N_13653,N_12149);
nand U16693 (N_16693,N_12679,N_11452);
or U16694 (N_16694,N_13268,N_13187);
nand U16695 (N_16695,N_14256,N_14842);
or U16696 (N_16696,N_10197,N_14981);
xor U16697 (N_16697,N_14607,N_11062);
xor U16698 (N_16698,N_10179,N_10742);
nor U16699 (N_16699,N_11740,N_11173);
xnor U16700 (N_16700,N_10133,N_10301);
or U16701 (N_16701,N_13733,N_12593);
nor U16702 (N_16702,N_12555,N_10368);
nand U16703 (N_16703,N_10653,N_11928);
xor U16704 (N_16704,N_14865,N_10427);
and U16705 (N_16705,N_14443,N_13328);
xnor U16706 (N_16706,N_13855,N_12834);
nand U16707 (N_16707,N_12880,N_12412);
nand U16708 (N_16708,N_10461,N_12265);
nand U16709 (N_16709,N_11286,N_12813);
or U16710 (N_16710,N_13686,N_12911);
and U16711 (N_16711,N_10980,N_11247);
nor U16712 (N_16712,N_11589,N_11584);
xor U16713 (N_16713,N_12171,N_12670);
nand U16714 (N_16714,N_11295,N_11823);
xnor U16715 (N_16715,N_14444,N_14451);
xor U16716 (N_16716,N_14080,N_13724);
or U16717 (N_16717,N_14596,N_13914);
nor U16718 (N_16718,N_11661,N_12075);
nand U16719 (N_16719,N_12323,N_11139);
or U16720 (N_16720,N_12930,N_11636);
or U16721 (N_16721,N_12456,N_14973);
and U16722 (N_16722,N_11902,N_13138);
and U16723 (N_16723,N_13765,N_11960);
nor U16724 (N_16724,N_14760,N_12746);
and U16725 (N_16725,N_12239,N_13932);
nand U16726 (N_16726,N_13529,N_12943);
xor U16727 (N_16727,N_13839,N_13891);
and U16728 (N_16728,N_14368,N_11195);
nand U16729 (N_16729,N_14592,N_10071);
and U16730 (N_16730,N_11432,N_10117);
nor U16731 (N_16731,N_12077,N_13058);
nor U16732 (N_16732,N_13250,N_11777);
and U16733 (N_16733,N_10621,N_11873);
nand U16734 (N_16734,N_13900,N_12076);
or U16735 (N_16735,N_10216,N_14645);
nor U16736 (N_16736,N_11206,N_11118);
nor U16737 (N_16737,N_13664,N_10892);
or U16738 (N_16738,N_10244,N_14841);
and U16739 (N_16739,N_12795,N_14696);
xor U16740 (N_16740,N_10237,N_14528);
or U16741 (N_16741,N_14436,N_14183);
nor U16742 (N_16742,N_12876,N_14133);
nand U16743 (N_16743,N_13303,N_14594);
or U16744 (N_16744,N_14827,N_13904);
and U16745 (N_16745,N_13033,N_13190);
nor U16746 (N_16746,N_14656,N_10069);
and U16747 (N_16747,N_11151,N_13876);
xnor U16748 (N_16748,N_10535,N_14588);
and U16749 (N_16749,N_13255,N_13285);
xor U16750 (N_16750,N_13149,N_11444);
nor U16751 (N_16751,N_10764,N_13182);
nor U16752 (N_16752,N_11274,N_13581);
nor U16753 (N_16753,N_12390,N_14835);
and U16754 (N_16754,N_11188,N_14137);
or U16755 (N_16755,N_10777,N_11822);
nand U16756 (N_16756,N_12604,N_11847);
nor U16757 (N_16757,N_12696,N_10497);
and U16758 (N_16758,N_12718,N_13629);
nand U16759 (N_16759,N_12084,N_14103);
xnor U16760 (N_16760,N_13469,N_14005);
nand U16761 (N_16761,N_13805,N_12376);
nand U16762 (N_16762,N_13730,N_11571);
xor U16763 (N_16763,N_11767,N_13446);
or U16764 (N_16764,N_13569,N_11185);
or U16765 (N_16765,N_12329,N_14784);
xor U16766 (N_16766,N_10733,N_13854);
nand U16767 (N_16767,N_10858,N_14364);
or U16768 (N_16768,N_14156,N_14094);
xnor U16769 (N_16769,N_11310,N_10775);
nor U16770 (N_16770,N_12127,N_14045);
or U16771 (N_16771,N_12611,N_14377);
nand U16772 (N_16772,N_10296,N_11443);
nor U16773 (N_16773,N_11595,N_11117);
or U16774 (N_16774,N_10879,N_10027);
and U16775 (N_16775,N_10664,N_10173);
nand U16776 (N_16776,N_10351,N_13010);
and U16777 (N_16777,N_11338,N_14426);
nand U16778 (N_16778,N_12695,N_13069);
or U16779 (N_16779,N_11634,N_12086);
nor U16780 (N_16780,N_14698,N_14539);
or U16781 (N_16781,N_14504,N_14761);
or U16782 (N_16782,N_14851,N_12651);
and U16783 (N_16783,N_10947,N_10864);
nor U16784 (N_16784,N_14721,N_13520);
nand U16785 (N_16785,N_14255,N_13968);
xnor U16786 (N_16786,N_11688,N_12916);
or U16787 (N_16787,N_10156,N_11037);
or U16788 (N_16788,N_10209,N_14212);
nand U16789 (N_16789,N_10985,N_13264);
nor U16790 (N_16790,N_13031,N_14050);
and U16791 (N_16791,N_12649,N_12972);
nand U16792 (N_16792,N_14999,N_10138);
xnor U16793 (N_16793,N_13179,N_13630);
xor U16794 (N_16794,N_13866,N_14207);
nand U16795 (N_16795,N_13899,N_14742);
nand U16796 (N_16796,N_10516,N_11034);
or U16797 (N_16797,N_10726,N_11043);
and U16798 (N_16798,N_10630,N_13843);
and U16799 (N_16799,N_14489,N_10860);
nand U16800 (N_16800,N_14744,N_13170);
or U16801 (N_16801,N_14772,N_14294);
nand U16802 (N_16802,N_12979,N_13731);
nor U16803 (N_16803,N_14714,N_10095);
xor U16804 (N_16804,N_11878,N_14293);
and U16805 (N_16805,N_13771,N_12242);
xnor U16806 (N_16806,N_14317,N_10073);
or U16807 (N_16807,N_13084,N_12863);
nor U16808 (N_16808,N_13066,N_13072);
nor U16809 (N_16809,N_14598,N_12897);
nand U16810 (N_16810,N_10002,N_12561);
and U16811 (N_16811,N_11727,N_14988);
nand U16812 (N_16812,N_10545,N_11794);
or U16813 (N_16813,N_12048,N_10546);
nand U16814 (N_16814,N_10362,N_13297);
nor U16815 (N_16815,N_13712,N_14178);
nand U16816 (N_16816,N_10529,N_11896);
and U16817 (N_16817,N_12520,N_14318);
xnor U16818 (N_16818,N_11585,N_13077);
xnor U16819 (N_16819,N_11531,N_14701);
and U16820 (N_16820,N_12882,N_11724);
and U16821 (N_16821,N_12365,N_11638);
nor U16822 (N_16822,N_14860,N_11583);
xor U16823 (N_16823,N_14099,N_11150);
nor U16824 (N_16824,N_14048,N_12449);
and U16825 (N_16825,N_10350,N_12689);
nand U16826 (N_16826,N_12385,N_14682);
xnor U16827 (N_16827,N_13319,N_12978);
xor U16828 (N_16828,N_10383,N_14845);
nor U16829 (N_16829,N_11138,N_12193);
xnor U16830 (N_16830,N_11682,N_11508);
nand U16831 (N_16831,N_13822,N_14723);
nor U16832 (N_16832,N_13153,N_13504);
nand U16833 (N_16833,N_10880,N_10128);
and U16834 (N_16834,N_11870,N_13209);
nand U16835 (N_16835,N_14569,N_13717);
nor U16836 (N_16836,N_10172,N_14478);
and U16837 (N_16837,N_13977,N_10340);
xor U16838 (N_16838,N_14993,N_13516);
nand U16839 (N_16839,N_11049,N_10440);
or U16840 (N_16840,N_12002,N_12282);
nand U16841 (N_16841,N_10600,N_10496);
and U16842 (N_16842,N_13677,N_12150);
and U16843 (N_16843,N_14709,N_14510);
nand U16844 (N_16844,N_13050,N_12563);
and U16845 (N_16845,N_11692,N_13955);
nand U16846 (N_16846,N_12446,N_13374);
nand U16847 (N_16847,N_12668,N_14322);
or U16848 (N_16848,N_13160,N_12073);
nand U16849 (N_16849,N_10412,N_14378);
xor U16850 (N_16850,N_12700,N_10211);
and U16851 (N_16851,N_11405,N_10055);
and U16852 (N_16852,N_10175,N_12612);
and U16853 (N_16853,N_12234,N_10431);
nor U16854 (N_16854,N_14513,N_10238);
or U16855 (N_16855,N_11581,N_10220);
and U16856 (N_16856,N_10874,N_12128);
or U16857 (N_16857,N_12186,N_12021);
nand U16858 (N_16858,N_10782,N_12153);
nand U16859 (N_16859,N_14641,N_11292);
xor U16860 (N_16860,N_11613,N_11351);
and U16861 (N_16861,N_11732,N_14873);
nor U16862 (N_16862,N_14316,N_13092);
nor U16863 (N_16863,N_11144,N_11889);
xor U16864 (N_16864,N_13492,N_13812);
nor U16865 (N_16865,N_14373,N_10502);
nand U16866 (N_16866,N_13082,N_14140);
nand U16867 (N_16867,N_10869,N_13468);
and U16868 (N_16868,N_10225,N_12035);
nand U16869 (N_16869,N_10581,N_13144);
and U16870 (N_16870,N_11624,N_10236);
nor U16871 (N_16871,N_14924,N_13424);
or U16872 (N_16872,N_12135,N_11382);
nor U16873 (N_16873,N_13406,N_14392);
xnor U16874 (N_16874,N_13613,N_10712);
or U16875 (N_16875,N_14722,N_11014);
nor U16876 (N_16876,N_11391,N_11448);
and U16877 (N_16877,N_13410,N_10578);
xnor U16878 (N_16878,N_10882,N_10426);
nor U16879 (N_16879,N_10531,N_14695);
nand U16880 (N_16880,N_14078,N_10946);
or U16881 (N_16881,N_12778,N_10958);
and U16882 (N_16882,N_13095,N_10018);
nand U16883 (N_16883,N_14508,N_13324);
or U16884 (N_16884,N_12823,N_13593);
nand U16885 (N_16885,N_13201,N_13886);
nor U16886 (N_16886,N_14274,N_10622);
nand U16887 (N_16887,N_13976,N_10976);
or U16888 (N_16888,N_14283,N_13833);
and U16889 (N_16889,N_12258,N_14732);
and U16890 (N_16890,N_14422,N_14549);
nor U16891 (N_16891,N_14705,N_11922);
and U16892 (N_16892,N_11153,N_13294);
xor U16893 (N_16893,N_12888,N_11856);
nand U16894 (N_16894,N_11203,N_14348);
nor U16895 (N_16895,N_13566,N_14174);
nand U16896 (N_16896,N_14372,N_10451);
or U16897 (N_16897,N_12008,N_10295);
nor U16898 (N_16898,N_13039,N_10394);
nand U16899 (N_16899,N_10861,N_13296);
xnor U16900 (N_16900,N_13965,N_10893);
nand U16901 (N_16901,N_13466,N_13139);
xnor U16902 (N_16902,N_14473,N_11271);
nand U16903 (N_16903,N_10901,N_11680);
and U16904 (N_16904,N_13038,N_11586);
or U16905 (N_16905,N_13444,N_10022);
and U16906 (N_16906,N_11833,N_10984);
or U16907 (N_16907,N_10702,N_13508);
nor U16908 (N_16908,N_10981,N_14623);
nand U16909 (N_16909,N_13195,N_10589);
nand U16910 (N_16910,N_10913,N_12655);
and U16911 (N_16911,N_10291,N_13913);
xnor U16912 (N_16912,N_12163,N_14896);
xnor U16913 (N_16913,N_13742,N_12312);
nor U16914 (N_16914,N_13067,N_12678);
and U16915 (N_16915,N_10429,N_11990);
nor U16916 (N_16916,N_12860,N_12842);
xnor U16917 (N_16917,N_11893,N_10191);
or U16918 (N_16918,N_10832,N_13343);
nor U16919 (N_16919,N_10166,N_12764);
nor U16920 (N_16920,N_12351,N_12466);
or U16921 (N_16921,N_12680,N_10396);
nand U16922 (N_16922,N_11551,N_11001);
and U16923 (N_16923,N_13585,N_13071);
xnor U16924 (N_16924,N_10347,N_13764);
xnor U16925 (N_16925,N_14658,N_13816);
or U16926 (N_16926,N_10070,N_14455);
xnor U16927 (N_16927,N_13434,N_14600);
or U16928 (N_16928,N_11623,N_12967);
xor U16929 (N_16929,N_11170,N_13785);
nor U16930 (N_16930,N_10476,N_11417);
or U16931 (N_16931,N_12502,N_13428);
or U16932 (N_16932,N_12579,N_13881);
nand U16933 (N_16933,N_11120,N_11086);
nor U16934 (N_16934,N_10324,N_11776);
or U16935 (N_16935,N_10251,N_10164);
nor U16936 (N_16936,N_13584,N_11579);
xnor U16937 (N_16937,N_14169,N_11494);
and U16938 (N_16938,N_12998,N_14633);
nor U16939 (N_16939,N_11715,N_12990);
xor U16940 (N_16940,N_13835,N_12199);
nor U16941 (N_16941,N_11312,N_14471);
nor U16942 (N_16942,N_10749,N_13933);
nand U16943 (N_16943,N_12610,N_10036);
or U16944 (N_16944,N_14375,N_12303);
xor U16945 (N_16945,N_10654,N_14162);
or U16946 (N_16946,N_11275,N_10547);
nor U16947 (N_16947,N_14526,N_10217);
or U16948 (N_16948,N_10338,N_12454);
nand U16949 (N_16949,N_13442,N_11348);
and U16950 (N_16950,N_10514,N_10483);
and U16951 (N_16951,N_11765,N_11921);
nor U16952 (N_16952,N_14110,N_11392);
or U16953 (N_16953,N_13605,N_12498);
or U16954 (N_16954,N_14729,N_12056);
nor U16955 (N_16955,N_11214,N_13543);
nor U16956 (N_16956,N_10088,N_13721);
nand U16957 (N_16957,N_11507,N_11820);
nor U16958 (N_16958,N_12496,N_10178);
nor U16959 (N_16959,N_14201,N_11516);
xor U16960 (N_16960,N_10793,N_12095);
and U16961 (N_16961,N_12676,N_13824);
nand U16962 (N_16962,N_13284,N_11189);
nor U16963 (N_16963,N_10077,N_14192);
xor U16964 (N_16964,N_11084,N_11152);
or U16965 (N_16965,N_13969,N_10212);
and U16966 (N_16966,N_14735,N_10498);
or U16967 (N_16967,N_11790,N_11121);
or U16968 (N_16968,N_11839,N_10231);
xnor U16969 (N_16969,N_11826,N_10593);
or U16970 (N_16970,N_13426,N_14923);
nor U16971 (N_16971,N_13719,N_12925);
and U16972 (N_16972,N_14561,N_14419);
nand U16973 (N_16973,N_13118,N_13060);
and U16974 (N_16974,N_13754,N_11245);
xor U16975 (N_16975,N_13147,N_14727);
nand U16976 (N_16976,N_12467,N_14970);
and U16977 (N_16977,N_12216,N_11394);
nand U16978 (N_16978,N_11815,N_12797);
nor U16979 (N_16979,N_10032,N_11251);
or U16980 (N_16980,N_13128,N_10881);
nor U16981 (N_16981,N_12783,N_14286);
or U16982 (N_16982,N_11287,N_10834);
nor U16983 (N_16983,N_11594,N_13841);
xnor U16984 (N_16984,N_12406,N_13947);
nand U16985 (N_16985,N_11713,N_13341);
or U16986 (N_16986,N_12708,N_12530);
nor U16987 (N_16987,N_12274,N_13054);
nor U16988 (N_16988,N_10234,N_11534);
nand U16989 (N_16989,N_13896,N_10620);
nand U16990 (N_16990,N_12762,N_14297);
nor U16991 (N_16991,N_11552,N_10604);
nand U16992 (N_16992,N_14800,N_12807);
nor U16993 (N_16993,N_13612,N_11083);
and U16994 (N_16994,N_13745,N_13495);
nor U16995 (N_16995,N_14193,N_13723);
and U16996 (N_16996,N_14947,N_14341);
xor U16997 (N_16997,N_11402,N_11015);
nand U16998 (N_16998,N_13631,N_13844);
xnor U16999 (N_16999,N_11099,N_13522);
nor U17000 (N_17000,N_11007,N_14885);
or U17001 (N_17001,N_11178,N_13051);
or U17002 (N_17002,N_14214,N_13042);
nand U17003 (N_17003,N_14187,N_12752);
xnor U17004 (N_17004,N_10300,N_11076);
or U17005 (N_17005,N_12832,N_10361);
and U17006 (N_17006,N_11415,N_14768);
xnor U17007 (N_17007,N_13815,N_12769);
xnor U17008 (N_17008,N_14725,N_13505);
and U17009 (N_17009,N_10326,N_14699);
nand U17010 (N_17010,N_13658,N_13880);
or U17011 (N_17011,N_10950,N_13484);
and U17012 (N_17012,N_14595,N_14158);
nor U17013 (N_17013,N_10334,N_11728);
xnor U17014 (N_17014,N_11966,N_11837);
nor U17015 (N_17015,N_11509,N_14869);
nor U17016 (N_17016,N_14799,N_13361);
nor U17017 (N_17017,N_11560,N_11734);
and U17018 (N_17018,N_13193,N_10577);
nor U17019 (N_17019,N_13556,N_10651);
or U17020 (N_17020,N_11860,N_11672);
nor U17021 (N_17021,N_13137,N_10454);
xor U17022 (N_17022,N_10907,N_13980);
or U17023 (N_17023,N_12356,N_10267);
or U17024 (N_17024,N_13796,N_11167);
nor U17025 (N_17025,N_11647,N_14743);
nand U17026 (N_17026,N_12846,N_12092);
nand U17027 (N_17027,N_13510,N_11526);
or U17028 (N_17028,N_10906,N_10475);
or U17029 (N_17029,N_13215,N_11025);
xnor U17030 (N_17030,N_11277,N_11629);
and U17031 (N_17031,N_14389,N_13248);
nand U17032 (N_17032,N_11163,N_11858);
xor U17033 (N_17033,N_10048,N_12806);
xor U17034 (N_17034,N_12845,N_10355);
nor U17035 (N_17035,N_11145,N_14878);
and U17036 (N_17036,N_10811,N_12078);
nand U17037 (N_17037,N_13776,N_13872);
xnor U17038 (N_17038,N_10152,N_12210);
or U17039 (N_17039,N_13315,N_14073);
nor U17040 (N_17040,N_13836,N_10570);
xor U17041 (N_17041,N_13271,N_14538);
nand U17042 (N_17042,N_10971,N_11318);
nand U17043 (N_17043,N_14948,N_12685);
or U17044 (N_17044,N_11559,N_11263);
nor U17045 (N_17045,N_11917,N_11619);
and U17046 (N_17046,N_12066,N_12733);
xnor U17047 (N_17047,N_13578,N_14394);
and U17048 (N_17048,N_12951,N_11997);
xor U17049 (N_17049,N_10751,N_13792);
or U17050 (N_17050,N_13897,N_12297);
nor U17051 (N_17051,N_14380,N_13165);
or U17052 (N_17052,N_12851,N_14260);
and U17053 (N_17053,N_12310,N_11296);
nor U17054 (N_17054,N_10618,N_14233);
or U17055 (N_17055,N_14511,N_14277);
or U17056 (N_17056,N_14335,N_11674);
nand U17057 (N_17057,N_12808,N_13415);
nand U17058 (N_17058,N_13936,N_11273);
or U17059 (N_17059,N_11575,N_14872);
or U17060 (N_17060,N_14712,N_12389);
nand U17061 (N_17061,N_12233,N_10970);
xnor U17062 (N_17062,N_14880,N_11269);
or U17063 (N_17063,N_14194,N_11479);
or U17064 (N_17064,N_13941,N_11111);
or U17065 (N_17065,N_11316,N_13868);
and U17066 (N_17066,N_11401,N_14353);
and U17067 (N_17067,N_10781,N_13146);
or U17068 (N_17068,N_10258,N_12055);
and U17069 (N_17069,N_12589,N_13239);
xor U17070 (N_17070,N_12450,N_10008);
nand U17071 (N_17071,N_13521,N_10928);
xor U17072 (N_17072,N_13648,N_12115);
nor U17073 (N_17073,N_10555,N_11176);
and U17074 (N_17074,N_13709,N_12675);
and U17075 (N_17075,N_10942,N_12288);
nand U17076 (N_17076,N_14786,N_10663);
xnor U17077 (N_17077,N_12883,N_13915);
nand U17078 (N_17078,N_13670,N_12505);
and U17079 (N_17079,N_13181,N_12694);
nand U17080 (N_17080,N_14980,N_14145);
xnor U17081 (N_17081,N_14854,N_14371);
nand U17082 (N_17082,N_12551,N_13659);
xnor U17083 (N_17083,N_12855,N_11961);
and U17084 (N_17084,N_11332,N_14669);
nand U17085 (N_17085,N_13883,N_14660);
or U17086 (N_17086,N_13610,N_12912);
and U17087 (N_17087,N_11563,N_10715);
or U17088 (N_17088,N_12988,N_11887);
or U17089 (N_17089,N_10270,N_10051);
nor U17090 (N_17090,N_13435,N_10279);
nand U17091 (N_17091,N_12182,N_11910);
nand U17092 (N_17092,N_11344,N_11562);
and U17093 (N_17093,N_11670,N_10115);
xnor U17094 (N_17094,N_12436,N_12574);
or U17095 (N_17095,N_11398,N_10259);
nand U17096 (N_17096,N_14068,N_10510);
xnor U17097 (N_17097,N_13053,N_10493);
xnor U17098 (N_17098,N_10619,N_13389);
and U17099 (N_17099,N_10741,N_11130);
nor U17100 (N_17100,N_10890,N_10460);
or U17101 (N_17101,N_14147,N_10325);
nor U17102 (N_17102,N_11895,N_13022);
and U17103 (N_17103,N_11373,N_14313);
xor U17104 (N_17104,N_12161,N_12603);
nor U17105 (N_17105,N_13597,N_13837);
and U17106 (N_17106,N_12588,N_12792);
xor U17107 (N_17107,N_13119,N_10597);
or U17108 (N_17108,N_10800,N_10538);
or U17109 (N_17109,N_12480,N_10453);
xor U17110 (N_17110,N_11857,N_12088);
nand U17111 (N_17111,N_10423,N_13825);
and U17112 (N_17112,N_10634,N_10438);
nor U17113 (N_17113,N_14636,N_10842);
nor U17114 (N_17114,N_11000,N_10464);
nor U17115 (N_17115,N_14689,N_13780);
or U17116 (N_17116,N_13869,N_13330);
xnor U17117 (N_17117,N_10490,N_11518);
nor U17118 (N_17118,N_14967,N_10999);
xnor U17119 (N_17119,N_10011,N_13043);
nand U17120 (N_17120,N_11210,N_11939);
nor U17121 (N_17121,N_12690,N_14016);
xor U17122 (N_17122,N_10960,N_11950);
or U17123 (N_17123,N_12370,N_11293);
or U17124 (N_17124,N_14683,N_11513);
and U17125 (N_17125,N_13411,N_13265);
or U17126 (N_17126,N_10576,N_14534);
nor U17127 (N_17127,N_14365,N_12814);
nand U17128 (N_17128,N_12411,N_13331);
xnor U17129 (N_17129,N_12527,N_12222);
or U17130 (N_17130,N_12940,N_14864);
nand U17131 (N_17131,N_13115,N_12803);
nand U17132 (N_17132,N_12567,N_10532);
xnor U17133 (N_17133,N_11886,N_12550);
xnor U17134 (N_17134,N_13532,N_13606);
or U17135 (N_17135,N_11809,N_10723);
nand U17136 (N_17136,N_10316,N_13935);
or U17137 (N_17137,N_12512,N_12497);
nor U17138 (N_17138,N_10061,N_12536);
or U17139 (N_17139,N_11830,N_11220);
nand U17140 (N_17140,N_13169,N_12264);
and U17141 (N_17141,N_10050,N_13944);
or U17142 (N_17142,N_14084,N_14223);
nor U17143 (N_17143,N_13587,N_11416);
nand U17144 (N_17144,N_12734,N_10344);
xnor U17145 (N_17145,N_13827,N_13829);
and U17146 (N_17146,N_13507,N_13727);
or U17147 (N_17147,N_14770,N_11468);
nor U17148 (N_17148,N_13902,N_14337);
nand U17149 (N_17149,N_13496,N_13109);
or U17150 (N_17150,N_10536,N_11229);
nor U17151 (N_17151,N_14963,N_14918);
xnor U17152 (N_17152,N_11087,N_12724);
nand U17153 (N_17153,N_14586,N_12471);
nand U17154 (N_17154,N_13333,N_13894);
nor U17155 (N_17155,N_13946,N_11681);
nand U17156 (N_17156,N_14671,N_14618);
nor U17157 (N_17157,N_12090,N_11912);
or U17158 (N_17158,N_13738,N_10143);
xnor U17159 (N_17159,N_12138,N_13081);
nor U17160 (N_17160,N_12244,N_13634);
and U17161 (N_17161,N_10904,N_11538);
nor U17162 (N_17162,N_12656,N_11249);
xor U17163 (N_17163,N_13478,N_14271);
or U17164 (N_17164,N_14643,N_12259);
xor U17165 (N_17165,N_13272,N_14847);
xor U17166 (N_17166,N_13448,N_11164);
or U17167 (N_17167,N_12114,N_13306);
nor U17168 (N_17168,N_11222,N_13267);
xor U17169 (N_17169,N_10305,N_11561);
nand U17170 (N_17170,N_10282,N_13813);
nand U17171 (N_17171,N_14467,N_14439);
nand U17172 (N_17172,N_13598,N_13555);
nor U17173 (N_17173,N_12627,N_11578);
and U17174 (N_17174,N_11125,N_13951);
nand U17175 (N_17175,N_14447,N_12905);
or U17176 (N_17176,N_13666,N_11459);
xor U17177 (N_17177,N_13596,N_14844);
nand U17178 (N_17178,N_10122,N_14149);
or U17179 (N_17179,N_10643,N_13086);
xor U17180 (N_17180,N_12333,N_10956);
nand U17181 (N_17181,N_13441,N_11489);
xor U17182 (N_17182,N_13818,N_13070);
or U17183 (N_17183,N_11819,N_14202);
xnor U17184 (N_17184,N_12097,N_10797);
and U17185 (N_17185,N_11055,N_12126);
xnor U17186 (N_17186,N_14211,N_10116);
xnor U17187 (N_17187,N_11285,N_14889);
xnor U17188 (N_17188,N_12324,N_10968);
and U17189 (N_17189,N_11707,N_11353);
nor U17190 (N_17190,N_12529,N_11442);
xnor U17191 (N_17191,N_12793,N_11781);
xnor U17192 (N_17192,N_11975,N_10964);
nand U17193 (N_17193,N_12903,N_13940);
nand U17194 (N_17194,N_10151,N_13436);
nor U17195 (N_17195,N_12915,N_14853);
and U17196 (N_17196,N_11861,N_12961);
and U17197 (N_17197,N_12874,N_11635);
nor U17198 (N_17198,N_13572,N_10873);
and U17199 (N_17199,N_11704,N_12838);
xor U17200 (N_17200,N_11648,N_10524);
or U17201 (N_17201,N_12169,N_13783);
and U17202 (N_17202,N_11590,N_12522);
or U17203 (N_17203,N_12552,N_13548);
nand U17204 (N_17204,N_10924,N_12873);
nand U17205 (N_17205,N_11769,N_10759);
or U17206 (N_17206,N_14794,N_14917);
or U17207 (N_17207,N_14257,N_14693);
nand U17208 (N_17208,N_14648,N_12141);
nand U17209 (N_17209,N_12628,N_14234);
or U17210 (N_17210,N_11843,N_13124);
or U17211 (N_17211,N_11646,N_11663);
or U17212 (N_17212,N_14930,N_13545);
and U17213 (N_17213,N_12155,N_10583);
xnor U17214 (N_17214,N_10714,N_14486);
or U17215 (N_17215,N_10557,N_11337);
nor U17216 (N_17216,N_12993,N_14733);
or U17217 (N_17217,N_11235,N_10393);
xor U17218 (N_17218,N_13888,N_13753);
nor U17219 (N_17219,N_13749,N_12291);
and U17220 (N_17220,N_10224,N_11503);
nand U17221 (N_17221,N_11460,N_12722);
nor U17222 (N_17222,N_13254,N_11871);
nand U17223 (N_17223,N_11863,N_13908);
nor U17224 (N_17224,N_11127,N_10057);
nand U17225 (N_17225,N_11607,N_13609);
nor U17226 (N_17226,N_14057,N_13421);
and U17227 (N_17227,N_14251,N_11965);
and U17228 (N_17228,N_13219,N_14655);
xnor U17229 (N_17229,N_10074,N_11684);
and U17230 (N_17230,N_11126,N_14190);
or U17231 (N_17231,N_11478,N_13799);
xnor U17232 (N_17232,N_13773,N_14191);
and U17233 (N_17233,N_12195,N_12422);
nand U17234 (N_17234,N_12394,N_11490);
and U17235 (N_17235,N_13650,N_13692);
xor U17236 (N_17236,N_13074,N_10841);
or U17237 (N_17237,N_12087,N_13395);
nand U17238 (N_17238,N_12111,N_13047);
and U17239 (N_17239,N_14232,N_10222);
nand U17240 (N_17240,N_14170,N_13684);
and U17241 (N_17241,N_14412,N_10488);
and U17242 (N_17242,N_10263,N_10052);
nand U17243 (N_17243,N_13506,N_14613);
nor U17244 (N_17244,N_10507,N_12340);
or U17245 (N_17245,N_11656,N_14562);
nand U17246 (N_17246,N_14114,N_14989);
xor U17247 (N_17247,N_11016,N_12861);
nand U17248 (N_17248,N_12710,N_11652);
and U17249 (N_17249,N_13638,N_12129);
or U17250 (N_17250,N_10738,N_12609);
or U17251 (N_17251,N_10883,N_13621);
or U17252 (N_17252,N_11082,N_13270);
and U17253 (N_17253,N_13360,N_12631);
and U17254 (N_17254,N_11808,N_12902);
nor U17255 (N_17255,N_14927,N_10925);
and U17256 (N_17256,N_11510,N_14387);
nor U17257 (N_17257,N_13794,N_14717);
nor U17258 (N_17258,N_12545,N_13120);
nor U17259 (N_17259,N_11451,N_14497);
nor U17260 (N_17260,N_11089,N_11710);
nand U17261 (N_17261,N_12608,N_13059);
nor U17262 (N_17262,N_10734,N_10673);
and U17263 (N_17263,N_11396,N_13871);
or U17264 (N_17264,N_11998,N_10028);
xnor U17265 (N_17265,N_11060,N_11810);
or U17266 (N_17266,N_13948,N_12759);
nor U17267 (N_17267,N_12181,N_12698);
nand U17268 (N_17268,N_10031,N_12183);
and U17269 (N_17269,N_13739,N_13643);
or U17270 (N_17270,N_13852,N_13901);
nor U17271 (N_17271,N_14129,N_11288);
and U17272 (N_17272,N_14333,N_14340);
nor U17273 (N_17273,N_10711,N_10905);
or U17274 (N_17274,N_13024,N_12945);
nand U17275 (N_17275,N_11454,N_13752);
or U17276 (N_17276,N_10810,N_14954);
or U17277 (N_17277,N_10784,N_11365);
nor U17278 (N_17278,N_14900,N_10080);
and U17279 (N_17279,N_12189,N_11143);
nand U17280 (N_17280,N_10275,N_10356);
and U17281 (N_17281,N_14767,N_13989);
nand U17282 (N_17282,N_14519,N_12958);
or U17283 (N_17283,N_14358,N_14060);
and U17284 (N_17284,N_12843,N_11458);
nand U17285 (N_17285,N_11795,N_11564);
nand U17286 (N_17286,N_11799,N_12768);
nand U17287 (N_17287,N_11186,N_13877);
and U17288 (N_17288,N_11698,N_14407);
and U17289 (N_17289,N_12534,N_13909);
xnor U17290 (N_17290,N_10571,N_13236);
nor U17291 (N_17291,N_13336,N_10769);
and U17292 (N_17292,N_14111,N_10407);
nand U17293 (N_17293,N_12854,N_13299);
and U17294 (N_17294,N_13180,N_13784);
xnor U17295 (N_17295,N_14891,N_12247);
xor U17296 (N_17296,N_11838,N_11731);
and U17297 (N_17297,N_13322,N_13238);
and U17298 (N_17298,N_10903,N_11227);
or U17299 (N_17299,N_11785,N_14448);
xor U17300 (N_17300,N_10799,N_14716);
or U17301 (N_17301,N_14642,N_13800);
nor U17302 (N_17302,N_14217,N_10794);
and U17303 (N_17303,N_11994,N_12745);
and U17304 (N_17304,N_12515,N_11104);
nor U17305 (N_17305,N_13707,N_11331);
nand U17306 (N_17306,N_11948,N_11324);
and U17307 (N_17307,N_10900,N_12501);
nor U17308 (N_17308,N_10366,N_14985);
and U17309 (N_17309,N_14328,N_12521);
nand U17310 (N_17310,N_14796,N_10335);
nor U17311 (N_17311,N_11903,N_12033);
xnor U17312 (N_17312,N_11547,N_13565);
nand U17313 (N_17313,N_13019,N_11511);
nor U17314 (N_17314,N_11092,N_12867);
or U17315 (N_17315,N_11098,N_14476);
or U17316 (N_17316,N_11311,N_12172);
or U17317 (N_17317,N_11774,N_13810);
xnor U17318 (N_17318,N_10506,N_12064);
nand U17319 (N_17319,N_13020,N_14279);
xor U17320 (N_17320,N_11197,N_12240);
nand U17321 (N_17321,N_10233,N_10395);
and U17322 (N_17322,N_10786,N_12162);
and U17323 (N_17323,N_12788,N_11841);
or U17324 (N_17324,N_13027,N_11546);
nand U17325 (N_17325,N_11737,N_12503);
nand U17326 (N_17326,N_14871,N_14173);
xnor U17327 (N_17327,N_13307,N_12336);
xnor U17328 (N_17328,N_10289,N_10120);
nor U17329 (N_17329,N_14463,N_10836);
or U17330 (N_17330,N_14433,N_12043);
xnor U17331 (N_17331,N_11340,N_10411);
or U17332 (N_17332,N_12495,N_13911);
and U17333 (N_17333,N_14250,N_10271);
nor U17334 (N_17334,N_14472,N_11717);
nor U17335 (N_17335,N_11747,N_14625);
nand U17336 (N_17336,N_14056,N_13769);
nand U17337 (N_17337,N_12533,N_13064);
and U17338 (N_17338,N_14577,N_13379);
nor U17339 (N_17339,N_13893,N_11660);
and U17340 (N_17340,N_14172,N_11056);
nand U17341 (N_17341,N_13798,N_10941);
and U17342 (N_17342,N_12927,N_10094);
or U17343 (N_17343,N_12119,N_14326);
and U17344 (N_17344,N_13034,N_12962);
nand U17345 (N_17345,N_10406,N_10568);
nor U17346 (N_17346,N_13538,N_10805);
nor U17347 (N_17347,N_14792,N_13363);
or U17348 (N_17348,N_12206,N_13823);
nand U17349 (N_17349,N_10352,N_10791);
and U17350 (N_17350,N_12334,N_12211);
nand U17351 (N_17351,N_14776,N_12595);
nor U17352 (N_17352,N_12197,N_12091);
or U17353 (N_17353,N_11610,N_12372);
nor U17354 (N_17354,N_13574,N_10005);
and U17355 (N_17355,N_14700,N_12157);
nand U17356 (N_17356,N_10482,N_13300);
and U17357 (N_17357,N_11488,N_11080);
and U17358 (N_17358,N_14167,N_13274);
nor U17359 (N_17359,N_12131,N_12215);
or U17360 (N_17360,N_13025,N_11248);
or U17361 (N_17361,N_10997,N_10196);
and U17362 (N_17362,N_13246,N_14839);
xor U17363 (N_17363,N_12770,N_12185);
or U17364 (N_17364,N_14343,N_11242);
and U17365 (N_17365,N_14524,N_14789);
nor U17366 (N_17366,N_14920,N_11424);
nand U17367 (N_17367,N_11307,N_11683);
nand U17368 (N_17368,N_10239,N_13462);
nor U17369 (N_17369,N_14082,N_11941);
or U17370 (N_17370,N_10961,N_14226);
nand U17371 (N_17371,N_12015,N_14249);
or U17372 (N_17372,N_14001,N_14545);
and U17373 (N_17373,N_12641,N_13526);
xor U17374 (N_17374,N_11974,N_10378);
nand U17375 (N_17375,N_10730,N_12547);
xor U17376 (N_17376,N_10803,N_10227);
xnor U17377 (N_17377,N_13476,N_13744);
or U17378 (N_17378,N_11350,N_13396);
nand U17379 (N_17379,N_14780,N_11572);
xor U17380 (N_17380,N_13061,N_10647);
nand U17381 (N_17381,N_11780,N_14163);
or U17382 (N_17382,N_12443,N_13633);
or U17383 (N_17383,N_14354,N_13642);
nand U17384 (N_17384,N_14215,N_10629);
xnor U17385 (N_17385,N_14678,N_12388);
nor U17386 (N_17386,N_13640,N_11695);
nor U17387 (N_17387,N_11678,N_10939);
xor U17388 (N_17388,N_10494,N_12632);
nand U17389 (N_17389,N_10814,N_10358);
nand U17390 (N_17390,N_12750,N_13831);
or U17391 (N_17391,N_12300,N_10499);
and U17392 (N_17392,N_13113,N_11256);
and U17393 (N_17393,N_14758,N_10299);
and U17394 (N_17394,N_14859,N_11261);
xor U17395 (N_17395,N_14230,N_11596);
and U17396 (N_17396,N_10974,N_11805);
xor U17397 (N_17397,N_14741,N_12730);
or U17398 (N_17398,N_11029,N_10528);
nand U17399 (N_17399,N_14783,N_11005);
xor U17400 (N_17400,N_12504,N_13151);
nand U17401 (N_17401,N_14943,N_11212);
and U17402 (N_17402,N_14122,N_10768);
nand U17403 (N_17403,N_11236,N_10635);
nor U17404 (N_17404,N_14978,N_13223);
nand U17405 (N_17405,N_13402,N_10875);
nor U17406 (N_17406,N_14003,N_13536);
or U17407 (N_17407,N_11943,N_14063);
nor U17408 (N_17408,N_12026,N_10330);
xnor U17409 (N_17409,N_12616,N_14263);
or U17410 (N_17410,N_14138,N_13347);
or U17411 (N_17411,N_12546,N_14514);
or U17412 (N_17412,N_13287,N_11908);
nand U17413 (N_17413,N_10311,N_11134);
nand U17414 (N_17414,N_14034,N_14824);
and U17415 (N_17415,N_10933,N_13667);
xor U17416 (N_17416,N_14021,N_13559);
or U17417 (N_17417,N_11465,N_10284);
nor U17418 (N_17418,N_14276,N_11631);
xor U17419 (N_17419,N_14719,N_10748);
xnor U17420 (N_17420,N_13477,N_14934);
nand U17421 (N_17421,N_12437,N_10180);
nand U17422 (N_17422,N_13275,N_10530);
nor U17423 (N_17423,N_10147,N_12535);
nand U17424 (N_17424,N_13550,N_11357);
or U17425 (N_17425,N_10364,N_10219);
or U17426 (N_17426,N_13646,N_11693);
and U17427 (N_17427,N_11013,N_14996);
nand U17428 (N_17428,N_10822,N_11484);
xnor U17429 (N_17429,N_11336,N_13327);
nand U17430 (N_17430,N_11797,N_12755);
xor U17431 (N_17431,N_14054,N_11745);
nor U17432 (N_17432,N_14490,N_11933);
xor U17433 (N_17433,N_14568,N_11983);
or U17434 (N_17434,N_11154,N_10518);
and U17435 (N_17435,N_11384,N_14206);
and U17436 (N_17436,N_12478,N_10843);
nor U17437 (N_17437,N_13244,N_12713);
nand U17438 (N_17438,N_13171,N_10750);
nand U17439 (N_17439,N_14105,N_14144);
or U17440 (N_17440,N_14529,N_12335);
and U17441 (N_17441,N_10086,N_11467);
or U17442 (N_17442,N_10995,N_12429);
nand U17443 (N_17443,N_12057,N_12960);
and U17444 (N_17444,N_14560,N_12262);
nand U17445 (N_17445,N_13847,N_14610);
nand U17446 (N_17446,N_10944,N_11557);
nor U17447 (N_17447,N_12599,N_11689);
xnor U17448 (N_17448,N_12736,N_11345);
xor U17449 (N_17449,N_12889,N_12844);
nor U17450 (N_17450,N_11855,N_13186);
and U17451 (N_17451,N_14797,N_13364);
xor U17452 (N_17452,N_10888,N_13934);
xnor U17453 (N_17453,N_13635,N_11616);
or U17454 (N_17454,N_11260,N_13892);
nor U17455 (N_17455,N_13583,N_12637);
nand U17456 (N_17456,N_11280,N_13392);
nor U17457 (N_17457,N_12014,N_13511);
nand U17458 (N_17458,N_10444,N_14737);
xor U17459 (N_17459,N_10010,N_12287);
nor U17460 (N_17460,N_13217,N_10203);
nor U17461 (N_17461,N_14505,N_12420);
nor U17462 (N_17462,N_11063,N_13895);
xor U17463 (N_17463,N_12191,N_11630);
nor U17464 (N_17464,N_14634,N_11147);
xor U17465 (N_17465,N_11476,N_11339);
nor U17466 (N_17466,N_12010,N_11609);
nor U17467 (N_17467,N_12691,N_12709);
nor U17468 (N_17468,N_12007,N_14621);
or U17469 (N_17469,N_12660,N_10923);
nand U17470 (N_17470,N_14363,N_14470);
nand U17471 (N_17471,N_12934,N_11057);
nand U17472 (N_17472,N_12352,N_11527);
xnor U17473 (N_17473,N_13622,N_14522);
nand U17474 (N_17474,N_10572,N_12901);
and U17475 (N_17475,N_10029,N_10082);
xor U17476 (N_17476,N_14926,N_12243);
and U17477 (N_17477,N_12364,N_11486);
and U17478 (N_17478,N_12926,N_12869);
or U17479 (N_17479,N_10512,N_10868);
or U17480 (N_17480,N_14134,N_10479);
or U17481 (N_17481,N_11131,N_10762);
nand U17482 (N_17482,N_11193,N_10717);
xnor U17483 (N_17483,N_12772,N_10449);
or U17484 (N_17484,N_10058,N_11915);
and U17485 (N_17485,N_13298,N_10592);
nand U17486 (N_17486,N_11783,N_10452);
nor U17487 (N_17487,N_11851,N_14617);
and U17488 (N_17488,N_11876,N_11845);
nand U17489 (N_17489,N_12896,N_12442);
and U17490 (N_17490,N_13993,N_12121);
or U17491 (N_17491,N_13826,N_12113);
nor U17492 (N_17492,N_14291,N_10287);
nor U17493 (N_17493,N_14047,N_14840);
nand U17494 (N_17494,N_11880,N_11407);
nor U17495 (N_17495,N_14067,N_10020);
nor U17496 (N_17496,N_12633,N_13858);
nor U17497 (N_17497,N_13432,N_11215);
or U17498 (N_17498,N_11400,N_10409);
nor U17499 (N_17499,N_10763,N_12899);
or U17500 (N_17500,N_10009,N_13487);
and U17501 (N_17501,N_14717,N_14970);
nand U17502 (N_17502,N_13665,N_13459);
nor U17503 (N_17503,N_11369,N_13387);
or U17504 (N_17504,N_13981,N_14961);
nand U17505 (N_17505,N_14343,N_12836);
or U17506 (N_17506,N_13107,N_14436);
nand U17507 (N_17507,N_13961,N_14189);
xor U17508 (N_17508,N_13987,N_14406);
or U17509 (N_17509,N_12712,N_12100);
or U17510 (N_17510,N_12610,N_13341);
nor U17511 (N_17511,N_10102,N_12560);
nor U17512 (N_17512,N_12738,N_14180);
nand U17513 (N_17513,N_10420,N_13469);
and U17514 (N_17514,N_10238,N_10511);
and U17515 (N_17515,N_11297,N_14765);
nor U17516 (N_17516,N_12627,N_10734);
nor U17517 (N_17517,N_12733,N_11052);
nor U17518 (N_17518,N_14053,N_14193);
and U17519 (N_17519,N_12079,N_11270);
and U17520 (N_17520,N_13504,N_14372);
xnor U17521 (N_17521,N_10461,N_10317);
or U17522 (N_17522,N_13701,N_13042);
nand U17523 (N_17523,N_14512,N_14616);
nor U17524 (N_17524,N_14874,N_14045);
nand U17525 (N_17525,N_13211,N_11046);
or U17526 (N_17526,N_10694,N_14127);
nor U17527 (N_17527,N_11085,N_14268);
nand U17528 (N_17528,N_11948,N_10289);
or U17529 (N_17529,N_13547,N_13531);
or U17530 (N_17530,N_13214,N_11404);
nand U17531 (N_17531,N_10470,N_13480);
or U17532 (N_17532,N_11114,N_10390);
or U17533 (N_17533,N_11791,N_14306);
and U17534 (N_17534,N_12963,N_14570);
nor U17535 (N_17535,N_12660,N_11335);
and U17536 (N_17536,N_10439,N_11383);
nor U17537 (N_17537,N_13291,N_13899);
nor U17538 (N_17538,N_14375,N_14169);
or U17539 (N_17539,N_13861,N_12018);
nor U17540 (N_17540,N_14131,N_14357);
or U17541 (N_17541,N_10734,N_10112);
nor U17542 (N_17542,N_12209,N_12824);
and U17543 (N_17543,N_10257,N_13050);
nor U17544 (N_17544,N_14480,N_12277);
xor U17545 (N_17545,N_13395,N_12783);
xnor U17546 (N_17546,N_12458,N_14729);
xor U17547 (N_17547,N_11215,N_14110);
nand U17548 (N_17548,N_12186,N_14363);
nor U17549 (N_17549,N_13269,N_13494);
or U17550 (N_17550,N_11604,N_11622);
and U17551 (N_17551,N_12879,N_14838);
nor U17552 (N_17552,N_14459,N_12210);
nor U17553 (N_17553,N_10917,N_14788);
nand U17554 (N_17554,N_11804,N_10613);
nor U17555 (N_17555,N_14884,N_14467);
xor U17556 (N_17556,N_11375,N_13069);
or U17557 (N_17557,N_14524,N_10487);
or U17558 (N_17558,N_13076,N_14963);
and U17559 (N_17559,N_14363,N_13027);
xor U17560 (N_17560,N_12431,N_12484);
and U17561 (N_17561,N_11311,N_12102);
xor U17562 (N_17562,N_11751,N_13973);
and U17563 (N_17563,N_10056,N_11614);
nor U17564 (N_17564,N_10265,N_14662);
and U17565 (N_17565,N_13354,N_11992);
or U17566 (N_17566,N_11609,N_13069);
and U17567 (N_17567,N_12079,N_12799);
nand U17568 (N_17568,N_12270,N_13992);
or U17569 (N_17569,N_14417,N_13476);
nor U17570 (N_17570,N_14130,N_14974);
xor U17571 (N_17571,N_14621,N_14071);
and U17572 (N_17572,N_14296,N_13251);
or U17573 (N_17573,N_10085,N_10897);
xnor U17574 (N_17574,N_13464,N_13088);
nand U17575 (N_17575,N_14708,N_13873);
xnor U17576 (N_17576,N_11807,N_10183);
and U17577 (N_17577,N_12369,N_12609);
nor U17578 (N_17578,N_11635,N_14796);
or U17579 (N_17579,N_11893,N_10162);
and U17580 (N_17580,N_11683,N_11625);
nor U17581 (N_17581,N_13681,N_14727);
xor U17582 (N_17582,N_11757,N_10414);
or U17583 (N_17583,N_11999,N_12137);
nor U17584 (N_17584,N_13342,N_14342);
nor U17585 (N_17585,N_10873,N_14389);
or U17586 (N_17586,N_14054,N_13740);
or U17587 (N_17587,N_14118,N_14431);
nand U17588 (N_17588,N_10905,N_14723);
nand U17589 (N_17589,N_10967,N_14532);
nand U17590 (N_17590,N_14065,N_12501);
and U17591 (N_17591,N_10398,N_10331);
nor U17592 (N_17592,N_14349,N_14252);
xnor U17593 (N_17593,N_13956,N_12128);
nand U17594 (N_17594,N_14573,N_13162);
xor U17595 (N_17595,N_10614,N_13773);
xnor U17596 (N_17596,N_10510,N_10649);
or U17597 (N_17597,N_10000,N_11952);
or U17598 (N_17598,N_11040,N_10891);
nand U17599 (N_17599,N_13456,N_12060);
nand U17600 (N_17600,N_14885,N_11053);
xnor U17601 (N_17601,N_13137,N_13309);
nand U17602 (N_17602,N_10423,N_12666);
nand U17603 (N_17603,N_12852,N_14299);
xnor U17604 (N_17604,N_11894,N_11257);
or U17605 (N_17605,N_11827,N_10009);
xor U17606 (N_17606,N_10432,N_11388);
and U17607 (N_17607,N_10878,N_10962);
nand U17608 (N_17608,N_14300,N_13545);
or U17609 (N_17609,N_14783,N_10431);
nand U17610 (N_17610,N_10438,N_10724);
nand U17611 (N_17611,N_13744,N_11808);
xnor U17612 (N_17612,N_14167,N_14031);
or U17613 (N_17613,N_11454,N_12925);
nand U17614 (N_17614,N_12001,N_12670);
or U17615 (N_17615,N_14025,N_10389);
or U17616 (N_17616,N_14650,N_14951);
nand U17617 (N_17617,N_14622,N_12287);
and U17618 (N_17618,N_14983,N_12240);
or U17619 (N_17619,N_10054,N_11979);
nor U17620 (N_17620,N_14661,N_14899);
or U17621 (N_17621,N_11152,N_11544);
nand U17622 (N_17622,N_10691,N_14576);
nor U17623 (N_17623,N_11311,N_11564);
nand U17624 (N_17624,N_10296,N_14215);
nand U17625 (N_17625,N_10780,N_13689);
or U17626 (N_17626,N_10933,N_10731);
nor U17627 (N_17627,N_10585,N_11165);
nand U17628 (N_17628,N_13413,N_10500);
nor U17629 (N_17629,N_11191,N_13488);
nand U17630 (N_17630,N_13263,N_12812);
xor U17631 (N_17631,N_10352,N_10163);
xnor U17632 (N_17632,N_13297,N_14653);
or U17633 (N_17633,N_11500,N_12033);
xnor U17634 (N_17634,N_12230,N_12907);
xnor U17635 (N_17635,N_11990,N_10974);
xnor U17636 (N_17636,N_10123,N_10986);
nand U17637 (N_17637,N_13759,N_10558);
xor U17638 (N_17638,N_13013,N_14930);
xor U17639 (N_17639,N_11950,N_10251);
nand U17640 (N_17640,N_10610,N_14709);
nand U17641 (N_17641,N_12176,N_13239);
or U17642 (N_17642,N_11246,N_12853);
or U17643 (N_17643,N_11577,N_12776);
and U17644 (N_17644,N_10298,N_11713);
and U17645 (N_17645,N_11249,N_11667);
nor U17646 (N_17646,N_11468,N_13645);
nand U17647 (N_17647,N_11955,N_14653);
xor U17648 (N_17648,N_13531,N_14399);
or U17649 (N_17649,N_12394,N_11614);
and U17650 (N_17650,N_13487,N_11046);
nor U17651 (N_17651,N_10817,N_14818);
or U17652 (N_17652,N_14591,N_11506);
or U17653 (N_17653,N_14150,N_11804);
or U17654 (N_17654,N_14380,N_14543);
nand U17655 (N_17655,N_11327,N_10532);
nor U17656 (N_17656,N_10068,N_10702);
or U17657 (N_17657,N_12192,N_14937);
or U17658 (N_17658,N_12854,N_13462);
nand U17659 (N_17659,N_10513,N_12988);
or U17660 (N_17660,N_10552,N_10385);
and U17661 (N_17661,N_14371,N_11735);
nor U17662 (N_17662,N_13313,N_11673);
nand U17663 (N_17663,N_14937,N_10123);
or U17664 (N_17664,N_12076,N_11828);
or U17665 (N_17665,N_10449,N_13621);
nand U17666 (N_17666,N_10568,N_10843);
nor U17667 (N_17667,N_10798,N_10976);
nor U17668 (N_17668,N_10321,N_12884);
xnor U17669 (N_17669,N_13512,N_11782);
or U17670 (N_17670,N_12148,N_13062);
nand U17671 (N_17671,N_12409,N_13206);
and U17672 (N_17672,N_13872,N_10936);
xnor U17673 (N_17673,N_11395,N_13505);
and U17674 (N_17674,N_11245,N_13163);
and U17675 (N_17675,N_14896,N_12404);
xor U17676 (N_17676,N_13883,N_13798);
xnor U17677 (N_17677,N_14407,N_12053);
or U17678 (N_17678,N_14645,N_14053);
and U17679 (N_17679,N_12597,N_10042);
nor U17680 (N_17680,N_10458,N_13912);
and U17681 (N_17681,N_11725,N_14811);
and U17682 (N_17682,N_12350,N_10641);
and U17683 (N_17683,N_11832,N_14169);
nand U17684 (N_17684,N_14789,N_12934);
nor U17685 (N_17685,N_13716,N_12027);
and U17686 (N_17686,N_14020,N_11246);
nand U17687 (N_17687,N_13422,N_14702);
xnor U17688 (N_17688,N_12239,N_10879);
xor U17689 (N_17689,N_10139,N_14896);
and U17690 (N_17690,N_14565,N_10804);
nand U17691 (N_17691,N_14328,N_13948);
or U17692 (N_17692,N_14157,N_12806);
and U17693 (N_17693,N_14806,N_10176);
nor U17694 (N_17694,N_14716,N_13254);
nand U17695 (N_17695,N_12123,N_11067);
and U17696 (N_17696,N_10417,N_12359);
nand U17697 (N_17697,N_12514,N_14069);
nand U17698 (N_17698,N_12700,N_12911);
or U17699 (N_17699,N_14569,N_14297);
nor U17700 (N_17700,N_10330,N_13660);
and U17701 (N_17701,N_10984,N_14271);
nand U17702 (N_17702,N_10331,N_12860);
or U17703 (N_17703,N_12651,N_12637);
and U17704 (N_17704,N_12313,N_10930);
or U17705 (N_17705,N_13502,N_11919);
or U17706 (N_17706,N_11708,N_11876);
nor U17707 (N_17707,N_13091,N_11928);
nor U17708 (N_17708,N_14931,N_14568);
nor U17709 (N_17709,N_12260,N_14066);
and U17710 (N_17710,N_14445,N_13094);
nor U17711 (N_17711,N_11633,N_10062);
nand U17712 (N_17712,N_10580,N_13857);
and U17713 (N_17713,N_10387,N_11718);
nand U17714 (N_17714,N_14715,N_10518);
nor U17715 (N_17715,N_14939,N_13588);
nand U17716 (N_17716,N_11186,N_13952);
and U17717 (N_17717,N_12172,N_12876);
and U17718 (N_17718,N_11646,N_12602);
or U17719 (N_17719,N_13144,N_14311);
or U17720 (N_17720,N_10187,N_13807);
xnor U17721 (N_17721,N_12279,N_10874);
nand U17722 (N_17722,N_10179,N_12344);
or U17723 (N_17723,N_14427,N_12949);
or U17724 (N_17724,N_13134,N_13887);
nand U17725 (N_17725,N_14211,N_14841);
and U17726 (N_17726,N_11788,N_13522);
xor U17727 (N_17727,N_12348,N_13467);
xnor U17728 (N_17728,N_14264,N_13170);
xnor U17729 (N_17729,N_12001,N_11656);
xnor U17730 (N_17730,N_12011,N_11231);
and U17731 (N_17731,N_11370,N_14547);
xor U17732 (N_17732,N_10383,N_13750);
and U17733 (N_17733,N_10683,N_12872);
nand U17734 (N_17734,N_12089,N_12452);
or U17735 (N_17735,N_11102,N_12749);
nor U17736 (N_17736,N_11184,N_11158);
or U17737 (N_17737,N_13601,N_10257);
xor U17738 (N_17738,N_11987,N_12861);
and U17739 (N_17739,N_14855,N_11551);
and U17740 (N_17740,N_12353,N_12585);
nor U17741 (N_17741,N_11176,N_10282);
nand U17742 (N_17742,N_10676,N_12349);
or U17743 (N_17743,N_10172,N_13262);
xor U17744 (N_17744,N_10209,N_12216);
nand U17745 (N_17745,N_10588,N_12633);
or U17746 (N_17746,N_13134,N_14873);
and U17747 (N_17747,N_13157,N_11639);
or U17748 (N_17748,N_13052,N_12110);
nor U17749 (N_17749,N_11153,N_14378);
and U17750 (N_17750,N_11707,N_14228);
nand U17751 (N_17751,N_14996,N_12852);
or U17752 (N_17752,N_13293,N_14113);
nand U17753 (N_17753,N_13850,N_11451);
nor U17754 (N_17754,N_10638,N_11414);
or U17755 (N_17755,N_13402,N_12569);
nand U17756 (N_17756,N_11563,N_12628);
or U17757 (N_17757,N_12150,N_13833);
xnor U17758 (N_17758,N_10810,N_10980);
xor U17759 (N_17759,N_12125,N_12347);
nand U17760 (N_17760,N_11515,N_12951);
nand U17761 (N_17761,N_10140,N_10856);
nor U17762 (N_17762,N_13843,N_13053);
xnor U17763 (N_17763,N_12101,N_14451);
nand U17764 (N_17764,N_12858,N_12475);
nand U17765 (N_17765,N_10756,N_13336);
and U17766 (N_17766,N_10544,N_10493);
nand U17767 (N_17767,N_13565,N_10141);
nor U17768 (N_17768,N_13659,N_14697);
xor U17769 (N_17769,N_13210,N_11188);
or U17770 (N_17770,N_13519,N_14270);
or U17771 (N_17771,N_12756,N_13635);
or U17772 (N_17772,N_12947,N_11602);
and U17773 (N_17773,N_14355,N_10636);
or U17774 (N_17774,N_11649,N_10314);
xnor U17775 (N_17775,N_11626,N_12250);
and U17776 (N_17776,N_13431,N_14964);
or U17777 (N_17777,N_14664,N_11735);
and U17778 (N_17778,N_11748,N_14478);
nand U17779 (N_17779,N_10320,N_11619);
nand U17780 (N_17780,N_10464,N_12102);
nand U17781 (N_17781,N_11206,N_12083);
nand U17782 (N_17782,N_13039,N_12279);
nor U17783 (N_17783,N_11513,N_13450);
and U17784 (N_17784,N_10708,N_13262);
and U17785 (N_17785,N_12767,N_14251);
and U17786 (N_17786,N_12684,N_14631);
nand U17787 (N_17787,N_11601,N_11520);
and U17788 (N_17788,N_14077,N_12310);
and U17789 (N_17789,N_10695,N_14696);
and U17790 (N_17790,N_13984,N_12912);
nor U17791 (N_17791,N_13913,N_12029);
or U17792 (N_17792,N_12885,N_13007);
nor U17793 (N_17793,N_14226,N_12799);
and U17794 (N_17794,N_13886,N_12440);
nand U17795 (N_17795,N_14869,N_11322);
xor U17796 (N_17796,N_13297,N_10850);
nor U17797 (N_17797,N_13281,N_14053);
nor U17798 (N_17798,N_12304,N_12448);
and U17799 (N_17799,N_14221,N_12932);
xor U17800 (N_17800,N_10783,N_10552);
nand U17801 (N_17801,N_11033,N_13362);
nor U17802 (N_17802,N_14564,N_12053);
nand U17803 (N_17803,N_10768,N_12560);
or U17804 (N_17804,N_13757,N_11373);
nand U17805 (N_17805,N_13844,N_13565);
nor U17806 (N_17806,N_10028,N_10101);
nand U17807 (N_17807,N_13995,N_14024);
xnor U17808 (N_17808,N_10748,N_12458);
nor U17809 (N_17809,N_11602,N_14721);
xnor U17810 (N_17810,N_12491,N_11271);
nor U17811 (N_17811,N_14996,N_11348);
nand U17812 (N_17812,N_14760,N_11794);
xnor U17813 (N_17813,N_13658,N_13523);
or U17814 (N_17814,N_13709,N_10107);
and U17815 (N_17815,N_14128,N_14140);
xor U17816 (N_17816,N_14542,N_12719);
xor U17817 (N_17817,N_11505,N_12936);
xor U17818 (N_17818,N_12348,N_10476);
and U17819 (N_17819,N_14635,N_11081);
and U17820 (N_17820,N_14790,N_10621);
nor U17821 (N_17821,N_10227,N_11485);
xnor U17822 (N_17822,N_10085,N_10119);
xor U17823 (N_17823,N_13091,N_10456);
xnor U17824 (N_17824,N_13255,N_11442);
or U17825 (N_17825,N_10770,N_14761);
xnor U17826 (N_17826,N_11553,N_10675);
and U17827 (N_17827,N_14738,N_14103);
nor U17828 (N_17828,N_11885,N_12155);
and U17829 (N_17829,N_12823,N_13191);
and U17830 (N_17830,N_11358,N_14108);
nor U17831 (N_17831,N_11944,N_10730);
nor U17832 (N_17832,N_11988,N_14918);
or U17833 (N_17833,N_13050,N_12686);
or U17834 (N_17834,N_14669,N_14904);
nor U17835 (N_17835,N_13044,N_13238);
or U17836 (N_17836,N_14098,N_12324);
or U17837 (N_17837,N_13575,N_12918);
or U17838 (N_17838,N_10214,N_14515);
xor U17839 (N_17839,N_13143,N_10772);
xor U17840 (N_17840,N_13416,N_11449);
nor U17841 (N_17841,N_14171,N_12325);
xnor U17842 (N_17842,N_11539,N_10681);
or U17843 (N_17843,N_10460,N_12038);
nor U17844 (N_17844,N_11983,N_10574);
nand U17845 (N_17845,N_12360,N_12179);
or U17846 (N_17846,N_11854,N_11699);
nor U17847 (N_17847,N_11766,N_10274);
and U17848 (N_17848,N_10927,N_13613);
nand U17849 (N_17849,N_13144,N_11304);
or U17850 (N_17850,N_10053,N_12143);
or U17851 (N_17851,N_10940,N_10201);
or U17852 (N_17852,N_13751,N_14360);
or U17853 (N_17853,N_12701,N_12695);
and U17854 (N_17854,N_12896,N_13734);
xor U17855 (N_17855,N_10519,N_13031);
or U17856 (N_17856,N_13177,N_14970);
or U17857 (N_17857,N_13205,N_10387);
xor U17858 (N_17858,N_14177,N_11842);
nand U17859 (N_17859,N_10508,N_10160);
nand U17860 (N_17860,N_14668,N_14107);
or U17861 (N_17861,N_14130,N_13756);
and U17862 (N_17862,N_10283,N_11136);
and U17863 (N_17863,N_11114,N_13931);
and U17864 (N_17864,N_13923,N_11923);
nor U17865 (N_17865,N_12412,N_14887);
xor U17866 (N_17866,N_13805,N_10231);
nand U17867 (N_17867,N_12886,N_10567);
nor U17868 (N_17868,N_12364,N_10050);
nand U17869 (N_17869,N_12012,N_10309);
and U17870 (N_17870,N_13004,N_10200);
or U17871 (N_17871,N_11645,N_14859);
and U17872 (N_17872,N_11123,N_10069);
and U17873 (N_17873,N_12790,N_10694);
or U17874 (N_17874,N_10571,N_10022);
xor U17875 (N_17875,N_14123,N_13378);
nor U17876 (N_17876,N_13175,N_13062);
nand U17877 (N_17877,N_12223,N_10341);
nand U17878 (N_17878,N_12843,N_13529);
or U17879 (N_17879,N_10125,N_14048);
or U17880 (N_17880,N_11504,N_10744);
or U17881 (N_17881,N_11291,N_12220);
or U17882 (N_17882,N_12723,N_11744);
and U17883 (N_17883,N_13937,N_10357);
nand U17884 (N_17884,N_12871,N_14290);
xnor U17885 (N_17885,N_11129,N_14706);
and U17886 (N_17886,N_14383,N_10493);
nand U17887 (N_17887,N_13987,N_14575);
or U17888 (N_17888,N_13327,N_13754);
nand U17889 (N_17889,N_13278,N_13797);
nand U17890 (N_17890,N_14552,N_12533);
nor U17891 (N_17891,N_12917,N_10404);
and U17892 (N_17892,N_14024,N_12161);
or U17893 (N_17893,N_12382,N_14697);
and U17894 (N_17894,N_11889,N_14746);
nor U17895 (N_17895,N_14042,N_11094);
or U17896 (N_17896,N_13825,N_10956);
and U17897 (N_17897,N_10632,N_14845);
and U17898 (N_17898,N_10905,N_12869);
xor U17899 (N_17899,N_10085,N_12705);
xor U17900 (N_17900,N_12792,N_13499);
or U17901 (N_17901,N_13781,N_10405);
nand U17902 (N_17902,N_10762,N_11204);
xnor U17903 (N_17903,N_10573,N_11276);
or U17904 (N_17904,N_10969,N_14809);
or U17905 (N_17905,N_11037,N_14403);
xor U17906 (N_17906,N_12841,N_12953);
nor U17907 (N_17907,N_10716,N_11947);
xor U17908 (N_17908,N_12929,N_11901);
xnor U17909 (N_17909,N_10027,N_10993);
nor U17910 (N_17910,N_10979,N_13213);
and U17911 (N_17911,N_14350,N_10461);
and U17912 (N_17912,N_13842,N_14148);
or U17913 (N_17913,N_14939,N_10352);
nor U17914 (N_17914,N_12399,N_12842);
nor U17915 (N_17915,N_10346,N_12303);
and U17916 (N_17916,N_11743,N_11302);
nand U17917 (N_17917,N_14217,N_13808);
nor U17918 (N_17918,N_11496,N_10683);
and U17919 (N_17919,N_14192,N_11696);
xnor U17920 (N_17920,N_12863,N_12827);
nor U17921 (N_17921,N_14885,N_14998);
and U17922 (N_17922,N_11260,N_10598);
nor U17923 (N_17923,N_12615,N_11085);
and U17924 (N_17924,N_13391,N_12017);
xor U17925 (N_17925,N_11873,N_10707);
nor U17926 (N_17926,N_14713,N_10792);
nand U17927 (N_17927,N_10355,N_10291);
or U17928 (N_17928,N_12666,N_13850);
nor U17929 (N_17929,N_12279,N_12568);
and U17930 (N_17930,N_14269,N_11982);
xnor U17931 (N_17931,N_12606,N_14362);
nor U17932 (N_17932,N_14204,N_13038);
nor U17933 (N_17933,N_13415,N_10368);
nor U17934 (N_17934,N_12244,N_11882);
nand U17935 (N_17935,N_12362,N_14094);
xnor U17936 (N_17936,N_11789,N_12086);
or U17937 (N_17937,N_14975,N_14762);
and U17938 (N_17938,N_12560,N_11201);
or U17939 (N_17939,N_13599,N_12221);
nand U17940 (N_17940,N_12018,N_13106);
nor U17941 (N_17941,N_13882,N_10990);
nor U17942 (N_17942,N_10996,N_13480);
or U17943 (N_17943,N_10691,N_12325);
nor U17944 (N_17944,N_10593,N_10614);
xnor U17945 (N_17945,N_13492,N_11355);
nor U17946 (N_17946,N_10368,N_10148);
xnor U17947 (N_17947,N_11192,N_11066);
and U17948 (N_17948,N_10719,N_10672);
nand U17949 (N_17949,N_12312,N_14698);
xnor U17950 (N_17950,N_10850,N_11653);
and U17951 (N_17951,N_14557,N_14245);
or U17952 (N_17952,N_12562,N_10446);
nor U17953 (N_17953,N_11461,N_10344);
xnor U17954 (N_17954,N_14308,N_10521);
and U17955 (N_17955,N_14140,N_14229);
xor U17956 (N_17956,N_11201,N_10833);
nor U17957 (N_17957,N_10108,N_10077);
nor U17958 (N_17958,N_13090,N_14420);
xnor U17959 (N_17959,N_11574,N_11471);
and U17960 (N_17960,N_12053,N_12801);
nor U17961 (N_17961,N_14801,N_14802);
nand U17962 (N_17962,N_12409,N_13794);
nor U17963 (N_17963,N_10300,N_14918);
or U17964 (N_17964,N_10995,N_12980);
nand U17965 (N_17965,N_14115,N_14926);
nor U17966 (N_17966,N_12501,N_12116);
xor U17967 (N_17967,N_11273,N_12152);
and U17968 (N_17968,N_11484,N_10671);
and U17969 (N_17969,N_10370,N_12721);
nand U17970 (N_17970,N_13995,N_11907);
or U17971 (N_17971,N_14038,N_13579);
xor U17972 (N_17972,N_13186,N_10254);
nand U17973 (N_17973,N_12266,N_14807);
nand U17974 (N_17974,N_11324,N_14574);
xor U17975 (N_17975,N_10589,N_11982);
and U17976 (N_17976,N_12626,N_10419);
nor U17977 (N_17977,N_12559,N_10270);
nand U17978 (N_17978,N_13565,N_13869);
or U17979 (N_17979,N_12545,N_13840);
nand U17980 (N_17980,N_10617,N_12988);
nor U17981 (N_17981,N_11945,N_13550);
or U17982 (N_17982,N_13148,N_10335);
nor U17983 (N_17983,N_14096,N_10506);
nand U17984 (N_17984,N_12371,N_10141);
xnor U17985 (N_17985,N_11486,N_10617);
or U17986 (N_17986,N_12946,N_11944);
nand U17987 (N_17987,N_14971,N_12823);
nor U17988 (N_17988,N_14266,N_12784);
or U17989 (N_17989,N_14506,N_14637);
nor U17990 (N_17990,N_14400,N_12366);
or U17991 (N_17991,N_11576,N_14331);
nand U17992 (N_17992,N_11691,N_13880);
xor U17993 (N_17993,N_12039,N_13078);
nand U17994 (N_17994,N_14175,N_11301);
nor U17995 (N_17995,N_10108,N_12125);
or U17996 (N_17996,N_13460,N_11681);
xor U17997 (N_17997,N_11579,N_14202);
or U17998 (N_17998,N_14458,N_14676);
and U17999 (N_17999,N_14687,N_14307);
nor U18000 (N_18000,N_10703,N_10550);
xor U18001 (N_18001,N_13034,N_12460);
xor U18002 (N_18002,N_13455,N_12139);
nand U18003 (N_18003,N_12080,N_13058);
or U18004 (N_18004,N_10738,N_11696);
and U18005 (N_18005,N_10148,N_13342);
and U18006 (N_18006,N_10943,N_13399);
xnor U18007 (N_18007,N_10741,N_12652);
nor U18008 (N_18008,N_12930,N_11663);
nand U18009 (N_18009,N_12998,N_11744);
nand U18010 (N_18010,N_13214,N_12087);
xor U18011 (N_18011,N_12113,N_12511);
nor U18012 (N_18012,N_12501,N_14353);
nand U18013 (N_18013,N_12034,N_11983);
nor U18014 (N_18014,N_13061,N_13224);
and U18015 (N_18015,N_14308,N_12301);
or U18016 (N_18016,N_10056,N_11896);
nand U18017 (N_18017,N_11728,N_11702);
or U18018 (N_18018,N_13468,N_14612);
or U18019 (N_18019,N_12701,N_10945);
and U18020 (N_18020,N_13390,N_10763);
nor U18021 (N_18021,N_10881,N_14389);
or U18022 (N_18022,N_10443,N_12854);
nor U18023 (N_18023,N_12705,N_11108);
xor U18024 (N_18024,N_11182,N_11156);
xor U18025 (N_18025,N_13436,N_14857);
xnor U18026 (N_18026,N_14586,N_10705);
and U18027 (N_18027,N_11583,N_12423);
and U18028 (N_18028,N_11222,N_12024);
or U18029 (N_18029,N_12027,N_14144);
and U18030 (N_18030,N_12185,N_11537);
nand U18031 (N_18031,N_14073,N_11026);
and U18032 (N_18032,N_13917,N_11731);
nor U18033 (N_18033,N_11742,N_14031);
and U18034 (N_18034,N_13554,N_14871);
or U18035 (N_18035,N_10920,N_14050);
xor U18036 (N_18036,N_13970,N_13176);
nor U18037 (N_18037,N_11842,N_12707);
or U18038 (N_18038,N_10422,N_14214);
xor U18039 (N_18039,N_14834,N_11419);
xor U18040 (N_18040,N_12673,N_12122);
nand U18041 (N_18041,N_13558,N_12701);
nand U18042 (N_18042,N_12061,N_13998);
or U18043 (N_18043,N_14696,N_13124);
nand U18044 (N_18044,N_13894,N_14859);
and U18045 (N_18045,N_14803,N_12655);
xor U18046 (N_18046,N_12261,N_12782);
and U18047 (N_18047,N_12536,N_12877);
or U18048 (N_18048,N_13549,N_13532);
and U18049 (N_18049,N_10991,N_11893);
and U18050 (N_18050,N_13818,N_11715);
xnor U18051 (N_18051,N_12437,N_13857);
nand U18052 (N_18052,N_14816,N_12731);
nor U18053 (N_18053,N_13421,N_14817);
and U18054 (N_18054,N_13119,N_11313);
nand U18055 (N_18055,N_11190,N_11676);
nand U18056 (N_18056,N_14567,N_14690);
or U18057 (N_18057,N_13593,N_10038);
and U18058 (N_18058,N_14849,N_12896);
nand U18059 (N_18059,N_12522,N_12068);
and U18060 (N_18060,N_11362,N_10925);
or U18061 (N_18061,N_14027,N_10223);
and U18062 (N_18062,N_14104,N_13298);
xor U18063 (N_18063,N_12330,N_13373);
xnor U18064 (N_18064,N_13864,N_10229);
or U18065 (N_18065,N_14085,N_11030);
and U18066 (N_18066,N_13886,N_14409);
and U18067 (N_18067,N_10027,N_13402);
or U18068 (N_18068,N_12531,N_10914);
nand U18069 (N_18069,N_11012,N_12224);
or U18070 (N_18070,N_11287,N_10148);
nor U18071 (N_18071,N_13663,N_10945);
xor U18072 (N_18072,N_10985,N_11701);
nor U18073 (N_18073,N_11099,N_11708);
nor U18074 (N_18074,N_10916,N_14542);
xnor U18075 (N_18075,N_13123,N_13552);
xnor U18076 (N_18076,N_13468,N_14352);
xor U18077 (N_18077,N_12940,N_13387);
and U18078 (N_18078,N_13526,N_10389);
nand U18079 (N_18079,N_10672,N_11438);
xor U18080 (N_18080,N_12204,N_10279);
nand U18081 (N_18081,N_10012,N_12811);
xor U18082 (N_18082,N_14360,N_12402);
nor U18083 (N_18083,N_13898,N_12484);
xnor U18084 (N_18084,N_12075,N_12587);
nor U18085 (N_18085,N_12158,N_14707);
nand U18086 (N_18086,N_14246,N_12140);
xor U18087 (N_18087,N_10303,N_11757);
nand U18088 (N_18088,N_14183,N_12632);
nor U18089 (N_18089,N_10427,N_11982);
xnor U18090 (N_18090,N_10568,N_10802);
xor U18091 (N_18091,N_13840,N_11089);
nand U18092 (N_18092,N_13253,N_12590);
and U18093 (N_18093,N_13429,N_13182);
nor U18094 (N_18094,N_13613,N_11472);
or U18095 (N_18095,N_10082,N_12908);
nor U18096 (N_18096,N_10211,N_12305);
nand U18097 (N_18097,N_10623,N_11164);
and U18098 (N_18098,N_14314,N_11439);
and U18099 (N_18099,N_13464,N_14611);
and U18100 (N_18100,N_11816,N_11488);
nor U18101 (N_18101,N_14454,N_11657);
xnor U18102 (N_18102,N_12243,N_13719);
nor U18103 (N_18103,N_13583,N_10261);
nor U18104 (N_18104,N_11657,N_11738);
xor U18105 (N_18105,N_13011,N_13861);
xor U18106 (N_18106,N_10419,N_13239);
and U18107 (N_18107,N_13865,N_11679);
or U18108 (N_18108,N_12140,N_14263);
and U18109 (N_18109,N_12341,N_10618);
and U18110 (N_18110,N_12004,N_10993);
nand U18111 (N_18111,N_14080,N_14504);
or U18112 (N_18112,N_13177,N_13800);
xnor U18113 (N_18113,N_14185,N_11569);
nor U18114 (N_18114,N_10294,N_13238);
and U18115 (N_18115,N_13814,N_13371);
xor U18116 (N_18116,N_10958,N_13200);
or U18117 (N_18117,N_14053,N_12388);
nand U18118 (N_18118,N_14895,N_14132);
nor U18119 (N_18119,N_13141,N_10801);
nor U18120 (N_18120,N_10680,N_14108);
or U18121 (N_18121,N_10744,N_14887);
nor U18122 (N_18122,N_10134,N_11260);
nor U18123 (N_18123,N_11560,N_11503);
nor U18124 (N_18124,N_14440,N_12528);
nand U18125 (N_18125,N_12092,N_12177);
or U18126 (N_18126,N_11548,N_11137);
and U18127 (N_18127,N_12901,N_13733);
nand U18128 (N_18128,N_10595,N_14461);
or U18129 (N_18129,N_11145,N_11908);
nand U18130 (N_18130,N_10347,N_13774);
nor U18131 (N_18131,N_14386,N_13642);
xnor U18132 (N_18132,N_14885,N_12547);
and U18133 (N_18133,N_14608,N_10785);
and U18134 (N_18134,N_14238,N_11623);
nor U18135 (N_18135,N_13688,N_13004);
and U18136 (N_18136,N_10061,N_11301);
nor U18137 (N_18137,N_11505,N_14868);
nor U18138 (N_18138,N_12041,N_14869);
or U18139 (N_18139,N_10774,N_13278);
and U18140 (N_18140,N_12015,N_14578);
or U18141 (N_18141,N_10048,N_11619);
nand U18142 (N_18142,N_14277,N_10743);
xor U18143 (N_18143,N_11605,N_11842);
xnor U18144 (N_18144,N_10239,N_10628);
xor U18145 (N_18145,N_10074,N_13249);
and U18146 (N_18146,N_11337,N_12787);
and U18147 (N_18147,N_13322,N_10596);
or U18148 (N_18148,N_12421,N_13649);
or U18149 (N_18149,N_14797,N_14716);
and U18150 (N_18150,N_14205,N_10296);
or U18151 (N_18151,N_12291,N_13517);
nor U18152 (N_18152,N_13440,N_10929);
xnor U18153 (N_18153,N_10848,N_14969);
or U18154 (N_18154,N_13804,N_12264);
nand U18155 (N_18155,N_10029,N_11727);
nor U18156 (N_18156,N_13125,N_14652);
nor U18157 (N_18157,N_10169,N_11417);
xnor U18158 (N_18158,N_10099,N_13268);
or U18159 (N_18159,N_13798,N_11775);
and U18160 (N_18160,N_10577,N_12192);
nor U18161 (N_18161,N_13340,N_14023);
nor U18162 (N_18162,N_10558,N_10419);
xor U18163 (N_18163,N_10263,N_10676);
xor U18164 (N_18164,N_13139,N_13108);
xnor U18165 (N_18165,N_11847,N_11644);
and U18166 (N_18166,N_10230,N_12308);
and U18167 (N_18167,N_11020,N_14142);
or U18168 (N_18168,N_14801,N_13032);
xor U18169 (N_18169,N_14393,N_12060);
nand U18170 (N_18170,N_10339,N_14689);
nand U18171 (N_18171,N_10714,N_13877);
nor U18172 (N_18172,N_13652,N_11368);
or U18173 (N_18173,N_14624,N_12248);
nor U18174 (N_18174,N_12313,N_12446);
nand U18175 (N_18175,N_13486,N_12818);
nor U18176 (N_18176,N_13666,N_11815);
nand U18177 (N_18177,N_12114,N_11110);
and U18178 (N_18178,N_11067,N_13845);
nor U18179 (N_18179,N_13004,N_13892);
nand U18180 (N_18180,N_10978,N_11504);
nor U18181 (N_18181,N_12876,N_12846);
xor U18182 (N_18182,N_10381,N_11736);
nor U18183 (N_18183,N_11027,N_12217);
nand U18184 (N_18184,N_13303,N_11513);
or U18185 (N_18185,N_12330,N_10011);
nand U18186 (N_18186,N_10649,N_13606);
xnor U18187 (N_18187,N_10337,N_12009);
or U18188 (N_18188,N_10003,N_14060);
and U18189 (N_18189,N_13990,N_11981);
or U18190 (N_18190,N_14789,N_10811);
nand U18191 (N_18191,N_11608,N_12217);
or U18192 (N_18192,N_12967,N_12143);
nor U18193 (N_18193,N_13966,N_11252);
or U18194 (N_18194,N_10332,N_10441);
or U18195 (N_18195,N_13310,N_14692);
and U18196 (N_18196,N_12238,N_11660);
xor U18197 (N_18197,N_14033,N_12611);
nor U18198 (N_18198,N_13330,N_14295);
xnor U18199 (N_18199,N_12366,N_14554);
xor U18200 (N_18200,N_13124,N_13385);
nand U18201 (N_18201,N_12099,N_12193);
xor U18202 (N_18202,N_11195,N_10723);
and U18203 (N_18203,N_14985,N_10727);
nor U18204 (N_18204,N_14426,N_13483);
nor U18205 (N_18205,N_11281,N_13424);
nor U18206 (N_18206,N_12924,N_11427);
nand U18207 (N_18207,N_11467,N_14230);
nor U18208 (N_18208,N_13269,N_11680);
and U18209 (N_18209,N_11700,N_13212);
nand U18210 (N_18210,N_14334,N_12519);
nor U18211 (N_18211,N_10421,N_13421);
xnor U18212 (N_18212,N_13769,N_11881);
xnor U18213 (N_18213,N_14304,N_11277);
and U18214 (N_18214,N_10958,N_10893);
nor U18215 (N_18215,N_13848,N_11038);
or U18216 (N_18216,N_11578,N_14832);
or U18217 (N_18217,N_10478,N_14757);
or U18218 (N_18218,N_13721,N_11612);
xnor U18219 (N_18219,N_11587,N_11211);
and U18220 (N_18220,N_10977,N_13378);
xnor U18221 (N_18221,N_14729,N_13325);
and U18222 (N_18222,N_14591,N_11390);
nor U18223 (N_18223,N_10535,N_10019);
or U18224 (N_18224,N_12921,N_10173);
and U18225 (N_18225,N_12724,N_13631);
nor U18226 (N_18226,N_12976,N_11857);
nor U18227 (N_18227,N_14548,N_14509);
nand U18228 (N_18228,N_12884,N_11076);
or U18229 (N_18229,N_14604,N_12889);
or U18230 (N_18230,N_14665,N_11121);
and U18231 (N_18231,N_13763,N_10971);
nor U18232 (N_18232,N_14779,N_10125);
or U18233 (N_18233,N_13814,N_13199);
xor U18234 (N_18234,N_12183,N_13124);
or U18235 (N_18235,N_11044,N_11426);
xnor U18236 (N_18236,N_14014,N_12541);
nor U18237 (N_18237,N_12938,N_11138);
nor U18238 (N_18238,N_12045,N_14320);
and U18239 (N_18239,N_12954,N_12807);
nand U18240 (N_18240,N_13909,N_12934);
xnor U18241 (N_18241,N_13513,N_12739);
nand U18242 (N_18242,N_11336,N_10629);
and U18243 (N_18243,N_12185,N_12103);
nand U18244 (N_18244,N_13425,N_10485);
xnor U18245 (N_18245,N_11688,N_12861);
and U18246 (N_18246,N_14721,N_14536);
or U18247 (N_18247,N_11026,N_11046);
and U18248 (N_18248,N_12617,N_10876);
and U18249 (N_18249,N_12335,N_12827);
nand U18250 (N_18250,N_12678,N_12564);
nor U18251 (N_18251,N_14196,N_14700);
or U18252 (N_18252,N_12565,N_10904);
nand U18253 (N_18253,N_11973,N_13735);
and U18254 (N_18254,N_11311,N_12581);
nor U18255 (N_18255,N_14118,N_11003);
xnor U18256 (N_18256,N_12066,N_13091);
xor U18257 (N_18257,N_10158,N_14076);
nand U18258 (N_18258,N_14570,N_12412);
nand U18259 (N_18259,N_13322,N_10933);
and U18260 (N_18260,N_11428,N_11534);
nand U18261 (N_18261,N_13627,N_10833);
and U18262 (N_18262,N_13167,N_10531);
xor U18263 (N_18263,N_10991,N_10803);
and U18264 (N_18264,N_13783,N_10485);
nand U18265 (N_18265,N_12643,N_11707);
xnor U18266 (N_18266,N_10236,N_14465);
xnor U18267 (N_18267,N_11805,N_11886);
xnor U18268 (N_18268,N_13019,N_13360);
or U18269 (N_18269,N_11493,N_10371);
or U18270 (N_18270,N_10335,N_13345);
or U18271 (N_18271,N_13450,N_14325);
nand U18272 (N_18272,N_12541,N_11808);
and U18273 (N_18273,N_10745,N_11260);
xor U18274 (N_18274,N_14387,N_13686);
and U18275 (N_18275,N_14152,N_13957);
nor U18276 (N_18276,N_12807,N_13668);
nor U18277 (N_18277,N_10534,N_12884);
xnor U18278 (N_18278,N_14548,N_12748);
or U18279 (N_18279,N_12603,N_14203);
or U18280 (N_18280,N_10013,N_12202);
nand U18281 (N_18281,N_14941,N_13287);
xnor U18282 (N_18282,N_10788,N_11715);
and U18283 (N_18283,N_10828,N_12262);
and U18284 (N_18284,N_12729,N_11028);
or U18285 (N_18285,N_12139,N_10548);
xnor U18286 (N_18286,N_11460,N_11428);
nor U18287 (N_18287,N_14228,N_12525);
nor U18288 (N_18288,N_10400,N_11574);
and U18289 (N_18289,N_10723,N_13463);
nand U18290 (N_18290,N_13553,N_13900);
nor U18291 (N_18291,N_12723,N_11420);
and U18292 (N_18292,N_11934,N_10782);
and U18293 (N_18293,N_11901,N_12559);
and U18294 (N_18294,N_12447,N_14969);
xnor U18295 (N_18295,N_11746,N_14437);
xor U18296 (N_18296,N_14066,N_12168);
nor U18297 (N_18297,N_10477,N_13301);
nor U18298 (N_18298,N_12296,N_10795);
or U18299 (N_18299,N_13667,N_10552);
or U18300 (N_18300,N_11155,N_11696);
or U18301 (N_18301,N_12446,N_14099);
xnor U18302 (N_18302,N_13962,N_14365);
and U18303 (N_18303,N_12894,N_10038);
nor U18304 (N_18304,N_14704,N_12520);
or U18305 (N_18305,N_12093,N_14930);
nor U18306 (N_18306,N_10833,N_11415);
nand U18307 (N_18307,N_14692,N_14981);
nor U18308 (N_18308,N_11705,N_12079);
nand U18309 (N_18309,N_12146,N_14982);
xor U18310 (N_18310,N_13829,N_10157);
nand U18311 (N_18311,N_12732,N_11122);
and U18312 (N_18312,N_14443,N_12779);
or U18313 (N_18313,N_13362,N_12796);
nand U18314 (N_18314,N_11796,N_11637);
nor U18315 (N_18315,N_14899,N_12127);
xnor U18316 (N_18316,N_11340,N_13077);
xor U18317 (N_18317,N_12712,N_12205);
and U18318 (N_18318,N_10600,N_12045);
or U18319 (N_18319,N_12789,N_12078);
or U18320 (N_18320,N_14524,N_14715);
nor U18321 (N_18321,N_10418,N_12780);
or U18322 (N_18322,N_12303,N_14619);
nand U18323 (N_18323,N_14311,N_10200);
nor U18324 (N_18324,N_13003,N_10385);
nand U18325 (N_18325,N_14940,N_14730);
xnor U18326 (N_18326,N_14871,N_11669);
or U18327 (N_18327,N_13491,N_11947);
xor U18328 (N_18328,N_12056,N_11694);
xnor U18329 (N_18329,N_14671,N_11868);
nand U18330 (N_18330,N_14745,N_14111);
and U18331 (N_18331,N_12915,N_12339);
xor U18332 (N_18332,N_10653,N_10336);
nand U18333 (N_18333,N_14952,N_11324);
nand U18334 (N_18334,N_13589,N_13592);
or U18335 (N_18335,N_11124,N_12816);
and U18336 (N_18336,N_13952,N_10718);
or U18337 (N_18337,N_10303,N_12106);
nand U18338 (N_18338,N_12590,N_14731);
or U18339 (N_18339,N_11870,N_10098);
or U18340 (N_18340,N_10870,N_10574);
and U18341 (N_18341,N_11107,N_11875);
xnor U18342 (N_18342,N_12977,N_14543);
xnor U18343 (N_18343,N_10015,N_12224);
or U18344 (N_18344,N_12740,N_14659);
and U18345 (N_18345,N_10235,N_14240);
nor U18346 (N_18346,N_11386,N_11414);
or U18347 (N_18347,N_13524,N_13796);
nor U18348 (N_18348,N_13377,N_12861);
nand U18349 (N_18349,N_14297,N_10862);
and U18350 (N_18350,N_14520,N_11744);
and U18351 (N_18351,N_13861,N_14283);
nor U18352 (N_18352,N_13153,N_13214);
xor U18353 (N_18353,N_13170,N_10822);
nor U18354 (N_18354,N_14859,N_11134);
nand U18355 (N_18355,N_11858,N_11517);
and U18356 (N_18356,N_13885,N_11214);
nand U18357 (N_18357,N_12230,N_13356);
xnor U18358 (N_18358,N_14596,N_14024);
or U18359 (N_18359,N_14958,N_14963);
and U18360 (N_18360,N_14910,N_14467);
nor U18361 (N_18361,N_11532,N_11299);
nand U18362 (N_18362,N_12578,N_12188);
or U18363 (N_18363,N_11309,N_14206);
or U18364 (N_18364,N_14842,N_10454);
nor U18365 (N_18365,N_11221,N_14207);
and U18366 (N_18366,N_11869,N_10050);
xnor U18367 (N_18367,N_10342,N_14735);
or U18368 (N_18368,N_14788,N_11927);
and U18369 (N_18369,N_14390,N_10039);
and U18370 (N_18370,N_10702,N_11161);
nand U18371 (N_18371,N_14741,N_11438);
nor U18372 (N_18372,N_13951,N_14690);
nand U18373 (N_18373,N_10126,N_11315);
xor U18374 (N_18374,N_14929,N_14139);
and U18375 (N_18375,N_11205,N_14746);
nand U18376 (N_18376,N_12898,N_12865);
or U18377 (N_18377,N_13828,N_11536);
xnor U18378 (N_18378,N_10451,N_11334);
nand U18379 (N_18379,N_10084,N_12020);
or U18380 (N_18380,N_10574,N_10797);
nand U18381 (N_18381,N_10823,N_10733);
or U18382 (N_18382,N_10583,N_10009);
or U18383 (N_18383,N_10993,N_14195);
and U18384 (N_18384,N_10871,N_13895);
or U18385 (N_18385,N_12544,N_14858);
nand U18386 (N_18386,N_10140,N_12310);
nand U18387 (N_18387,N_14415,N_12730);
nor U18388 (N_18388,N_11603,N_12296);
xor U18389 (N_18389,N_12601,N_10524);
nand U18390 (N_18390,N_12956,N_13046);
xnor U18391 (N_18391,N_11729,N_10720);
and U18392 (N_18392,N_10504,N_13700);
nand U18393 (N_18393,N_13273,N_11396);
nand U18394 (N_18394,N_14890,N_14627);
nand U18395 (N_18395,N_11973,N_14696);
nand U18396 (N_18396,N_14053,N_14352);
nor U18397 (N_18397,N_12970,N_14256);
nor U18398 (N_18398,N_14595,N_11987);
and U18399 (N_18399,N_11131,N_14566);
nor U18400 (N_18400,N_14047,N_14002);
xnor U18401 (N_18401,N_12059,N_10731);
nor U18402 (N_18402,N_11080,N_12150);
nor U18403 (N_18403,N_11427,N_14602);
xnor U18404 (N_18404,N_11225,N_10048);
and U18405 (N_18405,N_10959,N_14713);
nand U18406 (N_18406,N_10077,N_11894);
or U18407 (N_18407,N_11810,N_10227);
xor U18408 (N_18408,N_14783,N_13038);
and U18409 (N_18409,N_12012,N_13841);
or U18410 (N_18410,N_10489,N_13345);
nand U18411 (N_18411,N_13179,N_14319);
or U18412 (N_18412,N_14557,N_12459);
nand U18413 (N_18413,N_11405,N_14405);
xnor U18414 (N_18414,N_11103,N_10948);
nor U18415 (N_18415,N_13881,N_13868);
xor U18416 (N_18416,N_14953,N_10523);
xnor U18417 (N_18417,N_11400,N_13308);
nor U18418 (N_18418,N_12878,N_13083);
nor U18419 (N_18419,N_12308,N_14248);
or U18420 (N_18420,N_10878,N_10193);
nand U18421 (N_18421,N_11125,N_11934);
nor U18422 (N_18422,N_10445,N_14959);
or U18423 (N_18423,N_12635,N_10487);
or U18424 (N_18424,N_12044,N_13173);
nor U18425 (N_18425,N_14286,N_14500);
xor U18426 (N_18426,N_10905,N_11578);
or U18427 (N_18427,N_11137,N_11700);
xor U18428 (N_18428,N_14354,N_13700);
and U18429 (N_18429,N_12888,N_12788);
and U18430 (N_18430,N_12284,N_11272);
xnor U18431 (N_18431,N_13261,N_10035);
and U18432 (N_18432,N_10194,N_10176);
or U18433 (N_18433,N_13584,N_11370);
nor U18434 (N_18434,N_13275,N_10735);
and U18435 (N_18435,N_12572,N_10056);
nand U18436 (N_18436,N_12581,N_11867);
and U18437 (N_18437,N_11518,N_10956);
nand U18438 (N_18438,N_10670,N_12317);
nor U18439 (N_18439,N_10773,N_12976);
or U18440 (N_18440,N_11062,N_13750);
nor U18441 (N_18441,N_12970,N_11755);
nand U18442 (N_18442,N_12121,N_13738);
xor U18443 (N_18443,N_10381,N_13762);
nand U18444 (N_18444,N_11850,N_13892);
and U18445 (N_18445,N_14346,N_12474);
nor U18446 (N_18446,N_13400,N_13336);
nor U18447 (N_18447,N_13765,N_14768);
or U18448 (N_18448,N_13742,N_13504);
xnor U18449 (N_18449,N_12162,N_14443);
or U18450 (N_18450,N_12840,N_14320);
nand U18451 (N_18451,N_12700,N_13748);
xor U18452 (N_18452,N_14122,N_12838);
and U18453 (N_18453,N_11446,N_10636);
nor U18454 (N_18454,N_11212,N_14705);
and U18455 (N_18455,N_14814,N_13592);
xnor U18456 (N_18456,N_10698,N_11871);
or U18457 (N_18457,N_12697,N_10382);
xor U18458 (N_18458,N_12402,N_12084);
and U18459 (N_18459,N_12876,N_13477);
and U18460 (N_18460,N_12646,N_14975);
nor U18461 (N_18461,N_14725,N_13963);
xnor U18462 (N_18462,N_10321,N_11740);
xor U18463 (N_18463,N_13044,N_11699);
and U18464 (N_18464,N_11341,N_13857);
nand U18465 (N_18465,N_14931,N_13495);
nor U18466 (N_18466,N_14352,N_11085);
nand U18467 (N_18467,N_11999,N_14515);
and U18468 (N_18468,N_10813,N_13376);
xor U18469 (N_18469,N_14045,N_14145);
nor U18470 (N_18470,N_14388,N_11275);
nor U18471 (N_18471,N_10212,N_14257);
xor U18472 (N_18472,N_10101,N_13953);
and U18473 (N_18473,N_14857,N_11628);
nor U18474 (N_18474,N_14396,N_12062);
nand U18475 (N_18475,N_11853,N_14734);
xor U18476 (N_18476,N_12883,N_14415);
nand U18477 (N_18477,N_10996,N_12723);
nand U18478 (N_18478,N_11804,N_11144);
nand U18479 (N_18479,N_10768,N_10278);
nor U18480 (N_18480,N_12897,N_13778);
xnor U18481 (N_18481,N_10162,N_12417);
and U18482 (N_18482,N_13096,N_14811);
nand U18483 (N_18483,N_12946,N_13051);
or U18484 (N_18484,N_14686,N_11189);
nor U18485 (N_18485,N_10408,N_14356);
and U18486 (N_18486,N_12338,N_11244);
or U18487 (N_18487,N_11777,N_11462);
xor U18488 (N_18488,N_11403,N_11775);
nor U18489 (N_18489,N_11718,N_14152);
nand U18490 (N_18490,N_11548,N_10466);
nor U18491 (N_18491,N_13926,N_13907);
nor U18492 (N_18492,N_14176,N_10540);
xor U18493 (N_18493,N_13772,N_11659);
or U18494 (N_18494,N_14717,N_11085);
and U18495 (N_18495,N_13044,N_14635);
and U18496 (N_18496,N_12048,N_14421);
nor U18497 (N_18497,N_14062,N_12903);
xnor U18498 (N_18498,N_13872,N_10174);
xor U18499 (N_18499,N_11930,N_12988);
xnor U18500 (N_18500,N_13342,N_14487);
nand U18501 (N_18501,N_14781,N_14754);
xnor U18502 (N_18502,N_10108,N_11941);
or U18503 (N_18503,N_11106,N_13799);
nor U18504 (N_18504,N_13190,N_11083);
nor U18505 (N_18505,N_10034,N_12605);
and U18506 (N_18506,N_11623,N_12143);
and U18507 (N_18507,N_11282,N_12908);
or U18508 (N_18508,N_12183,N_14766);
nor U18509 (N_18509,N_14386,N_12500);
or U18510 (N_18510,N_11001,N_11462);
or U18511 (N_18511,N_11227,N_11199);
xnor U18512 (N_18512,N_13504,N_12451);
and U18513 (N_18513,N_12779,N_11302);
or U18514 (N_18514,N_13070,N_12406);
xor U18515 (N_18515,N_11432,N_13488);
or U18516 (N_18516,N_12676,N_11604);
or U18517 (N_18517,N_12972,N_14500);
nand U18518 (N_18518,N_12364,N_12511);
nand U18519 (N_18519,N_12641,N_10446);
and U18520 (N_18520,N_11034,N_14385);
or U18521 (N_18521,N_14719,N_13638);
and U18522 (N_18522,N_11163,N_10442);
xnor U18523 (N_18523,N_13969,N_10468);
or U18524 (N_18524,N_13002,N_11561);
and U18525 (N_18525,N_14086,N_13454);
and U18526 (N_18526,N_14219,N_10954);
xor U18527 (N_18527,N_12769,N_12869);
xnor U18528 (N_18528,N_13692,N_11569);
or U18529 (N_18529,N_13579,N_14985);
nand U18530 (N_18530,N_13492,N_10116);
nand U18531 (N_18531,N_12554,N_11517);
nand U18532 (N_18532,N_11021,N_11367);
xnor U18533 (N_18533,N_10744,N_12122);
xnor U18534 (N_18534,N_12938,N_12444);
nor U18535 (N_18535,N_11995,N_13034);
nor U18536 (N_18536,N_11610,N_14481);
xor U18537 (N_18537,N_10637,N_10287);
or U18538 (N_18538,N_11039,N_12241);
xnor U18539 (N_18539,N_12615,N_10462);
nand U18540 (N_18540,N_14267,N_12444);
nor U18541 (N_18541,N_11583,N_10579);
xor U18542 (N_18542,N_14548,N_13531);
nand U18543 (N_18543,N_10023,N_11136);
or U18544 (N_18544,N_10434,N_12572);
xor U18545 (N_18545,N_10725,N_13291);
nand U18546 (N_18546,N_13701,N_12427);
nor U18547 (N_18547,N_14684,N_11656);
nor U18548 (N_18548,N_13750,N_12264);
nand U18549 (N_18549,N_13229,N_10778);
or U18550 (N_18550,N_12064,N_13151);
xnor U18551 (N_18551,N_10973,N_10355);
and U18552 (N_18552,N_12038,N_10677);
nand U18553 (N_18553,N_10942,N_10715);
nand U18554 (N_18554,N_12454,N_10942);
nor U18555 (N_18555,N_13292,N_13372);
nand U18556 (N_18556,N_14360,N_12489);
and U18557 (N_18557,N_14521,N_11194);
nand U18558 (N_18558,N_14755,N_14979);
nor U18559 (N_18559,N_14533,N_14796);
nand U18560 (N_18560,N_14412,N_14846);
nor U18561 (N_18561,N_13405,N_12661);
nor U18562 (N_18562,N_12224,N_11535);
nand U18563 (N_18563,N_12531,N_11206);
or U18564 (N_18564,N_12026,N_14264);
or U18565 (N_18565,N_11732,N_13758);
and U18566 (N_18566,N_12691,N_13305);
or U18567 (N_18567,N_12392,N_10040);
nand U18568 (N_18568,N_12269,N_11633);
or U18569 (N_18569,N_10051,N_12610);
nor U18570 (N_18570,N_14675,N_11220);
nand U18571 (N_18571,N_12369,N_14095);
nand U18572 (N_18572,N_13264,N_13073);
and U18573 (N_18573,N_12867,N_10067);
xor U18574 (N_18574,N_14829,N_11196);
xnor U18575 (N_18575,N_13295,N_13984);
nand U18576 (N_18576,N_12266,N_11258);
nor U18577 (N_18577,N_14755,N_12663);
or U18578 (N_18578,N_11182,N_10346);
nand U18579 (N_18579,N_13322,N_14628);
nor U18580 (N_18580,N_14691,N_12053);
and U18581 (N_18581,N_13627,N_12185);
nor U18582 (N_18582,N_14068,N_10417);
xnor U18583 (N_18583,N_12258,N_13244);
xor U18584 (N_18584,N_11660,N_14196);
xor U18585 (N_18585,N_11582,N_11161);
xnor U18586 (N_18586,N_10122,N_14565);
xor U18587 (N_18587,N_11471,N_10067);
nor U18588 (N_18588,N_13401,N_13062);
nand U18589 (N_18589,N_14583,N_13575);
nand U18590 (N_18590,N_10462,N_13297);
and U18591 (N_18591,N_14841,N_11708);
and U18592 (N_18592,N_12387,N_14500);
or U18593 (N_18593,N_10817,N_14732);
nand U18594 (N_18594,N_13684,N_12976);
or U18595 (N_18595,N_12581,N_13646);
or U18596 (N_18596,N_12595,N_12203);
xor U18597 (N_18597,N_10204,N_13500);
nor U18598 (N_18598,N_13436,N_10924);
or U18599 (N_18599,N_14384,N_10552);
or U18600 (N_18600,N_12508,N_13584);
and U18601 (N_18601,N_10047,N_10018);
nor U18602 (N_18602,N_10753,N_11014);
xnor U18603 (N_18603,N_12924,N_10720);
xnor U18604 (N_18604,N_13259,N_10149);
xor U18605 (N_18605,N_13326,N_10767);
xnor U18606 (N_18606,N_10192,N_11107);
and U18607 (N_18607,N_12708,N_13292);
nand U18608 (N_18608,N_10251,N_12137);
xor U18609 (N_18609,N_14321,N_14848);
or U18610 (N_18610,N_13361,N_13427);
nor U18611 (N_18611,N_13026,N_13178);
xor U18612 (N_18612,N_13438,N_12057);
nand U18613 (N_18613,N_11184,N_11663);
or U18614 (N_18614,N_10884,N_11946);
and U18615 (N_18615,N_12337,N_13425);
or U18616 (N_18616,N_12360,N_11854);
nor U18617 (N_18617,N_14224,N_10507);
or U18618 (N_18618,N_13842,N_13872);
and U18619 (N_18619,N_11518,N_11752);
or U18620 (N_18620,N_13141,N_11736);
or U18621 (N_18621,N_10488,N_13295);
nand U18622 (N_18622,N_14380,N_10308);
and U18623 (N_18623,N_12196,N_13803);
xor U18624 (N_18624,N_12577,N_14854);
and U18625 (N_18625,N_14061,N_12610);
nand U18626 (N_18626,N_10058,N_11659);
or U18627 (N_18627,N_14531,N_11668);
xnor U18628 (N_18628,N_13302,N_12871);
nor U18629 (N_18629,N_12138,N_10336);
xor U18630 (N_18630,N_11414,N_10543);
nand U18631 (N_18631,N_11190,N_11188);
and U18632 (N_18632,N_10253,N_12746);
and U18633 (N_18633,N_13475,N_10229);
nand U18634 (N_18634,N_14885,N_14712);
or U18635 (N_18635,N_12483,N_10341);
nand U18636 (N_18636,N_11139,N_13016);
or U18637 (N_18637,N_11309,N_10020);
or U18638 (N_18638,N_13437,N_10600);
and U18639 (N_18639,N_11921,N_14075);
and U18640 (N_18640,N_13738,N_14869);
xor U18641 (N_18641,N_10494,N_12213);
or U18642 (N_18642,N_13190,N_10911);
xor U18643 (N_18643,N_12256,N_14899);
or U18644 (N_18644,N_10051,N_13689);
or U18645 (N_18645,N_13658,N_12270);
or U18646 (N_18646,N_14995,N_13256);
and U18647 (N_18647,N_10156,N_10494);
or U18648 (N_18648,N_14478,N_10379);
and U18649 (N_18649,N_11704,N_11159);
and U18650 (N_18650,N_14659,N_14510);
and U18651 (N_18651,N_11474,N_12382);
nor U18652 (N_18652,N_11261,N_13236);
nand U18653 (N_18653,N_13977,N_13349);
and U18654 (N_18654,N_10430,N_13579);
or U18655 (N_18655,N_13309,N_14731);
nand U18656 (N_18656,N_13294,N_11264);
and U18657 (N_18657,N_10320,N_11917);
nor U18658 (N_18658,N_10716,N_14959);
nor U18659 (N_18659,N_14341,N_12033);
nor U18660 (N_18660,N_13842,N_10142);
and U18661 (N_18661,N_12893,N_13620);
nor U18662 (N_18662,N_14922,N_10608);
nor U18663 (N_18663,N_14058,N_14285);
or U18664 (N_18664,N_12170,N_11646);
or U18665 (N_18665,N_12458,N_10687);
or U18666 (N_18666,N_12322,N_12316);
or U18667 (N_18667,N_12219,N_12320);
and U18668 (N_18668,N_14269,N_10986);
or U18669 (N_18669,N_10221,N_13644);
nand U18670 (N_18670,N_11006,N_14093);
and U18671 (N_18671,N_11449,N_11867);
and U18672 (N_18672,N_11816,N_12593);
or U18673 (N_18673,N_12304,N_14453);
nor U18674 (N_18674,N_11399,N_10245);
nor U18675 (N_18675,N_12825,N_13790);
or U18676 (N_18676,N_10592,N_14724);
nor U18677 (N_18677,N_12120,N_10343);
xor U18678 (N_18678,N_14729,N_12077);
xor U18679 (N_18679,N_14856,N_11662);
nand U18680 (N_18680,N_14683,N_14932);
nor U18681 (N_18681,N_12464,N_13261);
nor U18682 (N_18682,N_12405,N_10668);
nor U18683 (N_18683,N_12512,N_11009);
xor U18684 (N_18684,N_12976,N_14109);
and U18685 (N_18685,N_10321,N_12550);
and U18686 (N_18686,N_13066,N_14332);
nor U18687 (N_18687,N_10411,N_10814);
xnor U18688 (N_18688,N_11138,N_12574);
nand U18689 (N_18689,N_10465,N_11924);
or U18690 (N_18690,N_10991,N_11153);
nand U18691 (N_18691,N_10160,N_10830);
or U18692 (N_18692,N_10064,N_11516);
and U18693 (N_18693,N_12543,N_11142);
xnor U18694 (N_18694,N_10950,N_12998);
nor U18695 (N_18695,N_14639,N_12493);
and U18696 (N_18696,N_10388,N_10122);
nor U18697 (N_18697,N_13548,N_14889);
and U18698 (N_18698,N_13968,N_10102);
or U18699 (N_18699,N_10165,N_14654);
or U18700 (N_18700,N_13441,N_11587);
and U18701 (N_18701,N_12805,N_14856);
and U18702 (N_18702,N_10825,N_13572);
nor U18703 (N_18703,N_11629,N_10327);
and U18704 (N_18704,N_13439,N_11283);
nor U18705 (N_18705,N_14314,N_10917);
xnor U18706 (N_18706,N_13628,N_12320);
or U18707 (N_18707,N_10601,N_14833);
or U18708 (N_18708,N_14961,N_14190);
xnor U18709 (N_18709,N_13190,N_11576);
and U18710 (N_18710,N_11614,N_14701);
nor U18711 (N_18711,N_11789,N_11276);
and U18712 (N_18712,N_14369,N_10932);
nor U18713 (N_18713,N_10263,N_12417);
or U18714 (N_18714,N_11372,N_14362);
xor U18715 (N_18715,N_12834,N_14710);
or U18716 (N_18716,N_12656,N_11218);
nand U18717 (N_18717,N_14518,N_11026);
nand U18718 (N_18718,N_10875,N_10170);
or U18719 (N_18719,N_14259,N_13416);
xnor U18720 (N_18720,N_12487,N_10026);
and U18721 (N_18721,N_14713,N_14879);
nand U18722 (N_18722,N_12674,N_10820);
or U18723 (N_18723,N_14851,N_11108);
xnor U18724 (N_18724,N_13324,N_12309);
nor U18725 (N_18725,N_14172,N_10291);
nand U18726 (N_18726,N_10136,N_10532);
nand U18727 (N_18727,N_10345,N_13758);
nand U18728 (N_18728,N_14540,N_14692);
or U18729 (N_18729,N_11176,N_11442);
and U18730 (N_18730,N_10543,N_11527);
nand U18731 (N_18731,N_11916,N_10750);
nor U18732 (N_18732,N_12273,N_12574);
nor U18733 (N_18733,N_13761,N_13310);
or U18734 (N_18734,N_10485,N_12914);
or U18735 (N_18735,N_11378,N_11596);
xor U18736 (N_18736,N_13006,N_10244);
or U18737 (N_18737,N_14383,N_13824);
and U18738 (N_18738,N_11955,N_12898);
xor U18739 (N_18739,N_12176,N_10436);
and U18740 (N_18740,N_13562,N_10153);
or U18741 (N_18741,N_12096,N_12090);
nor U18742 (N_18742,N_10396,N_13069);
nor U18743 (N_18743,N_10689,N_10361);
nor U18744 (N_18744,N_10924,N_12366);
xor U18745 (N_18745,N_12524,N_12845);
or U18746 (N_18746,N_11552,N_14682);
nand U18747 (N_18747,N_10320,N_14071);
nor U18748 (N_18748,N_13331,N_11228);
or U18749 (N_18749,N_13290,N_11412);
or U18750 (N_18750,N_11644,N_10136);
nand U18751 (N_18751,N_13391,N_13461);
nand U18752 (N_18752,N_10730,N_10710);
and U18753 (N_18753,N_14257,N_14957);
and U18754 (N_18754,N_10751,N_13043);
nor U18755 (N_18755,N_12453,N_13856);
xnor U18756 (N_18756,N_13034,N_12409);
or U18757 (N_18757,N_14964,N_10454);
or U18758 (N_18758,N_12662,N_12597);
nor U18759 (N_18759,N_14498,N_11671);
nand U18760 (N_18760,N_13125,N_14842);
nand U18761 (N_18761,N_10354,N_13092);
and U18762 (N_18762,N_10506,N_13607);
nor U18763 (N_18763,N_12411,N_13668);
xor U18764 (N_18764,N_14730,N_14003);
nand U18765 (N_18765,N_14910,N_11788);
xor U18766 (N_18766,N_10440,N_11601);
nor U18767 (N_18767,N_10545,N_12456);
or U18768 (N_18768,N_14716,N_13769);
nand U18769 (N_18769,N_11506,N_11668);
and U18770 (N_18770,N_11469,N_12648);
nor U18771 (N_18771,N_12405,N_13994);
xnor U18772 (N_18772,N_14110,N_13489);
and U18773 (N_18773,N_12809,N_13093);
xnor U18774 (N_18774,N_14702,N_12219);
or U18775 (N_18775,N_10828,N_11991);
nor U18776 (N_18776,N_14764,N_11086);
xor U18777 (N_18777,N_10356,N_13519);
nor U18778 (N_18778,N_12754,N_12894);
and U18779 (N_18779,N_12881,N_11521);
xnor U18780 (N_18780,N_10083,N_13075);
or U18781 (N_18781,N_14009,N_12509);
and U18782 (N_18782,N_11470,N_14739);
or U18783 (N_18783,N_11294,N_11104);
nand U18784 (N_18784,N_11974,N_11219);
nor U18785 (N_18785,N_14998,N_12445);
nor U18786 (N_18786,N_12030,N_12039);
nor U18787 (N_18787,N_14604,N_12817);
xnor U18788 (N_18788,N_12158,N_10254);
or U18789 (N_18789,N_12744,N_12896);
and U18790 (N_18790,N_12370,N_11619);
xnor U18791 (N_18791,N_14467,N_11244);
nand U18792 (N_18792,N_11473,N_11782);
xnor U18793 (N_18793,N_14050,N_13305);
and U18794 (N_18794,N_14182,N_10928);
nor U18795 (N_18795,N_10469,N_11181);
xor U18796 (N_18796,N_11205,N_11813);
nand U18797 (N_18797,N_14995,N_13891);
nor U18798 (N_18798,N_12466,N_14558);
nand U18799 (N_18799,N_13945,N_11867);
or U18800 (N_18800,N_14962,N_13971);
nor U18801 (N_18801,N_13557,N_13730);
or U18802 (N_18802,N_14410,N_12090);
nand U18803 (N_18803,N_13232,N_11822);
and U18804 (N_18804,N_13622,N_13341);
nor U18805 (N_18805,N_12931,N_13657);
nor U18806 (N_18806,N_11440,N_13614);
nor U18807 (N_18807,N_11630,N_11066);
or U18808 (N_18808,N_11673,N_10365);
nor U18809 (N_18809,N_11034,N_11777);
and U18810 (N_18810,N_12166,N_14071);
or U18811 (N_18811,N_14202,N_10224);
nor U18812 (N_18812,N_11013,N_13867);
or U18813 (N_18813,N_13308,N_14590);
nand U18814 (N_18814,N_10469,N_10214);
xor U18815 (N_18815,N_14210,N_14652);
xnor U18816 (N_18816,N_14425,N_11269);
or U18817 (N_18817,N_12610,N_11883);
and U18818 (N_18818,N_10064,N_10872);
xnor U18819 (N_18819,N_12317,N_11222);
nor U18820 (N_18820,N_12945,N_12903);
nor U18821 (N_18821,N_14880,N_10711);
nand U18822 (N_18822,N_12278,N_13450);
and U18823 (N_18823,N_14807,N_12676);
nand U18824 (N_18824,N_12162,N_10465);
xor U18825 (N_18825,N_11519,N_12074);
nand U18826 (N_18826,N_10833,N_14239);
nand U18827 (N_18827,N_14724,N_10378);
or U18828 (N_18828,N_13586,N_12218);
xnor U18829 (N_18829,N_14743,N_14972);
nor U18830 (N_18830,N_13222,N_11660);
xor U18831 (N_18831,N_10671,N_13322);
or U18832 (N_18832,N_13192,N_12916);
nand U18833 (N_18833,N_12497,N_11502);
or U18834 (N_18834,N_14452,N_13216);
or U18835 (N_18835,N_12398,N_12561);
or U18836 (N_18836,N_11919,N_12377);
and U18837 (N_18837,N_13603,N_14121);
nor U18838 (N_18838,N_10366,N_10952);
or U18839 (N_18839,N_14639,N_13925);
and U18840 (N_18840,N_12568,N_14443);
xnor U18841 (N_18841,N_14278,N_14484);
and U18842 (N_18842,N_10066,N_14251);
nand U18843 (N_18843,N_12130,N_11778);
nand U18844 (N_18844,N_11522,N_13793);
and U18845 (N_18845,N_11230,N_12248);
and U18846 (N_18846,N_13525,N_11392);
nand U18847 (N_18847,N_10513,N_11132);
xor U18848 (N_18848,N_11534,N_12339);
and U18849 (N_18849,N_12006,N_13687);
xnor U18850 (N_18850,N_14790,N_10088);
nor U18851 (N_18851,N_10802,N_10295);
nand U18852 (N_18852,N_14401,N_12999);
xnor U18853 (N_18853,N_13282,N_11977);
nor U18854 (N_18854,N_12162,N_14839);
or U18855 (N_18855,N_11452,N_10029);
nor U18856 (N_18856,N_11743,N_13077);
nor U18857 (N_18857,N_10385,N_11101);
and U18858 (N_18858,N_14361,N_11637);
nand U18859 (N_18859,N_12663,N_13562);
or U18860 (N_18860,N_13926,N_14253);
xor U18861 (N_18861,N_12898,N_12814);
nor U18862 (N_18862,N_10810,N_13202);
xnor U18863 (N_18863,N_14887,N_10565);
or U18864 (N_18864,N_12494,N_10398);
nor U18865 (N_18865,N_13806,N_14341);
or U18866 (N_18866,N_10193,N_11846);
nand U18867 (N_18867,N_14268,N_12931);
nand U18868 (N_18868,N_14677,N_12393);
nor U18869 (N_18869,N_12022,N_11310);
and U18870 (N_18870,N_11858,N_14623);
nand U18871 (N_18871,N_10841,N_13793);
xor U18872 (N_18872,N_10281,N_11941);
nand U18873 (N_18873,N_13344,N_13296);
nand U18874 (N_18874,N_12748,N_12726);
xnor U18875 (N_18875,N_14513,N_14823);
and U18876 (N_18876,N_10378,N_10066);
and U18877 (N_18877,N_10330,N_14456);
nand U18878 (N_18878,N_11083,N_12287);
or U18879 (N_18879,N_13295,N_14309);
or U18880 (N_18880,N_14274,N_14156);
and U18881 (N_18881,N_11949,N_11281);
nand U18882 (N_18882,N_13197,N_14623);
nand U18883 (N_18883,N_10625,N_11885);
xor U18884 (N_18884,N_10342,N_14796);
nand U18885 (N_18885,N_13812,N_11698);
or U18886 (N_18886,N_11920,N_10648);
and U18887 (N_18887,N_11868,N_11758);
or U18888 (N_18888,N_12613,N_10696);
nand U18889 (N_18889,N_14636,N_13097);
nor U18890 (N_18890,N_11137,N_13609);
nand U18891 (N_18891,N_11871,N_13562);
and U18892 (N_18892,N_10551,N_12141);
nand U18893 (N_18893,N_13922,N_11821);
nand U18894 (N_18894,N_12334,N_12619);
nor U18895 (N_18895,N_10407,N_14779);
nor U18896 (N_18896,N_10515,N_10317);
or U18897 (N_18897,N_10887,N_10099);
nand U18898 (N_18898,N_11314,N_14865);
nor U18899 (N_18899,N_10943,N_14054);
nor U18900 (N_18900,N_13907,N_10344);
xnor U18901 (N_18901,N_10734,N_14279);
nor U18902 (N_18902,N_14402,N_10491);
xor U18903 (N_18903,N_12234,N_11212);
or U18904 (N_18904,N_11860,N_11074);
xnor U18905 (N_18905,N_12838,N_12834);
xnor U18906 (N_18906,N_11896,N_13679);
or U18907 (N_18907,N_12648,N_11949);
nor U18908 (N_18908,N_13929,N_12993);
nor U18909 (N_18909,N_13783,N_14147);
or U18910 (N_18910,N_10850,N_11146);
and U18911 (N_18911,N_14099,N_12560);
xor U18912 (N_18912,N_14810,N_14405);
nor U18913 (N_18913,N_13360,N_13224);
or U18914 (N_18914,N_14072,N_12985);
nand U18915 (N_18915,N_13651,N_14808);
nor U18916 (N_18916,N_13330,N_14174);
nand U18917 (N_18917,N_10416,N_11825);
xnor U18918 (N_18918,N_11453,N_11054);
xnor U18919 (N_18919,N_12631,N_11341);
nor U18920 (N_18920,N_12537,N_14711);
nand U18921 (N_18921,N_13799,N_11610);
or U18922 (N_18922,N_13012,N_13268);
xnor U18923 (N_18923,N_10840,N_10035);
xor U18924 (N_18924,N_14965,N_11739);
nand U18925 (N_18925,N_12220,N_10951);
nand U18926 (N_18926,N_11808,N_14436);
nand U18927 (N_18927,N_13828,N_11227);
nand U18928 (N_18928,N_14709,N_14583);
and U18929 (N_18929,N_12721,N_12742);
nand U18930 (N_18930,N_10954,N_14170);
xnor U18931 (N_18931,N_12684,N_13433);
or U18932 (N_18932,N_14340,N_12856);
nand U18933 (N_18933,N_12671,N_12814);
xor U18934 (N_18934,N_12360,N_13838);
and U18935 (N_18935,N_12447,N_12352);
nand U18936 (N_18936,N_10615,N_11115);
xnor U18937 (N_18937,N_10771,N_12564);
nor U18938 (N_18938,N_10879,N_13337);
or U18939 (N_18939,N_12687,N_14371);
and U18940 (N_18940,N_12997,N_10123);
xor U18941 (N_18941,N_14219,N_14438);
nor U18942 (N_18942,N_11192,N_10459);
nor U18943 (N_18943,N_13343,N_10739);
and U18944 (N_18944,N_13088,N_10769);
nand U18945 (N_18945,N_13497,N_11869);
nor U18946 (N_18946,N_14618,N_13096);
or U18947 (N_18947,N_12620,N_13666);
and U18948 (N_18948,N_10735,N_14214);
nor U18949 (N_18949,N_13533,N_12599);
or U18950 (N_18950,N_13089,N_13319);
xor U18951 (N_18951,N_11988,N_13140);
or U18952 (N_18952,N_12076,N_10775);
and U18953 (N_18953,N_12119,N_11229);
or U18954 (N_18954,N_10511,N_14770);
nor U18955 (N_18955,N_10672,N_10900);
xnor U18956 (N_18956,N_11468,N_12203);
xor U18957 (N_18957,N_11722,N_12306);
and U18958 (N_18958,N_13273,N_12124);
or U18959 (N_18959,N_10425,N_14812);
or U18960 (N_18960,N_11874,N_11157);
nor U18961 (N_18961,N_12030,N_12395);
and U18962 (N_18962,N_10355,N_14740);
nand U18963 (N_18963,N_13060,N_11877);
xnor U18964 (N_18964,N_11955,N_12032);
xnor U18965 (N_18965,N_13589,N_11768);
or U18966 (N_18966,N_14583,N_10986);
and U18967 (N_18967,N_12184,N_14791);
and U18968 (N_18968,N_10551,N_14468);
or U18969 (N_18969,N_10368,N_13990);
xnor U18970 (N_18970,N_13468,N_12455);
xor U18971 (N_18971,N_12540,N_14185);
xor U18972 (N_18972,N_13515,N_12380);
and U18973 (N_18973,N_11935,N_14882);
and U18974 (N_18974,N_13785,N_14958);
and U18975 (N_18975,N_12483,N_14964);
or U18976 (N_18976,N_13657,N_12634);
and U18977 (N_18977,N_13629,N_12134);
xnor U18978 (N_18978,N_13817,N_12702);
or U18979 (N_18979,N_12874,N_10999);
or U18980 (N_18980,N_14672,N_11534);
or U18981 (N_18981,N_13419,N_13290);
and U18982 (N_18982,N_13151,N_12115);
nor U18983 (N_18983,N_14411,N_13311);
or U18984 (N_18984,N_11539,N_12684);
and U18985 (N_18985,N_12397,N_10809);
nand U18986 (N_18986,N_11650,N_14175);
nor U18987 (N_18987,N_12376,N_10428);
nand U18988 (N_18988,N_13150,N_14703);
xnor U18989 (N_18989,N_13853,N_10186);
nor U18990 (N_18990,N_12374,N_13538);
and U18991 (N_18991,N_10362,N_11437);
nor U18992 (N_18992,N_13626,N_13355);
or U18993 (N_18993,N_11159,N_11441);
xnor U18994 (N_18994,N_11469,N_12240);
nor U18995 (N_18995,N_14315,N_10758);
nand U18996 (N_18996,N_13486,N_10665);
and U18997 (N_18997,N_14776,N_11544);
and U18998 (N_18998,N_11865,N_13030);
xor U18999 (N_18999,N_13649,N_12534);
xor U19000 (N_19000,N_10938,N_13588);
and U19001 (N_19001,N_14157,N_11647);
nor U19002 (N_19002,N_11834,N_14391);
nor U19003 (N_19003,N_12400,N_11030);
nor U19004 (N_19004,N_10217,N_12482);
xor U19005 (N_19005,N_12666,N_13068);
xor U19006 (N_19006,N_12348,N_11768);
nor U19007 (N_19007,N_13626,N_10953);
xor U19008 (N_19008,N_14737,N_12504);
and U19009 (N_19009,N_11399,N_10919);
nor U19010 (N_19010,N_10113,N_10598);
xnor U19011 (N_19011,N_11143,N_10336);
nor U19012 (N_19012,N_11833,N_10432);
and U19013 (N_19013,N_12666,N_11456);
nand U19014 (N_19014,N_13672,N_12565);
nand U19015 (N_19015,N_11672,N_14132);
xnor U19016 (N_19016,N_12564,N_13208);
or U19017 (N_19017,N_12986,N_14604);
and U19018 (N_19018,N_10216,N_13846);
nor U19019 (N_19019,N_11924,N_13085);
or U19020 (N_19020,N_13907,N_10613);
nand U19021 (N_19021,N_11476,N_11498);
xor U19022 (N_19022,N_14072,N_10976);
or U19023 (N_19023,N_13943,N_12213);
nor U19024 (N_19024,N_13064,N_12481);
nand U19025 (N_19025,N_10405,N_14052);
or U19026 (N_19026,N_11228,N_11901);
nor U19027 (N_19027,N_11900,N_11755);
nor U19028 (N_19028,N_14808,N_10700);
and U19029 (N_19029,N_10134,N_12649);
and U19030 (N_19030,N_14510,N_13217);
nor U19031 (N_19031,N_10365,N_14251);
nand U19032 (N_19032,N_10879,N_14533);
nand U19033 (N_19033,N_14774,N_11815);
nand U19034 (N_19034,N_10800,N_13771);
nand U19035 (N_19035,N_12040,N_10135);
xnor U19036 (N_19036,N_13714,N_13819);
nor U19037 (N_19037,N_14766,N_11230);
nand U19038 (N_19038,N_12582,N_10392);
xnor U19039 (N_19039,N_12310,N_13583);
and U19040 (N_19040,N_10426,N_10055);
nand U19041 (N_19041,N_10273,N_13429);
and U19042 (N_19042,N_10639,N_11918);
nor U19043 (N_19043,N_13747,N_12166);
and U19044 (N_19044,N_13845,N_10613);
and U19045 (N_19045,N_10848,N_14930);
nor U19046 (N_19046,N_14190,N_14014);
nand U19047 (N_19047,N_14996,N_11897);
nor U19048 (N_19048,N_12256,N_12473);
and U19049 (N_19049,N_14187,N_12590);
nand U19050 (N_19050,N_13031,N_10630);
xnor U19051 (N_19051,N_12804,N_11766);
nor U19052 (N_19052,N_14986,N_12720);
xor U19053 (N_19053,N_11398,N_12188);
xor U19054 (N_19054,N_14964,N_10839);
or U19055 (N_19055,N_11247,N_10779);
nand U19056 (N_19056,N_14531,N_13660);
and U19057 (N_19057,N_13715,N_10458);
or U19058 (N_19058,N_12447,N_12182);
xor U19059 (N_19059,N_14582,N_13822);
or U19060 (N_19060,N_12702,N_10015);
and U19061 (N_19061,N_10984,N_14211);
nor U19062 (N_19062,N_12437,N_11768);
nand U19063 (N_19063,N_11326,N_10838);
nor U19064 (N_19064,N_13893,N_13283);
nor U19065 (N_19065,N_12478,N_14798);
xor U19066 (N_19066,N_13258,N_14516);
nand U19067 (N_19067,N_11200,N_10553);
and U19068 (N_19068,N_12838,N_10460);
nor U19069 (N_19069,N_13457,N_10702);
nor U19070 (N_19070,N_12299,N_10634);
xnor U19071 (N_19071,N_14658,N_10545);
nor U19072 (N_19072,N_10332,N_14170);
and U19073 (N_19073,N_10359,N_12685);
xor U19074 (N_19074,N_14906,N_11857);
and U19075 (N_19075,N_11347,N_14035);
xor U19076 (N_19076,N_11438,N_12046);
xnor U19077 (N_19077,N_10533,N_11482);
xnor U19078 (N_19078,N_14582,N_14494);
xor U19079 (N_19079,N_10560,N_11154);
nor U19080 (N_19080,N_10531,N_10226);
nand U19081 (N_19081,N_13168,N_11630);
or U19082 (N_19082,N_10007,N_11091);
nand U19083 (N_19083,N_13261,N_14457);
or U19084 (N_19084,N_14423,N_10797);
nand U19085 (N_19085,N_11227,N_10496);
and U19086 (N_19086,N_14770,N_13528);
xor U19087 (N_19087,N_14954,N_10007);
nor U19088 (N_19088,N_12894,N_12186);
nand U19089 (N_19089,N_12987,N_10985);
or U19090 (N_19090,N_14977,N_12479);
and U19091 (N_19091,N_10986,N_10838);
or U19092 (N_19092,N_12800,N_13077);
xnor U19093 (N_19093,N_11478,N_12350);
and U19094 (N_19094,N_10428,N_11539);
nand U19095 (N_19095,N_14907,N_13421);
nor U19096 (N_19096,N_11455,N_13719);
or U19097 (N_19097,N_10650,N_11436);
nor U19098 (N_19098,N_13020,N_11081);
xor U19099 (N_19099,N_12449,N_14289);
xor U19100 (N_19100,N_11992,N_10252);
nor U19101 (N_19101,N_12799,N_13887);
xnor U19102 (N_19102,N_10785,N_12300);
nor U19103 (N_19103,N_10812,N_14477);
or U19104 (N_19104,N_11046,N_13250);
xnor U19105 (N_19105,N_10845,N_13284);
nor U19106 (N_19106,N_11473,N_12918);
nor U19107 (N_19107,N_14537,N_11499);
or U19108 (N_19108,N_12471,N_10788);
nand U19109 (N_19109,N_10510,N_11157);
and U19110 (N_19110,N_10092,N_13560);
nor U19111 (N_19111,N_14793,N_12670);
xnor U19112 (N_19112,N_13851,N_12110);
and U19113 (N_19113,N_13051,N_10783);
or U19114 (N_19114,N_14805,N_12023);
or U19115 (N_19115,N_11913,N_11832);
or U19116 (N_19116,N_10882,N_12370);
or U19117 (N_19117,N_11982,N_11371);
nand U19118 (N_19118,N_13575,N_12595);
or U19119 (N_19119,N_12983,N_12432);
xor U19120 (N_19120,N_10882,N_14180);
or U19121 (N_19121,N_12675,N_12228);
xnor U19122 (N_19122,N_13349,N_12186);
nand U19123 (N_19123,N_10275,N_10887);
nor U19124 (N_19124,N_14580,N_12034);
nor U19125 (N_19125,N_12541,N_11064);
nand U19126 (N_19126,N_10398,N_10877);
nor U19127 (N_19127,N_13728,N_12152);
nand U19128 (N_19128,N_14858,N_10209);
xnor U19129 (N_19129,N_10284,N_13077);
nand U19130 (N_19130,N_13173,N_12315);
and U19131 (N_19131,N_11141,N_10168);
xnor U19132 (N_19132,N_10822,N_13805);
xor U19133 (N_19133,N_12916,N_12374);
xor U19134 (N_19134,N_14589,N_13221);
xor U19135 (N_19135,N_10991,N_14071);
xnor U19136 (N_19136,N_11492,N_14181);
nor U19137 (N_19137,N_14017,N_13089);
nand U19138 (N_19138,N_11621,N_10109);
nor U19139 (N_19139,N_11329,N_10201);
and U19140 (N_19140,N_11988,N_12917);
xnor U19141 (N_19141,N_14357,N_14737);
and U19142 (N_19142,N_12761,N_12941);
and U19143 (N_19143,N_11833,N_12081);
and U19144 (N_19144,N_14748,N_10575);
nand U19145 (N_19145,N_11937,N_10706);
nor U19146 (N_19146,N_10245,N_14350);
nor U19147 (N_19147,N_14630,N_10641);
nor U19148 (N_19148,N_11594,N_13108);
nand U19149 (N_19149,N_13630,N_10945);
nand U19150 (N_19150,N_13717,N_13106);
nor U19151 (N_19151,N_14287,N_11051);
and U19152 (N_19152,N_10916,N_12801);
xor U19153 (N_19153,N_11695,N_12979);
xor U19154 (N_19154,N_12754,N_12779);
nor U19155 (N_19155,N_10693,N_11224);
and U19156 (N_19156,N_12695,N_11426);
nand U19157 (N_19157,N_11013,N_14983);
nand U19158 (N_19158,N_10680,N_13359);
xnor U19159 (N_19159,N_11801,N_11636);
or U19160 (N_19160,N_10602,N_11176);
xor U19161 (N_19161,N_14178,N_10477);
nand U19162 (N_19162,N_11431,N_14120);
and U19163 (N_19163,N_12069,N_12454);
and U19164 (N_19164,N_10118,N_12524);
nor U19165 (N_19165,N_12631,N_13929);
xnor U19166 (N_19166,N_11314,N_10911);
nor U19167 (N_19167,N_11163,N_10453);
nor U19168 (N_19168,N_13208,N_11166);
xnor U19169 (N_19169,N_13110,N_13153);
nor U19170 (N_19170,N_13702,N_13208);
and U19171 (N_19171,N_13755,N_13049);
or U19172 (N_19172,N_13891,N_10553);
and U19173 (N_19173,N_12828,N_14224);
nand U19174 (N_19174,N_12814,N_13585);
and U19175 (N_19175,N_13545,N_12941);
nand U19176 (N_19176,N_12546,N_12074);
or U19177 (N_19177,N_12442,N_13702);
and U19178 (N_19178,N_12276,N_12976);
xnor U19179 (N_19179,N_14143,N_11563);
and U19180 (N_19180,N_13359,N_14309);
and U19181 (N_19181,N_11677,N_13768);
nand U19182 (N_19182,N_11079,N_14274);
xor U19183 (N_19183,N_14934,N_12156);
nand U19184 (N_19184,N_12692,N_11888);
or U19185 (N_19185,N_10440,N_12391);
nor U19186 (N_19186,N_11750,N_11388);
nor U19187 (N_19187,N_11426,N_10960);
nand U19188 (N_19188,N_13458,N_12062);
xnor U19189 (N_19189,N_11058,N_10723);
nor U19190 (N_19190,N_14695,N_13704);
nand U19191 (N_19191,N_14814,N_12193);
nor U19192 (N_19192,N_10632,N_13148);
and U19193 (N_19193,N_11963,N_12973);
xor U19194 (N_19194,N_11638,N_11397);
or U19195 (N_19195,N_12826,N_11667);
nand U19196 (N_19196,N_13025,N_14589);
nor U19197 (N_19197,N_12110,N_13006);
nand U19198 (N_19198,N_12028,N_10027);
nor U19199 (N_19199,N_14889,N_11720);
nor U19200 (N_19200,N_11846,N_13897);
and U19201 (N_19201,N_10793,N_12118);
xnor U19202 (N_19202,N_13900,N_11537);
nor U19203 (N_19203,N_14800,N_10206);
nor U19204 (N_19204,N_13982,N_11075);
xnor U19205 (N_19205,N_13786,N_10849);
and U19206 (N_19206,N_11515,N_11136);
and U19207 (N_19207,N_10405,N_11714);
nor U19208 (N_19208,N_12687,N_14495);
xnor U19209 (N_19209,N_14306,N_10883);
xnor U19210 (N_19210,N_11256,N_10240);
and U19211 (N_19211,N_13025,N_14078);
xor U19212 (N_19212,N_10328,N_10502);
nand U19213 (N_19213,N_12117,N_14827);
nor U19214 (N_19214,N_12853,N_12577);
or U19215 (N_19215,N_14176,N_12261);
nor U19216 (N_19216,N_13517,N_11467);
xnor U19217 (N_19217,N_14270,N_11021);
nor U19218 (N_19218,N_12576,N_11930);
nor U19219 (N_19219,N_13472,N_10407);
xor U19220 (N_19220,N_11345,N_13286);
nor U19221 (N_19221,N_13047,N_13125);
nand U19222 (N_19222,N_12103,N_13551);
or U19223 (N_19223,N_14300,N_12898);
nand U19224 (N_19224,N_13593,N_10057);
nand U19225 (N_19225,N_13394,N_11853);
or U19226 (N_19226,N_10903,N_14082);
or U19227 (N_19227,N_12878,N_12696);
and U19228 (N_19228,N_10589,N_11606);
nand U19229 (N_19229,N_14044,N_10282);
or U19230 (N_19230,N_14488,N_13630);
or U19231 (N_19231,N_10465,N_10086);
or U19232 (N_19232,N_12376,N_13570);
xor U19233 (N_19233,N_11194,N_12271);
xnor U19234 (N_19234,N_10961,N_13839);
nor U19235 (N_19235,N_10116,N_14024);
nor U19236 (N_19236,N_10655,N_14329);
or U19237 (N_19237,N_14884,N_10695);
nand U19238 (N_19238,N_11725,N_14088);
nand U19239 (N_19239,N_10589,N_10169);
nor U19240 (N_19240,N_13065,N_11196);
xor U19241 (N_19241,N_10435,N_12072);
nor U19242 (N_19242,N_10305,N_13658);
nand U19243 (N_19243,N_11814,N_13071);
or U19244 (N_19244,N_11806,N_13947);
and U19245 (N_19245,N_12454,N_11847);
or U19246 (N_19246,N_11223,N_12685);
or U19247 (N_19247,N_10827,N_12821);
nand U19248 (N_19248,N_14758,N_11141);
nand U19249 (N_19249,N_13534,N_11832);
nand U19250 (N_19250,N_10627,N_13388);
or U19251 (N_19251,N_14446,N_13676);
and U19252 (N_19252,N_12324,N_10871);
nand U19253 (N_19253,N_13566,N_10709);
nor U19254 (N_19254,N_13035,N_10946);
or U19255 (N_19255,N_10908,N_11216);
and U19256 (N_19256,N_12246,N_12696);
nor U19257 (N_19257,N_11151,N_13264);
nor U19258 (N_19258,N_12503,N_11166);
and U19259 (N_19259,N_10183,N_13827);
and U19260 (N_19260,N_12738,N_13233);
nor U19261 (N_19261,N_14258,N_12312);
xor U19262 (N_19262,N_13869,N_10470);
nand U19263 (N_19263,N_14828,N_12058);
and U19264 (N_19264,N_14733,N_12379);
and U19265 (N_19265,N_12171,N_13159);
xor U19266 (N_19266,N_12307,N_14405);
or U19267 (N_19267,N_11628,N_13250);
and U19268 (N_19268,N_14517,N_10500);
nand U19269 (N_19269,N_13317,N_14263);
xor U19270 (N_19270,N_11949,N_11304);
and U19271 (N_19271,N_12871,N_10566);
xnor U19272 (N_19272,N_12255,N_10053);
and U19273 (N_19273,N_13141,N_12408);
xor U19274 (N_19274,N_12259,N_14940);
and U19275 (N_19275,N_12785,N_13127);
and U19276 (N_19276,N_12222,N_13386);
and U19277 (N_19277,N_12487,N_13190);
nand U19278 (N_19278,N_11672,N_14601);
or U19279 (N_19279,N_14606,N_11704);
nor U19280 (N_19280,N_14808,N_11518);
xor U19281 (N_19281,N_11778,N_10798);
xnor U19282 (N_19282,N_14725,N_11233);
nand U19283 (N_19283,N_13738,N_10344);
nand U19284 (N_19284,N_10891,N_14908);
nor U19285 (N_19285,N_14308,N_13939);
and U19286 (N_19286,N_10891,N_11633);
or U19287 (N_19287,N_14601,N_12787);
or U19288 (N_19288,N_13367,N_13616);
nor U19289 (N_19289,N_11895,N_10535);
xnor U19290 (N_19290,N_13804,N_12247);
nand U19291 (N_19291,N_12314,N_10375);
nand U19292 (N_19292,N_14014,N_13919);
or U19293 (N_19293,N_12375,N_13949);
nand U19294 (N_19294,N_13227,N_13955);
nor U19295 (N_19295,N_11474,N_13174);
xnor U19296 (N_19296,N_13948,N_14070);
nand U19297 (N_19297,N_11422,N_11185);
or U19298 (N_19298,N_12179,N_10407);
and U19299 (N_19299,N_12682,N_11851);
nand U19300 (N_19300,N_13213,N_12971);
nand U19301 (N_19301,N_11514,N_12319);
and U19302 (N_19302,N_10311,N_13491);
xor U19303 (N_19303,N_14923,N_10534);
or U19304 (N_19304,N_10190,N_14160);
or U19305 (N_19305,N_14020,N_13570);
or U19306 (N_19306,N_13675,N_11844);
nor U19307 (N_19307,N_14343,N_14010);
xor U19308 (N_19308,N_10646,N_14453);
or U19309 (N_19309,N_10218,N_13231);
xor U19310 (N_19310,N_14020,N_11880);
nor U19311 (N_19311,N_12091,N_11070);
and U19312 (N_19312,N_12715,N_13391);
and U19313 (N_19313,N_14104,N_12164);
nor U19314 (N_19314,N_14354,N_11960);
and U19315 (N_19315,N_10242,N_12047);
nor U19316 (N_19316,N_11888,N_10897);
and U19317 (N_19317,N_14967,N_14234);
xor U19318 (N_19318,N_12488,N_11105);
nor U19319 (N_19319,N_14568,N_12540);
and U19320 (N_19320,N_12740,N_13945);
nor U19321 (N_19321,N_12197,N_14540);
nand U19322 (N_19322,N_14766,N_10269);
xor U19323 (N_19323,N_12710,N_11482);
xnor U19324 (N_19324,N_10855,N_10958);
xor U19325 (N_19325,N_14956,N_10553);
nor U19326 (N_19326,N_12192,N_11322);
or U19327 (N_19327,N_11618,N_13996);
and U19328 (N_19328,N_11614,N_12299);
xnor U19329 (N_19329,N_14295,N_10711);
nor U19330 (N_19330,N_12362,N_12035);
nor U19331 (N_19331,N_14429,N_12290);
and U19332 (N_19332,N_13888,N_13496);
nand U19333 (N_19333,N_14129,N_10442);
xnor U19334 (N_19334,N_14942,N_11319);
xnor U19335 (N_19335,N_12473,N_14264);
nand U19336 (N_19336,N_11865,N_14572);
or U19337 (N_19337,N_14316,N_13125);
nor U19338 (N_19338,N_11422,N_12305);
or U19339 (N_19339,N_12735,N_13855);
nor U19340 (N_19340,N_13432,N_13231);
xor U19341 (N_19341,N_14420,N_14645);
nor U19342 (N_19342,N_10726,N_14313);
nor U19343 (N_19343,N_12512,N_14016);
nand U19344 (N_19344,N_11397,N_11396);
and U19345 (N_19345,N_13394,N_10754);
xor U19346 (N_19346,N_14505,N_10624);
nor U19347 (N_19347,N_14176,N_13605);
or U19348 (N_19348,N_12865,N_13381);
nor U19349 (N_19349,N_11928,N_11033);
or U19350 (N_19350,N_10433,N_10930);
xor U19351 (N_19351,N_11117,N_11181);
xnor U19352 (N_19352,N_13191,N_12263);
or U19353 (N_19353,N_10108,N_11998);
and U19354 (N_19354,N_13991,N_11194);
and U19355 (N_19355,N_14224,N_10710);
nand U19356 (N_19356,N_10445,N_10713);
or U19357 (N_19357,N_10012,N_10992);
or U19358 (N_19358,N_10082,N_12205);
and U19359 (N_19359,N_12412,N_13489);
or U19360 (N_19360,N_10139,N_11251);
and U19361 (N_19361,N_11353,N_11314);
xnor U19362 (N_19362,N_12142,N_11317);
or U19363 (N_19363,N_12583,N_14606);
or U19364 (N_19364,N_11392,N_12692);
xnor U19365 (N_19365,N_14358,N_11311);
xnor U19366 (N_19366,N_12461,N_12014);
nor U19367 (N_19367,N_13018,N_13320);
xnor U19368 (N_19368,N_10878,N_11874);
xnor U19369 (N_19369,N_14060,N_11268);
nand U19370 (N_19370,N_10016,N_14900);
or U19371 (N_19371,N_10162,N_13467);
and U19372 (N_19372,N_13772,N_13885);
and U19373 (N_19373,N_11838,N_10951);
nor U19374 (N_19374,N_11729,N_12718);
and U19375 (N_19375,N_11729,N_11387);
and U19376 (N_19376,N_14642,N_13132);
and U19377 (N_19377,N_11944,N_14455);
nor U19378 (N_19378,N_13022,N_13057);
and U19379 (N_19379,N_14165,N_14907);
xnor U19380 (N_19380,N_13837,N_10930);
and U19381 (N_19381,N_13617,N_10573);
nand U19382 (N_19382,N_12269,N_11332);
or U19383 (N_19383,N_14487,N_11333);
or U19384 (N_19384,N_10607,N_10253);
nor U19385 (N_19385,N_13458,N_12315);
nor U19386 (N_19386,N_14370,N_12573);
xnor U19387 (N_19387,N_14269,N_13369);
and U19388 (N_19388,N_12898,N_14671);
and U19389 (N_19389,N_10013,N_10695);
nand U19390 (N_19390,N_10147,N_13141);
xor U19391 (N_19391,N_14743,N_12128);
nor U19392 (N_19392,N_13348,N_13224);
or U19393 (N_19393,N_10558,N_13121);
xnor U19394 (N_19394,N_11827,N_10637);
nand U19395 (N_19395,N_11171,N_10335);
and U19396 (N_19396,N_13545,N_13260);
nand U19397 (N_19397,N_11226,N_10815);
nand U19398 (N_19398,N_14393,N_10859);
or U19399 (N_19399,N_13278,N_12695);
nor U19400 (N_19400,N_14381,N_10073);
nand U19401 (N_19401,N_11860,N_13142);
nor U19402 (N_19402,N_12150,N_12870);
xor U19403 (N_19403,N_14022,N_14220);
xnor U19404 (N_19404,N_12047,N_11861);
nor U19405 (N_19405,N_10883,N_13040);
nor U19406 (N_19406,N_11327,N_13688);
xnor U19407 (N_19407,N_14236,N_14227);
xnor U19408 (N_19408,N_10998,N_11553);
nor U19409 (N_19409,N_14161,N_14033);
nand U19410 (N_19410,N_11908,N_12982);
nand U19411 (N_19411,N_10487,N_10953);
and U19412 (N_19412,N_14154,N_12529);
and U19413 (N_19413,N_11091,N_12041);
nand U19414 (N_19414,N_13186,N_13485);
or U19415 (N_19415,N_14778,N_14702);
nand U19416 (N_19416,N_14627,N_10234);
and U19417 (N_19417,N_14979,N_11771);
xnor U19418 (N_19418,N_14837,N_13779);
and U19419 (N_19419,N_14852,N_11741);
and U19420 (N_19420,N_10908,N_14638);
xor U19421 (N_19421,N_14787,N_10198);
xor U19422 (N_19422,N_13631,N_10131);
xnor U19423 (N_19423,N_10436,N_11274);
nor U19424 (N_19424,N_11888,N_12861);
and U19425 (N_19425,N_11367,N_13299);
xor U19426 (N_19426,N_14012,N_12059);
and U19427 (N_19427,N_10235,N_12499);
nand U19428 (N_19428,N_11361,N_11074);
or U19429 (N_19429,N_10105,N_12932);
and U19430 (N_19430,N_10812,N_14807);
and U19431 (N_19431,N_13183,N_12273);
and U19432 (N_19432,N_13440,N_13357);
nand U19433 (N_19433,N_12379,N_11382);
nor U19434 (N_19434,N_13373,N_12960);
xnor U19435 (N_19435,N_14398,N_11465);
nand U19436 (N_19436,N_13119,N_12880);
nand U19437 (N_19437,N_12527,N_14767);
nor U19438 (N_19438,N_14439,N_12428);
or U19439 (N_19439,N_14184,N_10547);
and U19440 (N_19440,N_14168,N_14039);
or U19441 (N_19441,N_12889,N_12818);
nand U19442 (N_19442,N_10866,N_10076);
nor U19443 (N_19443,N_11932,N_13597);
or U19444 (N_19444,N_10526,N_11055);
or U19445 (N_19445,N_11465,N_14732);
nand U19446 (N_19446,N_12793,N_13524);
nand U19447 (N_19447,N_10217,N_12243);
nand U19448 (N_19448,N_11616,N_10756);
xnor U19449 (N_19449,N_11028,N_14845);
or U19450 (N_19450,N_14944,N_12935);
nor U19451 (N_19451,N_14920,N_10140);
nor U19452 (N_19452,N_10908,N_12833);
nor U19453 (N_19453,N_14668,N_13323);
xnor U19454 (N_19454,N_14947,N_13236);
nor U19455 (N_19455,N_13983,N_14842);
nor U19456 (N_19456,N_10450,N_10532);
nand U19457 (N_19457,N_11811,N_12024);
or U19458 (N_19458,N_14400,N_14982);
nor U19459 (N_19459,N_14567,N_13577);
xor U19460 (N_19460,N_14773,N_12219);
and U19461 (N_19461,N_13851,N_14190);
or U19462 (N_19462,N_12920,N_13723);
and U19463 (N_19463,N_10761,N_12900);
xnor U19464 (N_19464,N_13980,N_14831);
xor U19465 (N_19465,N_10071,N_14557);
xnor U19466 (N_19466,N_12304,N_10218);
or U19467 (N_19467,N_11163,N_12687);
xnor U19468 (N_19468,N_14144,N_13554);
or U19469 (N_19469,N_14847,N_13454);
nand U19470 (N_19470,N_10074,N_11638);
and U19471 (N_19471,N_12634,N_10821);
nor U19472 (N_19472,N_12176,N_14505);
nand U19473 (N_19473,N_14702,N_10394);
nor U19474 (N_19474,N_10491,N_10539);
or U19475 (N_19475,N_14785,N_11972);
or U19476 (N_19476,N_13221,N_14596);
or U19477 (N_19477,N_11665,N_11240);
xor U19478 (N_19478,N_10269,N_12447);
xor U19479 (N_19479,N_14118,N_12449);
nor U19480 (N_19480,N_14765,N_14295);
and U19481 (N_19481,N_14432,N_10540);
nor U19482 (N_19482,N_14255,N_10811);
xnor U19483 (N_19483,N_10357,N_13325);
nand U19484 (N_19484,N_12466,N_10491);
xor U19485 (N_19485,N_10344,N_11941);
and U19486 (N_19486,N_10263,N_11004);
or U19487 (N_19487,N_11610,N_12793);
or U19488 (N_19488,N_12774,N_12053);
xor U19489 (N_19489,N_12886,N_14520);
nor U19490 (N_19490,N_14126,N_13516);
nand U19491 (N_19491,N_11084,N_10448);
and U19492 (N_19492,N_10387,N_13004);
nor U19493 (N_19493,N_10056,N_14180);
nor U19494 (N_19494,N_12211,N_12865);
nor U19495 (N_19495,N_13639,N_13040);
nor U19496 (N_19496,N_12234,N_12188);
nor U19497 (N_19497,N_12221,N_13248);
nor U19498 (N_19498,N_11990,N_13778);
nor U19499 (N_19499,N_10535,N_11287);
nand U19500 (N_19500,N_14028,N_14607);
or U19501 (N_19501,N_13547,N_10749);
nor U19502 (N_19502,N_14604,N_11644);
xnor U19503 (N_19503,N_13140,N_12761);
xor U19504 (N_19504,N_11557,N_10429);
or U19505 (N_19505,N_12099,N_13966);
xor U19506 (N_19506,N_13745,N_14664);
nand U19507 (N_19507,N_12389,N_12938);
and U19508 (N_19508,N_10138,N_12321);
xnor U19509 (N_19509,N_11968,N_11509);
or U19510 (N_19510,N_13214,N_14610);
and U19511 (N_19511,N_14542,N_13145);
or U19512 (N_19512,N_11536,N_11686);
and U19513 (N_19513,N_14887,N_13054);
and U19514 (N_19514,N_14417,N_11682);
or U19515 (N_19515,N_11490,N_13598);
nand U19516 (N_19516,N_14119,N_12689);
and U19517 (N_19517,N_14081,N_14354);
nor U19518 (N_19518,N_14026,N_10583);
nand U19519 (N_19519,N_12071,N_10862);
or U19520 (N_19520,N_11411,N_11591);
xnor U19521 (N_19521,N_12223,N_14328);
xor U19522 (N_19522,N_10685,N_11924);
nor U19523 (N_19523,N_12030,N_10569);
and U19524 (N_19524,N_11878,N_14949);
xnor U19525 (N_19525,N_10277,N_14564);
xor U19526 (N_19526,N_12187,N_10043);
xnor U19527 (N_19527,N_13201,N_11312);
xor U19528 (N_19528,N_10183,N_14514);
or U19529 (N_19529,N_10918,N_10587);
nand U19530 (N_19530,N_13680,N_10016);
xnor U19531 (N_19531,N_12552,N_10625);
or U19532 (N_19532,N_10289,N_12495);
nand U19533 (N_19533,N_11380,N_13210);
and U19534 (N_19534,N_11634,N_13888);
nor U19535 (N_19535,N_12611,N_13779);
nor U19536 (N_19536,N_11000,N_14548);
nor U19537 (N_19537,N_11225,N_14862);
xnor U19538 (N_19538,N_11297,N_13091);
nor U19539 (N_19539,N_13150,N_14619);
xor U19540 (N_19540,N_11666,N_10271);
or U19541 (N_19541,N_12797,N_14167);
nand U19542 (N_19542,N_11261,N_10390);
nor U19543 (N_19543,N_11842,N_11873);
or U19544 (N_19544,N_14887,N_12052);
nand U19545 (N_19545,N_10944,N_12437);
nor U19546 (N_19546,N_11708,N_13442);
nand U19547 (N_19547,N_14763,N_14711);
nor U19548 (N_19548,N_10321,N_12084);
or U19549 (N_19549,N_10504,N_11004);
nor U19550 (N_19550,N_14105,N_11399);
nand U19551 (N_19551,N_14452,N_14148);
nand U19552 (N_19552,N_12398,N_10291);
nor U19553 (N_19553,N_11582,N_14556);
nor U19554 (N_19554,N_14400,N_13293);
nand U19555 (N_19555,N_14307,N_11082);
and U19556 (N_19556,N_13033,N_12334);
nand U19557 (N_19557,N_14886,N_12679);
or U19558 (N_19558,N_12738,N_13589);
or U19559 (N_19559,N_11355,N_13217);
or U19560 (N_19560,N_13727,N_13222);
nand U19561 (N_19561,N_11263,N_12719);
nand U19562 (N_19562,N_10512,N_10627);
xnor U19563 (N_19563,N_14239,N_11655);
or U19564 (N_19564,N_14110,N_12368);
xor U19565 (N_19565,N_13710,N_11166);
xor U19566 (N_19566,N_12393,N_13226);
or U19567 (N_19567,N_12352,N_10953);
nand U19568 (N_19568,N_11428,N_11646);
xnor U19569 (N_19569,N_12739,N_11568);
and U19570 (N_19570,N_14214,N_10471);
and U19571 (N_19571,N_14458,N_12099);
nor U19572 (N_19572,N_10916,N_12394);
xnor U19573 (N_19573,N_13735,N_14628);
nor U19574 (N_19574,N_10834,N_11843);
xor U19575 (N_19575,N_11308,N_14203);
nand U19576 (N_19576,N_10212,N_13927);
or U19577 (N_19577,N_12848,N_10430);
and U19578 (N_19578,N_14764,N_10371);
nor U19579 (N_19579,N_10654,N_10588);
and U19580 (N_19580,N_14720,N_12570);
xnor U19581 (N_19581,N_14003,N_11948);
or U19582 (N_19582,N_11912,N_14067);
or U19583 (N_19583,N_10606,N_12271);
and U19584 (N_19584,N_11554,N_14418);
nor U19585 (N_19585,N_10485,N_11820);
xor U19586 (N_19586,N_14312,N_14033);
nor U19587 (N_19587,N_10454,N_14303);
and U19588 (N_19588,N_14312,N_10115);
and U19589 (N_19589,N_10031,N_13345);
or U19590 (N_19590,N_13699,N_12642);
nor U19591 (N_19591,N_10812,N_14134);
and U19592 (N_19592,N_12677,N_14630);
and U19593 (N_19593,N_13787,N_13730);
nand U19594 (N_19594,N_10387,N_14247);
nor U19595 (N_19595,N_11662,N_11237);
or U19596 (N_19596,N_12845,N_10067);
nand U19597 (N_19597,N_14055,N_11520);
nand U19598 (N_19598,N_10627,N_11263);
xor U19599 (N_19599,N_11520,N_11898);
or U19600 (N_19600,N_13846,N_10659);
xnor U19601 (N_19601,N_13931,N_11810);
nand U19602 (N_19602,N_12591,N_10705);
nor U19603 (N_19603,N_13550,N_13267);
and U19604 (N_19604,N_13698,N_11516);
nand U19605 (N_19605,N_14843,N_13109);
xnor U19606 (N_19606,N_12502,N_10132);
nor U19607 (N_19607,N_14825,N_13321);
or U19608 (N_19608,N_12800,N_11153);
xnor U19609 (N_19609,N_14746,N_13593);
nor U19610 (N_19610,N_12259,N_11846);
and U19611 (N_19611,N_12930,N_12376);
nand U19612 (N_19612,N_10739,N_12513);
nand U19613 (N_19613,N_14245,N_10235);
xnor U19614 (N_19614,N_13942,N_10099);
nand U19615 (N_19615,N_14922,N_11815);
or U19616 (N_19616,N_13663,N_13821);
nor U19617 (N_19617,N_10327,N_11150);
nand U19618 (N_19618,N_13752,N_12097);
or U19619 (N_19619,N_11683,N_13572);
nor U19620 (N_19620,N_12853,N_10644);
nand U19621 (N_19621,N_10544,N_10284);
nand U19622 (N_19622,N_14547,N_10346);
xor U19623 (N_19623,N_12620,N_10088);
or U19624 (N_19624,N_11121,N_10832);
xnor U19625 (N_19625,N_12761,N_13424);
or U19626 (N_19626,N_13093,N_12334);
nand U19627 (N_19627,N_10196,N_14779);
nand U19628 (N_19628,N_12685,N_13931);
and U19629 (N_19629,N_11906,N_10889);
nand U19630 (N_19630,N_14592,N_11508);
or U19631 (N_19631,N_12407,N_12265);
or U19632 (N_19632,N_12094,N_11680);
and U19633 (N_19633,N_12697,N_14852);
or U19634 (N_19634,N_12533,N_11531);
xor U19635 (N_19635,N_13744,N_12264);
nand U19636 (N_19636,N_13679,N_14517);
xor U19637 (N_19637,N_13895,N_14562);
or U19638 (N_19638,N_12851,N_10032);
and U19639 (N_19639,N_10247,N_13954);
xor U19640 (N_19640,N_12761,N_14392);
and U19641 (N_19641,N_11229,N_11822);
xnor U19642 (N_19642,N_14798,N_13792);
nor U19643 (N_19643,N_11458,N_14679);
xnor U19644 (N_19644,N_13991,N_13230);
and U19645 (N_19645,N_13801,N_14851);
or U19646 (N_19646,N_10357,N_13345);
xnor U19647 (N_19647,N_13102,N_14988);
xnor U19648 (N_19648,N_12775,N_13955);
or U19649 (N_19649,N_11763,N_14924);
xor U19650 (N_19650,N_11291,N_12325);
and U19651 (N_19651,N_14611,N_10854);
xnor U19652 (N_19652,N_13404,N_12441);
nand U19653 (N_19653,N_11091,N_11851);
nor U19654 (N_19654,N_12958,N_12903);
nor U19655 (N_19655,N_13122,N_14360);
and U19656 (N_19656,N_10645,N_11186);
nor U19657 (N_19657,N_12450,N_10130);
or U19658 (N_19658,N_14984,N_11128);
nand U19659 (N_19659,N_12728,N_13664);
nor U19660 (N_19660,N_12921,N_10800);
xor U19661 (N_19661,N_11262,N_10488);
nor U19662 (N_19662,N_14522,N_11339);
nand U19663 (N_19663,N_12776,N_13647);
nor U19664 (N_19664,N_14349,N_14305);
xnor U19665 (N_19665,N_10666,N_10043);
nand U19666 (N_19666,N_13873,N_12890);
xnor U19667 (N_19667,N_13167,N_10093);
nor U19668 (N_19668,N_13382,N_10854);
or U19669 (N_19669,N_13496,N_12581);
xor U19670 (N_19670,N_10605,N_10057);
nor U19671 (N_19671,N_13358,N_13198);
xnor U19672 (N_19672,N_14264,N_10728);
nand U19673 (N_19673,N_11631,N_10960);
or U19674 (N_19674,N_13692,N_14011);
xor U19675 (N_19675,N_13655,N_11360);
or U19676 (N_19676,N_11051,N_13480);
and U19677 (N_19677,N_11112,N_10059);
nand U19678 (N_19678,N_12244,N_11484);
or U19679 (N_19679,N_13343,N_12521);
and U19680 (N_19680,N_14397,N_13324);
nor U19681 (N_19681,N_11373,N_13258);
xor U19682 (N_19682,N_13626,N_14062);
nor U19683 (N_19683,N_13798,N_14899);
nand U19684 (N_19684,N_10886,N_14042);
xor U19685 (N_19685,N_14954,N_11900);
or U19686 (N_19686,N_14582,N_13994);
or U19687 (N_19687,N_13194,N_11384);
nand U19688 (N_19688,N_12552,N_10432);
and U19689 (N_19689,N_11486,N_13446);
nor U19690 (N_19690,N_10110,N_14193);
xor U19691 (N_19691,N_13284,N_14888);
and U19692 (N_19692,N_12988,N_10730);
nand U19693 (N_19693,N_10862,N_11702);
nand U19694 (N_19694,N_12557,N_10768);
nor U19695 (N_19695,N_10664,N_10167);
and U19696 (N_19696,N_10619,N_10270);
nand U19697 (N_19697,N_11763,N_13760);
or U19698 (N_19698,N_10699,N_11602);
nor U19699 (N_19699,N_12805,N_13995);
xnor U19700 (N_19700,N_10445,N_12588);
xnor U19701 (N_19701,N_11749,N_10797);
nor U19702 (N_19702,N_10002,N_13144);
or U19703 (N_19703,N_10376,N_14549);
nand U19704 (N_19704,N_13856,N_12812);
or U19705 (N_19705,N_14625,N_12714);
nor U19706 (N_19706,N_11829,N_12017);
nand U19707 (N_19707,N_11432,N_13031);
xnor U19708 (N_19708,N_14873,N_11329);
nor U19709 (N_19709,N_11538,N_14021);
or U19710 (N_19710,N_12420,N_12326);
nand U19711 (N_19711,N_14085,N_13105);
nor U19712 (N_19712,N_13283,N_12290);
and U19713 (N_19713,N_10501,N_13073);
and U19714 (N_19714,N_13447,N_10235);
or U19715 (N_19715,N_12505,N_13303);
and U19716 (N_19716,N_10007,N_14985);
nand U19717 (N_19717,N_10355,N_13007);
xor U19718 (N_19718,N_12389,N_12572);
or U19719 (N_19719,N_14669,N_12311);
nand U19720 (N_19720,N_14384,N_14865);
nor U19721 (N_19721,N_13652,N_10527);
nand U19722 (N_19722,N_13164,N_11742);
or U19723 (N_19723,N_14052,N_10078);
and U19724 (N_19724,N_12545,N_10020);
nand U19725 (N_19725,N_10565,N_10376);
or U19726 (N_19726,N_14305,N_11449);
and U19727 (N_19727,N_11961,N_11947);
xor U19728 (N_19728,N_10942,N_12980);
nor U19729 (N_19729,N_11008,N_13537);
or U19730 (N_19730,N_14902,N_11061);
nand U19731 (N_19731,N_12156,N_13289);
xor U19732 (N_19732,N_12185,N_11681);
nand U19733 (N_19733,N_11648,N_12315);
nand U19734 (N_19734,N_13533,N_14180);
nor U19735 (N_19735,N_10972,N_11051);
xor U19736 (N_19736,N_14046,N_11285);
xnor U19737 (N_19737,N_14206,N_14442);
nor U19738 (N_19738,N_12216,N_12607);
or U19739 (N_19739,N_11089,N_12382);
nand U19740 (N_19740,N_11202,N_14112);
or U19741 (N_19741,N_13684,N_11720);
nand U19742 (N_19742,N_14295,N_13604);
xnor U19743 (N_19743,N_14637,N_11454);
and U19744 (N_19744,N_11490,N_11661);
and U19745 (N_19745,N_14639,N_11140);
xnor U19746 (N_19746,N_11439,N_12550);
xnor U19747 (N_19747,N_14232,N_13541);
xor U19748 (N_19748,N_11944,N_14734);
and U19749 (N_19749,N_14188,N_12990);
and U19750 (N_19750,N_11666,N_12732);
xor U19751 (N_19751,N_13818,N_13679);
nand U19752 (N_19752,N_11771,N_10842);
or U19753 (N_19753,N_14259,N_13468);
nor U19754 (N_19754,N_13221,N_14592);
nor U19755 (N_19755,N_10148,N_10009);
nor U19756 (N_19756,N_11601,N_11563);
nand U19757 (N_19757,N_11208,N_10042);
or U19758 (N_19758,N_10654,N_11235);
or U19759 (N_19759,N_14065,N_11466);
and U19760 (N_19760,N_11469,N_10272);
nand U19761 (N_19761,N_11513,N_10146);
nor U19762 (N_19762,N_13083,N_12857);
nor U19763 (N_19763,N_10155,N_11997);
nor U19764 (N_19764,N_11022,N_11312);
or U19765 (N_19765,N_10920,N_12870);
nor U19766 (N_19766,N_14684,N_11850);
xor U19767 (N_19767,N_10471,N_14500);
and U19768 (N_19768,N_12910,N_12198);
nand U19769 (N_19769,N_12510,N_10998);
nand U19770 (N_19770,N_13459,N_14150);
and U19771 (N_19771,N_10174,N_11126);
or U19772 (N_19772,N_12669,N_10088);
xnor U19773 (N_19773,N_13304,N_13278);
and U19774 (N_19774,N_10071,N_11020);
nor U19775 (N_19775,N_11243,N_13313);
nor U19776 (N_19776,N_11203,N_14196);
xnor U19777 (N_19777,N_10685,N_10182);
or U19778 (N_19778,N_13940,N_12243);
or U19779 (N_19779,N_14093,N_13100);
and U19780 (N_19780,N_12034,N_14227);
xnor U19781 (N_19781,N_10303,N_13140);
or U19782 (N_19782,N_11713,N_13926);
or U19783 (N_19783,N_14079,N_10204);
or U19784 (N_19784,N_12476,N_11879);
nor U19785 (N_19785,N_12618,N_14643);
xnor U19786 (N_19786,N_11854,N_12885);
nand U19787 (N_19787,N_12962,N_13072);
nand U19788 (N_19788,N_10179,N_13514);
and U19789 (N_19789,N_11560,N_10549);
or U19790 (N_19790,N_14313,N_14451);
nor U19791 (N_19791,N_12263,N_12231);
nor U19792 (N_19792,N_11481,N_10446);
or U19793 (N_19793,N_12965,N_13958);
nand U19794 (N_19794,N_10796,N_14562);
and U19795 (N_19795,N_13327,N_13355);
nor U19796 (N_19796,N_11086,N_10911);
or U19797 (N_19797,N_11042,N_10381);
nor U19798 (N_19798,N_13485,N_11044);
or U19799 (N_19799,N_10596,N_12634);
xor U19800 (N_19800,N_14116,N_13368);
nor U19801 (N_19801,N_14020,N_10119);
xor U19802 (N_19802,N_11106,N_10554);
nand U19803 (N_19803,N_13206,N_10120);
xnor U19804 (N_19804,N_13682,N_11755);
or U19805 (N_19805,N_14881,N_11200);
xor U19806 (N_19806,N_11933,N_14204);
nand U19807 (N_19807,N_12979,N_12101);
nor U19808 (N_19808,N_11401,N_14009);
xnor U19809 (N_19809,N_11611,N_14339);
and U19810 (N_19810,N_12293,N_10971);
xor U19811 (N_19811,N_14908,N_14852);
and U19812 (N_19812,N_12909,N_13826);
nand U19813 (N_19813,N_14105,N_12433);
xor U19814 (N_19814,N_12171,N_13729);
and U19815 (N_19815,N_11055,N_13129);
nor U19816 (N_19816,N_11156,N_12272);
or U19817 (N_19817,N_12458,N_13737);
or U19818 (N_19818,N_14699,N_11833);
or U19819 (N_19819,N_11114,N_12470);
nor U19820 (N_19820,N_10004,N_10842);
nand U19821 (N_19821,N_14377,N_13636);
nor U19822 (N_19822,N_11245,N_10445);
and U19823 (N_19823,N_14765,N_14945);
xor U19824 (N_19824,N_12275,N_14568);
xor U19825 (N_19825,N_14924,N_10284);
or U19826 (N_19826,N_14547,N_11834);
xor U19827 (N_19827,N_11761,N_12108);
xor U19828 (N_19828,N_12786,N_11432);
and U19829 (N_19829,N_12300,N_13806);
nand U19830 (N_19830,N_11094,N_11816);
nand U19831 (N_19831,N_12431,N_12690);
nor U19832 (N_19832,N_14482,N_13995);
xor U19833 (N_19833,N_12838,N_10999);
nor U19834 (N_19834,N_12908,N_14187);
nand U19835 (N_19835,N_12324,N_10156);
xor U19836 (N_19836,N_12456,N_10910);
or U19837 (N_19837,N_13081,N_12789);
and U19838 (N_19838,N_13765,N_10855);
and U19839 (N_19839,N_12074,N_10306);
nor U19840 (N_19840,N_14024,N_14113);
nand U19841 (N_19841,N_13636,N_12489);
and U19842 (N_19842,N_13826,N_13616);
or U19843 (N_19843,N_10244,N_13604);
xor U19844 (N_19844,N_12801,N_14871);
xor U19845 (N_19845,N_10568,N_14637);
nand U19846 (N_19846,N_10634,N_10425);
nor U19847 (N_19847,N_13094,N_12690);
or U19848 (N_19848,N_11853,N_13157);
nand U19849 (N_19849,N_10531,N_14094);
or U19850 (N_19850,N_13090,N_11928);
and U19851 (N_19851,N_11133,N_13394);
nor U19852 (N_19852,N_13209,N_13216);
xnor U19853 (N_19853,N_11110,N_10729);
xor U19854 (N_19854,N_12702,N_10215);
or U19855 (N_19855,N_12329,N_12237);
and U19856 (N_19856,N_14473,N_11164);
and U19857 (N_19857,N_10316,N_12693);
nand U19858 (N_19858,N_10960,N_13012);
or U19859 (N_19859,N_12813,N_14773);
nand U19860 (N_19860,N_11774,N_14522);
nor U19861 (N_19861,N_12332,N_10689);
or U19862 (N_19862,N_10737,N_14059);
and U19863 (N_19863,N_14842,N_10280);
nor U19864 (N_19864,N_13394,N_13269);
or U19865 (N_19865,N_14170,N_11344);
or U19866 (N_19866,N_14072,N_10625);
xnor U19867 (N_19867,N_11619,N_11539);
and U19868 (N_19868,N_12074,N_10570);
nor U19869 (N_19869,N_12924,N_10994);
nand U19870 (N_19870,N_14792,N_14448);
nand U19871 (N_19871,N_11854,N_14422);
and U19872 (N_19872,N_11165,N_14564);
and U19873 (N_19873,N_13204,N_12409);
nand U19874 (N_19874,N_11517,N_13463);
and U19875 (N_19875,N_11280,N_14854);
nand U19876 (N_19876,N_10374,N_11326);
xor U19877 (N_19877,N_13714,N_13352);
or U19878 (N_19878,N_13292,N_13756);
and U19879 (N_19879,N_13831,N_13973);
or U19880 (N_19880,N_14679,N_13740);
nor U19881 (N_19881,N_14302,N_11488);
and U19882 (N_19882,N_14110,N_11269);
nand U19883 (N_19883,N_11512,N_12816);
and U19884 (N_19884,N_12113,N_12171);
nand U19885 (N_19885,N_13095,N_11792);
nor U19886 (N_19886,N_13787,N_14934);
or U19887 (N_19887,N_13082,N_11956);
nand U19888 (N_19888,N_12564,N_11388);
nor U19889 (N_19889,N_10030,N_14338);
nor U19890 (N_19890,N_14859,N_14810);
nand U19891 (N_19891,N_12702,N_14281);
or U19892 (N_19892,N_12145,N_11445);
nand U19893 (N_19893,N_11949,N_13749);
or U19894 (N_19894,N_13628,N_11264);
nand U19895 (N_19895,N_13032,N_10756);
and U19896 (N_19896,N_11815,N_11342);
xor U19897 (N_19897,N_13410,N_10510);
nand U19898 (N_19898,N_14408,N_13653);
nand U19899 (N_19899,N_14328,N_12064);
xor U19900 (N_19900,N_10935,N_11171);
nor U19901 (N_19901,N_13170,N_12275);
or U19902 (N_19902,N_12628,N_12035);
xor U19903 (N_19903,N_14576,N_14084);
nor U19904 (N_19904,N_10438,N_11956);
nor U19905 (N_19905,N_10782,N_12192);
xor U19906 (N_19906,N_13934,N_12722);
or U19907 (N_19907,N_12613,N_14288);
xnor U19908 (N_19908,N_14533,N_10267);
nor U19909 (N_19909,N_10039,N_11749);
or U19910 (N_19910,N_14546,N_11942);
nand U19911 (N_19911,N_14801,N_10796);
or U19912 (N_19912,N_12554,N_14498);
nor U19913 (N_19913,N_12389,N_11852);
xor U19914 (N_19914,N_12976,N_14396);
or U19915 (N_19915,N_14948,N_11717);
nor U19916 (N_19916,N_10806,N_11512);
and U19917 (N_19917,N_14746,N_11136);
and U19918 (N_19918,N_13768,N_13356);
and U19919 (N_19919,N_10210,N_10777);
xor U19920 (N_19920,N_13177,N_11101);
xnor U19921 (N_19921,N_14009,N_13512);
nor U19922 (N_19922,N_13544,N_13421);
xor U19923 (N_19923,N_10206,N_11335);
or U19924 (N_19924,N_10813,N_13531);
nand U19925 (N_19925,N_12683,N_11148);
and U19926 (N_19926,N_10165,N_11476);
and U19927 (N_19927,N_14842,N_11674);
and U19928 (N_19928,N_14714,N_11430);
or U19929 (N_19929,N_14163,N_14913);
and U19930 (N_19930,N_11107,N_13944);
xor U19931 (N_19931,N_11225,N_13253);
nand U19932 (N_19932,N_11292,N_13980);
and U19933 (N_19933,N_12701,N_10216);
nor U19934 (N_19934,N_14946,N_10165);
or U19935 (N_19935,N_13349,N_10919);
or U19936 (N_19936,N_10271,N_10403);
xnor U19937 (N_19937,N_12689,N_13925);
xnor U19938 (N_19938,N_11464,N_13265);
nand U19939 (N_19939,N_12204,N_12057);
and U19940 (N_19940,N_13311,N_14313);
or U19941 (N_19941,N_14302,N_10433);
or U19942 (N_19942,N_10686,N_14322);
nand U19943 (N_19943,N_14902,N_12027);
nand U19944 (N_19944,N_12240,N_14607);
nor U19945 (N_19945,N_10316,N_12015);
and U19946 (N_19946,N_10293,N_13602);
xnor U19947 (N_19947,N_13548,N_13263);
nand U19948 (N_19948,N_12717,N_13850);
or U19949 (N_19949,N_11720,N_12425);
or U19950 (N_19950,N_14405,N_13909);
and U19951 (N_19951,N_14709,N_12226);
nor U19952 (N_19952,N_14959,N_11676);
nor U19953 (N_19953,N_13831,N_14148);
nand U19954 (N_19954,N_11207,N_13754);
xnor U19955 (N_19955,N_13209,N_13125);
or U19956 (N_19956,N_13840,N_12695);
and U19957 (N_19957,N_14757,N_11114);
xnor U19958 (N_19958,N_11124,N_12501);
and U19959 (N_19959,N_13894,N_12909);
nand U19960 (N_19960,N_12957,N_12305);
xnor U19961 (N_19961,N_10359,N_13778);
nor U19962 (N_19962,N_10181,N_12109);
and U19963 (N_19963,N_14012,N_10314);
xor U19964 (N_19964,N_14110,N_13927);
xor U19965 (N_19965,N_10365,N_14105);
nand U19966 (N_19966,N_14665,N_12188);
xor U19967 (N_19967,N_13413,N_13623);
nor U19968 (N_19968,N_14876,N_12617);
and U19969 (N_19969,N_10755,N_12891);
nand U19970 (N_19970,N_12261,N_11038);
and U19971 (N_19971,N_11347,N_12400);
nand U19972 (N_19972,N_10421,N_11331);
nand U19973 (N_19973,N_13112,N_10026);
or U19974 (N_19974,N_12437,N_10859);
nor U19975 (N_19975,N_10970,N_12084);
xnor U19976 (N_19976,N_14865,N_13564);
xnor U19977 (N_19977,N_12420,N_13583);
and U19978 (N_19978,N_14187,N_10131);
and U19979 (N_19979,N_11942,N_13411);
xor U19980 (N_19980,N_13207,N_13645);
or U19981 (N_19981,N_12893,N_12527);
or U19982 (N_19982,N_10487,N_11877);
nand U19983 (N_19983,N_11346,N_13911);
or U19984 (N_19984,N_11510,N_11263);
or U19985 (N_19985,N_14442,N_12416);
and U19986 (N_19986,N_11009,N_10244);
xnor U19987 (N_19987,N_14577,N_11499);
and U19988 (N_19988,N_12097,N_12270);
xnor U19989 (N_19989,N_10899,N_10443);
xor U19990 (N_19990,N_12074,N_12847);
nand U19991 (N_19991,N_13193,N_14493);
nand U19992 (N_19992,N_11498,N_14012);
or U19993 (N_19993,N_13180,N_13273);
or U19994 (N_19994,N_10966,N_10291);
nand U19995 (N_19995,N_10658,N_14596);
xor U19996 (N_19996,N_13155,N_14619);
and U19997 (N_19997,N_12212,N_14836);
xnor U19998 (N_19998,N_10992,N_12039);
nor U19999 (N_19999,N_12143,N_11740);
nand U20000 (N_20000,N_16720,N_18105);
xor U20001 (N_20001,N_17229,N_15648);
nand U20002 (N_20002,N_19106,N_16467);
and U20003 (N_20003,N_15924,N_19495);
nor U20004 (N_20004,N_16649,N_16672);
or U20005 (N_20005,N_19821,N_15259);
and U20006 (N_20006,N_16851,N_17697);
or U20007 (N_20007,N_17676,N_18098);
nor U20008 (N_20008,N_16784,N_16984);
or U20009 (N_20009,N_15512,N_18380);
xnor U20010 (N_20010,N_15515,N_16268);
or U20011 (N_20011,N_16075,N_18495);
nand U20012 (N_20012,N_16226,N_17209);
nand U20013 (N_20013,N_19746,N_16455);
nor U20014 (N_20014,N_19778,N_16880);
and U20015 (N_20015,N_17200,N_16449);
nand U20016 (N_20016,N_16735,N_17234);
nand U20017 (N_20017,N_16648,N_17900);
nor U20018 (N_20018,N_15246,N_15170);
xnor U20019 (N_20019,N_19665,N_15151);
or U20020 (N_20020,N_19058,N_16955);
nor U20021 (N_20021,N_16386,N_16956);
xor U20022 (N_20022,N_19517,N_19274);
nand U20023 (N_20023,N_19296,N_18843);
and U20024 (N_20024,N_19994,N_15289);
and U20025 (N_20025,N_18154,N_18860);
nand U20026 (N_20026,N_18075,N_19595);
or U20027 (N_20027,N_18285,N_17553);
xor U20028 (N_20028,N_15478,N_19742);
xor U20029 (N_20029,N_18073,N_17595);
xor U20030 (N_20030,N_16829,N_19151);
and U20031 (N_20031,N_15461,N_19945);
xor U20032 (N_20032,N_16764,N_19620);
and U20033 (N_20033,N_18251,N_18517);
xor U20034 (N_20034,N_17404,N_16964);
or U20035 (N_20035,N_19524,N_17581);
or U20036 (N_20036,N_15665,N_16323);
and U20037 (N_20037,N_18120,N_17632);
nand U20038 (N_20038,N_18097,N_19811);
nor U20039 (N_20039,N_17945,N_19010);
xnor U20040 (N_20040,N_18276,N_17348);
nand U20041 (N_20041,N_19139,N_17092);
or U20042 (N_20042,N_15396,N_19919);
nor U20043 (N_20043,N_15467,N_18686);
nor U20044 (N_20044,N_19732,N_19067);
xor U20045 (N_20045,N_18823,N_19861);
or U20046 (N_20046,N_16145,N_19553);
and U20047 (N_20047,N_16980,N_18630);
xnor U20048 (N_20048,N_17197,N_18773);
and U20049 (N_20049,N_18347,N_16523);
and U20050 (N_20050,N_17809,N_19483);
nor U20051 (N_20051,N_19364,N_18513);
or U20052 (N_20052,N_18752,N_16532);
or U20053 (N_20053,N_15118,N_15325);
nor U20054 (N_20054,N_19030,N_17417);
xnor U20055 (N_20055,N_15321,N_16883);
nand U20056 (N_20056,N_16103,N_19249);
nor U20057 (N_20057,N_18050,N_16727);
and U20058 (N_20058,N_19458,N_18086);
or U20059 (N_20059,N_16387,N_18137);
xnor U20060 (N_20060,N_15197,N_15141);
xor U20061 (N_20061,N_16834,N_15200);
and U20062 (N_20062,N_19178,N_19282);
and U20063 (N_20063,N_17052,N_17452);
nand U20064 (N_20064,N_18564,N_17338);
xor U20065 (N_20065,N_17969,N_17248);
xor U20066 (N_20066,N_16379,N_17614);
nor U20067 (N_20067,N_19651,N_15481);
and U20068 (N_20068,N_19488,N_18508);
xnor U20069 (N_20069,N_15416,N_16334);
nand U20070 (N_20070,N_17874,N_17635);
nand U20071 (N_20071,N_15212,N_19774);
nor U20072 (N_20072,N_18440,N_17571);
and U20073 (N_20073,N_18943,N_19117);
nand U20074 (N_20074,N_18775,N_15057);
nor U20075 (N_20075,N_19963,N_16412);
nand U20076 (N_20076,N_16465,N_19463);
nor U20077 (N_20077,N_18881,N_18963);
nor U20078 (N_20078,N_19528,N_15641);
nand U20079 (N_20079,N_19535,N_19461);
or U20080 (N_20080,N_19242,N_19940);
nand U20081 (N_20081,N_17165,N_16017);
nand U20082 (N_20082,N_18465,N_15875);
and U20083 (N_20083,N_16314,N_15109);
or U20084 (N_20084,N_15821,N_18806);
and U20085 (N_20085,N_17817,N_16256);
nor U20086 (N_20086,N_15620,N_15016);
xnor U20087 (N_20087,N_16651,N_16916);
nor U20088 (N_20088,N_16786,N_19158);
nand U20089 (N_20089,N_16442,N_15868);
and U20090 (N_20090,N_15097,N_19478);
xor U20091 (N_20091,N_15703,N_19453);
and U20092 (N_20092,N_16495,N_15638);
and U20093 (N_20093,N_19239,N_18287);
and U20094 (N_20094,N_16933,N_18448);
xnor U20095 (N_20095,N_17266,N_15407);
nor U20096 (N_20096,N_19074,N_16437);
xnor U20097 (N_20097,N_19812,N_16349);
nor U20098 (N_20098,N_19878,N_17527);
xor U20099 (N_20099,N_19934,N_15856);
or U20100 (N_20100,N_18520,N_19137);
nor U20101 (N_20101,N_19638,N_19307);
xnor U20102 (N_20102,N_17685,N_15587);
xnor U20103 (N_20103,N_16677,N_17956);
and U20104 (N_20104,N_17115,N_17392);
nand U20105 (N_20105,N_17419,N_19897);
or U20106 (N_20106,N_19924,N_19741);
nand U20107 (N_20107,N_16042,N_15981);
nand U20108 (N_20108,N_18556,N_17739);
and U20109 (N_20109,N_16634,N_15230);
nor U20110 (N_20110,N_17469,N_17625);
nand U20111 (N_20111,N_18559,N_18900);
nor U20112 (N_20112,N_16587,N_17296);
and U20113 (N_20113,N_15299,N_16190);
nor U20114 (N_20114,N_19283,N_15253);
xnor U20115 (N_20115,N_15140,N_17299);
xnor U20116 (N_20116,N_19673,N_15082);
or U20117 (N_20117,N_15329,N_17645);
nor U20118 (N_20118,N_16547,N_19246);
xor U20119 (N_20119,N_16741,N_16111);
xor U20120 (N_20120,N_17374,N_18712);
or U20121 (N_20121,N_19554,N_18210);
and U20122 (N_20122,N_15031,N_17465);
xnor U20123 (N_20123,N_15672,N_16207);
nor U20124 (N_20124,N_17378,N_19747);
or U20125 (N_20125,N_18064,N_17649);
and U20126 (N_20126,N_19346,N_19698);
and U20127 (N_20127,N_17481,N_16596);
and U20128 (N_20128,N_15208,N_17307);
nand U20129 (N_20129,N_15406,N_18572);
nor U20130 (N_20130,N_16492,N_19988);
nand U20131 (N_20131,N_19550,N_18614);
nor U20132 (N_20132,N_15549,N_18703);
or U20133 (N_20133,N_19072,N_16557);
or U20134 (N_20134,N_18986,N_16912);
nand U20135 (N_20135,N_16223,N_18979);
or U20136 (N_20136,N_16678,N_17932);
nand U20137 (N_20137,N_16011,N_15881);
or U20138 (N_20138,N_16030,N_19708);
or U20139 (N_20139,N_19704,N_16280);
nor U20140 (N_20140,N_17004,N_18011);
nor U20141 (N_20141,N_16036,N_16163);
xnor U20142 (N_20142,N_18461,N_15844);
nor U20143 (N_20143,N_18557,N_15182);
and U20144 (N_20144,N_16925,N_19331);
or U20145 (N_20145,N_18263,N_18000);
and U20146 (N_20146,N_15931,N_17716);
or U20147 (N_20147,N_19906,N_15571);
xnor U20148 (N_20148,N_17198,N_17023);
nor U20149 (N_20149,N_18204,N_19567);
xor U20150 (N_20150,N_16884,N_17498);
xnor U20151 (N_20151,N_19252,N_19454);
or U20152 (N_20152,N_18407,N_15829);
nand U20153 (N_20153,N_16553,N_17416);
nor U20154 (N_20154,N_18340,N_19599);
or U20155 (N_20155,N_16019,N_19764);
xor U20156 (N_20156,N_18230,N_17997);
xor U20157 (N_20157,N_17844,N_16087);
nor U20158 (N_20158,N_16270,N_19925);
or U20159 (N_20159,N_18087,N_18476);
and U20160 (N_20160,N_15945,N_15417);
or U20161 (N_20161,N_15566,N_16689);
or U20162 (N_20162,N_17896,N_16541);
nor U20163 (N_20163,N_18953,N_17841);
nand U20164 (N_20164,N_19352,N_16643);
nand U20165 (N_20165,N_15846,N_16679);
nand U20166 (N_20166,N_17174,N_19536);
nand U20167 (N_20167,N_18092,N_19088);
nor U20168 (N_20168,N_19890,N_17184);
xnor U20169 (N_20169,N_16767,N_15813);
and U20170 (N_20170,N_16718,N_16468);
nor U20171 (N_20171,N_19179,N_17497);
or U20172 (N_20172,N_18727,N_17077);
nor U20173 (N_20173,N_15483,N_18084);
or U20174 (N_20174,N_16257,N_19722);
xor U20175 (N_20175,N_17759,N_16125);
or U20176 (N_20176,N_15893,N_15780);
nor U20177 (N_20177,N_18725,N_18139);
nor U20178 (N_20178,N_16774,N_15536);
nand U20179 (N_20179,N_16792,N_16115);
or U20180 (N_20180,N_15840,N_19970);
nand U20181 (N_20181,N_19689,N_17974);
or U20182 (N_20182,N_16262,N_16065);
or U20183 (N_20183,N_18027,N_18936);
nor U20184 (N_20184,N_16475,N_15500);
and U20185 (N_20185,N_19586,N_15775);
nand U20186 (N_20186,N_17070,N_19926);
or U20187 (N_20187,N_15317,N_18008);
or U20188 (N_20188,N_17479,N_18776);
and U20189 (N_20189,N_16133,N_18372);
nand U20190 (N_20190,N_16488,N_18149);
nand U20191 (N_20191,N_17923,N_19201);
or U20192 (N_20192,N_15534,N_15801);
or U20193 (N_20193,N_16135,N_16534);
nor U20194 (N_20194,N_15996,N_16084);
and U20195 (N_20195,N_19777,N_17935);
and U20196 (N_20196,N_17083,N_19204);
nand U20197 (N_20197,N_17866,N_18598);
nor U20198 (N_20198,N_16775,N_16242);
xnor U20199 (N_20199,N_16358,N_17142);
xnor U20200 (N_20200,N_18275,N_18700);
or U20201 (N_20201,N_15726,N_19218);
or U20202 (N_20202,N_19455,N_15282);
xor U20203 (N_20203,N_18709,N_15514);
nand U20204 (N_20204,N_15697,N_15979);
and U20205 (N_20205,N_18262,N_16776);
or U20206 (N_20206,N_19782,N_15838);
or U20207 (N_20207,N_19266,N_16005);
or U20208 (N_20208,N_17563,N_16580);
and U20209 (N_20209,N_16150,N_16188);
nand U20210 (N_20210,N_16875,N_16791);
nand U20211 (N_20211,N_15916,N_18470);
nor U20212 (N_20212,N_18715,N_17233);
xnor U20213 (N_20213,N_18152,N_18730);
nand U20214 (N_20214,N_17987,N_18278);
nand U20215 (N_20215,N_17045,N_19448);
xnor U20216 (N_20216,N_19789,N_15210);
xor U20217 (N_20217,N_18056,N_15088);
or U20218 (N_20218,N_17977,N_15696);
xnor U20219 (N_20219,N_16430,N_16804);
xor U20220 (N_20220,N_17770,N_17407);
or U20221 (N_20221,N_19631,N_16470);
xor U20222 (N_20222,N_16441,N_17836);
nand U20223 (N_20223,N_17855,N_19557);
nor U20224 (N_20224,N_19836,N_19501);
or U20225 (N_20225,N_19691,N_17801);
and U20226 (N_20226,N_15387,N_16800);
nand U20227 (N_20227,N_18885,N_19976);
xor U20228 (N_20228,N_18910,N_17017);
nor U20229 (N_20229,N_16899,N_18761);
nor U20230 (N_20230,N_15800,N_15578);
xnor U20231 (N_20231,N_15626,N_17838);
nor U20232 (N_20232,N_18221,N_15508);
nor U20233 (N_20233,N_17710,N_16151);
nand U20234 (N_20234,N_16514,N_19587);
nor U20235 (N_20235,N_16865,N_19412);
xor U20236 (N_20236,N_15589,N_19422);
nor U20237 (N_20237,N_15181,N_17193);
and U20238 (N_20238,N_17424,N_18672);
nand U20239 (N_20239,N_19061,N_17210);
and U20240 (N_20240,N_19669,N_19735);
nand U20241 (N_20241,N_17704,N_19039);
xnor U20242 (N_20242,N_15306,N_18496);
nand U20243 (N_20243,N_15449,N_16566);
nand U20244 (N_20244,N_16723,N_16813);
and U20245 (N_20245,N_15788,N_16069);
nor U20246 (N_20246,N_15643,N_17068);
nand U20247 (N_20247,N_17090,N_18122);
nand U20248 (N_20248,N_16225,N_18988);
xnor U20249 (N_20249,N_17274,N_17080);
nand U20250 (N_20250,N_17166,N_15733);
and U20251 (N_20251,N_15437,N_17689);
nand U20252 (N_20252,N_19687,N_15843);
nor U20253 (N_20253,N_17871,N_15388);
xor U20254 (N_20254,N_19080,N_17908);
xnor U20255 (N_20255,N_15802,N_15487);
and U20256 (N_20256,N_19024,N_19995);
nor U20257 (N_20257,N_15929,N_15137);
or U20258 (N_20258,N_17413,N_15267);
or U20259 (N_20259,N_15691,N_17062);
nor U20260 (N_20260,N_17602,N_18466);
xnor U20261 (N_20261,N_17321,N_15466);
and U20262 (N_20262,N_17095,N_19614);
nand U20263 (N_20263,N_16335,N_19357);
nand U20264 (N_20264,N_19748,N_18786);
or U20265 (N_20265,N_19949,N_18311);
xnor U20266 (N_20266,N_18897,N_16604);
and U20267 (N_20267,N_15926,N_16760);
xor U20268 (N_20268,N_18892,N_19593);
nand U20269 (N_20269,N_17385,N_15166);
and U20270 (N_20270,N_19472,N_15271);
or U20271 (N_20271,N_19028,N_15921);
nor U20272 (N_20272,N_15614,N_15211);
and U20273 (N_20273,N_18198,N_15535);
and U20274 (N_20274,N_16288,N_18416);
nand U20275 (N_20275,N_17798,N_18101);
nand U20276 (N_20276,N_17214,N_17010);
nand U20277 (N_20277,N_17201,N_16212);
nand U20278 (N_20278,N_17705,N_15784);
xor U20279 (N_20279,N_18216,N_16932);
and U20280 (N_20280,N_18303,N_19892);
and U20281 (N_20281,N_19378,N_18151);
or U20282 (N_20282,N_17258,N_19788);
nor U20283 (N_20283,N_17679,N_18615);
xnor U20284 (N_20284,N_19180,N_18049);
nor U20285 (N_20285,N_19914,N_17403);
xor U20286 (N_20286,N_19308,N_16239);
nand U20287 (N_20287,N_15824,N_19409);
xnor U20288 (N_20288,N_15600,N_17402);
xor U20289 (N_20289,N_18121,N_15982);
nor U20290 (N_20290,N_19414,N_19690);
xor U20291 (N_20291,N_18296,N_19016);
nand U20292 (N_20292,N_16204,N_16165);
or U20293 (N_20293,N_19645,N_18434);
and U20294 (N_20294,N_17101,N_19092);
or U20295 (N_20295,N_18225,N_15865);
nand U20296 (N_20296,N_15489,N_16330);
nand U20297 (N_20297,N_18778,N_18159);
nand U20298 (N_20298,N_15002,N_15090);
xnor U20299 (N_20299,N_15073,N_18035);
nand U20300 (N_20300,N_15000,N_19834);
and U20301 (N_20301,N_18270,N_16699);
or U20302 (N_20302,N_16007,N_18504);
xor U20303 (N_20303,N_16729,N_18501);
or U20304 (N_20304,N_19041,N_16370);
and U20305 (N_20305,N_15202,N_15007);
nand U20306 (N_20306,N_15792,N_17509);
and U20307 (N_20307,N_17930,N_17192);
nor U20308 (N_20308,N_18985,N_17875);
nor U20309 (N_20309,N_15443,N_18037);
xnor U20310 (N_20310,N_16321,N_17160);
nand U20311 (N_20311,N_19600,N_15193);
or U20312 (N_20312,N_15542,N_18991);
and U20313 (N_20313,N_17121,N_18315);
nand U20314 (N_20314,N_16605,N_18660);
nor U20315 (N_20315,N_17910,N_15080);
xor U20316 (N_20316,N_15906,N_15532);
and U20317 (N_20317,N_17957,N_17703);
nand U20318 (N_20318,N_18415,N_16014);
xnor U20319 (N_20319,N_15992,N_19841);
or U20320 (N_20320,N_19290,N_15569);
or U20321 (N_20321,N_19993,N_19157);
and U20322 (N_20322,N_15652,N_17096);
nor U20323 (N_20323,N_15330,N_16653);
and U20324 (N_20324,N_19664,N_16160);
and U20325 (N_20325,N_17973,N_19739);
and U20326 (N_20326,N_19056,N_16578);
xnor U20327 (N_20327,N_15234,N_19957);
xnor U20328 (N_20328,N_17250,N_15344);
or U20329 (N_20329,N_16333,N_18560);
nor U20330 (N_20330,N_19358,N_15959);
or U20331 (N_20331,N_18076,N_17122);
nand U20332 (N_20332,N_15591,N_15660);
nand U20333 (N_20333,N_15831,N_17484);
nor U20334 (N_20334,N_17332,N_16486);
nor U20335 (N_20335,N_18391,N_15971);
nor U20336 (N_20336,N_18932,N_19539);
nand U20337 (N_20337,N_19267,N_15447);
nand U20338 (N_20338,N_16783,N_15662);
xor U20339 (N_20339,N_19477,N_17130);
or U20340 (N_20340,N_19733,N_16588);
nor U20341 (N_20341,N_18882,N_15173);
nand U20342 (N_20342,N_17661,N_16259);
xnor U20343 (N_20343,N_19470,N_15608);
nor U20344 (N_20344,N_17050,N_15869);
xor U20345 (N_20345,N_19862,N_15889);
nand U20346 (N_20346,N_15415,N_15540);
nand U20347 (N_20347,N_17447,N_16736);
and U20348 (N_20348,N_18147,N_19416);
and U20349 (N_20349,N_17252,N_17267);
xor U20350 (N_20350,N_15596,N_18866);
and U20351 (N_20351,N_19336,N_19941);
or U20352 (N_20352,N_17333,N_15872);
xor U20353 (N_20353,N_15106,N_16568);
and U20354 (N_20354,N_18327,N_18929);
and U20355 (N_20355,N_18845,N_18418);
and U20356 (N_20356,N_16291,N_17837);
nand U20357 (N_20357,N_17864,N_15991);
and U20358 (N_20358,N_17828,N_19577);
nor U20359 (N_20359,N_15134,N_17899);
nor U20360 (N_20360,N_18942,N_17822);
xnor U20361 (N_20361,N_16975,N_15286);
and U20362 (N_20362,N_16232,N_15133);
xor U20363 (N_20363,N_18544,N_15562);
nand U20364 (N_20364,N_16616,N_16406);
nor U20365 (N_20365,N_19351,N_16181);
or U20366 (N_20366,N_19224,N_18197);
and U20367 (N_20367,N_17780,N_16051);
or U20368 (N_20368,N_19728,N_18279);
xor U20369 (N_20369,N_16098,N_16336);
xor U20370 (N_20370,N_19173,N_19814);
nand U20371 (N_20371,N_17708,N_18694);
and U20372 (N_20372,N_17372,N_16373);
xnor U20373 (N_20373,N_16461,N_17736);
nor U20374 (N_20374,N_19226,N_16083);
nor U20375 (N_20375,N_18474,N_19601);
xnor U20376 (N_20376,N_16116,N_19276);
and U20377 (N_20377,N_18078,N_15264);
and U20378 (N_20378,N_16445,N_18981);
nor U20379 (N_20379,N_19435,N_15324);
xor U20380 (N_20380,N_16743,N_16569);
nor U20381 (N_20381,N_18665,N_15730);
and U20382 (N_20382,N_15884,N_19775);
nand U20383 (N_20383,N_15805,N_17763);
and U20384 (N_20384,N_18489,N_17019);
and U20385 (N_20385,N_18048,N_18609);
nor U20386 (N_20386,N_15086,N_18928);
nand U20387 (N_20387,N_19624,N_18144);
and U20388 (N_20388,N_15891,N_16419);
nor U20389 (N_20389,N_15948,N_19543);
nor U20390 (N_20390,N_18511,N_18247);
nor U20391 (N_20391,N_18102,N_15539);
nand U20392 (N_20392,N_18529,N_17756);
nor U20393 (N_20393,N_18768,N_16620);
and U20394 (N_20394,N_17651,N_18431);
xnor U20395 (N_20395,N_17304,N_15568);
nand U20396 (N_20396,N_18926,N_16402);
nand U20397 (N_20397,N_15998,N_15341);
nor U20398 (N_20398,N_16369,N_15607);
nand U20399 (N_20399,N_18451,N_15625);
and U20400 (N_20400,N_16854,N_16624);
or U20401 (N_20401,N_17768,N_17520);
nand U20402 (N_20402,N_16529,N_18631);
and U20403 (N_20403,N_15342,N_16444);
or U20404 (N_20404,N_17721,N_15474);
or U20405 (N_20405,N_18873,N_15492);
nor U20406 (N_20406,N_15072,N_16926);
nor U20407 (N_20407,N_16996,N_16099);
xor U20408 (N_20408,N_18293,N_18211);
nand U20409 (N_20409,N_15867,N_18411);
and U20410 (N_20410,N_18153,N_19508);
nand U20411 (N_20411,N_19618,N_17883);
nor U20412 (N_20412,N_17499,N_16598);
nor U20413 (N_20413,N_16848,N_18189);
xnor U20414 (N_20414,N_18993,N_15834);
xnor U20415 (N_20415,N_19717,N_15204);
or U20416 (N_20416,N_19724,N_15419);
nor U20417 (N_20417,N_16585,N_19426);
or U20418 (N_20418,N_19858,N_19216);
nor U20419 (N_20419,N_18369,N_16606);
or U20420 (N_20420,N_17349,N_15135);
and U20421 (N_20421,N_15630,N_15276);
and U20422 (N_20422,N_17196,N_17706);
and U20423 (N_20423,N_17021,N_17047);
or U20424 (N_20424,N_18414,N_19082);
and U20425 (N_20425,N_17642,N_17513);
nand U20426 (N_20426,N_17851,N_18600);
or U20427 (N_20427,N_18980,N_19663);
xnor U20428 (N_20428,N_19922,N_16092);
and U20429 (N_20429,N_17558,N_15669);
and U20430 (N_20430,N_19983,N_16673);
xnor U20431 (N_20431,N_19032,N_19496);
nor U20432 (N_20432,N_16560,N_17470);
nand U20433 (N_20433,N_16998,N_17016);
xor U20434 (N_20434,N_16429,N_17217);
nor U20435 (N_20435,N_18478,N_17510);
or U20436 (N_20436,N_19584,N_16101);
xor U20437 (N_20437,N_17297,N_18760);
and U20438 (N_20438,N_18023,N_18819);
nand U20439 (N_20439,N_15559,N_15089);
nor U20440 (N_20440,N_16853,N_15601);
nand U20441 (N_20441,N_16746,N_15556);
nor U20442 (N_20442,N_16733,N_17126);
or U20443 (N_20443,N_17580,N_18379);
xor U20444 (N_20444,N_17972,N_18780);
nor U20445 (N_20445,N_17226,N_19150);
nor U20446 (N_20446,N_16091,N_18844);
or U20447 (N_20447,N_19660,N_15668);
and U20448 (N_20448,N_16417,N_17639);
xnor U20449 (N_20449,N_19817,N_17291);
or U20450 (N_20450,N_15796,N_16617);
xor U20451 (N_20451,N_18758,N_16176);
and U20452 (N_20452,N_15414,N_16765);
nand U20453 (N_20453,N_19705,N_17055);
nor U20454 (N_20454,N_15736,N_19098);
nand U20455 (N_20455,N_19966,N_16027);
xnor U20456 (N_20456,N_15093,N_16408);
xor U20457 (N_20457,N_16272,N_15942);
xor U20458 (N_20458,N_15303,N_15919);
nor U20459 (N_20459,N_16658,N_19090);
nor U20460 (N_20460,N_17711,N_18063);
and U20461 (N_20461,N_18133,N_16613);
and U20462 (N_20462,N_15168,N_19084);
and U20463 (N_20463,N_19279,N_18803);
or U20464 (N_20464,N_15520,N_17787);
or U20465 (N_20465,N_19191,N_16346);
and U20466 (N_20466,N_15338,N_16337);
or U20467 (N_20467,N_17389,N_18740);
or U20468 (N_20468,N_16351,N_18518);
and U20469 (N_20469,N_15604,N_17432);
or U20470 (N_20470,N_16622,N_18692);
nor U20471 (N_20471,N_15319,N_19161);
nand U20472 (N_20472,N_18624,N_17980);
nand U20473 (N_20473,N_17501,N_16218);
or U20474 (N_20474,N_18455,N_18487);
and U20475 (N_20475,N_19652,N_15275);
xor U20476 (N_20476,N_17948,N_15766);
and U20477 (N_20477,N_19367,N_16022);
xnor U20478 (N_20478,N_16196,N_17604);
and U20479 (N_20479,N_16384,N_17037);
nand U20480 (N_20480,N_15076,N_19001);
xor U20481 (N_20481,N_17748,N_17001);
or U20482 (N_20482,N_15244,N_19286);
or U20483 (N_20483,N_17671,N_17819);
xor U20484 (N_20484,N_18041,N_17251);
and U20485 (N_20485,N_15195,N_17993);
nor U20486 (N_20486,N_16361,N_17556);
xor U20487 (N_20487,N_18729,N_16206);
xor U20488 (N_20488,N_19604,N_16201);
nand U20489 (N_20489,N_15293,N_16282);
nand U20490 (N_20490,N_19324,N_16454);
nand U20491 (N_20491,N_19240,N_17207);
and U20492 (N_20492,N_17680,N_16021);
nor U20493 (N_20493,N_15313,N_19129);
xnor U20494 (N_20494,N_19002,N_15110);
or U20495 (N_20495,N_15836,N_18813);
xnor U20496 (N_20496,N_16589,N_17597);
or U20497 (N_20497,N_19128,N_16787);
or U20498 (N_20498,N_19159,N_19939);
nor U20499 (N_20499,N_19189,N_16586);
xnor U20500 (N_20500,N_17537,N_17100);
xor U20501 (N_20501,N_15157,N_18696);
and U20502 (N_20502,N_18417,N_18743);
xnor U20503 (N_20503,N_15285,N_16768);
xor U20504 (N_20504,N_19019,N_19177);
and U20505 (N_20505,N_18958,N_17444);
or U20506 (N_20506,N_16001,N_18833);
nor U20507 (N_20507,N_16790,N_17970);
nor U20508 (N_20508,N_17849,N_16615);
and U20509 (N_20509,N_18720,N_17655);
nor U20510 (N_20510,N_15354,N_17256);
nor U20511 (N_20511,N_19511,N_15028);
nor U20512 (N_20512,N_17346,N_19648);
or U20513 (N_20513,N_17766,N_18003);
or U20514 (N_20514,N_17793,N_15394);
xnor U20515 (N_20515,N_18267,N_15126);
and U20516 (N_20516,N_18542,N_18264);
xnor U20517 (N_20517,N_18838,N_16003);
nor U20518 (N_20518,N_17827,N_16399);
or U20519 (N_20519,N_17495,N_16702);
nand U20520 (N_20520,N_16513,N_17125);
or U20521 (N_20521,N_15383,N_18563);
xnor U20522 (N_20522,N_18044,N_17776);
and U20523 (N_20523,N_16505,N_15222);
nand U20524 (N_20524,N_17636,N_16882);
nor U20525 (N_20525,N_19532,N_16059);
xor U20526 (N_20526,N_16796,N_19806);
nand U20527 (N_20527,N_17933,N_17779);
nor U20528 (N_20528,N_19977,N_16697);
or U20529 (N_20529,N_18238,N_17088);
and U20530 (N_20530,N_18922,N_17729);
and U20531 (N_20531,N_15724,N_17205);
or U20532 (N_20532,N_17707,N_18540);
or U20533 (N_20533,N_16973,N_19315);
and U20534 (N_20534,N_15751,N_19864);
or U20535 (N_20535,N_16104,N_18046);
nand U20536 (N_20536,N_19529,N_19837);
and U20537 (N_20537,N_19217,N_15904);
nor U20538 (N_20538,N_16205,N_16599);
nand U20539 (N_20539,N_16551,N_18574);
xor U20540 (N_20540,N_19382,N_15729);
or U20541 (N_20541,N_15145,N_18155);
nand U20542 (N_20542,N_15526,N_19561);
nand U20543 (N_20543,N_17545,N_15769);
or U20544 (N_20544,N_16010,N_19238);
and U20545 (N_20545,N_19445,N_19633);
xnor U20546 (N_20546,N_18213,N_15890);
nand U20547 (N_20547,N_17752,N_18338);
nor U20548 (N_20548,N_16418,N_18310);
xor U20549 (N_20549,N_19264,N_16930);
and U20550 (N_20550,N_15862,N_17223);
xnor U20551 (N_20551,N_18337,N_15099);
nand U20552 (N_20552,N_16832,N_15887);
and U20553 (N_20553,N_15032,N_18397);
nor U20554 (N_20554,N_17025,N_18090);
xnor U20555 (N_20555,N_15162,N_17590);
xnor U20556 (N_20556,N_18581,N_19744);
xor U20557 (N_20557,N_16364,N_18750);
nor U20558 (N_20558,N_19562,N_19653);
nand U20559 (N_20559,N_15547,N_17727);
or U20560 (N_20560,N_15918,N_19127);
and U20561 (N_20561,N_18714,N_18736);
nor U20562 (N_20562,N_15795,N_15019);
nand U20563 (N_20563,N_15714,N_19492);
or U20564 (N_20564,N_17049,N_17542);
xnor U20565 (N_20565,N_18423,N_16564);
nor U20566 (N_20566,N_18438,N_15155);
nor U20567 (N_20567,N_19273,N_18356);
nand U20568 (N_20568,N_15132,N_15873);
nand U20569 (N_20569,N_17461,N_15357);
xnor U20570 (N_20570,N_16552,N_16986);
and U20571 (N_20571,N_17861,N_17303);
and U20572 (N_20572,N_19752,N_17412);
or U20573 (N_20573,N_18012,N_16397);
xor U20574 (N_20574,N_15221,N_18430);
nand U20575 (N_20575,N_18412,N_17528);
and U20576 (N_20576,N_17343,N_19526);
nor U20577 (N_20577,N_15167,N_16357);
xor U20578 (N_20578,N_19112,N_18601);
and U20579 (N_20579,N_18976,N_15974);
or U20580 (N_20580,N_17998,N_17583);
and U20581 (N_20581,N_18918,N_15190);
nand U20582 (N_20582,N_17504,N_15312);
and U20583 (N_20583,N_16519,N_19873);
and U20584 (N_20584,N_16000,N_19182);
or U20585 (N_20585,N_16817,N_19345);
nor U20586 (N_20586,N_15042,N_19964);
xor U20587 (N_20587,N_16877,N_17123);
xnor U20588 (N_20588,N_15619,N_19985);
or U20589 (N_20589,N_19506,N_17104);
and U20590 (N_20590,N_17087,N_16403);
nor U20591 (N_20591,N_18158,N_17134);
xnor U20592 (N_20592,N_15092,N_18856);
and U20593 (N_20593,N_15832,N_16456);
xor U20594 (N_20594,N_16183,N_19447);
or U20595 (N_20595,N_18923,N_18006);
nor U20596 (N_20596,N_17700,N_18812);
xnor U20597 (N_20597,N_18867,N_19473);
xnor U20598 (N_20598,N_15579,N_19485);
nand U20599 (N_20599,N_19927,N_15586);
nand U20600 (N_20600,N_18755,N_16891);
xor U20601 (N_20601,N_16863,N_16920);
nand U20602 (N_20602,N_17186,N_18410);
nor U20603 (N_20603,N_19255,N_19089);
or U20604 (N_20604,N_19231,N_19237);
or U20605 (N_20605,N_19679,N_16725);
nand U20606 (N_20606,N_16166,N_18650);
nor U20607 (N_20607,N_18591,N_17139);
and U20608 (N_20608,N_15350,N_15713);
nand U20609 (N_20609,N_17902,N_15983);
nor U20610 (N_20610,N_18134,N_18662);
xnor U20611 (N_20611,N_16426,N_19973);
and U20612 (N_20612,N_18783,N_18717);
and U20613 (N_20613,N_18182,N_19556);
xor U20614 (N_20614,N_16661,N_17147);
nor U20615 (N_20615,N_18571,N_16601);
nor U20616 (N_20616,N_16324,N_17044);
and U20617 (N_20617,N_17958,N_18840);
and U20618 (N_20618,N_18047,N_17487);
or U20619 (N_20619,N_18785,N_19396);
and U20620 (N_20620,N_18208,N_15980);
nor U20621 (N_20621,N_15731,N_17526);
nand U20622 (N_20622,N_16458,N_15624);
or U20623 (N_20623,N_16177,N_19236);
nor U20624 (N_20624,N_16489,N_19980);
or U20625 (N_20625,N_17681,N_17936);
nor U20626 (N_20626,N_15927,N_19813);
and U20627 (N_20627,N_15243,N_16843);
xor U20628 (N_20628,N_16577,N_16758);
or U20629 (N_20629,N_15315,N_17013);
nand U20630 (N_20630,N_16801,N_19542);
and U20631 (N_20631,N_15049,N_19316);
nor U20632 (N_20632,N_17792,N_16047);
or U20633 (N_20633,N_18880,N_17852);
xnor U20634 (N_20634,N_15465,N_16316);
xor U20635 (N_20635,N_17734,N_18799);
nor U20636 (N_20636,N_19670,N_15018);
nand U20637 (N_20637,N_15590,N_16846);
and U20638 (N_20638,N_17543,N_19816);
xnor U20639 (N_20639,N_16913,N_18565);
or U20640 (N_20640,N_16706,N_17867);
nor U20641 (N_20641,N_17337,N_18567);
nor U20642 (N_20642,N_18184,N_17622);
and U20643 (N_20643,N_19613,N_16731);
nor U20644 (N_20644,N_16210,N_19605);
nor U20645 (N_20645,N_16473,N_16670);
nand U20646 (N_20646,N_19850,N_18471);
nor U20647 (N_20647,N_17112,N_18863);
nor U20648 (N_20648,N_17788,N_16527);
nor U20649 (N_20649,N_18148,N_17003);
nand U20650 (N_20650,N_17667,N_16730);
or U20651 (N_20651,N_15176,N_15810);
xor U20652 (N_20652,N_17955,N_18691);
and U20653 (N_20653,N_15030,N_16982);
nand U20654 (N_20654,N_15239,N_15544);
and U20655 (N_20655,N_19840,N_18009);
nand U20656 (N_20656,N_15504,N_19854);
and U20657 (N_20657,N_19799,N_17746);
or U20658 (N_20658,N_18790,N_18911);
and U20659 (N_20659,N_17245,N_19134);
or U20660 (N_20660,N_19736,N_18846);
and U20661 (N_20661,N_17659,N_17063);
nand U20662 (N_20662,N_18872,N_18118);
nor U20663 (N_20663,N_18592,N_19608);
or U20664 (N_20664,N_18641,N_18534);
or U20665 (N_20665,N_18959,N_19243);
and U20666 (N_20666,N_17559,N_17796);
nand U20667 (N_20667,N_18177,N_18516);
nand U20668 (N_20668,N_19655,N_15616);
and U20669 (N_20669,N_16915,N_16963);
or U20670 (N_20670,N_19323,N_16388);
and U20671 (N_20671,N_16401,N_17220);
nor U20672 (N_20672,N_16640,N_15746);
or U20673 (N_20673,N_18099,N_17228);
nand U20674 (N_20674,N_15382,N_19046);
or U20675 (N_20675,N_16048,N_16438);
nor U20676 (N_20676,N_15242,N_19374);
or U20677 (N_20677,N_19417,N_19935);
or U20678 (N_20678,N_15876,N_19695);
nor U20679 (N_20679,N_18401,N_17034);
nor U20680 (N_20680,N_16570,N_18757);
and U20681 (N_20681,N_15794,N_19711);
xnor U20682 (N_20682,N_18722,N_15305);
xor U20683 (N_20683,N_15252,N_19701);
nor U20684 (N_20684,N_16528,N_16825);
or U20685 (N_20685,N_19441,N_15227);
or U20686 (N_20686,N_19184,N_16342);
or U20687 (N_20687,N_19078,N_15782);
and U20688 (N_20688,N_16328,N_16994);
nor U20689 (N_20689,N_18320,N_16737);
or U20690 (N_20690,N_15215,N_15175);
and U20691 (N_20691,N_19391,N_18052);
and U20692 (N_20692,N_18906,N_17694);
and U20693 (N_20693,N_17127,N_18355);
and U20694 (N_20694,N_16147,N_16782);
and U20695 (N_20695,N_17665,N_17799);
or U20696 (N_20696,N_16434,N_18088);
nand U20697 (N_20697,N_19942,N_17138);
nor U20698 (N_20698,N_15010,N_17536);
nand U20699 (N_20699,N_16420,N_18202);
nand U20700 (N_20700,N_18506,N_18222);
or U20701 (N_20701,N_19199,N_16378);
nor U20702 (N_20702,N_16701,N_18297);
xor U20703 (N_20703,N_19931,N_18237);
xor U20704 (N_20704,N_16818,N_15480);
xor U20705 (N_20705,N_18483,N_15395);
nand U20706 (N_20706,N_17326,N_15819);
and U20707 (N_20707,N_18475,N_17946);
and U20708 (N_20708,N_15250,N_17638);
nand U20709 (N_20709,N_17213,N_19027);
or U20710 (N_20710,N_15811,N_17675);
or U20711 (N_20711,N_18317,N_17640);
xnor U20712 (N_20712,N_18488,N_15013);
nand U20713 (N_20713,N_17995,N_15119);
nand U20714 (N_20714,N_19761,N_19305);
nand U20715 (N_20715,N_15015,N_16062);
nand U20716 (N_20716,N_17375,N_17568);
nand U20717 (N_20717,N_18854,N_17552);
xor U20718 (N_20718,N_17185,N_19057);
or U20719 (N_20719,N_17606,N_16018);
nand U20720 (N_20720,N_19154,N_16812);
nor U20721 (N_20721,N_15320,N_16944);
nor U20722 (N_20722,N_15987,N_16669);
xor U20723 (N_20723,N_17359,N_19910);
nor U20724 (N_20724,N_16343,N_19641);
xnor U20725 (N_20725,N_17925,N_17380);
or U20726 (N_20726,N_19013,N_19114);
nand U20727 (N_20727,N_19206,N_16861);
or U20728 (N_20728,N_16876,N_18234);
and U20729 (N_20729,N_16411,N_18348);
nor U20730 (N_20730,N_19619,N_18248);
xor U20731 (N_20731,N_17975,N_18473);
xor U20732 (N_20732,N_18436,N_15278);
and U20733 (N_20733,N_16058,N_17391);
or U20734 (N_20734,N_19311,N_17187);
or U20735 (N_20735,N_16497,N_16549);
nand U20736 (N_20736,N_15950,N_16506);
and U20737 (N_20737,N_17425,N_19967);
and U20738 (N_20738,N_15491,N_18684);
or U20739 (N_20739,N_19497,N_17728);
xor U20740 (N_20740,N_16515,N_19415);
or U20741 (N_20741,N_15949,N_19997);
xnor U20742 (N_20742,N_17954,N_19397);
or U20743 (N_20743,N_16802,N_18062);
nand U20744 (N_20744,N_16777,N_15177);
xor U20745 (N_20745,N_18301,N_15859);
nor U20746 (N_20746,N_17753,N_17931);
or U20747 (N_20747,N_15634,N_16844);
xor U20748 (N_20748,N_17181,N_19575);
nor U20749 (N_20749,N_17369,N_19773);
nor U20750 (N_20750,N_18469,N_17312);
nand U20751 (N_20751,N_16102,N_16770);
nor U20752 (N_20752,N_17949,N_18404);
and U20753 (N_20753,N_17206,N_15255);
and U20754 (N_20754,N_18316,N_16472);
and U20755 (N_20755,N_16793,N_16744);
nor U20756 (N_20756,N_19716,N_18580);
nand U20757 (N_20757,N_18362,N_16200);
nor U20758 (N_20758,N_15635,N_19737);
or U20759 (N_20759,N_18666,N_18289);
and U20760 (N_20760,N_18635,N_18094);
xor U20761 (N_20761,N_19063,N_16779);
and U20762 (N_20762,N_17005,N_17227);
or U20763 (N_20763,N_16347,N_17271);
and U20764 (N_20764,N_19221,N_19152);
nor U20765 (N_20765,N_19355,N_17075);
and U20766 (N_20766,N_15462,N_16958);
and U20767 (N_20767,N_19000,N_16345);
xor U20768 (N_20768,N_19186,N_18294);
nor U20769 (N_20769,N_17491,N_16319);
or U20770 (N_20770,N_16498,N_16254);
and U20771 (N_20771,N_16807,N_19696);
nor U20772 (N_20772,N_17750,N_17449);
or U20773 (N_20773,N_15725,N_17554);
xor U20774 (N_20774,N_19839,N_16381);
nor U20775 (N_20775,N_17182,N_17097);
nor U20776 (N_20776,N_18553,N_16531);
nand U20777 (N_20777,N_17212,N_17984);
nor U20778 (N_20778,N_19138,N_15611);
nor U20779 (N_20779,N_15291,N_19131);
nor U20780 (N_20780,N_15937,N_17493);
nand U20781 (N_20781,N_18502,N_18933);
or U20782 (N_20782,N_17131,N_16903);
or U20783 (N_20783,N_17246,N_15355);
and U20784 (N_20784,N_19710,N_19787);
and U20785 (N_20785,N_19004,N_16902);
and U20786 (N_20786,N_15418,N_17843);
xnor U20787 (N_20787,N_18255,N_16910);
or U20788 (N_20788,N_17656,N_16747);
nand U20789 (N_20789,N_16788,N_16038);
and U20790 (N_20790,N_19847,N_18537);
and U20791 (N_20791,N_16501,N_19457);
xor U20792 (N_20792,N_17440,N_18724);
and U20793 (N_20793,N_19868,N_16096);
and U20794 (N_20794,N_18302,N_15943);
or U20795 (N_20795,N_15380,N_16948);
or U20796 (N_20796,N_15656,N_17323);
or U20797 (N_20797,N_18500,N_18753);
xnor U20798 (N_20798,N_16646,N_16922);
xnor U20799 (N_20799,N_17968,N_16929);
and U20800 (N_20800,N_16076,N_16603);
nand U20801 (N_20801,N_16045,N_18808);
or U20802 (N_20802,N_16692,N_17662);
nor U20803 (N_20803,N_19531,N_16088);
and U20804 (N_20804,N_18680,N_17725);
xnor U20805 (N_20805,N_17450,N_18123);
and U20806 (N_20806,N_18336,N_17254);
xnor U20807 (N_20807,N_18007,N_18655);
or U20808 (N_20808,N_18150,N_15196);
nor U20809 (N_20809,N_18349,N_15349);
xnor U20810 (N_20810,N_17399,N_17539);
or U20811 (N_20811,N_16186,N_17191);
nand U20812 (N_20812,N_16079,N_17564);
or U20813 (N_20813,N_17760,N_19790);
nand U20814 (N_20814,N_18206,N_15815);
nand U20815 (N_20815,N_15294,N_15266);
nor U20816 (N_20816,N_17802,N_19917);
xor U20817 (N_20817,N_17573,N_15327);
xnor U20818 (N_20818,N_15240,N_16409);
and U20819 (N_20819,N_17991,N_15933);
xnor U20820 (N_20820,N_18031,N_17959);
or U20821 (N_20821,N_16693,N_16404);
and U20822 (N_20822,N_15280,N_16376);
nor U20823 (N_20823,N_19928,N_18203);
or U20824 (N_20824,N_15524,N_15025);
xor U20825 (N_20825,N_18663,N_19827);
nand U20826 (N_20826,N_15518,N_17051);
nor U20827 (N_20827,N_17907,N_18025);
or U20828 (N_20828,N_18460,N_16655);
and U20829 (N_20829,N_17887,N_17445);
xor U20830 (N_20830,N_19849,N_16995);
nor U20831 (N_20831,N_17008,N_16241);
nor U20832 (N_20832,N_15694,N_16536);
xnor U20833 (N_20833,N_15144,N_15989);
xor U20834 (N_20834,N_18288,N_16439);
nor U20835 (N_20835,N_18325,N_15249);
xnor U20836 (N_20836,N_15541,N_15143);
and U20837 (N_20837,N_18021,N_17377);
nand U20838 (N_20838,N_18326,N_17442);
or U20839 (N_20839,N_17870,N_16660);
and U20840 (N_20840,N_17731,N_18399);
and U20841 (N_20841,N_16987,N_16198);
nand U20842 (N_20842,N_19667,N_15262);
or U20843 (N_20843,N_16484,N_19882);
nor U20844 (N_20844,N_18667,N_17897);
xor U20845 (N_20845,N_18904,N_16847);
nor U20846 (N_20846,N_16650,N_15457);
and U20847 (N_20847,N_18286,N_19411);
nand U20848 (N_20848,N_16631,N_16656);
or U20849 (N_20849,N_18820,N_16517);
and U20850 (N_20850,N_17778,N_18857);
xor U20851 (N_20851,N_19911,N_18428);
nand U20852 (N_20852,N_17506,N_16097);
xnor U20853 (N_20853,N_19729,N_19388);
or U20854 (N_20854,N_15642,N_16974);
nor U20855 (N_20855,N_19419,N_18333);
nor U20856 (N_20856,N_17532,N_15675);
nand U20857 (N_20857,N_16881,N_19763);
nand U20858 (N_20858,N_17818,N_18427);
xor U20859 (N_20859,N_15727,N_16972);
nor U20860 (N_20860,N_16187,N_15951);
and U20861 (N_20861,N_19330,N_19694);
nor U20862 (N_20862,N_19100,N_19110);
xnor U20863 (N_20863,N_16667,N_19794);
xnor U20864 (N_20864,N_17464,N_18457);
nor U20865 (N_20865,N_18029,N_17488);
nand U20866 (N_20866,N_16537,N_18697);
and U20867 (N_20867,N_17058,N_15165);
nor U20868 (N_20868,N_15905,N_18413);
xnor U20869 (N_20869,N_18917,N_19225);
nand U20870 (N_20870,N_15226,N_16938);
nor U20871 (N_20871,N_17585,N_18283);
nand U20872 (N_20872,N_17145,N_17886);
nor U20873 (N_20873,N_16039,N_19213);
nor U20874 (N_20874,N_19932,N_19842);
nand U20875 (N_20875,N_15748,N_15994);
and U20876 (N_20876,N_16144,N_18026);
xnor U20877 (N_20877,N_16540,N_19630);
or U20878 (N_20878,N_17643,N_19034);
xor U20879 (N_20879,N_16350,N_15201);
or U20880 (N_20880,N_19487,N_15678);
and U20881 (N_20881,N_15521,N_17411);
xor U20882 (N_20882,N_15848,N_19025);
xnor U20883 (N_20883,N_17305,N_19784);
xor U20884 (N_20884,N_16367,N_18818);
nor U20885 (N_20885,N_19202,N_15223);
xnor U20886 (N_20886,N_15258,N_15046);
nand U20887 (N_20887,N_19810,N_19099);
or U20888 (N_20888,N_18896,N_17678);
xnor U20889 (N_20889,N_19423,N_18930);
nand U20890 (N_20890,N_17938,N_15011);
nor U20891 (N_20891,N_18138,N_17666);
xor U20892 (N_20892,N_16009,N_19688);
nand U20893 (N_20893,N_16962,N_17634);
nand U20894 (N_20894,N_18252,N_16911);
or U20895 (N_20895,N_15645,N_16742);
or U20896 (N_20896,N_16143,N_19792);
xnor U20897 (N_20897,N_17259,N_16331);
nand U20898 (N_20898,N_19031,N_15522);
nand U20899 (N_20899,N_15426,N_17784);
or U20900 (N_20900,N_19087,N_15946);
or U20901 (N_20901,N_19756,N_19146);
and U20902 (N_20902,N_18322,N_15899);
and U20903 (N_20903,N_18458,N_18527);
or U20904 (N_20904,N_16315,N_17043);
or U20905 (N_20905,N_18835,N_17879);
nor U20906 (N_20906,N_19263,N_19885);
xnor U20907 (N_20907,N_17775,N_19400);
and U20908 (N_20908,N_17148,N_17027);
xor U20909 (N_20909,N_15673,N_18108);
nor U20910 (N_20910,N_16063,N_18389);
or U20911 (N_20911,N_15283,N_19281);
xor U20912 (N_20912,N_16688,N_16004);
xor U20913 (N_20913,N_16739,N_16940);
and U20914 (N_20914,N_19521,N_16738);
nor U20915 (N_20915,N_15740,N_17533);
xnor U20916 (N_20916,N_19405,N_15702);
or U20917 (N_20917,N_19650,N_16873);
and U20918 (N_20918,N_18579,N_15424);
and U20919 (N_20919,N_18329,N_15771);
nor U20920 (N_20920,N_15400,N_18842);
or U20921 (N_20921,N_16178,N_18607);
nand U20922 (N_20922,N_18091,N_16503);
and U20923 (N_20923,N_19809,N_17713);
or U20924 (N_20924,N_17888,N_19144);
or U20925 (N_20925,N_19430,N_17771);
and U20926 (N_20926,N_17572,N_16901);
nand U20927 (N_20927,N_15798,N_18996);
nor U20928 (N_20928,N_19384,N_19153);
nor U20929 (N_20929,N_19442,N_16753);
xnor U20930 (N_20930,N_19334,N_18935);
nand U20931 (N_20931,N_19681,N_18861);
nor U20932 (N_20932,N_15454,N_17472);
or U20933 (N_20933,N_18670,N_19684);
xnor U20934 (N_20934,N_18723,N_19996);
or U20935 (N_20935,N_19163,N_19909);
and U20936 (N_20936,N_19632,N_17790);
nand U20937 (N_20937,N_16571,N_16396);
nor U20938 (N_20938,N_19828,N_16683);
nand U20939 (N_20939,N_17566,N_16772);
nand U20940 (N_20940,N_15537,N_17422);
nand U20941 (N_20941,N_15583,N_17575);
or U20942 (N_20942,N_17953,N_18711);
nand U20943 (N_20943,N_18970,N_19354);
xnor U20944 (N_20944,N_19479,N_19527);
or U20945 (N_20945,N_19889,N_19254);
nand U20946 (N_20946,N_16253,N_17398);
nand U20947 (N_20947,N_15545,N_15653);
nor U20948 (N_20948,N_19750,N_18509);
or U20949 (N_20949,N_16180,N_17690);
or U20950 (N_20950,N_19259,N_16093);
nand U20951 (N_20951,N_17821,N_19625);
or U20952 (N_20952,N_15823,N_19621);
xor U20953 (N_20953,N_19647,N_16248);
nand U20954 (N_20954,N_15914,N_19793);
or U20955 (N_20955,N_18168,N_18022);
nand U20956 (N_20956,N_16671,N_15337);
or U20957 (N_20957,N_17839,N_15563);
or U20958 (N_20958,N_15198,N_15886);
or U20959 (N_20959,N_17847,N_19167);
and U20960 (N_20960,N_17594,N_16780);
nor U20961 (N_20961,N_16255,N_18490);
xor U20962 (N_20962,N_17331,N_15318);
or U20963 (N_20963,N_17190,N_16008);
nand U20964 (N_20964,N_19278,N_16785);
xor U20965 (N_20965,N_16629,N_17686);
or U20966 (N_20966,N_18903,N_16769);
or U20967 (N_20967,N_18173,N_17073);
nor U20968 (N_20968,N_15761,N_17467);
xnor U20969 (N_20969,N_19338,N_19175);
and U20970 (N_20970,N_19376,N_15045);
nor U20971 (N_20971,N_16690,N_18532);
nand U20972 (N_20972,N_19171,N_16806);
and U20973 (N_20973,N_15188,N_15610);
or U20974 (N_20974,N_17988,N_16594);
xor U20975 (N_20975,N_16593,N_17277);
or U20976 (N_20976,N_15707,N_18888);
nand U20977 (N_20977,N_15399,N_18346);
and U20978 (N_20978,N_19335,N_19103);
nor U20979 (N_20979,N_18737,N_18802);
and U20980 (N_20980,N_19569,N_17803);
nor U20981 (N_20981,N_16756,N_15358);
nand U20982 (N_20982,N_16339,N_17093);
and U20983 (N_20983,N_16173,N_18330);
or U20984 (N_20984,N_18646,N_18795);
xnor U20985 (N_20985,N_19721,N_17319);
xnor U20986 (N_20986,N_15827,N_17439);
nor U20987 (N_20987,N_17061,N_16611);
and U20988 (N_20988,N_19295,N_19594);
and U20989 (N_20989,N_18398,N_19306);
and U20990 (N_20990,N_18862,N_17872);
or U20991 (N_20991,N_18083,N_15693);
nor U20992 (N_20992,N_17489,N_16459);
nor U20993 (N_20993,N_18744,N_17719);
nor U20994 (N_20994,N_15498,N_16563);
nor U20995 (N_20995,N_19318,N_15343);
and U20996 (N_20996,N_19325,N_15174);
xnor U20997 (N_20997,N_15666,N_16657);
nor U20998 (N_20998,N_15256,N_17565);
nand U20999 (N_20999,N_19033,N_15001);
or U21000 (N_21000,N_18161,N_15063);
nand U21001 (N_21001,N_19611,N_17831);
nor U21002 (N_21002,N_17529,N_16216);
or U21003 (N_21003,N_17757,N_15391);
or U21004 (N_21004,N_17505,N_15968);
nand U21005 (N_21005,N_19389,N_17113);
or U21006 (N_21006,N_18479,N_15314);
nand U21007 (N_21007,N_16466,N_16904);
nand U21008 (N_21008,N_19071,N_17835);
or U21009 (N_21009,N_17657,N_15692);
or U21010 (N_21010,N_16591,N_16794);
nor U21011 (N_21011,N_18875,N_17356);
and U21012 (N_21012,N_15687,N_17812);
xnor U21013 (N_21013,N_19612,N_15427);
or U21014 (N_21014,N_17696,N_18829);
xor U21015 (N_21015,N_19697,N_17868);
nor U21016 (N_21016,N_18447,N_16893);
and U21017 (N_21017,N_16895,N_15218);
and U21018 (N_21018,N_17918,N_18292);
nand U21019 (N_21019,N_17820,N_19852);
and U21020 (N_21020,N_19954,N_18165);
nand U21021 (N_21021,N_18566,N_17502);
xnor U21022 (N_21022,N_17937,N_15684);
or U21023 (N_21023,N_18368,N_18235);
nand U21024 (N_21024,N_19271,N_18383);
and U21025 (N_21025,N_16542,N_15156);
xnor U21026 (N_21026,N_15954,N_16502);
nand U21027 (N_21027,N_15421,N_19820);
xor U21028 (N_21028,N_15580,N_19077);
or U21029 (N_21029,N_17941,N_19749);
xor U21030 (N_21030,N_15923,N_16122);
xor U21031 (N_21031,N_16524,N_17270);
nand U21032 (N_21032,N_15557,N_16977);
xor U21033 (N_21033,N_16482,N_16140);
nor U21034 (N_21034,N_19682,N_16582);
or U21035 (N_21035,N_15737,N_18754);
or U21036 (N_21036,N_15472,N_16961);
nand U21037 (N_21037,N_17648,N_16837);
and U21038 (N_21038,N_19053,N_16383);
and U21039 (N_21039,N_16835,N_18104);
or U21040 (N_21040,N_18215,N_17257);
and U21041 (N_21041,N_15401,N_15367);
and U21042 (N_21042,N_17177,N_15014);
nand U21043 (N_21043,N_17738,N_17901);
nor U21044 (N_21044,N_16708,N_18886);
nand U21045 (N_21045,N_19835,N_18381);
xnor U21046 (N_21046,N_18745,N_19843);
nand U21047 (N_21047,N_17519,N_19165);
nand U21048 (N_21048,N_17451,N_15699);
or U21049 (N_21049,N_15482,N_19476);
nor U21050 (N_21050,N_17963,N_16141);
nand U21051 (N_21051,N_17494,N_16309);
nand U21052 (N_21052,N_15340,N_19297);
xor U21053 (N_21053,N_17805,N_18273);
xnor U21054 (N_21054,N_19819,N_18351);
and U21055 (N_21055,N_19603,N_15900);
nand U21056 (N_21056,N_15124,N_17846);
or U21057 (N_21057,N_17726,N_15961);
xor U21058 (N_21058,N_19055,N_17943);
nand U21059 (N_21059,N_17408,N_18272);
nand U21060 (N_21060,N_17589,N_18246);
or U21061 (N_21061,N_18656,N_15352);
nor U21062 (N_21062,N_16644,N_15689);
xor U21063 (N_21063,N_15316,N_15304);
xnor U21064 (N_21064,N_18281,N_16748);
xor U21065 (N_21065,N_17971,N_16795);
nor U21066 (N_21066,N_15420,N_16023);
and U21067 (N_21067,N_18787,N_19832);
nor U21068 (N_21068,N_19265,N_16539);
and U21069 (N_21069,N_19947,N_17368);
or U21070 (N_21070,N_19899,N_17032);
or U21071 (N_21071,N_17094,N_19181);
or U21072 (N_21072,N_16652,N_17199);
nor U21073 (N_21073,N_17215,N_18358);
nand U21074 (N_21074,N_18055,N_18924);
and U21075 (N_21075,N_19943,N_16561);
nor U21076 (N_21076,N_19469,N_17247);
and U21077 (N_21077,N_17951,N_19235);
and U21078 (N_21078,N_15854,N_19304);
and U21079 (N_21079,N_15627,N_18766);
xnor U21080 (N_21080,N_15393,N_15444);
or U21081 (N_21081,N_17524,N_19105);
nand U21082 (N_21082,N_19936,N_15295);
nand U21083 (N_21083,N_19219,N_17324);
or U21084 (N_21084,N_18370,N_16407);
xnor U21085 (N_21085,N_16976,N_16400);
nand U21086 (N_21086,N_17631,N_19293);
xnor U21087 (N_21087,N_15003,N_17650);
and U21088 (N_21088,N_16674,N_16170);
xnor U21089 (N_21089,N_15269,N_16887);
xnor U21090 (N_21090,N_18117,N_17476);
xor U21091 (N_21091,N_15517,N_16778);
or U21092 (N_21092,N_16474,N_18548);
nand U21093 (N_21093,N_16665,N_17588);
or U21094 (N_21094,N_18798,N_17992);
or U21095 (N_21095,N_17203,N_17260);
nand U21096 (N_21096,N_15438,N_17124);
nand U21097 (N_21097,N_15623,N_18067);
or U21098 (N_21098,N_15062,N_17106);
nand U21099 (N_21099,N_19195,N_15938);
or U21100 (N_21100,N_15229,N_19680);
nand U21101 (N_21101,N_17854,N_16273);
nor U21102 (N_21102,N_18321,N_15377);
xnor U21103 (N_21103,N_18637,N_17903);
and U21104 (N_21104,N_18710,N_15425);
nor U21105 (N_21105,N_15364,N_15857);
xor U21106 (N_21106,N_17990,N_16798);
nor U21107 (N_21107,N_17420,N_18191);
xor U21108 (N_21108,N_17829,N_17912);
nand U21109 (N_21109,N_18967,N_17749);
or U21110 (N_21110,N_17807,N_15732);
and U21111 (N_21111,N_18728,N_18334);
nor U21112 (N_21112,N_17546,N_17362);
nand U21113 (N_21113,N_15069,N_15621);
and U21114 (N_21114,N_16338,N_16635);
nand U21115 (N_21115,N_18997,N_18747);
or U21116 (N_21116,N_15047,N_18378);
or U21117 (N_21117,N_15962,N_19884);
nand U21118 (N_21118,N_15371,N_17966);
xor U21119 (N_21119,N_17627,N_19446);
or U21120 (N_21120,N_16044,N_18898);
nor U21121 (N_21121,N_18912,N_16012);
nand U21122 (N_21122,N_15493,N_19965);
xnor U21123 (N_21123,N_19475,N_17599);
nand U21124 (N_21124,N_16202,N_17054);
nand U21125 (N_21125,N_18195,N_16164);
nor U21126 (N_21126,N_17929,N_19375);
or U21127 (N_21127,N_16898,N_19160);
xor U21128 (N_21128,N_15161,N_16341);
nor U21129 (N_21129,N_18157,N_19404);
and U21130 (N_21130,N_17175,N_19802);
and U21131 (N_21131,N_17624,N_19859);
or U21132 (N_21132,N_16243,N_15148);
nor U21133 (N_21133,N_16700,N_16630);
or U21134 (N_21134,N_18015,N_16840);
nor U21135 (N_21135,N_19313,N_15490);
or U21136 (N_21136,N_18620,N_18551);
and U21137 (N_21137,N_17183,N_15910);
nor U21138 (N_21138,N_19546,N_16453);
and U21139 (N_21139,N_17664,N_18602);
or U21140 (N_21140,N_15913,N_16968);
nor U21141 (N_21141,N_19026,N_16749);
xnor U21142 (N_21142,N_15102,N_17547);
and U21143 (N_21143,N_15958,N_17249);
or U21144 (N_21144,N_16392,N_19780);
nor U21145 (N_21145,N_18300,N_18290);
xor U21146 (N_21146,N_18318,N_16344);
xnor U21147 (N_21147,N_15453,N_17500);
nand U21148 (N_21148,N_18491,N_17085);
or U21149 (N_21149,N_18794,N_19205);
nand U21150 (N_21150,N_17028,N_18188);
xnor U21151 (N_21151,N_16191,N_17889);
nand U21152 (N_21152,N_15754,N_19826);
or U21153 (N_21153,N_15728,N_18170);
and U21154 (N_21154,N_16950,N_19121);
xor U21155 (N_21155,N_16032,N_16805);
xor U21156 (N_21156,N_16500,N_15525);
or U21157 (N_21157,N_15888,N_19830);
and U21158 (N_21158,N_18952,N_17415);
nor U21159 (N_21159,N_15903,N_17682);
or U21160 (N_21160,N_16511,N_15682);
and U21161 (N_21161,N_19320,N_17352);
nand U21162 (N_21162,N_15068,N_18595);
and U21163 (N_21163,N_19581,N_15964);
xor U21164 (N_21164,N_17783,N_17285);
and U21165 (N_21165,N_18130,N_19700);
nand U21166 (N_21166,N_15050,N_17482);
xnor U21167 (N_21167,N_16425,N_16368);
nor U21168 (N_21168,N_16592,N_17180);
nand U21169 (N_21169,N_16934,N_18217);
nand U21170 (N_21170,N_18716,N_18377);
or U21171 (N_21171,N_19075,N_15440);
or U21172 (N_21172,N_19326,N_15774);
xor U21173 (N_21173,N_18938,N_15976);
and U21174 (N_21174,N_19824,N_16354);
nand U21175 (N_21175,N_16123,N_15059);
and U21176 (N_21176,N_15237,N_18541);
xor U21177 (N_21177,N_18625,N_16073);
or U21178 (N_21178,N_16627,N_15362);
xor U21179 (N_21179,N_15288,N_17549);
and U21180 (N_21180,N_18683,N_17446);
nand U21181 (N_21181,N_19658,N_18253);
and U21182 (N_21182,N_17745,N_19096);
and U21183 (N_21183,N_15034,N_18359);
and U21184 (N_21184,N_15822,N_17040);
and U21185 (N_21185,N_17584,N_19248);
or U21186 (N_21186,N_19860,N_18116);
nor U21187 (N_21187,N_16639,N_18593);
nor U21188 (N_21188,N_19383,N_19022);
nand U21189 (N_21189,N_15435,N_15445);
and U21190 (N_21190,N_16249,N_15502);
and U21191 (N_21191,N_18764,N_16132);
xnor U21192 (N_21192,N_17342,N_15431);
nor U21193 (N_21193,N_16558,N_18841);
or U21194 (N_21194,N_19005,N_16174);
xor U21195 (N_21195,N_15966,N_15781);
nand U21196 (N_21196,N_15755,N_18733);
or U21197 (N_21197,N_17660,N_18575);
nand U21198 (N_21198,N_19895,N_16897);
xor U21199 (N_21199,N_15458,N_16221);
xnor U21200 (N_21200,N_17264,N_16312);
and U21201 (N_21201,N_17386,N_19714);
xor U21202 (N_21202,N_16440,N_15947);
or U21203 (N_21203,N_17433,N_18960);
nand U21204 (N_21204,N_15441,N_18525);
nand U21205 (N_21205,N_15235,N_19386);
xnor U21206 (N_21206,N_17426,N_16352);
nand U21207 (N_21207,N_15033,N_16476);
nand U21208 (N_21208,N_19989,N_19615);
xor U21209 (N_21209,N_18651,N_19328);
nor U21210 (N_21210,N_18931,N_16828);
or U21211 (N_21211,N_19373,N_18110);
nand U21212 (N_21212,N_15037,N_19726);
nor U21213 (N_21213,N_18077,N_19505);
and U21214 (N_21214,N_15451,N_19253);
nand U21215 (N_21215,N_15469,N_17548);
or U21216 (N_21216,N_16831,N_17344);
nor U21217 (N_21217,N_19628,N_16548);
and U21218 (N_21218,N_17579,N_18421);
nand U21219 (N_21219,N_19523,N_17143);
xor U21220 (N_21220,N_17741,N_18126);
xnor U21221 (N_21221,N_15486,N_17390);
nand U21222 (N_21222,N_18454,N_17534);
or U21223 (N_21223,N_16923,N_19952);
xnor U21224 (N_21224,N_17146,N_17860);
or U21225 (N_21225,N_15528,N_19343);
or U21226 (N_21226,N_17236,N_18654);
nand U21227 (N_21227,N_15723,N_15373);
and U21228 (N_21228,N_16687,N_15786);
xor U21229 (N_21229,N_17109,N_19617);
xor U21230 (N_21230,N_17255,N_15456);
or U21231 (N_21231,N_15999,N_16608);
and U21232 (N_21232,N_15027,N_16279);
xnor U21233 (N_21233,N_18245,N_16546);
xnor U21234 (N_21234,N_18494,N_17102);
xor U21235 (N_21235,N_19891,N_15260);
nor U21236 (N_21236,N_18816,N_19955);
or U21237 (N_21237,N_15351,N_16719);
or U21238 (N_21238,N_15302,N_17268);
xnor U21239 (N_21239,N_15405,N_15392);
or U21240 (N_21240,N_18061,N_17460);
xnor U21241 (N_21241,N_15189,N_18142);
and U21242 (N_21242,N_19499,N_15812);
xnor U21243 (N_21243,N_16247,N_19552);
xnor U21244 (N_21244,N_17762,N_16965);
or U21245 (N_21245,N_18307,N_16516);
nor U21246 (N_21246,N_18180,N_19155);
nor U21247 (N_21247,N_16182,N_19547);
nor U21248 (N_21248,N_18045,N_15153);
nand U21249 (N_21249,N_18849,N_18341);
or U21250 (N_21250,N_18828,N_19982);
or U21251 (N_21251,N_16245,N_19738);
or U21252 (N_21252,N_17747,N_17284);
xnor U21253 (N_21253,N_15247,N_18894);
nor U21254 (N_21254,N_18441,N_15985);
xor U21255 (N_21255,N_17238,N_16988);
nor U21256 (N_21256,N_16618,N_15021);
and U21257 (N_21257,N_16981,N_16308);
or U21258 (N_21258,N_19432,N_16478);
nor U21259 (N_21259,N_19559,N_15957);
xnor U21260 (N_21260,N_18735,N_16213);
nor U21261 (N_21261,N_19197,N_19109);
and U21262 (N_21262,N_18831,N_18392);
or U21263 (N_21263,N_16130,N_18990);
nor U21264 (N_21264,N_19915,N_19699);
nand U21265 (N_21265,N_17035,N_19269);
and U21266 (N_21266,N_16246,N_19049);
or U21267 (N_21267,N_18763,N_16110);
nand U21268 (N_21268,N_15081,N_17610);
or U21269 (N_21269,N_19431,N_16161);
nand U21270 (N_21270,N_17615,N_15390);
nand U21271 (N_21271,N_18259,N_15695);
nand U21272 (N_21272,N_18877,N_16584);
nand U21273 (N_21273,N_19148,N_16433);
and U21274 (N_21274,N_18895,N_18612);
nand U21275 (N_21275,N_17485,N_15849);
or U21276 (N_21276,N_19563,N_17979);
or U21277 (N_21277,N_18181,N_15432);
nand U21278 (N_21278,N_19251,N_17587);
xor U21279 (N_21279,N_16645,N_17480);
nor U21280 (N_21280,N_17151,N_16072);
and U21281 (N_21281,N_17172,N_19020);
and U21282 (N_21282,N_16220,N_18112);
or U21283 (N_21283,N_19912,N_16724);
and U21284 (N_21284,N_16139,N_16761);
nand U21285 (N_21285,N_19300,N_19168);
nand U21286 (N_21286,N_17904,N_18420);
nor U21287 (N_21287,N_15460,N_16077);
and U21288 (N_21288,N_17281,N_16085);
nor U21289 (N_21289,N_15129,N_17406);
nor U21290 (N_21290,N_15706,N_16999);
xor U21291 (N_21291,N_18779,N_18385);
or U21292 (N_21292,N_16056,N_19456);
or U21293 (N_21293,N_17965,N_19578);
and U21294 (N_21294,N_15231,N_18668);
and U21295 (N_21295,N_17535,N_17156);
and U21296 (N_21296,N_18664,N_19893);
nand U21297 (N_21297,N_15094,N_17132);
nor U21298 (N_21298,N_16067,N_16809);
nand U21299 (N_21299,N_15654,N_18852);
xor U21300 (N_21300,N_19392,N_17009);
nand U21301 (N_21301,N_17014,N_18080);
xor U21302 (N_21302,N_15972,N_17423);
or U21303 (N_21303,N_16971,N_19640);
xor U21304 (N_21304,N_17617,N_15232);
and U21305 (N_21305,N_15499,N_15029);
nor U21306 (N_21306,N_16390,N_16810);
and U21307 (N_21307,N_15333,N_19450);
nand U21308 (N_21308,N_15411,N_17717);
or U21309 (N_21309,N_16838,N_19875);
or U21310 (N_21310,N_18343,N_16050);
nor U21311 (N_21311,N_15661,N_15172);
and U21312 (N_21312,N_16879,N_16855);
xnor U21313 (N_21313,N_17591,N_17507);
and U21314 (N_21314,N_16026,N_19064);
xnor U21315 (N_21315,N_18597,N_17873);
nor U21316 (N_21316,N_19344,N_18965);
or U21317 (N_21317,N_18577,N_16696);
or U21318 (N_21318,N_18242,N_16959);
xnor U21319 (N_21319,N_17334,N_19244);
and U21320 (N_21320,N_15576,N_19579);
nand U21321 (N_21321,N_18987,N_17986);
or U21322 (N_21322,N_19359,N_15413);
or U21323 (N_21323,N_16808,N_19962);
nand U21324 (N_21324,N_17144,N_16685);
nor U21325 (N_21325,N_18284,N_17364);
or U21326 (N_21326,N_19484,N_16298);
or U21327 (N_21327,N_15552,N_15058);
nand U21328 (N_21328,N_18944,N_17455);
nor U21329 (N_21329,N_17926,N_15932);
and U21330 (N_21330,N_17620,N_18769);
nor U21331 (N_21331,N_16979,N_16295);
xnor U21332 (N_21332,N_19803,N_19933);
and U21333 (N_21333,N_15265,N_18220);
nor U21334 (N_21334,N_19574,N_19101);
and U21335 (N_21335,N_19795,N_19923);
and U21336 (N_21336,N_18741,N_19870);
nand U21337 (N_21337,N_18128,N_16485);
or U21338 (N_21338,N_19200,N_18919);
xor U21339 (N_21339,N_17078,N_15908);
nand U21340 (N_21340,N_17076,N_19951);
and U21341 (N_21341,N_19626,N_15048);
or U21342 (N_21342,N_16375,N_18583);
xor U21343 (N_21343,N_19866,N_18749);
and U21344 (N_21344,N_18966,N_17373);
nor U21345 (N_21345,N_16927,N_18331);
xnor U21346 (N_21346,N_15238,N_19014);
or U21347 (N_21347,N_15087,N_19361);
xor U21348 (N_21348,N_17178,N_17613);
or U21349 (N_21349,N_15839,N_17273);
nand U21350 (N_21350,N_16137,N_18533);
nand U21351 (N_21351,N_17616,N_18435);
or U21352 (N_21352,N_19194,N_18558);
or U21353 (N_21353,N_17289,N_15085);
nand U21354 (N_21354,N_16208,N_15209);
or U21355 (N_21355,N_15442,N_15509);
nand U21356 (N_21356,N_19634,N_18408);
nand U21357 (N_21357,N_16713,N_19003);
and U21358 (N_21358,N_18698,N_17743);
nor U21359 (N_21359,N_17347,N_15043);
and U21360 (N_21360,N_16305,N_19091);
xor U21361 (N_21361,N_18937,N_18801);
or U21362 (N_21362,N_19755,N_16483);
and U21363 (N_21363,N_16153,N_16251);
nor U21364 (N_21364,N_18493,N_17434);
nand U21365 (N_21365,N_16951,N_15531);
and U21366 (N_21366,N_19223,N_15920);
nand U21367 (N_21367,N_15756,N_19865);
nand U21368 (N_21368,N_15622,N_19258);
xnor U21369 (N_21369,N_18350,N_15816);
nor U21370 (N_21370,N_17318,N_15690);
nand U21371 (N_21371,N_15850,N_15651);
xnor U21372 (N_21372,N_16914,N_17118);
nand U21373 (N_21373,N_16870,N_18539);
nand U21374 (N_21374,N_17431,N_18268);
xnor U21375 (N_21375,N_18249,N_15039);
nor U21376 (N_21376,N_16874,N_18955);
nor U21377 (N_21377,N_19073,N_17026);
xor U21378 (N_21378,N_17239,N_17039);
xnor U21379 (N_21379,N_16595,N_15901);
xnor U21380 (N_21380,N_19188,N_15436);
nand U21381 (N_21381,N_15308,N_18185);
nor U21382 (N_21382,N_15768,N_16289);
xnor U21383 (N_21383,N_19533,N_15745);
xor U21384 (N_21384,N_15005,N_18260);
or U21385 (N_21385,N_17086,N_16090);
and U21386 (N_21386,N_17262,N_19108);
nor U21387 (N_21387,N_18588,N_19518);
nand U21388 (N_21388,N_19509,N_15067);
nand U21389 (N_21389,N_18477,N_18205);
xor U21390 (N_21390,N_19280,N_18893);
or U21391 (N_21391,N_19818,N_18669);
nor U21392 (N_21392,N_19452,N_15763);
xor U21393 (N_21393,N_15122,N_18363);
and U21394 (N_21394,N_15473,N_17188);
nand U21395 (N_21395,N_15307,N_16450);
nand U21396 (N_21396,N_17562,N_19771);
or U21397 (N_21397,N_18132,N_15261);
and U21398 (N_21398,N_16095,N_19029);
xnor U21399 (N_21399,N_15575,N_19040);
or U21400 (N_21400,N_16155,N_18732);
xor U21401 (N_21401,N_17996,N_16909);
or U21402 (N_21402,N_16686,N_17724);
xnor U21403 (N_21403,N_16680,N_19076);
and U21404 (N_21404,N_17561,N_15346);
xnor U21405 (N_21405,N_16803,N_15248);
nand U21406 (N_21406,N_19398,N_15988);
nand U21407 (N_21407,N_19853,N_19393);
or U21408 (N_21408,N_17179,N_19727);
xor U21409 (N_21409,N_19758,N_19261);
and U21410 (N_21410,N_16427,N_19474);
and U21411 (N_21411,N_19288,N_15128);
or U21412 (N_21412,N_19132,N_18800);
nand U21413 (N_21413,N_19959,N_17755);
and U21414 (N_21414,N_19418,N_16389);
or U21415 (N_21415,N_16641,N_18212);
and U21416 (N_21416,N_18030,N_17623);
xor U21417 (N_21417,N_18618,N_15071);
xor U21418 (N_21418,N_17397,N_18826);
xnor U21419 (N_21419,N_17232,N_17384);
and U21420 (N_21420,N_19319,N_17167);
or U21421 (N_21421,N_18163,N_19902);
or U21422 (N_21422,N_19036,N_15558);
or U21423 (N_21423,N_16949,N_17744);
nor U21424 (N_21424,N_19366,N_18033);
and U21425 (N_21425,N_16238,N_16332);
nand U21426 (N_21426,N_19047,N_15709);
xor U21427 (N_21427,N_18973,N_15035);
or U21428 (N_21428,N_18271,N_19145);
nand U21429 (N_21429,N_15877,N_16306);
or U21430 (N_21430,N_15560,N_17677);
nor U21431 (N_21431,N_16074,N_18707);
or U21432 (N_21432,N_16296,N_17892);
nor U21433 (N_21433,N_17082,N_18426);
nand U21434 (N_21434,N_18850,N_18243);
nand U21435 (N_21435,N_19920,N_17646);
xor U21436 (N_21436,N_19541,N_19767);
and U21437 (N_21437,N_16889,N_17608);
or U21438 (N_21438,N_19427,N_16244);
or U21439 (N_21439,N_16841,N_15450);
nand U21440 (N_21440,N_17999,N_19990);
or U21441 (N_21441,N_18908,N_19115);
and U21442 (N_21442,N_19921,N_18057);
xor U21443 (N_21443,N_17950,N_15494);
and U21444 (N_21444,N_15990,N_18042);
and U21445 (N_21445,N_15671,N_17699);
xnor U21446 (N_21446,N_17216,N_19662);
or U21447 (N_21447,N_19953,N_19008);
or U21448 (N_21448,N_16707,N_15553);
and U21449 (N_21449,N_18902,N_16120);
xnor U21450 (N_21450,N_17275,N_16148);
or U21451 (N_21451,N_19410,N_19823);
and U21452 (N_21452,N_17059,N_15716);
nor U21453 (N_21453,N_18256,N_15717);
nor U21454 (N_21454,N_15065,N_18810);
or U21455 (N_21455,N_17154,N_18437);
and U21456 (N_21456,N_15613,N_16970);
nand U21457 (N_21457,N_19715,N_16131);
nor U21458 (N_21458,N_16471,N_15408);
and U21459 (N_21459,N_19583,N_15111);
nand U21460 (N_21460,N_15841,N_19371);
nor U21461 (N_21461,N_18920,N_18699);
nor U21462 (N_21462,N_19720,N_18573);
nor U21463 (N_21463,N_18194,N_15476);
xor U21464 (N_21464,N_16046,N_19576);
and U21465 (N_21465,N_17823,N_17149);
nand U21466 (N_21466,N_19460,N_17159);
or U21467 (N_21467,N_19768,N_19209);
nor U21468 (N_21468,N_16716,N_16146);
and U21469 (N_21469,N_16149,N_19969);
nand U21470 (N_21470,N_17367,N_15649);
nor U21471 (N_21471,N_18395,N_18228);
nor U21472 (N_21472,N_19570,N_17231);
xnor U21473 (N_21473,N_18788,N_15718);
nand U21474 (N_21474,N_15797,N_16329);
nand U21475 (N_21475,N_16572,N_15779);
and U21476 (N_21476,N_16535,N_17960);
or U21477 (N_21477,N_16931,N_19512);
xor U21478 (N_21478,N_18531,N_15593);
nor U21479 (N_21479,N_19903,N_19294);
and U21480 (N_21480,N_18871,N_16327);
xnor U21481 (N_21481,N_16508,N_19471);
or U21482 (N_21482,N_19685,N_17786);
or U21483 (N_21483,N_17895,N_15842);
nor U21484 (N_21484,N_15224,N_17577);
or U21485 (N_21485,N_17898,N_17358);
nand U21486 (N_21486,N_18590,N_17515);
nor U21487 (N_21487,N_15241,N_18295);
xor U21488 (N_21488,N_15907,N_18439);
nand U21489 (N_21489,N_17295,N_15565);
and U21490 (N_21490,N_16013,N_15104);
nand U21491 (N_21491,N_17320,N_16224);
nand U21492 (N_21492,N_19104,N_16106);
and U21493 (N_21493,N_17306,N_18036);
or U21494 (N_21494,N_19760,N_17742);
nand U21495 (N_21495,N_17672,N_15511);
or U21496 (N_21496,N_17490,N_15770);
and U21497 (N_21497,N_18817,N_16214);
xor U21498 (N_21498,N_19356,N_18782);
xor U21499 (N_21499,N_15790,N_19342);
xor U21500 (N_21500,N_16326,N_19133);
nand U21501 (N_21501,N_19394,N_18071);
or U21502 (N_21502,N_16302,N_18545);
or U21503 (N_21503,N_18113,N_19930);
xnor U21504 (N_21504,N_18319,N_15701);
and U21505 (N_21505,N_17629,N_19070);
and U21506 (N_21506,N_17098,N_17435);
nor U21507 (N_21507,N_17540,N_15206);
nand U21508 (N_21508,N_18679,N_19038);
nor U21509 (N_21509,N_17194,N_15871);
nand U21510 (N_21510,N_18393,N_15636);
nor U21511 (N_21511,N_16460,N_15078);
and U21512 (N_21512,N_15064,N_19009);
nor U21513 (N_21513,N_17630,N_16432);
nand U21514 (N_21514,N_15883,N_18940);
nand U21515 (N_21515,N_18962,N_16663);
xor U21516 (N_21516,N_18605,N_18328);
nor U21517 (N_21517,N_15825,N_17714);
and U21518 (N_21518,N_17308,N_17774);
nand U21519 (N_21519,N_17683,N_17038);
or U21520 (N_21520,N_17574,N_17394);
nor U21521 (N_21521,N_17496,N_18190);
xnor U21522 (N_21522,N_16274,N_15637);
and U21523 (N_21523,N_15245,N_18536);
and U21524 (N_21524,N_17327,N_17863);
and U21525 (N_21525,N_18562,N_16574);
nand U21526 (N_21526,N_17283,N_16301);
xor U21527 (N_21527,N_18507,N_19333);
nor U21528 (N_21528,N_18519,N_19905);
xnor U21529 (N_21529,N_18429,N_18673);
nand U21530 (N_21530,N_18640,N_19233);
nor U21531 (N_21531,N_19314,N_19671);
xor U21532 (N_21532,N_18916,N_15934);
or U21533 (N_21533,N_15739,N_17020);
xnor U21534 (N_21534,N_18514,N_16623);
nand U21535 (N_21535,N_15757,N_18059);
and U21536 (N_21536,N_19564,N_17376);
or U21537 (N_21537,N_15463,N_17400);
or U21538 (N_21538,N_19303,N_18954);
and U21539 (N_21539,N_19021,N_16423);
or U21540 (N_21540,N_17531,N_19590);
and U21541 (N_21541,N_16820,N_15738);
or U21542 (N_21542,N_18244,N_15105);
xnor U21543 (N_21543,N_17024,N_18594);
or U21544 (N_21544,N_16168,N_18459);
xor U21545 (N_21545,N_15708,N_18878);
nand U21546 (N_21546,N_19256,N_18058);
and U21547 (N_21547,N_19743,N_19164);
or U21548 (N_21548,N_17292,N_15676);
nor U21549 (N_21549,N_17825,N_19589);
and U21550 (N_21550,N_19170,N_15952);
nor U21551 (N_21551,N_18834,N_18040);
or U21552 (N_21552,N_18901,N_17382);
xor U21553 (N_21553,N_15609,N_15572);
nand U21554 (N_21554,N_18968,N_16113);
and U21555 (N_21555,N_17688,N_16969);
nand U21556 (N_21556,N_17663,N_18394);
or U21557 (N_21557,N_18726,N_19037);
and U21558 (N_21558,N_18167,N_16121);
and U21559 (N_21559,N_15554,N_17601);
nor U21560 (N_21560,N_18066,N_15356);
xnor U21561 (N_21561,N_17952,N_17353);
and U21562 (N_21562,N_16610,N_15897);
xor U21563 (N_21563,N_15564,N_18644);
nand U21564 (N_21564,N_15006,N_17477);
and U21565 (N_21565,N_18400,N_17845);
xor U21566 (N_21566,N_18626,N_18524);
nand U21567 (N_21567,N_18406,N_17355);
nor U21568 (N_21568,N_18576,N_16937);
nor U21569 (N_21569,N_17924,N_17740);
and U21570 (N_21570,N_17795,N_18661);
nor U21571 (N_21571,N_18001,N_16304);
nor U21572 (N_21572,N_17720,N_19677);
xnor U21573 (N_21573,N_15433,N_15503);
nand U21574 (N_21574,N_18277,N_18633);
nand U21575 (N_21575,N_17715,N_15715);
xnor U21576 (N_21576,N_19683,N_19974);
xor U21577 (N_21577,N_18839,N_19999);
or U21578 (N_21578,N_16842,N_17782);
and U21579 (N_21579,N_16960,N_15363);
and U21580 (N_21580,N_19560,N_15154);
and U21581 (N_21581,N_16576,N_18582);
xnor U21582 (N_21582,N_16952,N_19851);
nand U21583 (N_21583,N_19551,N_15711);
nand U21584 (N_21584,N_18807,N_19015);
nor U21585 (N_21585,N_15205,N_15581);
nand U21586 (N_21586,N_16954,N_18914);
or U21587 (N_21587,N_19880,N_17913);
nor U21588 (N_21588,N_15902,N_18160);
nand U21589 (N_21589,N_15628,N_15292);
xor U21590 (N_21590,N_16530,N_15911);
nor U21591 (N_21591,N_15365,N_18313);
and U21592 (N_21592,N_16763,N_19066);
nor U21593 (N_21593,N_16990,N_17698);
nand U21594 (N_21594,N_19643,N_15765);
xnor U21595 (N_21595,N_17340,N_18899);
nand U21596 (N_21596,N_18561,N_18339);
and U21597 (N_21597,N_15650,N_19437);
or U21598 (N_21598,N_19011,N_16124);
or U21599 (N_21599,N_19212,N_19975);
and U21600 (N_21600,N_17011,N_19668);
nor U21601 (N_21601,N_15024,N_18688);
nand U21602 (N_21602,N_18017,N_19622);
and U21603 (N_21603,N_16299,N_15772);
and U21604 (N_21604,N_16512,N_19519);
nand U21605 (N_21605,N_19291,N_16209);
xor U21606 (N_21606,N_18374,N_19054);
and U21607 (N_21607,N_19302,N_19678);
and U21608 (N_21608,N_17311,N_15310);
and U21609 (N_21609,N_19428,N_16374);
nand U21610 (N_21610,N_19017,N_18038);
or U21611 (N_21611,N_16040,N_18068);
or U21612 (N_21612,N_19395,N_15375);
nor U21613 (N_21613,N_15570,N_18613);
xor U21614 (N_21614,N_16900,N_19491);
nor U21615 (N_21615,N_16662,N_16638);
nor U21616 (N_21616,N_19018,N_18074);
or U21617 (N_21617,N_15207,N_16410);
nand U21618 (N_21618,N_16109,N_15468);
nor U21619 (N_21619,N_15720,N_16060);
xnor U21620 (N_21620,N_19482,N_15017);
nand U21621 (N_21621,N_19981,N_15187);
nor U21622 (N_21622,N_18734,N_17006);
or U21623 (N_21623,N_18616,N_19838);
nand U21624 (N_21624,N_15658,N_17478);
and U21625 (N_21625,N_19402,N_15573);
and U21626 (N_21626,N_18219,N_18870);
and U21627 (N_21627,N_15543,N_15764);
and U21628 (N_21628,N_17658,N_19363);
nand U21629 (N_21629,N_17692,N_18830);
or U21630 (N_21630,N_15861,N_15758);
nand U21631 (N_21631,N_16878,N_19403);
nor U21632 (N_21632,N_15597,N_16082);
nand U21633 (N_21633,N_18388,N_15359);
or U21634 (N_21634,N_15112,N_18569);
or U21635 (N_21635,N_18043,N_19048);
nor U21636 (N_21636,N_16325,N_15773);
and U21637 (N_21637,N_17350,N_18360);
nand U21638 (N_21638,N_19272,N_18192);
nand U21639 (N_21639,N_19867,N_16193);
and U21640 (N_21640,N_17551,N_18463);
nor U21641 (N_21641,N_16757,N_16185);
and U21642 (N_21642,N_15496,N_19596);
xnor U21643 (N_21643,N_16751,N_19135);
xnor U21644 (N_21644,N_19781,N_16016);
or U21645 (N_21645,N_16447,N_17668);
nand U21646 (N_21646,N_19407,N_18971);
or U21647 (N_21647,N_15582,N_18166);
or U21648 (N_21648,N_17702,N_15577);
xnor U21649 (N_21649,N_17626,N_19798);
nor U21650 (N_21650,N_15719,N_15507);
nor U21651 (N_21651,N_18100,N_18772);
nand U21652 (N_21652,N_17365,N_17140);
nand U21653 (N_21653,N_15023,N_18983);
or U21654 (N_21654,N_17806,N_15194);
nand U21655 (N_21655,N_19341,N_17429);
and U21656 (N_21656,N_17578,N_16265);
and U21657 (N_21657,N_17994,N_18510);
nand U21658 (N_21658,N_15603,N_16799);
and U21659 (N_21659,N_19944,N_18742);
or U21660 (N_21660,N_15159,N_15529);
and U21661 (N_21661,N_16633,N_15115);
nor U21662 (N_21662,N_16222,N_17865);
nand U21663 (N_21663,N_18824,N_18584);
xor U21664 (N_21664,N_18659,N_15114);
and U21665 (N_21665,N_16443,N_18060);
or U21666 (N_21666,N_19686,N_16619);
nor U21667 (N_21667,N_19299,N_19232);
xnor U21668 (N_21668,N_16167,N_19220);
nor U21669 (N_21669,N_19504,N_17117);
and U21670 (N_21670,N_16520,N_16573);
or U21671 (N_21671,N_19369,N_18649);
nand U21672 (N_21672,N_18627,N_18554);
nand U21673 (N_21673,N_15348,N_17313);
nand U21674 (N_21674,N_19703,N_16398);
nand U21675 (N_21675,N_19007,N_19872);
xnor U21676 (N_21676,N_16583,N_17237);
and U21677 (N_21677,N_15370,N_16567);
and U21678 (N_21678,N_17081,N_19097);
or U21679 (N_21679,N_19377,N_16543);
and U21680 (N_21680,N_17939,N_19555);
xnor U21681 (N_21681,N_15284,N_16935);
nor U21682 (N_21682,N_17840,N_15334);
nand U21683 (N_21683,N_16822,N_16868);
and U21684 (N_21684,N_18172,N_19466);
and U21685 (N_21685,N_16607,N_16771);
nand U21686 (N_21686,N_19979,N_19429);
nand U21687 (N_21687,N_16422,N_17856);
nand U21688 (N_21688,N_16219,N_19260);
xor U21689 (N_21689,N_15546,N_19480);
nand U21690 (N_21690,N_16550,N_18568);
xor U21691 (N_21691,N_16313,N_18767);
nor U21692 (N_21692,N_16797,N_16250);
nor U21693 (N_21693,N_19804,N_17018);
or U21694 (N_21694,N_16494,N_15863);
nand U21695 (N_21695,N_18065,N_19904);
or U21696 (N_21696,N_15548,N_18125);
xor U21697 (N_21697,N_17418,N_16184);
or U21698 (N_21698,N_16372,N_19498);
xor U21699 (N_21699,N_17224,N_16939);
nand U21700 (N_21700,N_19123,N_15584);
nand U21701 (N_21701,N_16156,N_17733);
xnor U21702 (N_21702,N_15452,N_15131);
xnor U21703 (N_21703,N_15777,N_18695);
or U21704 (N_21704,N_15530,N_19116);
xnor U21705 (N_21705,N_19883,N_19856);
and U21706 (N_21706,N_19515,N_19241);
nor U21707 (N_21707,N_16826,N_19950);
xor U21708 (N_21708,N_16348,N_18969);
and U21709 (N_21709,N_19381,N_19380);
and U21710 (N_21710,N_16117,N_17155);
nor U21711 (N_21711,N_17218,N_17859);
or U21712 (N_21712,N_16487,N_17136);
nor U21713 (N_21713,N_17797,N_18827);
and U21714 (N_21714,N_17328,N_17354);
or U21715 (N_21715,N_16726,N_17644);
nor U21716 (N_21716,N_15826,N_16228);
nand U21717 (N_21717,N_17670,N_15083);
nand U21718 (N_21718,N_16068,N_19916);
or U21719 (N_21719,N_19185,N_16281);
nor U21720 (N_21720,N_19730,N_18014);
nand U21721 (N_21721,N_17162,N_16267);
and U21722 (N_21722,N_19568,N_15040);
and U21723 (N_21723,N_17878,N_16992);
xnor U21724 (N_21724,N_15479,N_18748);
and U21725 (N_21725,N_19360,N_18354);
nor U21726 (N_21726,N_16905,N_17361);
nand U21727 (N_21727,N_19960,N_17609);
nand U21728 (N_21728,N_17053,N_17693);
or U21729 (N_21729,N_16684,N_17486);
and U21730 (N_21730,N_19062,N_17813);
nor U21731 (N_21731,N_19675,N_18114);
or U21732 (N_21732,N_15185,N_17448);
or U21733 (N_21733,N_17607,N_15044);
nor U21734 (N_21734,N_16252,N_18746);
and U21735 (N_21735,N_15767,N_15970);
nor U21736 (N_21736,N_19310,N_15410);
nand U21737 (N_21737,N_17983,N_19637);
nand U21738 (N_21738,N_17357,N_18596);
xnor U21739 (N_21739,N_16052,N_18941);
nor U21740 (N_21740,N_19639,N_17880);
and U21741 (N_21741,N_16179,N_16750);
nand U21742 (N_21742,N_15670,N_18883);
and U21743 (N_21743,N_19451,N_16860);
nor U21744 (N_21744,N_16227,N_17060);
nor U21745 (N_21745,N_16997,N_18586);
or U21746 (N_21746,N_17336,N_16230);
and U21747 (N_21747,N_15272,N_18497);
and U21748 (N_21748,N_19530,N_17876);
xnor U21749 (N_21749,N_18868,N_19449);
nor U21750 (N_21750,N_19192,N_17120);
or U21751 (N_21751,N_18546,N_19513);
xnor U21752 (N_21752,N_18977,N_19706);
nand U21753 (N_21753,N_17208,N_19379);
nor U21754 (N_21754,N_18685,N_15588);
and U21755 (N_21755,N_18109,N_18884);
and U21756 (N_21756,N_16839,N_18675);
or U21757 (N_21757,N_16654,N_18887);
xor U21758 (N_21758,N_15236,N_17091);
nand U21759 (N_21759,N_17794,N_18265);
nor U21760 (N_21760,N_17674,N_19707);
and U21761 (N_21761,N_16894,N_18879);
and U21762 (N_21762,N_15944,N_15612);
or U21763 (N_21763,N_19545,N_15681);
nand U21764 (N_21764,N_17335,N_19946);
or U21765 (N_21765,N_19769,N_19494);
or U21766 (N_21766,N_15136,N_18274);
xnor U21767 (N_21767,N_16211,N_16049);
and U21768 (N_21768,N_18608,N_19140);
or U21769 (N_21769,N_19215,N_18171);
or U21770 (N_21770,N_17243,N_17471);
xnor U21771 (N_21771,N_19372,N_18636);
xor U21772 (N_21772,N_15368,N_17695);
or U21773 (N_21773,N_16908,N_15360);
and U21774 (N_21774,N_18016,N_16666);
xor U21775 (N_21775,N_18512,N_16340);
nand U21776 (N_21776,N_19558,N_15969);
nand U21777 (N_21777,N_16134,N_18214);
nand U21778 (N_21778,N_16127,N_18913);
xor U21779 (N_21779,N_15817,N_15912);
and U21780 (N_21780,N_15789,N_17618);
or U21781 (N_21781,N_15009,N_18353);
xnor U21782 (N_21782,N_15361,N_18143);
nor U21783 (N_21783,N_18629,N_18456);
xor U21784 (N_21784,N_15169,N_15667);
nand U21785 (N_21785,N_19898,N_19929);
and U21786 (N_21786,N_16162,N_19169);
or U21787 (N_21787,N_19250,N_16945);
nand U21788 (N_21788,N_17315,N_17857);
xnor U21789 (N_21789,N_16533,N_18869);
nand U21790 (N_21790,N_16100,N_16261);
and U21791 (N_21791,N_18628,N_15378);
nor U21792 (N_21792,N_16436,N_16405);
xor U21793 (N_21793,N_16278,N_16237);
nand U21794 (N_21794,N_15806,N_16862);
xor U21795 (N_21795,N_17514,N_16236);
xnor U21796 (N_21796,N_16698,N_16154);
xor U21797 (N_21797,N_16983,N_17603);
nand U21798 (N_21798,N_17458,N_18070);
nor U21799 (N_21799,N_15592,N_19582);
nor U21800 (N_21800,N_17371,N_15251);
nand U21801 (N_21801,N_19871,N_18543);
and U21802 (N_21802,N_16556,N_16695);
xor U21803 (N_21803,N_18482,N_16628);
nor U21804 (N_21804,N_15677,N_16819);
nand U21805 (N_21805,N_18648,N_18890);
nand U21806 (N_21806,N_17468,N_19901);
nand U21807 (N_21807,N_18498,N_17915);
or U21808 (N_21808,N_15977,N_18085);
nand U21809 (N_21809,N_16682,N_17033);
and U21810 (N_21810,N_19805,N_19387);
nor U21811 (N_21811,N_19948,N_16991);
nor U21812 (N_21812,N_18433,N_17858);
nand U21813 (N_21813,N_15984,N_15053);
nor U21814 (N_21814,N_19052,N_17225);
or U21815 (N_21815,N_16234,N_17512);
or U21816 (N_21816,N_18606,N_19370);
and U21817 (N_21817,N_16269,N_17119);
nor U21818 (N_21818,N_19766,N_15434);
nor U21819 (N_21819,N_15455,N_18992);
and U21820 (N_21820,N_18054,N_17538);
and U21821 (N_21821,N_19093,N_19321);
or U21822 (N_21822,N_19385,N_16394);
nor U21823 (N_21823,N_17158,N_19085);
nor U21824 (N_21824,N_18486,N_18815);
and U21825 (N_21825,N_19606,N_19642);
xor U21826 (N_21826,N_19807,N_17316);
or U21827 (N_21827,N_18781,N_19489);
xor U21828 (N_21828,N_16833,N_15776);
nor U21829 (N_21829,N_15640,N_19268);
nand U21830 (N_21830,N_16711,N_15257);
and U21831 (N_21831,N_17322,N_15199);
nand U21832 (N_21832,N_15079,N_16199);
or U21833 (N_21833,N_19275,N_17474);
and U21834 (N_21834,N_16107,N_19666);
or U21835 (N_21835,N_17811,N_19301);
nor U21836 (N_21836,N_17569,N_17430);
or U21837 (N_21837,N_19894,N_18449);
nand U21838 (N_21838,N_18232,N_18352);
or U21839 (N_21839,N_17761,N_18224);
nor U21840 (N_21840,N_15973,N_16490);
nor U21841 (N_21841,N_18443,N_15331);
or U21842 (N_21842,N_15997,N_15615);
xor U21843 (N_21843,N_15213,N_18915);
nand U21844 (N_21844,N_18135,N_15533);
xnor U21845 (N_21845,N_15519,N_16856);
xor U21846 (N_21846,N_18306,N_17381);
or U21847 (N_21847,N_16555,N_18731);
xnor U21848 (N_21848,N_16691,N_16424);
and U21849 (N_21849,N_17523,N_18505);
and U21850 (N_21850,N_17129,N_18978);
nand U21851 (N_21851,N_18681,N_16157);
or U21852 (N_21852,N_15925,N_15398);
and U21853 (N_21853,N_18103,N_16355);
xor U21854 (N_21854,N_18549,N_19228);
and U21855 (N_21855,N_19887,N_17341);
or U21856 (N_21856,N_16393,N_17919);
or U21857 (N_21857,N_15602,N_15012);
xnor U21858 (N_21858,N_15225,N_17457);
nand U21859 (N_21859,N_19958,N_15311);
and U21860 (N_21860,N_18587,N_18851);
or U21861 (N_21861,N_18982,N_19094);
nand U21862 (N_21862,N_17976,N_17405);
and U21863 (N_21863,N_18266,N_18706);
xnor U21864 (N_21864,N_19991,N_19908);
xnor U21865 (N_21865,N_15066,N_16080);
nand U21866 (N_21866,N_16229,N_16921);
or U21867 (N_21867,N_18257,N_17673);
nand U21868 (N_21868,N_15753,N_17396);
and U21869 (N_21869,N_16105,N_17826);
xnor U21870 (N_21870,N_15402,N_15149);
xor U21871 (N_21871,N_18373,N_18909);
and U21872 (N_21872,N_16175,N_17598);
xnor U21873 (N_21873,N_19627,N_16055);
xor U21874 (N_21874,N_16581,N_17171);
and U21875 (N_21875,N_18759,N_15300);
or U21876 (N_21876,N_19118,N_19833);
or U21877 (N_21877,N_16632,N_18231);
xor U21878 (N_21878,N_17769,N_16554);
or U21879 (N_21879,N_18762,N_16499);
and U21880 (N_21880,N_15595,N_15787);
and U21881 (N_21881,N_16823,N_16626);
nor U21882 (N_21882,N_17041,N_19208);
or U21883 (N_21883,N_16194,N_15038);
and U21884 (N_21884,N_15550,N_15164);
nor U21885 (N_21885,N_16957,N_15860);
xnor U21886 (N_21886,N_15369,N_19211);
or U21887 (N_21887,N_19938,N_19745);
and U21888 (N_21888,N_17278,N_16015);
and U21889 (N_21889,N_17967,N_15935);
or U21890 (N_21890,N_19399,N_19051);
or U21891 (N_21891,N_16057,N_18639);
or U21892 (N_21892,N_18376,N_16989);
nand U21893 (N_21893,N_16481,N_15820);
xor U21894 (N_21894,N_17325,N_15298);
xor U21895 (N_21895,N_15121,N_16759);
nor U21896 (N_21896,N_15116,N_19347);
or U21897 (N_21897,N_15722,N_17922);
nand U21898 (N_21898,N_18622,N_16869);
xor U21899 (N_21899,N_18199,N_18521);
or U21900 (N_21900,N_15833,N_19353);
or U21901 (N_21901,N_19044,N_19538);
xor U21902 (N_21902,N_17437,N_18550);
or U21903 (N_21903,N_16451,N_18129);
nor U21904 (N_21904,N_17240,N_19591);
or U21905 (N_21905,N_16811,N_18947);
and U21906 (N_21906,N_15835,N_18136);
and U21907 (N_21907,N_17781,N_15146);
nand U21908 (N_21908,N_17576,N_19317);
or U21909 (N_21909,N_16464,N_16919);
nand U21910 (N_21910,N_16710,N_15993);
xor U21911 (N_21911,N_16415,N_16538);
and U21912 (N_21912,N_15639,N_19230);
xnor U21913 (N_21913,N_15664,N_17877);
nor U21914 (N_21914,N_18472,N_19776);
or U21915 (N_21915,N_18610,N_18619);
nand U21916 (N_21916,N_18424,N_16037);
nor U21917 (N_21917,N_17360,N_19961);
xor U21918 (N_21918,N_15663,N_15279);
nor U21919 (N_21919,N_15374,N_19610);
and U21920 (N_21920,N_19162,N_17942);
xor U21921 (N_21921,N_18946,N_17280);
and U21922 (N_21922,N_15585,N_15874);
nor U21923 (N_21923,N_16518,N_16712);
xnor U21924 (N_21924,N_17084,N_17276);
or U21925 (N_21925,N_15055,N_17483);
or U21926 (N_21926,N_15061,N_17767);
or U21927 (N_21927,N_18405,N_16024);
xnor U21928 (N_21928,N_17764,N_17421);
and U21929 (N_21929,N_18280,N_16192);
or U21930 (N_21930,N_18791,N_19709);
xnor U21931 (N_21931,N_19888,N_15052);
nor U21932 (N_21932,N_15470,N_18804);
xor U21933 (N_21933,N_18948,N_15179);
and U21934 (N_21934,N_17339,N_19174);
xor U21935 (N_21935,N_19156,N_15103);
nand U21936 (N_21936,N_18589,N_15879);
or U21937 (N_21937,N_17944,N_19086);
xor U21938 (N_21938,N_16307,N_18805);
xnor U21939 (N_21939,N_15939,N_16064);
nor U21940 (N_21940,N_17772,N_16871);
and U21941 (N_21941,N_16544,N_17286);
and U21942 (N_21942,N_19125,N_18677);
nor U21943 (N_21943,N_16126,N_15561);
nor U21944 (N_21944,N_19464,N_18657);
or U21945 (N_21945,N_19095,N_15339);
nand U21946 (N_21946,N_17810,N_19284);
nand U21947 (N_21947,N_19187,N_18227);
nand U21948 (N_21948,N_17036,N_18821);
nor U21949 (N_21949,N_15322,N_16463);
xor U21950 (N_21950,N_19855,N_16172);
and U21951 (N_21951,N_19406,N_16789);
nand U21952 (N_21952,N_18364,N_19420);
or U21953 (N_21953,N_19172,N_18774);
and U21954 (N_21954,N_19421,N_15008);
nand U21955 (N_21955,N_16479,N_15743);
nand U21956 (N_21956,N_17176,N_17410);
or U21957 (N_21957,N_18956,N_19598);
or U21958 (N_21958,N_17653,N_17351);
and U21959 (N_21959,N_16953,N_17684);
and U21960 (N_21960,N_17370,N_15882);
xor U21961 (N_21961,N_16867,N_17652);
or U21962 (N_21962,N_15353,N_18682);
nor U21963 (N_21963,N_16740,N_18409);
nor U21964 (N_21964,N_17379,N_18446);
xor U21965 (N_21965,N_15191,N_19900);
xor U21966 (N_21966,N_16294,N_18585);
nand U21967 (N_21967,N_19270,N_16152);
or U21968 (N_21968,N_18499,N_19434);
xor U21969 (N_21969,N_19198,N_19713);
and U21970 (N_21970,N_16086,N_18069);
nand U21971 (N_21971,N_15527,N_15051);
nor U21972 (N_21972,N_19876,N_16614);
and U21973 (N_21973,N_17989,N_17317);
and U21974 (N_21974,N_19537,N_17934);
and U21975 (N_21975,N_16054,N_19069);
or U21976 (N_21976,N_15464,N_19753);
and U21977 (N_21977,N_17917,N_15885);
nor U21978 (N_21978,N_19234,N_18124);
and U21979 (N_21979,N_15192,N_18481);
and U21980 (N_21980,N_15446,N_17961);
xnor U21981 (N_21981,N_19972,N_19566);
xor U21982 (N_21982,N_18822,N_17730);
nand U21983 (N_21983,N_19119,N_16158);
and U21984 (N_21984,N_18689,N_16029);
and U21985 (N_21985,N_17654,N_18989);
xor U21986 (N_21986,N_17031,N_16028);
nor U21987 (N_21987,N_15296,N_19585);
xnor U21988 (N_21988,N_18927,N_19845);
or U21989 (N_21989,N_17294,N_15785);
nor U21990 (N_21990,N_18704,N_16917);
or U21991 (N_21991,N_18638,N_15870);
nor U21992 (N_21992,N_19757,N_17466);
nand U21993 (N_21993,N_18018,N_19571);
and U21994 (N_21994,N_18179,N_18305);
or U21995 (N_21995,N_19712,N_18972);
and U21996 (N_21996,N_16946,N_15646);
nor U21997 (N_21997,N_19968,N_18809);
nor U21998 (N_21998,N_17928,N_19644);
nor U21999 (N_21999,N_17596,N_15953);
nor U22000 (N_22000,N_19102,N_19937);
and U22001 (N_22001,N_16762,N_18738);
and U22002 (N_22002,N_15555,N_15495);
xor U22003 (N_22003,N_19227,N_18765);
or U22004 (N_22004,N_17414,N_19913);
nor U22005 (N_22005,N_18344,N_15909);
xor U22006 (N_22006,N_15631,N_16850);
nor U22007 (N_22007,N_15347,N_16734);
xnor U22008 (N_22008,N_18678,N_18604);
nand U22009 (N_22009,N_17522,N_16395);
nor U22010 (N_22010,N_16452,N_19413);
nor U22011 (N_22011,N_19661,N_17211);
or U22012 (N_22012,N_16849,N_16233);
xor U22013 (N_22013,N_18403,N_17816);
xnor U22014 (N_22014,N_17314,N_18599);
nor U22015 (N_22015,N_16416,N_18291);
or U22016 (N_22016,N_16827,N_19444);
or U22017 (N_22017,N_17691,N_17833);
nand U22018 (N_22018,N_16664,N_18178);
nand U22019 (N_22019,N_15219,N_15752);
xnor U22020 (N_22020,N_19042,N_15685);
nand U22021 (N_22021,N_18442,N_18889);
and U22022 (N_22022,N_18382,N_17309);
xnor U22023 (N_22023,N_15698,N_18535);
xnor U22024 (N_22024,N_17288,N_15095);
nor U22025 (N_22025,N_18367,N_16565);
xor U22026 (N_22026,N_16283,N_16053);
nor U22027 (N_22027,N_18332,N_18705);
and U22028 (N_22028,N_18974,N_15928);
nor U22029 (N_22029,N_19149,N_19083);
or U22030 (N_22030,N_15430,N_17133);
nor U22031 (N_22031,N_17550,N_18771);
or U22032 (N_22032,N_16078,N_17301);
and U22033 (N_22033,N_15505,N_18141);
and U22034 (N_22034,N_19808,N_18671);
and U22035 (N_22035,N_19544,N_15852);
xor U22036 (N_22036,N_17628,N_15273);
nand U22037 (N_22037,N_15618,N_15323);
nor U22038 (N_22038,N_17884,N_19486);
or U22039 (N_22039,N_16118,N_16525);
xor U22040 (N_22040,N_19796,N_15606);
and U22041 (N_22041,N_18718,N_17814);
nand U22042 (N_22042,N_19588,N_19502);
xnor U22043 (N_22043,N_18784,N_17804);
and U22044 (N_22044,N_19309,N_15020);
nand U22045 (N_22045,N_19573,N_19348);
nor U22046 (N_22046,N_15026,N_17202);
or U22047 (N_22047,N_16002,N_19629);
nor U22048 (N_22048,N_16943,N_17475);
nor U22049 (N_22049,N_18701,N_17541);
and U22050 (N_22050,N_18250,N_16428);
nor U22051 (N_22051,N_15214,N_16907);
or U22052 (N_22052,N_17141,N_17456);
xnor U22053 (N_22053,N_19636,N_17842);
nand U22054 (N_22054,N_16285,N_19646);
xnor U22055 (N_22055,N_17300,N_15986);
and U22056 (N_22056,N_16636,N_16681);
or U22057 (N_22057,N_17056,N_17265);
nor U22058 (N_22058,N_15070,N_17204);
or U22059 (N_22059,N_16493,N_18342);
and U22060 (N_22060,N_17637,N_15896);
nand U22061 (N_22061,N_18876,N_18853);
nand U22062 (N_22062,N_15403,N_15700);
xnor U22063 (N_22063,N_16142,N_19337);
nand U22064 (N_22064,N_18570,N_17401);
and U22065 (N_22065,N_19493,N_19126);
or U22066 (N_22066,N_16448,N_18623);
nor U22067 (N_22067,N_19481,N_18002);
nand U22068 (N_22068,N_16642,N_17067);
or U22069 (N_22069,N_19829,N_18811);
or U22070 (N_22070,N_19879,N_17517);
and U22071 (N_22071,N_18371,N_17428);
nand U22072 (N_22072,N_19791,N_16659);
and U22073 (N_22073,N_19465,N_16892);
xor U22074 (N_22074,N_15917,N_15022);
nor U22075 (N_22075,N_19822,N_15513);
nor U22076 (N_22076,N_18169,N_19659);
nand U22077 (N_22077,N_18523,N_16025);
xnor U22078 (N_22078,N_15075,N_15686);
nor U22079 (N_22079,N_16773,N_15747);
or U22080 (N_22080,N_15922,N_18999);
and U22081 (N_22081,N_15799,N_19045);
xnor U22082 (N_22082,N_17718,N_15657);
xor U22083 (N_22083,N_18081,N_17985);
xnor U22084 (N_22084,N_18611,N_16936);
nor U22085 (N_22085,N_16203,N_16043);
and U22086 (N_22086,N_18739,N_17722);
xnor U22087 (N_22087,N_17253,N_15516);
xor U22088 (N_22088,N_15108,N_16271);
nand U22089 (N_22089,N_19292,N_18005);
and U22090 (N_22090,N_18269,N_18503);
nand U22091 (N_22091,N_17473,N_15429);
nand U22092 (N_22092,N_17222,N_15428);
or U22093 (N_22093,N_18480,N_16714);
or U22094 (N_22094,N_18223,N_15683);
or U22095 (N_22095,N_19772,N_15423);
xnor U22096 (N_22096,N_15216,N_15485);
or U22097 (N_22097,N_18299,N_16705);
xor U22098 (N_22098,N_17114,N_18072);
or U22099 (N_22099,N_16385,N_16830);
xnor U22100 (N_22100,N_15940,N_19147);
nor U22101 (N_22101,N_16717,N_18309);
xnor U22102 (N_22102,N_18183,N_16260);
or U22103 (N_22103,N_17940,N_16300);
or U22104 (N_22104,N_16709,N_19247);
nand U22105 (N_22105,N_19881,N_18445);
nor U22106 (N_22106,N_19831,N_18864);
and U22107 (N_22107,N_15160,N_15385);
xnor U22108 (N_22108,N_18236,N_17927);
and U22109 (N_22109,N_15384,N_17022);
nand U22110 (N_22110,N_18957,N_18859);
nand U22111 (N_22111,N_16637,N_18145);
nor U22112 (N_22112,N_15301,N_16621);
or U22113 (N_22113,N_15647,N_19754);
xnor U22114 (N_22114,N_17409,N_16521);
and U22115 (N_22115,N_18174,N_17462);
xnor U22116 (N_22116,N_18485,N_16526);
and U22117 (N_22117,N_17916,N_15277);
nand U22118 (N_22118,N_16597,N_19654);
nor U22119 (N_22119,N_18721,N_18004);
nand U22120 (N_22120,N_15142,N_15056);
nor U22121 (N_22121,N_17586,N_17525);
or U22122 (N_22122,N_17914,N_16317);
xor U22123 (N_22123,N_15471,N_15941);
nor U22124 (N_22124,N_18402,N_19490);
and U22125 (N_22125,N_15523,N_17882);
and U22126 (N_22126,N_16382,N_19229);
xor U22127 (N_22127,N_17920,N_16824);
and U22128 (N_22128,N_15475,N_19006);
nand U22129 (N_22129,N_16722,N_15152);
or U22130 (N_22130,N_15851,N_16858);
xor U22131 (N_22131,N_16715,N_16496);
or U22132 (N_22132,N_19443,N_15150);
and U22133 (N_22133,N_15742,N_19692);
xor U22134 (N_22134,N_19956,N_17765);
or U22135 (N_22135,N_19857,N_18464);
and U22136 (N_22136,N_19869,N_16362);
or U22137 (N_22137,N_18797,N_18079);
xnor U22138 (N_22138,N_17157,N_18994);
nand U22139 (N_22139,N_17002,N_17387);
nor U22140 (N_22140,N_15712,N_17830);
nor U22141 (N_22141,N_15130,N_16446);
nand U22142 (N_22142,N_18484,N_18146);
nor U22143 (N_22143,N_19723,N_18032);
xnor U22144 (N_22144,N_18462,N_19436);
and U22145 (N_22145,N_16231,N_17633);
or U22146 (N_22146,N_18643,N_17777);
nand U22147 (N_22147,N_15574,N_17808);
xnor U22148 (N_22148,N_15783,N_17592);
and U22149 (N_22149,N_17570,N_19440);
nand U22150 (N_22150,N_16035,N_16978);
nor U22151 (N_22151,N_17135,N_19035);
or U22152 (N_22152,N_15837,N_16857);
or U22153 (N_22153,N_19214,N_19635);
nand U22154 (N_22154,N_15125,N_16728);
nand U22155 (N_22155,N_15598,N_17815);
xnor U22156 (N_22156,N_17110,N_17891);
xor U22157 (N_22157,N_18187,N_15965);
nor U22158 (N_22158,N_19339,N_17921);
or U22159 (N_22159,N_15412,N_19510);
nand U22160 (N_22160,N_17195,N_18298);
and U22161 (N_22161,N_19079,N_15892);
xor U22162 (N_22162,N_16703,N_15864);
and U22163 (N_22163,N_17492,N_15704);
or U22164 (N_22164,N_18096,N_18526);
nand U22165 (N_22165,N_16318,N_17363);
xor U22166 (N_22166,N_18345,N_18865);
xor U22167 (N_22167,N_16852,N_15228);
nand U22168 (N_22168,N_17163,N_16006);
nand U22169 (N_22169,N_15936,N_17150);
or U22170 (N_22170,N_15004,N_18713);
nand U22171 (N_22171,N_18751,N_15328);
and U22172 (N_22172,N_15760,N_16462);
or U22173 (N_22173,N_15735,N_15930);
xnor U22174 (N_22174,N_18855,N_15506);
nor U22175 (N_22175,N_16391,N_18874);
nand U22176 (N_22176,N_17947,N_18095);
nand U22177 (N_22177,N_16119,N_19815);
xor U22178 (N_22178,N_19863,N_15791);
nor U22179 (N_22179,N_19142,N_17329);
or U22180 (N_22180,N_15477,N_17030);
nor U22181 (N_22181,N_17521,N_18452);
nand U22182 (N_22182,N_16941,N_16089);
nand U22183 (N_22183,N_17152,N_16906);
or U22184 (N_22184,N_15853,N_17128);
xor U22185 (N_22185,N_16031,N_15376);
xor U22186 (N_22186,N_19433,N_19196);
nor U22187 (N_22187,N_17894,N_19978);
nand U22188 (N_22188,N_19312,N_17012);
nor U22189 (N_22189,N_18051,N_19277);
or U22190 (N_22190,N_19770,N_15217);
nand U22191 (N_22191,N_16081,N_18522);
xor U22192 (N_22192,N_15808,N_15096);
or U22193 (N_22193,N_16491,N_15107);
or U22194 (N_22194,N_18647,N_15484);
nand U22195 (N_22195,N_19783,N_19525);
nor U22196 (N_22196,N_16297,N_19572);
nand U22197 (N_22197,N_17029,N_18950);
nand U22198 (N_22198,N_16752,N_15655);
nor U22199 (N_22199,N_18939,N_16647);
nor U22200 (N_22200,N_18039,N_17279);
and U22201 (N_22201,N_18312,N_18254);
or U22202 (N_22202,N_17503,N_16414);
nor U22203 (N_22203,N_18492,N_18053);
xnor U22204 (N_22204,N_17701,N_19765);
nand U22205 (N_22205,N_15345,N_15139);
or U22206 (N_22206,N_15975,N_18323);
or U22207 (N_22207,N_16562,N_17099);
nand U22208 (N_22208,N_19877,N_19050);
nor U22209 (N_22209,N_18949,N_18127);
xor U22210 (N_22210,N_19193,N_16510);
xnor U22211 (N_22211,N_15389,N_15594);
xor U22212 (N_22212,N_19886,N_18789);
and U22213 (N_22213,N_16600,N_18324);
nor U22214 (N_22214,N_15721,N_19065);
nor U22215 (N_22215,N_18396,N_17906);
nand U22216 (N_22216,N_17560,N_19210);
or U22217 (N_22217,N_18653,N_19207);
or U22218 (N_22218,N_17219,N_17116);
xnor U22219 (N_22219,N_16263,N_17046);
nand U22220 (N_22220,N_17057,N_16704);
and U22221 (N_22221,N_15915,N_17241);
nor U22222 (N_22222,N_19203,N_15750);
xor U22223 (N_22223,N_16380,N_17687);
and U22224 (N_22224,N_19130,N_19740);
and U22225 (N_22225,N_15163,N_16413);
and U22226 (N_22226,N_18690,N_17235);
xor U22227 (N_22227,N_18162,N_16504);
or U22228 (N_22228,N_19693,N_19462);
and U22229 (N_22229,N_15036,N_15409);
xor U22230 (N_22230,N_16745,N_15439);
xor U22231 (N_22231,N_17712,N_18357);
nand U22232 (N_22232,N_19287,N_16277);
or U22233 (N_22233,N_17605,N_17170);
and U22234 (N_22234,N_15510,N_17065);
xnor U22235 (N_22235,N_17454,N_16886);
nor U22236 (N_22236,N_19534,N_19514);
and U22237 (N_22237,N_19340,N_16609);
nand U22238 (N_22238,N_19676,N_19896);
xnor U22239 (N_22239,N_19825,N_17982);
nor U22240 (N_22240,N_19327,N_17530);
nand U22241 (N_22241,N_17647,N_17244);
xnor U22242 (N_22242,N_17330,N_15858);
xnor U22243 (N_22243,N_15372,N_18975);
or U22244 (N_22244,N_17137,N_17905);
nor U22245 (N_22245,N_17557,N_16928);
nand U22246 (N_22246,N_15422,N_16602);
or U22247 (N_22247,N_17962,N_17582);
or U22248 (N_22248,N_19350,N_15290);
nand U22249 (N_22249,N_15878,N_15617);
nor U22250 (N_22250,N_15895,N_15060);
or U22251 (N_22251,N_17111,N_15297);
and U22252 (N_22252,N_16845,N_16836);
xor U22253 (N_22253,N_15894,N_16676);
xnor U22254 (N_22254,N_19520,N_18719);
or U22255 (N_22255,N_19424,N_19725);
xnor U22256 (N_22256,N_19143,N_17834);
nor U22257 (N_22257,N_17298,N_17641);
nor U22258 (N_22258,N_16171,N_19540);
and U22259 (N_22259,N_17074,N_15960);
nor U22260 (N_22260,N_17709,N_17069);
nand U22261 (N_22261,N_19111,N_16189);
nand U22262 (N_22262,N_16477,N_19368);
nand U22263 (N_22263,N_18642,N_17567);
nand U22264 (N_22264,N_17272,N_15117);
xor U22265 (N_22265,N_19408,N_18814);
or U22266 (N_22266,N_19971,N_18218);
nand U22267 (N_22267,N_18836,N_18119);
xor U22268 (N_22268,N_16612,N_16754);
and U22269 (N_22269,N_16545,N_17287);
or U22270 (N_22270,N_15158,N_18796);
and U22271 (N_22271,N_15828,N_19649);
or U22272 (N_22272,N_19592,N_15171);
xor U22273 (N_22273,N_17909,N_16070);
and U22274 (N_22274,N_15366,N_16766);
nand U22275 (N_22275,N_17853,N_15710);
and U22276 (N_22276,N_17881,N_15404);
or U22277 (N_22277,N_19702,N_18107);
or U22278 (N_22278,N_19176,N_17518);
nand U22279 (N_22279,N_15113,N_15679);
or U22280 (N_22280,N_17443,N_16061);
nor U22281 (N_22281,N_18832,N_18193);
nand U22282 (N_22282,N_18645,N_19797);
nand U22283 (N_22283,N_17593,N_16918);
and U22284 (N_22284,N_16258,N_16864);
or U22285 (N_22285,N_17388,N_18925);
and U22286 (N_22286,N_17893,N_15898);
nor U22287 (N_22287,N_19918,N_16112);
or U22288 (N_22288,N_19390,N_18687);
nor U22289 (N_22289,N_18658,N_17221);
nand U22290 (N_22290,N_15807,N_16322);
nand U22291 (N_22291,N_19401,N_17089);
nor U22292 (N_22292,N_16431,N_15397);
and U22293 (N_22293,N_18825,N_18201);
or U22294 (N_22294,N_19012,N_16579);
xnor U22295 (N_22295,N_18010,N_19257);
xnor U22296 (N_22296,N_18847,N_18386);
nor U22297 (N_22297,N_17366,N_17463);
xor U22298 (N_22298,N_19987,N_16041);
nand U22299 (N_22299,N_19580,N_17890);
or U22300 (N_22300,N_19759,N_19786);
nor U22301 (N_22301,N_19549,N_17612);
and U22302 (N_22302,N_15978,N_19609);
xnor U22303 (N_22303,N_18676,N_15633);
or U22304 (N_22304,N_17261,N_19522);
nor U22305 (N_22305,N_15814,N_18196);
or U22306 (N_22306,N_19507,N_16366);
or U22307 (N_22307,N_17282,N_17383);
and U22308 (N_22308,N_15967,N_18450);
nor U22309 (N_22309,N_18419,N_17395);
or U22310 (N_22310,N_15332,N_19425);
xor U22311 (N_22311,N_19322,N_18365);
nand U22312 (N_22312,N_15186,N_18617);
xnor U22313 (N_22313,N_16814,N_17754);
or U22314 (N_22314,N_18793,N_18905);
nor U22315 (N_22315,N_19190,N_17105);
nand U22316 (N_22316,N_15659,N_19081);
xnor U22317 (N_22317,N_17310,N_18837);
and U22318 (N_22318,N_15123,N_17438);
xnor U22319 (N_22319,N_19332,N_15386);
nand U22320 (N_22320,N_17737,N_19329);
xnor U22321 (N_22321,N_18390,N_19060);
or U22322 (N_22322,N_17978,N_17751);
or U22323 (N_22323,N_19607,N_15963);
xor U22324 (N_22324,N_18984,N_16293);
or U22325 (N_22325,N_18792,N_18756);
nand U22326 (N_22326,N_19222,N_15233);
nor U22327 (N_22327,N_15274,N_19762);
or U22328 (N_22328,N_15183,N_17071);
or U22329 (N_22329,N_15381,N_19734);
nand U22330 (N_22330,N_16197,N_17544);
or U22331 (N_22331,N_15127,N_19068);
or U22332 (N_22332,N_19122,N_16195);
xor U22333 (N_22333,N_15270,N_19672);
or U22334 (N_22334,N_18361,N_16320);
nand U22335 (N_22335,N_16020,N_19023);
nor U22336 (N_22336,N_18366,N_16359);
xor U22337 (N_22337,N_17153,N_16169);
xnor U22338 (N_22338,N_18538,N_16240);
or U22339 (N_22339,N_17169,N_16377);
and U22340 (N_22340,N_16353,N_19801);
xor U22341 (N_22341,N_15254,N_18858);
or U22342 (N_22342,N_18028,N_18444);
xor U22343 (N_22343,N_17981,N_16694);
nand U22344 (N_22344,N_17042,N_15488);
and U22345 (N_22345,N_17964,N_15629);
nor U22346 (N_22346,N_17161,N_19468);
nand U22347 (N_22347,N_16859,N_17015);
or U22348 (N_22348,N_18425,N_18164);
xnor U22349 (N_22349,N_15263,N_16138);
xnor U22350 (N_22350,N_17511,N_17441);
xnor U22351 (N_22351,N_15100,N_17555);
nand U22352 (N_22352,N_15845,N_16668);
nor U22353 (N_22353,N_16290,N_18013);
xnor U22354 (N_22354,N_18530,N_17048);
nand U22355 (N_22355,N_16816,N_19548);
nand U22356 (N_22356,N_16821,N_17885);
xnor U22357 (N_22357,N_19298,N_19800);
xor U22358 (N_22358,N_17516,N_15538);
nand U22359 (N_22359,N_17453,N_19907);
and U22360 (N_22360,N_17436,N_18552);
nand U22361 (N_22361,N_17007,N_18093);
or U22362 (N_22362,N_18528,N_18282);
xor U22363 (N_22363,N_15551,N_15644);
nor U22364 (N_22364,N_17263,N_18632);
xor U22365 (N_22365,N_15632,N_18891);
xnor U22366 (N_22366,N_19467,N_17732);
nor U22367 (N_22367,N_15220,N_15336);
and U22368 (N_22368,N_17621,N_15041);
nand U22369 (N_22369,N_15091,N_18089);
or U22370 (N_22370,N_19656,N_16872);
nand U22371 (N_22371,N_17459,N_19846);
nand U22372 (N_22372,N_16114,N_17290);
nand U22373 (N_22373,N_16128,N_16066);
or U22374 (N_22374,N_16276,N_19113);
or U22375 (N_22375,N_19362,N_18621);
or U22376 (N_22376,N_16287,N_16363);
or U22377 (N_22377,N_19986,N_18652);
xnor U22378 (N_22378,N_17072,N_18961);
or U22379 (N_22379,N_18239,N_15184);
or U22380 (N_22380,N_16890,N_16365);
nand U22381 (N_22381,N_15098,N_19503);
xnor U22382 (N_22382,N_15309,N_16159);
nand U22383 (N_22383,N_16275,N_18229);
nor U22384 (N_22384,N_18115,N_16732);
nand U22385 (N_22385,N_18934,N_15335);
nand U22386 (N_22386,N_18034,N_15749);
xor U22387 (N_22387,N_17669,N_17791);
or U22388 (N_22388,N_17427,N_15744);
xnor U22389 (N_22389,N_19516,N_17508);
xor U22390 (N_22390,N_15120,N_16266);
xnor U22391 (N_22391,N_15847,N_16469);
nor U22392 (N_22392,N_17064,N_18106);
or U22393 (N_22393,N_18848,N_15830);
xor U22394 (N_22394,N_15804,N_16136);
and U22395 (N_22395,N_18207,N_19785);
xnor U22396 (N_22396,N_18708,N_18019);
and U22397 (N_22397,N_16034,N_15054);
nand U22398 (N_22398,N_18432,N_16942);
and U22399 (N_22399,N_17869,N_19262);
or U22400 (N_22400,N_19719,N_17723);
and U22401 (N_22401,N_18140,N_17293);
nor U22402 (N_22402,N_16215,N_19245);
or U22403 (N_22403,N_15138,N_15326);
xnor U22404 (N_22404,N_16371,N_15674);
nor U22405 (N_22405,N_17345,N_17269);
nand U22406 (N_22406,N_19059,N_18907);
nand U22407 (N_22407,N_18024,N_16284);
xor U22408 (N_22408,N_16781,N_18176);
or U22409 (N_22409,N_17832,N_18468);
or U22410 (N_22410,N_19731,N_15762);
nor U22411 (N_22411,N_18515,N_16235);
xnor U22412 (N_22412,N_17107,N_19779);
and U22413 (N_22413,N_15705,N_18964);
xnor U22414 (N_22414,N_19565,N_16311);
nand U22415 (N_22415,N_18335,N_16129);
nand U22416 (N_22416,N_17164,N_18082);
and U22417 (N_22417,N_19657,N_15803);
or U22418 (N_22418,N_16033,N_16985);
nor U22419 (N_22419,N_15074,N_15448);
nor U22420 (N_22420,N_16457,N_19166);
nand U22421 (N_22421,N_18422,N_15741);
or U22422 (N_22422,N_18693,N_18578);
nand U22423 (N_22423,N_18175,N_18233);
nand U22424 (N_22424,N_19992,N_18200);
and U22425 (N_22425,N_16094,N_15459);
nor U22426 (N_22426,N_16507,N_17302);
nand U22427 (N_22427,N_18111,N_17393);
xnor U22428 (N_22428,N_16310,N_18156);
nand U22429 (N_22429,N_17619,N_19141);
and U22430 (N_22430,N_16480,N_16625);
nor U22431 (N_22431,N_19124,N_18998);
nor U22432 (N_22432,N_19107,N_16590);
and U22433 (N_22433,N_16108,N_16675);
and U22434 (N_22434,N_15101,N_18314);
and U22435 (N_22435,N_17735,N_18995);
and U22436 (N_22436,N_15759,N_18702);
or U22437 (N_22437,N_19459,N_17000);
nand U22438 (N_22438,N_17066,N_17789);
nor U22439 (N_22439,N_16435,N_19874);
nor U22440 (N_22440,N_18226,N_18258);
and U22441 (N_22441,N_16866,N_15178);
nor U22442 (N_22442,N_17911,N_15281);
or U22443 (N_22443,N_18467,N_17242);
or U22444 (N_22444,N_19183,N_17862);
and U22445 (N_22445,N_18384,N_15866);
nand U22446 (N_22446,N_17824,N_19751);
or U22447 (N_22447,N_19349,N_16360);
nor U22448 (N_22448,N_15501,N_18951);
nor U22449 (N_22449,N_17173,N_19984);
nor U22450 (N_22450,N_19120,N_17103);
nor U22451 (N_22451,N_18674,N_17800);
nand U22452 (N_22452,N_15778,N_19365);
nor U22453 (N_22453,N_15203,N_15077);
or U22454 (N_22454,N_17189,N_15793);
xor U22455 (N_22455,N_19616,N_17168);
xnor U22456 (N_22456,N_19998,N_16303);
xnor U22457 (N_22457,N_15734,N_19674);
and U22458 (N_22458,N_18634,N_16966);
or U22459 (N_22459,N_16815,N_16575);
and U22460 (N_22460,N_15497,N_17758);
and U22461 (N_22461,N_19597,N_17773);
nor U22462 (N_22462,N_18387,N_15818);
and U22463 (N_22463,N_16522,N_15880);
xor U22464 (N_22464,N_19043,N_19500);
and U22465 (N_22465,N_15855,N_16509);
nor U22466 (N_22466,N_16721,N_19285);
nand U22467 (N_22467,N_15955,N_18020);
or U22468 (N_22468,N_17108,N_18603);
and U22469 (N_22469,N_19718,N_15287);
or U22470 (N_22470,N_15809,N_17230);
and U22471 (N_22471,N_16264,N_15995);
or U22472 (N_22472,N_18375,N_16217);
xnor U22473 (N_22473,N_17850,N_18921);
or U22474 (N_22474,N_15688,N_18241);
or U22475 (N_22475,N_18547,N_19289);
nor U22476 (N_22476,N_19438,N_16286);
or U22477 (N_22477,N_18209,N_18240);
xnor U22478 (N_22478,N_16292,N_17600);
and U22479 (N_22479,N_16993,N_16947);
xor U22480 (N_22480,N_15567,N_16755);
nor U22481 (N_22481,N_15599,N_16559);
or U22482 (N_22482,N_15379,N_16888);
nor U22483 (N_22483,N_16967,N_18304);
and U22484 (N_22484,N_18186,N_19623);
nand U22485 (N_22485,N_15956,N_15180);
and U22486 (N_22486,N_18777,N_18555);
xor U22487 (N_22487,N_16896,N_15147);
nor U22488 (N_22488,N_18308,N_16924);
nor U22489 (N_22489,N_16071,N_15605);
xor U22490 (N_22490,N_18945,N_19136);
nor U22491 (N_22491,N_16421,N_17611);
xor U22492 (N_22492,N_17848,N_19602);
nand U22493 (N_22493,N_16885,N_18261);
nor U22494 (N_22494,N_19439,N_18770);
or U22495 (N_22495,N_18453,N_15680);
or U22496 (N_22496,N_19844,N_17079);
or U22497 (N_22497,N_16356,N_15084);
nor U22498 (N_22498,N_17785,N_19848);
or U22499 (N_22499,N_18131,N_15268);
and U22500 (N_22500,N_19913,N_16873);
xnor U22501 (N_22501,N_18166,N_18930);
or U22502 (N_22502,N_16525,N_16446);
nor U22503 (N_22503,N_18893,N_17649);
nand U22504 (N_22504,N_15623,N_17634);
and U22505 (N_22505,N_15446,N_15254);
or U22506 (N_22506,N_18856,N_15070);
or U22507 (N_22507,N_15489,N_17029);
or U22508 (N_22508,N_17185,N_17912);
nand U22509 (N_22509,N_15932,N_17665);
nand U22510 (N_22510,N_19957,N_19997);
xor U22511 (N_22511,N_15181,N_16112);
and U22512 (N_22512,N_15672,N_18261);
or U22513 (N_22513,N_19023,N_19809);
nand U22514 (N_22514,N_17272,N_17671);
xnor U22515 (N_22515,N_18310,N_18359);
xnor U22516 (N_22516,N_15720,N_16406);
nor U22517 (N_22517,N_16652,N_16023);
xor U22518 (N_22518,N_18544,N_19708);
nand U22519 (N_22519,N_16677,N_16546);
nor U22520 (N_22520,N_18349,N_19612);
xnor U22521 (N_22521,N_16254,N_19455);
xor U22522 (N_22522,N_17866,N_19319);
nor U22523 (N_22523,N_15202,N_15432);
nand U22524 (N_22524,N_16626,N_15223);
nor U22525 (N_22525,N_19973,N_19201);
xor U22526 (N_22526,N_19264,N_15148);
nor U22527 (N_22527,N_19154,N_19991);
or U22528 (N_22528,N_19857,N_16263);
or U22529 (N_22529,N_15128,N_18436);
xnor U22530 (N_22530,N_18859,N_18756);
nor U22531 (N_22531,N_19937,N_15919);
xnor U22532 (N_22532,N_18710,N_16353);
xnor U22533 (N_22533,N_18705,N_16250);
xnor U22534 (N_22534,N_16630,N_17792);
nor U22535 (N_22535,N_16401,N_19103);
nor U22536 (N_22536,N_19693,N_19862);
nand U22537 (N_22537,N_15210,N_19474);
and U22538 (N_22538,N_15872,N_18969);
or U22539 (N_22539,N_16206,N_17316);
nor U22540 (N_22540,N_16795,N_17428);
and U22541 (N_22541,N_15377,N_19410);
nor U22542 (N_22542,N_18963,N_16959);
nand U22543 (N_22543,N_15617,N_15336);
nor U22544 (N_22544,N_17463,N_17410);
and U22545 (N_22545,N_19283,N_18695);
xnor U22546 (N_22546,N_17417,N_16417);
or U22547 (N_22547,N_15682,N_17115);
nor U22548 (N_22548,N_18593,N_15485);
nor U22549 (N_22549,N_18816,N_16069);
nor U22550 (N_22550,N_17456,N_19978);
nor U22551 (N_22551,N_15504,N_19981);
nor U22552 (N_22552,N_16152,N_15229);
xnor U22553 (N_22553,N_16855,N_15311);
or U22554 (N_22554,N_19952,N_15341);
or U22555 (N_22555,N_15803,N_15677);
nor U22556 (N_22556,N_18291,N_18301);
or U22557 (N_22557,N_18708,N_18173);
and U22558 (N_22558,N_18424,N_19332);
nand U22559 (N_22559,N_19020,N_16244);
and U22560 (N_22560,N_18822,N_19558);
nand U22561 (N_22561,N_16922,N_18015);
and U22562 (N_22562,N_17037,N_15484);
nand U22563 (N_22563,N_19577,N_16133);
nand U22564 (N_22564,N_19428,N_17644);
nand U22565 (N_22565,N_18279,N_19901);
or U22566 (N_22566,N_15365,N_19148);
nor U22567 (N_22567,N_16776,N_15543);
nor U22568 (N_22568,N_16191,N_19175);
or U22569 (N_22569,N_17967,N_16682);
nand U22570 (N_22570,N_18705,N_15260);
xnor U22571 (N_22571,N_19831,N_16450);
or U22572 (N_22572,N_17488,N_19603);
nand U22573 (N_22573,N_16321,N_18640);
or U22574 (N_22574,N_16874,N_16984);
and U22575 (N_22575,N_18613,N_17381);
nor U22576 (N_22576,N_17280,N_15320);
nor U22577 (N_22577,N_19588,N_18796);
xnor U22578 (N_22578,N_19383,N_15810);
nand U22579 (N_22579,N_18520,N_17390);
nor U22580 (N_22580,N_19879,N_19276);
nand U22581 (N_22581,N_19050,N_16560);
and U22582 (N_22582,N_15769,N_19093);
or U22583 (N_22583,N_18540,N_15507);
xnor U22584 (N_22584,N_18526,N_16967);
xnor U22585 (N_22585,N_18763,N_18228);
or U22586 (N_22586,N_18844,N_17806);
nor U22587 (N_22587,N_17193,N_18703);
or U22588 (N_22588,N_19914,N_15844);
xnor U22589 (N_22589,N_17455,N_15858);
or U22590 (N_22590,N_15688,N_16335);
xnor U22591 (N_22591,N_16870,N_17743);
xnor U22592 (N_22592,N_16186,N_15023);
or U22593 (N_22593,N_18788,N_19882);
nor U22594 (N_22594,N_15834,N_17474);
xor U22595 (N_22595,N_17849,N_17208);
xnor U22596 (N_22596,N_17142,N_19151);
or U22597 (N_22597,N_17208,N_18181);
nor U22598 (N_22598,N_18307,N_15489);
nor U22599 (N_22599,N_17267,N_16579);
or U22600 (N_22600,N_17188,N_16178);
xor U22601 (N_22601,N_18958,N_19095);
nor U22602 (N_22602,N_18521,N_18046);
and U22603 (N_22603,N_17753,N_17560);
nor U22604 (N_22604,N_18499,N_15699);
or U22605 (N_22605,N_19047,N_15796);
and U22606 (N_22606,N_17966,N_15930);
and U22607 (N_22607,N_18002,N_19220);
and U22608 (N_22608,N_15747,N_19951);
nand U22609 (N_22609,N_18435,N_18001);
or U22610 (N_22610,N_19147,N_19307);
xor U22611 (N_22611,N_18364,N_16347);
xnor U22612 (N_22612,N_17629,N_15214);
and U22613 (N_22613,N_16354,N_18772);
xnor U22614 (N_22614,N_15963,N_17564);
and U22615 (N_22615,N_15295,N_16252);
nand U22616 (N_22616,N_19272,N_15832);
xnor U22617 (N_22617,N_18147,N_17563);
nor U22618 (N_22618,N_17205,N_18888);
nor U22619 (N_22619,N_15252,N_16573);
nor U22620 (N_22620,N_16507,N_19893);
or U22621 (N_22621,N_19021,N_18053);
and U22622 (N_22622,N_19467,N_16261);
nand U22623 (N_22623,N_16953,N_15847);
nor U22624 (N_22624,N_17626,N_18391);
nor U22625 (N_22625,N_19026,N_19625);
and U22626 (N_22626,N_18712,N_17149);
or U22627 (N_22627,N_18243,N_15945);
and U22628 (N_22628,N_15958,N_17656);
or U22629 (N_22629,N_17430,N_16489);
and U22630 (N_22630,N_18259,N_17988);
and U22631 (N_22631,N_16758,N_18332);
and U22632 (N_22632,N_15568,N_19731);
nor U22633 (N_22633,N_19923,N_16661);
nor U22634 (N_22634,N_17801,N_19022);
xnor U22635 (N_22635,N_18672,N_15912);
and U22636 (N_22636,N_15854,N_19963);
nand U22637 (N_22637,N_18473,N_18334);
nand U22638 (N_22638,N_16687,N_18197);
or U22639 (N_22639,N_19149,N_15975);
and U22640 (N_22640,N_15420,N_15996);
xnor U22641 (N_22641,N_18787,N_15508);
nor U22642 (N_22642,N_15086,N_17163);
nor U22643 (N_22643,N_18719,N_15389);
or U22644 (N_22644,N_17580,N_15150);
or U22645 (N_22645,N_15658,N_18333);
or U22646 (N_22646,N_16738,N_15063);
xor U22647 (N_22647,N_17786,N_17084);
and U22648 (N_22648,N_19136,N_16743);
or U22649 (N_22649,N_19680,N_16257);
or U22650 (N_22650,N_18727,N_17582);
nand U22651 (N_22651,N_19386,N_17690);
nand U22652 (N_22652,N_19366,N_19647);
or U22653 (N_22653,N_17193,N_18926);
nor U22654 (N_22654,N_15602,N_19665);
nand U22655 (N_22655,N_18143,N_16358);
or U22656 (N_22656,N_17150,N_19840);
nand U22657 (N_22657,N_17720,N_15133);
nand U22658 (N_22658,N_16813,N_17173);
nand U22659 (N_22659,N_19020,N_19078);
or U22660 (N_22660,N_15575,N_16028);
and U22661 (N_22661,N_15374,N_15254);
and U22662 (N_22662,N_17676,N_18856);
nor U22663 (N_22663,N_19450,N_17022);
nand U22664 (N_22664,N_17535,N_19607);
or U22665 (N_22665,N_17723,N_19544);
nand U22666 (N_22666,N_16555,N_17412);
nand U22667 (N_22667,N_16737,N_18865);
nor U22668 (N_22668,N_15458,N_18044);
or U22669 (N_22669,N_19827,N_16811);
nand U22670 (N_22670,N_19327,N_17195);
nor U22671 (N_22671,N_19399,N_17061);
nor U22672 (N_22672,N_17740,N_17562);
nor U22673 (N_22673,N_16560,N_19394);
xor U22674 (N_22674,N_16807,N_19924);
and U22675 (N_22675,N_15783,N_16388);
and U22676 (N_22676,N_17420,N_17686);
nor U22677 (N_22677,N_18599,N_15603);
nand U22678 (N_22678,N_17476,N_18280);
nand U22679 (N_22679,N_15284,N_18081);
nor U22680 (N_22680,N_18058,N_18855);
xnor U22681 (N_22681,N_15295,N_15111);
xnor U22682 (N_22682,N_18046,N_18808);
nor U22683 (N_22683,N_16173,N_15192);
xnor U22684 (N_22684,N_19698,N_19746);
nand U22685 (N_22685,N_17188,N_15137);
xnor U22686 (N_22686,N_17794,N_18214);
nor U22687 (N_22687,N_17202,N_19116);
or U22688 (N_22688,N_19265,N_19130);
and U22689 (N_22689,N_18161,N_16501);
nor U22690 (N_22690,N_15176,N_15126);
nand U22691 (N_22691,N_15198,N_17795);
and U22692 (N_22692,N_19474,N_16357);
and U22693 (N_22693,N_19855,N_16655);
xor U22694 (N_22694,N_19402,N_19301);
nand U22695 (N_22695,N_18754,N_16063);
and U22696 (N_22696,N_18949,N_17402);
xor U22697 (N_22697,N_16976,N_19250);
and U22698 (N_22698,N_17345,N_15827);
nand U22699 (N_22699,N_15053,N_17001);
and U22700 (N_22700,N_19861,N_18863);
or U22701 (N_22701,N_16890,N_19591);
nor U22702 (N_22702,N_17146,N_18690);
nand U22703 (N_22703,N_19310,N_19957);
and U22704 (N_22704,N_15195,N_15956);
nor U22705 (N_22705,N_16018,N_17595);
xnor U22706 (N_22706,N_15935,N_18995);
nand U22707 (N_22707,N_18524,N_17976);
xnor U22708 (N_22708,N_16837,N_16691);
and U22709 (N_22709,N_15537,N_15361);
xor U22710 (N_22710,N_17174,N_18551);
or U22711 (N_22711,N_18446,N_16053);
and U22712 (N_22712,N_16103,N_17027);
and U22713 (N_22713,N_17239,N_16464);
xor U22714 (N_22714,N_19307,N_19978);
nor U22715 (N_22715,N_17710,N_17137);
nor U22716 (N_22716,N_19031,N_19192);
and U22717 (N_22717,N_16891,N_15302);
or U22718 (N_22718,N_16111,N_18935);
and U22719 (N_22719,N_19023,N_15912);
xor U22720 (N_22720,N_15223,N_15401);
xor U22721 (N_22721,N_15894,N_15446);
and U22722 (N_22722,N_17581,N_15434);
nor U22723 (N_22723,N_16612,N_15636);
and U22724 (N_22724,N_16423,N_15666);
xor U22725 (N_22725,N_18361,N_19502);
and U22726 (N_22726,N_19725,N_17848);
nor U22727 (N_22727,N_15001,N_17620);
or U22728 (N_22728,N_18349,N_15749);
and U22729 (N_22729,N_16436,N_17201);
nor U22730 (N_22730,N_16725,N_15932);
nand U22731 (N_22731,N_15895,N_18945);
xnor U22732 (N_22732,N_19408,N_19622);
nand U22733 (N_22733,N_17673,N_19757);
and U22734 (N_22734,N_19703,N_15666);
nor U22735 (N_22735,N_18186,N_19823);
or U22736 (N_22736,N_17037,N_16295);
nand U22737 (N_22737,N_16653,N_18530);
or U22738 (N_22738,N_16086,N_17591);
nor U22739 (N_22739,N_17500,N_19885);
or U22740 (N_22740,N_16419,N_18484);
and U22741 (N_22741,N_18028,N_15951);
xnor U22742 (N_22742,N_17315,N_18116);
or U22743 (N_22743,N_19123,N_18980);
or U22744 (N_22744,N_19103,N_17583);
nand U22745 (N_22745,N_16314,N_19737);
xor U22746 (N_22746,N_15815,N_15198);
nor U22747 (N_22747,N_16230,N_15048);
nand U22748 (N_22748,N_15531,N_17787);
nor U22749 (N_22749,N_19524,N_19818);
nor U22750 (N_22750,N_16992,N_16351);
nor U22751 (N_22751,N_17812,N_18971);
nand U22752 (N_22752,N_19688,N_15332);
xnor U22753 (N_22753,N_15155,N_19551);
nand U22754 (N_22754,N_17580,N_17539);
or U22755 (N_22755,N_19795,N_18830);
or U22756 (N_22756,N_17945,N_19837);
nand U22757 (N_22757,N_17228,N_15797);
nor U22758 (N_22758,N_19534,N_18174);
xor U22759 (N_22759,N_18258,N_16082);
or U22760 (N_22760,N_17342,N_18934);
and U22761 (N_22761,N_18666,N_15264);
xnor U22762 (N_22762,N_19121,N_15747);
or U22763 (N_22763,N_17300,N_18827);
and U22764 (N_22764,N_19078,N_19110);
nor U22765 (N_22765,N_16866,N_18897);
or U22766 (N_22766,N_16637,N_18282);
or U22767 (N_22767,N_16140,N_16184);
nand U22768 (N_22768,N_16926,N_16513);
nor U22769 (N_22769,N_19822,N_15185);
nor U22770 (N_22770,N_18483,N_18560);
or U22771 (N_22771,N_17443,N_16979);
xnor U22772 (N_22772,N_19274,N_19103);
nor U22773 (N_22773,N_16161,N_15079);
or U22774 (N_22774,N_16402,N_15859);
xnor U22775 (N_22775,N_17964,N_15431);
xor U22776 (N_22776,N_16167,N_18454);
xnor U22777 (N_22777,N_16923,N_19345);
or U22778 (N_22778,N_19069,N_15541);
nor U22779 (N_22779,N_18560,N_16078);
nor U22780 (N_22780,N_16516,N_18252);
nor U22781 (N_22781,N_18131,N_18394);
nor U22782 (N_22782,N_15948,N_18277);
nand U22783 (N_22783,N_19740,N_18620);
or U22784 (N_22784,N_16976,N_15299);
and U22785 (N_22785,N_15994,N_17507);
xnor U22786 (N_22786,N_15737,N_18489);
or U22787 (N_22787,N_19619,N_16390);
nor U22788 (N_22788,N_16351,N_15461);
nand U22789 (N_22789,N_15800,N_19172);
and U22790 (N_22790,N_18598,N_18952);
or U22791 (N_22791,N_16541,N_17437);
nor U22792 (N_22792,N_19806,N_15538);
nand U22793 (N_22793,N_18636,N_15751);
or U22794 (N_22794,N_19926,N_16743);
nor U22795 (N_22795,N_17081,N_16112);
nor U22796 (N_22796,N_15345,N_19798);
nand U22797 (N_22797,N_19388,N_19685);
xor U22798 (N_22798,N_15729,N_19990);
or U22799 (N_22799,N_17196,N_17242);
or U22800 (N_22800,N_17628,N_16095);
nor U22801 (N_22801,N_16302,N_16401);
or U22802 (N_22802,N_16547,N_15387);
nor U22803 (N_22803,N_16653,N_17816);
nor U22804 (N_22804,N_17527,N_19438);
nor U22805 (N_22805,N_18985,N_17216);
and U22806 (N_22806,N_16375,N_16867);
or U22807 (N_22807,N_18637,N_18420);
or U22808 (N_22808,N_16356,N_17063);
or U22809 (N_22809,N_17221,N_15332);
and U22810 (N_22810,N_18174,N_17988);
and U22811 (N_22811,N_17318,N_18856);
nor U22812 (N_22812,N_16362,N_17207);
xnor U22813 (N_22813,N_18460,N_17061);
or U22814 (N_22814,N_16261,N_16909);
xnor U22815 (N_22815,N_16397,N_19649);
xnor U22816 (N_22816,N_15934,N_18396);
xor U22817 (N_22817,N_16460,N_15674);
nand U22818 (N_22818,N_15596,N_15417);
nand U22819 (N_22819,N_18763,N_17506);
xnor U22820 (N_22820,N_18706,N_15296);
xor U22821 (N_22821,N_15016,N_16818);
xnor U22822 (N_22822,N_19940,N_17950);
xnor U22823 (N_22823,N_17919,N_17501);
nand U22824 (N_22824,N_16613,N_19888);
xnor U22825 (N_22825,N_16193,N_19619);
and U22826 (N_22826,N_19747,N_16940);
xnor U22827 (N_22827,N_15129,N_17837);
or U22828 (N_22828,N_18805,N_16327);
and U22829 (N_22829,N_18203,N_16927);
or U22830 (N_22830,N_19961,N_18153);
xnor U22831 (N_22831,N_17042,N_19199);
and U22832 (N_22832,N_19255,N_15120);
xnor U22833 (N_22833,N_18015,N_19369);
nand U22834 (N_22834,N_18553,N_18071);
or U22835 (N_22835,N_18970,N_17124);
nor U22836 (N_22836,N_19134,N_18336);
nand U22837 (N_22837,N_17956,N_15116);
or U22838 (N_22838,N_16898,N_19070);
xnor U22839 (N_22839,N_18384,N_17037);
nand U22840 (N_22840,N_15835,N_18094);
nor U22841 (N_22841,N_15781,N_16340);
nand U22842 (N_22842,N_19358,N_16372);
nand U22843 (N_22843,N_17677,N_19913);
xor U22844 (N_22844,N_19087,N_15378);
xnor U22845 (N_22845,N_15348,N_19866);
and U22846 (N_22846,N_17902,N_16163);
nand U22847 (N_22847,N_18711,N_15495);
nor U22848 (N_22848,N_17065,N_19914);
xor U22849 (N_22849,N_19101,N_16336);
or U22850 (N_22850,N_19440,N_17727);
nand U22851 (N_22851,N_16588,N_16235);
xor U22852 (N_22852,N_19221,N_19205);
xnor U22853 (N_22853,N_18333,N_19390);
or U22854 (N_22854,N_16226,N_17524);
or U22855 (N_22855,N_19699,N_16922);
xor U22856 (N_22856,N_16303,N_17887);
and U22857 (N_22857,N_16586,N_15795);
xor U22858 (N_22858,N_17708,N_15636);
nor U22859 (N_22859,N_17881,N_18378);
or U22860 (N_22860,N_17897,N_17444);
xnor U22861 (N_22861,N_15275,N_19782);
nor U22862 (N_22862,N_18310,N_16606);
nand U22863 (N_22863,N_19385,N_18347);
xnor U22864 (N_22864,N_15524,N_18479);
or U22865 (N_22865,N_18816,N_15685);
or U22866 (N_22866,N_17726,N_17442);
and U22867 (N_22867,N_18358,N_16942);
or U22868 (N_22868,N_17018,N_17107);
and U22869 (N_22869,N_16826,N_17688);
nand U22870 (N_22870,N_18644,N_16206);
xnor U22871 (N_22871,N_15035,N_15109);
and U22872 (N_22872,N_16826,N_18457);
nand U22873 (N_22873,N_18634,N_18901);
and U22874 (N_22874,N_19645,N_19598);
and U22875 (N_22875,N_19506,N_19885);
nand U22876 (N_22876,N_19665,N_18779);
or U22877 (N_22877,N_15255,N_16232);
nor U22878 (N_22878,N_16046,N_18868);
nor U22879 (N_22879,N_19998,N_15192);
or U22880 (N_22880,N_16259,N_18748);
nor U22881 (N_22881,N_18143,N_18712);
nor U22882 (N_22882,N_18266,N_15636);
and U22883 (N_22883,N_18672,N_19062);
nand U22884 (N_22884,N_19774,N_15749);
nand U22885 (N_22885,N_16124,N_16190);
or U22886 (N_22886,N_18019,N_17393);
xor U22887 (N_22887,N_16370,N_18559);
nand U22888 (N_22888,N_19403,N_15411);
nor U22889 (N_22889,N_18582,N_19101);
or U22890 (N_22890,N_17586,N_15284);
and U22891 (N_22891,N_18609,N_17918);
nand U22892 (N_22892,N_19102,N_16786);
or U22893 (N_22893,N_16396,N_16883);
or U22894 (N_22894,N_15966,N_16037);
nor U22895 (N_22895,N_16113,N_17106);
nor U22896 (N_22896,N_18771,N_17220);
nor U22897 (N_22897,N_19788,N_15330);
xor U22898 (N_22898,N_19749,N_18023);
nand U22899 (N_22899,N_17675,N_19174);
nor U22900 (N_22900,N_15554,N_15625);
nand U22901 (N_22901,N_15376,N_17436);
nor U22902 (N_22902,N_17836,N_16299);
nor U22903 (N_22903,N_19746,N_16352);
and U22904 (N_22904,N_17016,N_18563);
nor U22905 (N_22905,N_18551,N_18058);
nand U22906 (N_22906,N_19767,N_18007);
and U22907 (N_22907,N_16382,N_16003);
nor U22908 (N_22908,N_16971,N_18970);
nor U22909 (N_22909,N_18825,N_18556);
nor U22910 (N_22910,N_18041,N_16853);
or U22911 (N_22911,N_16683,N_18950);
or U22912 (N_22912,N_19753,N_19663);
xnor U22913 (N_22913,N_15464,N_16323);
and U22914 (N_22914,N_18277,N_18840);
nor U22915 (N_22915,N_18396,N_17004);
nor U22916 (N_22916,N_16018,N_17350);
nand U22917 (N_22917,N_17091,N_18048);
and U22918 (N_22918,N_19642,N_17101);
nand U22919 (N_22919,N_16842,N_18827);
nand U22920 (N_22920,N_17129,N_19840);
or U22921 (N_22921,N_15301,N_17656);
nor U22922 (N_22922,N_17410,N_16603);
xor U22923 (N_22923,N_19072,N_19684);
and U22924 (N_22924,N_19627,N_16188);
nand U22925 (N_22925,N_18655,N_18936);
and U22926 (N_22926,N_18529,N_15516);
or U22927 (N_22927,N_18836,N_17769);
xnor U22928 (N_22928,N_16192,N_17003);
or U22929 (N_22929,N_16342,N_19769);
and U22930 (N_22930,N_16083,N_16133);
nand U22931 (N_22931,N_16563,N_17661);
and U22932 (N_22932,N_18883,N_19258);
and U22933 (N_22933,N_16819,N_15235);
or U22934 (N_22934,N_17699,N_18066);
nor U22935 (N_22935,N_16406,N_17694);
and U22936 (N_22936,N_17450,N_15720);
xor U22937 (N_22937,N_16743,N_17686);
xor U22938 (N_22938,N_16127,N_18972);
nor U22939 (N_22939,N_15665,N_17474);
nand U22940 (N_22940,N_16792,N_16716);
and U22941 (N_22941,N_16692,N_16928);
nor U22942 (N_22942,N_15849,N_15110);
nand U22943 (N_22943,N_19346,N_19530);
nor U22944 (N_22944,N_19670,N_18871);
xor U22945 (N_22945,N_16675,N_19084);
xnor U22946 (N_22946,N_17175,N_15783);
nor U22947 (N_22947,N_19362,N_19206);
nor U22948 (N_22948,N_16120,N_18978);
xor U22949 (N_22949,N_17888,N_15159);
or U22950 (N_22950,N_19199,N_18950);
xnor U22951 (N_22951,N_17096,N_19217);
nand U22952 (N_22952,N_15808,N_18103);
nand U22953 (N_22953,N_16227,N_16051);
or U22954 (N_22954,N_16646,N_16938);
nand U22955 (N_22955,N_17899,N_15975);
nor U22956 (N_22956,N_18518,N_16745);
xnor U22957 (N_22957,N_19625,N_18007);
xnor U22958 (N_22958,N_18229,N_19897);
or U22959 (N_22959,N_17180,N_19876);
and U22960 (N_22960,N_17106,N_19591);
nand U22961 (N_22961,N_18023,N_16432);
xnor U22962 (N_22962,N_16444,N_18686);
nand U22963 (N_22963,N_18610,N_17664);
or U22964 (N_22964,N_15630,N_18438);
xnor U22965 (N_22965,N_18842,N_16018);
nor U22966 (N_22966,N_16455,N_17938);
xnor U22967 (N_22967,N_17047,N_17099);
or U22968 (N_22968,N_19436,N_15886);
xor U22969 (N_22969,N_18649,N_15946);
and U22970 (N_22970,N_18603,N_15033);
xnor U22971 (N_22971,N_18877,N_15553);
or U22972 (N_22972,N_15887,N_16500);
xor U22973 (N_22973,N_15708,N_19033);
nor U22974 (N_22974,N_17343,N_15168);
or U22975 (N_22975,N_15568,N_18471);
or U22976 (N_22976,N_15172,N_15755);
or U22977 (N_22977,N_17472,N_18570);
and U22978 (N_22978,N_16123,N_15826);
and U22979 (N_22979,N_18623,N_19776);
nand U22980 (N_22980,N_15987,N_15030);
nor U22981 (N_22981,N_15673,N_16457);
or U22982 (N_22982,N_18799,N_15627);
nand U22983 (N_22983,N_19557,N_17035);
nor U22984 (N_22984,N_19224,N_19178);
nand U22985 (N_22985,N_17190,N_17867);
nand U22986 (N_22986,N_15848,N_18256);
nor U22987 (N_22987,N_17829,N_16743);
and U22988 (N_22988,N_18093,N_15970);
or U22989 (N_22989,N_17901,N_17379);
nor U22990 (N_22990,N_18430,N_16002);
or U22991 (N_22991,N_19415,N_17991);
nor U22992 (N_22992,N_17849,N_18133);
and U22993 (N_22993,N_19291,N_19608);
and U22994 (N_22994,N_19530,N_18506);
and U22995 (N_22995,N_18459,N_19160);
nand U22996 (N_22996,N_18360,N_19412);
nand U22997 (N_22997,N_15437,N_19184);
xor U22998 (N_22998,N_16118,N_16911);
nand U22999 (N_22999,N_16082,N_16716);
and U23000 (N_23000,N_19811,N_19491);
nand U23001 (N_23001,N_15126,N_19708);
and U23002 (N_23002,N_17360,N_16457);
or U23003 (N_23003,N_15395,N_18352);
or U23004 (N_23004,N_19944,N_15238);
nor U23005 (N_23005,N_19999,N_16558);
xor U23006 (N_23006,N_19827,N_19602);
nor U23007 (N_23007,N_16509,N_18976);
or U23008 (N_23008,N_19745,N_15352);
and U23009 (N_23009,N_18724,N_15762);
or U23010 (N_23010,N_16944,N_18382);
or U23011 (N_23011,N_18751,N_19383);
nor U23012 (N_23012,N_16184,N_16625);
nor U23013 (N_23013,N_16387,N_16591);
xnor U23014 (N_23014,N_17039,N_15192);
nor U23015 (N_23015,N_17626,N_17686);
nor U23016 (N_23016,N_15119,N_15637);
nor U23017 (N_23017,N_15781,N_18516);
nor U23018 (N_23018,N_19127,N_19357);
and U23019 (N_23019,N_15464,N_19689);
and U23020 (N_23020,N_16546,N_17945);
nor U23021 (N_23021,N_19789,N_16210);
nand U23022 (N_23022,N_16478,N_15247);
and U23023 (N_23023,N_19247,N_15896);
or U23024 (N_23024,N_18727,N_19898);
nand U23025 (N_23025,N_15762,N_19656);
or U23026 (N_23026,N_15744,N_18732);
xnor U23027 (N_23027,N_17968,N_17576);
nand U23028 (N_23028,N_15401,N_16158);
nor U23029 (N_23029,N_17202,N_15816);
and U23030 (N_23030,N_17290,N_19659);
or U23031 (N_23031,N_17736,N_15308);
or U23032 (N_23032,N_15090,N_15637);
nand U23033 (N_23033,N_18011,N_17326);
nand U23034 (N_23034,N_16667,N_19449);
nor U23035 (N_23035,N_17017,N_16640);
nand U23036 (N_23036,N_15711,N_17439);
and U23037 (N_23037,N_15176,N_15920);
nor U23038 (N_23038,N_19005,N_19821);
xor U23039 (N_23039,N_16391,N_19337);
or U23040 (N_23040,N_15364,N_18586);
or U23041 (N_23041,N_16399,N_19423);
nand U23042 (N_23042,N_18497,N_18991);
or U23043 (N_23043,N_15543,N_17763);
nor U23044 (N_23044,N_16885,N_17678);
nand U23045 (N_23045,N_16720,N_17077);
nor U23046 (N_23046,N_15599,N_19984);
nand U23047 (N_23047,N_15530,N_18168);
nand U23048 (N_23048,N_18095,N_15379);
nand U23049 (N_23049,N_16265,N_18158);
or U23050 (N_23050,N_15085,N_15160);
nand U23051 (N_23051,N_18598,N_16335);
xor U23052 (N_23052,N_19700,N_18981);
or U23053 (N_23053,N_19090,N_19443);
xnor U23054 (N_23054,N_15309,N_15002);
or U23055 (N_23055,N_17745,N_16417);
nor U23056 (N_23056,N_19204,N_19654);
nand U23057 (N_23057,N_19942,N_16841);
nor U23058 (N_23058,N_18963,N_15978);
nand U23059 (N_23059,N_15454,N_16222);
xor U23060 (N_23060,N_17165,N_15553);
nand U23061 (N_23061,N_15326,N_15716);
and U23062 (N_23062,N_19766,N_16420);
xnor U23063 (N_23063,N_19300,N_15956);
nand U23064 (N_23064,N_16099,N_15994);
and U23065 (N_23065,N_18619,N_15526);
nand U23066 (N_23066,N_19755,N_15222);
and U23067 (N_23067,N_15958,N_19328);
and U23068 (N_23068,N_15276,N_16858);
or U23069 (N_23069,N_18981,N_16312);
nor U23070 (N_23070,N_16943,N_15484);
nor U23071 (N_23071,N_15114,N_16042);
nand U23072 (N_23072,N_16591,N_19447);
nand U23073 (N_23073,N_16332,N_15709);
nand U23074 (N_23074,N_19100,N_18412);
or U23075 (N_23075,N_16924,N_16055);
xor U23076 (N_23076,N_17124,N_19070);
or U23077 (N_23077,N_16688,N_16019);
and U23078 (N_23078,N_16268,N_16732);
nor U23079 (N_23079,N_17129,N_19592);
or U23080 (N_23080,N_19283,N_18950);
nor U23081 (N_23081,N_19618,N_15032);
or U23082 (N_23082,N_17039,N_19081);
xnor U23083 (N_23083,N_18801,N_16277);
nand U23084 (N_23084,N_19617,N_15616);
and U23085 (N_23085,N_17045,N_19955);
xor U23086 (N_23086,N_17875,N_17637);
nand U23087 (N_23087,N_15781,N_18309);
or U23088 (N_23088,N_15635,N_16165);
nor U23089 (N_23089,N_16598,N_15631);
nand U23090 (N_23090,N_17125,N_18631);
nand U23091 (N_23091,N_19728,N_19647);
or U23092 (N_23092,N_17160,N_15267);
xor U23093 (N_23093,N_15104,N_19363);
xor U23094 (N_23094,N_19998,N_15044);
xnor U23095 (N_23095,N_18705,N_16775);
nand U23096 (N_23096,N_18804,N_16199);
nand U23097 (N_23097,N_18870,N_18199);
or U23098 (N_23098,N_17012,N_17843);
xor U23099 (N_23099,N_18522,N_16770);
nor U23100 (N_23100,N_15164,N_17941);
nor U23101 (N_23101,N_17364,N_18366);
xnor U23102 (N_23102,N_15586,N_18893);
nor U23103 (N_23103,N_15037,N_15189);
and U23104 (N_23104,N_19631,N_18134);
and U23105 (N_23105,N_19574,N_17560);
and U23106 (N_23106,N_15652,N_15623);
nand U23107 (N_23107,N_19247,N_15860);
or U23108 (N_23108,N_19456,N_15021);
nor U23109 (N_23109,N_18498,N_19528);
nor U23110 (N_23110,N_17115,N_19454);
or U23111 (N_23111,N_18727,N_19188);
nand U23112 (N_23112,N_17674,N_16825);
nor U23113 (N_23113,N_18016,N_18372);
xor U23114 (N_23114,N_15314,N_16385);
or U23115 (N_23115,N_16868,N_15678);
and U23116 (N_23116,N_16755,N_18227);
and U23117 (N_23117,N_18552,N_19064);
xor U23118 (N_23118,N_16804,N_18357);
nand U23119 (N_23119,N_17106,N_15774);
and U23120 (N_23120,N_19384,N_17580);
nor U23121 (N_23121,N_17133,N_15646);
nand U23122 (N_23122,N_17522,N_17185);
nor U23123 (N_23123,N_18143,N_16003);
or U23124 (N_23124,N_16463,N_19281);
xnor U23125 (N_23125,N_18162,N_16930);
xor U23126 (N_23126,N_16286,N_16217);
or U23127 (N_23127,N_17969,N_19364);
nor U23128 (N_23128,N_19811,N_19278);
xor U23129 (N_23129,N_18166,N_17550);
nand U23130 (N_23130,N_18534,N_16502);
and U23131 (N_23131,N_18077,N_15649);
and U23132 (N_23132,N_16663,N_18176);
nand U23133 (N_23133,N_19198,N_17759);
nand U23134 (N_23134,N_17123,N_19914);
xor U23135 (N_23135,N_16502,N_17510);
xor U23136 (N_23136,N_15551,N_16998);
or U23137 (N_23137,N_18579,N_19631);
nor U23138 (N_23138,N_15109,N_17138);
and U23139 (N_23139,N_16999,N_18575);
nor U23140 (N_23140,N_16262,N_18892);
or U23141 (N_23141,N_19759,N_19721);
xor U23142 (N_23142,N_16828,N_18378);
xnor U23143 (N_23143,N_19603,N_16348);
or U23144 (N_23144,N_18985,N_19636);
nor U23145 (N_23145,N_16305,N_19120);
nor U23146 (N_23146,N_15986,N_16145);
nand U23147 (N_23147,N_17954,N_19229);
and U23148 (N_23148,N_19432,N_19252);
xnor U23149 (N_23149,N_17417,N_15681);
or U23150 (N_23150,N_19971,N_18161);
xor U23151 (N_23151,N_17720,N_17526);
nor U23152 (N_23152,N_17070,N_17637);
nand U23153 (N_23153,N_16902,N_19815);
and U23154 (N_23154,N_15135,N_17629);
or U23155 (N_23155,N_15407,N_17687);
or U23156 (N_23156,N_18741,N_18177);
xor U23157 (N_23157,N_16797,N_17999);
nor U23158 (N_23158,N_18126,N_19772);
xor U23159 (N_23159,N_18901,N_18885);
and U23160 (N_23160,N_19438,N_19666);
nor U23161 (N_23161,N_17806,N_15845);
nor U23162 (N_23162,N_16994,N_16535);
nor U23163 (N_23163,N_19875,N_16332);
nor U23164 (N_23164,N_15470,N_15975);
nor U23165 (N_23165,N_18643,N_15795);
and U23166 (N_23166,N_15647,N_15758);
and U23167 (N_23167,N_15966,N_17561);
nor U23168 (N_23168,N_19398,N_17817);
nor U23169 (N_23169,N_16014,N_15107);
or U23170 (N_23170,N_19662,N_17624);
or U23171 (N_23171,N_19884,N_18278);
nand U23172 (N_23172,N_19945,N_16214);
and U23173 (N_23173,N_15505,N_19371);
xor U23174 (N_23174,N_18577,N_19730);
nor U23175 (N_23175,N_15282,N_15322);
and U23176 (N_23176,N_19083,N_16655);
nand U23177 (N_23177,N_17415,N_15963);
nor U23178 (N_23178,N_17698,N_15042);
nand U23179 (N_23179,N_15265,N_15447);
and U23180 (N_23180,N_18138,N_19818);
nor U23181 (N_23181,N_15546,N_15177);
nand U23182 (N_23182,N_16498,N_18011);
or U23183 (N_23183,N_19631,N_19559);
xnor U23184 (N_23184,N_18151,N_16892);
and U23185 (N_23185,N_16427,N_15650);
nand U23186 (N_23186,N_18927,N_15900);
nand U23187 (N_23187,N_16783,N_18481);
xnor U23188 (N_23188,N_18639,N_17348);
nand U23189 (N_23189,N_18483,N_19916);
nand U23190 (N_23190,N_19987,N_19444);
or U23191 (N_23191,N_17937,N_16571);
or U23192 (N_23192,N_19370,N_18646);
xor U23193 (N_23193,N_16957,N_18583);
nor U23194 (N_23194,N_19434,N_17260);
nor U23195 (N_23195,N_16538,N_18432);
or U23196 (N_23196,N_18327,N_19351);
and U23197 (N_23197,N_15285,N_18057);
or U23198 (N_23198,N_19594,N_17743);
nand U23199 (N_23199,N_15646,N_18018);
nor U23200 (N_23200,N_18046,N_19773);
and U23201 (N_23201,N_16946,N_19012);
or U23202 (N_23202,N_16558,N_17270);
nand U23203 (N_23203,N_17671,N_15059);
nand U23204 (N_23204,N_17112,N_18263);
and U23205 (N_23205,N_19535,N_18105);
xor U23206 (N_23206,N_16393,N_18770);
nand U23207 (N_23207,N_17767,N_18508);
nand U23208 (N_23208,N_15594,N_16315);
nor U23209 (N_23209,N_19683,N_17282);
and U23210 (N_23210,N_16248,N_16665);
nor U23211 (N_23211,N_16973,N_18755);
or U23212 (N_23212,N_17578,N_19777);
and U23213 (N_23213,N_16456,N_15055);
and U23214 (N_23214,N_18042,N_17579);
nor U23215 (N_23215,N_19407,N_18306);
nor U23216 (N_23216,N_15841,N_16938);
and U23217 (N_23217,N_15969,N_17134);
xnor U23218 (N_23218,N_15847,N_18410);
nand U23219 (N_23219,N_16720,N_18967);
nand U23220 (N_23220,N_16271,N_18290);
and U23221 (N_23221,N_17187,N_19941);
xnor U23222 (N_23222,N_19147,N_15323);
or U23223 (N_23223,N_19445,N_19731);
nand U23224 (N_23224,N_19092,N_15769);
and U23225 (N_23225,N_17311,N_17053);
xnor U23226 (N_23226,N_15030,N_18960);
and U23227 (N_23227,N_19473,N_16173);
and U23228 (N_23228,N_18119,N_15456);
and U23229 (N_23229,N_18559,N_16231);
or U23230 (N_23230,N_18301,N_18084);
xnor U23231 (N_23231,N_18847,N_18835);
nor U23232 (N_23232,N_16218,N_15433);
and U23233 (N_23233,N_16067,N_19692);
nand U23234 (N_23234,N_18485,N_18012);
nor U23235 (N_23235,N_19334,N_19331);
or U23236 (N_23236,N_18032,N_19125);
or U23237 (N_23237,N_15299,N_17192);
nor U23238 (N_23238,N_18378,N_17403);
nand U23239 (N_23239,N_17907,N_17855);
or U23240 (N_23240,N_18423,N_18504);
or U23241 (N_23241,N_17454,N_16461);
xnor U23242 (N_23242,N_16784,N_19783);
nand U23243 (N_23243,N_17516,N_17530);
or U23244 (N_23244,N_19447,N_18456);
nor U23245 (N_23245,N_15258,N_18412);
or U23246 (N_23246,N_17409,N_19294);
xnor U23247 (N_23247,N_19376,N_16269);
xor U23248 (N_23248,N_17455,N_15427);
and U23249 (N_23249,N_19146,N_15449);
and U23250 (N_23250,N_19527,N_16160);
xor U23251 (N_23251,N_19837,N_18507);
or U23252 (N_23252,N_18218,N_15086);
xnor U23253 (N_23253,N_15618,N_15220);
or U23254 (N_23254,N_19138,N_19920);
nand U23255 (N_23255,N_17864,N_16534);
or U23256 (N_23256,N_16998,N_15414);
nand U23257 (N_23257,N_17106,N_18251);
nand U23258 (N_23258,N_19330,N_19002);
xnor U23259 (N_23259,N_19494,N_17532);
and U23260 (N_23260,N_16128,N_18639);
nor U23261 (N_23261,N_18293,N_16482);
xnor U23262 (N_23262,N_15952,N_15932);
xnor U23263 (N_23263,N_18353,N_17266);
and U23264 (N_23264,N_16503,N_16282);
or U23265 (N_23265,N_16284,N_19035);
xnor U23266 (N_23266,N_16960,N_15059);
nand U23267 (N_23267,N_15645,N_16260);
nand U23268 (N_23268,N_19443,N_17504);
nand U23269 (N_23269,N_15027,N_18336);
or U23270 (N_23270,N_16970,N_16759);
nand U23271 (N_23271,N_17330,N_18303);
nand U23272 (N_23272,N_16756,N_18607);
and U23273 (N_23273,N_19512,N_18205);
and U23274 (N_23274,N_15373,N_19073);
and U23275 (N_23275,N_16850,N_17128);
or U23276 (N_23276,N_18639,N_17210);
and U23277 (N_23277,N_19999,N_18617);
or U23278 (N_23278,N_19134,N_17868);
nor U23279 (N_23279,N_16142,N_17508);
xnor U23280 (N_23280,N_15226,N_18988);
nand U23281 (N_23281,N_16669,N_15140);
xnor U23282 (N_23282,N_17087,N_18530);
nand U23283 (N_23283,N_19113,N_15623);
and U23284 (N_23284,N_15643,N_16268);
xnor U23285 (N_23285,N_19578,N_15456);
nand U23286 (N_23286,N_19972,N_17685);
xor U23287 (N_23287,N_18811,N_15752);
nor U23288 (N_23288,N_18781,N_18626);
nor U23289 (N_23289,N_19781,N_15490);
nand U23290 (N_23290,N_19677,N_18482);
and U23291 (N_23291,N_17154,N_16675);
nand U23292 (N_23292,N_19366,N_18609);
nand U23293 (N_23293,N_19018,N_16754);
nor U23294 (N_23294,N_17829,N_17013);
and U23295 (N_23295,N_15830,N_17027);
and U23296 (N_23296,N_15788,N_17069);
nand U23297 (N_23297,N_18812,N_18206);
and U23298 (N_23298,N_17055,N_15625);
and U23299 (N_23299,N_16575,N_18058);
and U23300 (N_23300,N_17848,N_19629);
and U23301 (N_23301,N_16514,N_17858);
nor U23302 (N_23302,N_17531,N_17175);
nor U23303 (N_23303,N_18732,N_19015);
xor U23304 (N_23304,N_19910,N_17630);
and U23305 (N_23305,N_19124,N_17021);
xor U23306 (N_23306,N_18956,N_19544);
or U23307 (N_23307,N_17276,N_19975);
nand U23308 (N_23308,N_17537,N_15595);
or U23309 (N_23309,N_16218,N_16945);
nand U23310 (N_23310,N_17503,N_15649);
xor U23311 (N_23311,N_16263,N_19348);
nand U23312 (N_23312,N_17213,N_15744);
nand U23313 (N_23313,N_19905,N_15150);
or U23314 (N_23314,N_19625,N_18355);
and U23315 (N_23315,N_18519,N_16232);
nor U23316 (N_23316,N_19515,N_15750);
nor U23317 (N_23317,N_17546,N_17200);
or U23318 (N_23318,N_16323,N_18225);
and U23319 (N_23319,N_19182,N_16604);
nand U23320 (N_23320,N_16519,N_15527);
and U23321 (N_23321,N_17763,N_16282);
and U23322 (N_23322,N_19003,N_18730);
nor U23323 (N_23323,N_18683,N_18188);
or U23324 (N_23324,N_19025,N_19105);
xor U23325 (N_23325,N_19046,N_15351);
nand U23326 (N_23326,N_19135,N_17541);
xnor U23327 (N_23327,N_19450,N_19326);
nand U23328 (N_23328,N_16745,N_19853);
nand U23329 (N_23329,N_16393,N_18528);
xor U23330 (N_23330,N_19007,N_15688);
nand U23331 (N_23331,N_16050,N_16450);
nand U23332 (N_23332,N_18211,N_19947);
xor U23333 (N_23333,N_19820,N_15280);
nor U23334 (N_23334,N_18575,N_17529);
nor U23335 (N_23335,N_19970,N_15771);
nand U23336 (N_23336,N_19366,N_17071);
xnor U23337 (N_23337,N_19678,N_17262);
and U23338 (N_23338,N_18446,N_18991);
or U23339 (N_23339,N_17488,N_18248);
or U23340 (N_23340,N_18663,N_18022);
nand U23341 (N_23341,N_17202,N_17892);
xor U23342 (N_23342,N_18633,N_19128);
nor U23343 (N_23343,N_16861,N_18779);
and U23344 (N_23344,N_18411,N_17993);
nand U23345 (N_23345,N_16635,N_16941);
nor U23346 (N_23346,N_18306,N_18323);
nand U23347 (N_23347,N_16566,N_17151);
nand U23348 (N_23348,N_16551,N_16504);
and U23349 (N_23349,N_19601,N_15968);
nand U23350 (N_23350,N_18355,N_18375);
xnor U23351 (N_23351,N_15157,N_17104);
nand U23352 (N_23352,N_16201,N_17555);
xnor U23353 (N_23353,N_16223,N_16956);
nor U23354 (N_23354,N_15646,N_18527);
xor U23355 (N_23355,N_16341,N_18153);
xor U23356 (N_23356,N_16815,N_17666);
nand U23357 (N_23357,N_18310,N_15382);
xnor U23358 (N_23358,N_16709,N_15000);
nand U23359 (N_23359,N_18788,N_15231);
nor U23360 (N_23360,N_19189,N_19976);
nand U23361 (N_23361,N_19354,N_19271);
or U23362 (N_23362,N_16880,N_15250);
nor U23363 (N_23363,N_16297,N_16570);
nand U23364 (N_23364,N_15198,N_18973);
or U23365 (N_23365,N_18051,N_15788);
xnor U23366 (N_23366,N_19658,N_16445);
nor U23367 (N_23367,N_15729,N_17625);
or U23368 (N_23368,N_18125,N_18800);
nand U23369 (N_23369,N_18364,N_16256);
or U23370 (N_23370,N_19092,N_15368);
nor U23371 (N_23371,N_15049,N_16899);
nand U23372 (N_23372,N_16233,N_17430);
or U23373 (N_23373,N_19699,N_18353);
and U23374 (N_23374,N_19712,N_16574);
xnor U23375 (N_23375,N_15410,N_15074);
nor U23376 (N_23376,N_19284,N_16072);
xnor U23377 (N_23377,N_15573,N_16855);
and U23378 (N_23378,N_16892,N_17761);
and U23379 (N_23379,N_19013,N_17916);
nor U23380 (N_23380,N_15449,N_17697);
or U23381 (N_23381,N_17962,N_16324);
nand U23382 (N_23382,N_16829,N_15742);
xnor U23383 (N_23383,N_16432,N_17772);
nand U23384 (N_23384,N_15169,N_19171);
xnor U23385 (N_23385,N_15557,N_17022);
nor U23386 (N_23386,N_19196,N_15437);
xor U23387 (N_23387,N_17564,N_18492);
and U23388 (N_23388,N_18227,N_17471);
nand U23389 (N_23389,N_17493,N_16530);
nor U23390 (N_23390,N_18891,N_15210);
nor U23391 (N_23391,N_18888,N_16814);
nor U23392 (N_23392,N_16958,N_19174);
xnor U23393 (N_23393,N_16746,N_19248);
nor U23394 (N_23394,N_15145,N_19154);
nor U23395 (N_23395,N_16560,N_17227);
nor U23396 (N_23396,N_15699,N_17720);
xor U23397 (N_23397,N_16328,N_19333);
nand U23398 (N_23398,N_16805,N_16706);
nor U23399 (N_23399,N_16643,N_17051);
nor U23400 (N_23400,N_17237,N_18412);
nand U23401 (N_23401,N_18357,N_18398);
nand U23402 (N_23402,N_16680,N_19773);
or U23403 (N_23403,N_18709,N_18276);
nand U23404 (N_23404,N_16838,N_15073);
or U23405 (N_23405,N_16025,N_19220);
nor U23406 (N_23406,N_19130,N_19816);
nor U23407 (N_23407,N_17699,N_19481);
or U23408 (N_23408,N_18124,N_15344);
xnor U23409 (N_23409,N_16530,N_15239);
nand U23410 (N_23410,N_15819,N_16666);
xor U23411 (N_23411,N_15618,N_17274);
or U23412 (N_23412,N_16922,N_19713);
nor U23413 (N_23413,N_18116,N_19956);
xor U23414 (N_23414,N_17636,N_18900);
xnor U23415 (N_23415,N_17458,N_15526);
xnor U23416 (N_23416,N_19479,N_19569);
xnor U23417 (N_23417,N_19349,N_16496);
nand U23418 (N_23418,N_15664,N_15679);
and U23419 (N_23419,N_19191,N_18951);
and U23420 (N_23420,N_17813,N_19977);
and U23421 (N_23421,N_19116,N_17560);
xnor U23422 (N_23422,N_19637,N_17985);
nor U23423 (N_23423,N_15237,N_16437);
nand U23424 (N_23424,N_17642,N_16603);
nor U23425 (N_23425,N_19170,N_17481);
xor U23426 (N_23426,N_19233,N_17170);
or U23427 (N_23427,N_19327,N_17067);
or U23428 (N_23428,N_15926,N_17243);
nand U23429 (N_23429,N_19375,N_19901);
and U23430 (N_23430,N_18706,N_18070);
and U23431 (N_23431,N_19302,N_16494);
and U23432 (N_23432,N_17005,N_17436);
and U23433 (N_23433,N_19266,N_16607);
xnor U23434 (N_23434,N_16244,N_16282);
nor U23435 (N_23435,N_18022,N_18653);
and U23436 (N_23436,N_17388,N_15677);
xnor U23437 (N_23437,N_17798,N_18787);
xnor U23438 (N_23438,N_18522,N_17558);
nand U23439 (N_23439,N_17739,N_15095);
nand U23440 (N_23440,N_18334,N_18040);
nand U23441 (N_23441,N_18994,N_19514);
and U23442 (N_23442,N_16392,N_15045);
xor U23443 (N_23443,N_19927,N_16683);
nor U23444 (N_23444,N_16109,N_15550);
xor U23445 (N_23445,N_17299,N_16836);
and U23446 (N_23446,N_19974,N_17288);
xor U23447 (N_23447,N_15744,N_16507);
or U23448 (N_23448,N_19464,N_18379);
or U23449 (N_23449,N_15951,N_18462);
nor U23450 (N_23450,N_19705,N_19318);
or U23451 (N_23451,N_15696,N_15202);
nor U23452 (N_23452,N_15721,N_17772);
and U23453 (N_23453,N_18337,N_17084);
and U23454 (N_23454,N_19201,N_15297);
xnor U23455 (N_23455,N_18823,N_17297);
nand U23456 (N_23456,N_15996,N_18891);
nor U23457 (N_23457,N_15705,N_17302);
nand U23458 (N_23458,N_17527,N_18978);
nor U23459 (N_23459,N_16805,N_15196);
nand U23460 (N_23460,N_15825,N_16707);
and U23461 (N_23461,N_17680,N_15883);
and U23462 (N_23462,N_15216,N_17022);
nand U23463 (N_23463,N_16163,N_15942);
nand U23464 (N_23464,N_17942,N_17193);
and U23465 (N_23465,N_15053,N_16986);
xor U23466 (N_23466,N_16707,N_15034);
and U23467 (N_23467,N_18652,N_16392);
xnor U23468 (N_23468,N_16631,N_16616);
or U23469 (N_23469,N_15285,N_18243);
or U23470 (N_23470,N_18843,N_15122);
xor U23471 (N_23471,N_17960,N_15784);
or U23472 (N_23472,N_16203,N_15450);
and U23473 (N_23473,N_16546,N_17116);
or U23474 (N_23474,N_15636,N_19553);
or U23475 (N_23475,N_19402,N_17896);
nor U23476 (N_23476,N_15410,N_18449);
and U23477 (N_23477,N_16071,N_17593);
or U23478 (N_23478,N_18929,N_15805);
xor U23479 (N_23479,N_18272,N_18833);
and U23480 (N_23480,N_19518,N_16059);
xnor U23481 (N_23481,N_16250,N_18575);
nand U23482 (N_23482,N_16579,N_19398);
xnor U23483 (N_23483,N_18959,N_15055);
nor U23484 (N_23484,N_18997,N_18678);
nor U23485 (N_23485,N_16523,N_16153);
nor U23486 (N_23486,N_15640,N_15631);
and U23487 (N_23487,N_18688,N_17782);
xor U23488 (N_23488,N_16199,N_15138);
nand U23489 (N_23489,N_15645,N_16248);
or U23490 (N_23490,N_17416,N_17674);
nor U23491 (N_23491,N_16263,N_17595);
and U23492 (N_23492,N_19848,N_15025);
or U23493 (N_23493,N_17611,N_16621);
nand U23494 (N_23494,N_17193,N_17586);
xnor U23495 (N_23495,N_15628,N_18188);
nand U23496 (N_23496,N_15922,N_18814);
nand U23497 (N_23497,N_19556,N_16113);
and U23498 (N_23498,N_16023,N_16460);
or U23499 (N_23499,N_17844,N_15337);
xor U23500 (N_23500,N_15433,N_16145);
or U23501 (N_23501,N_16552,N_19701);
nand U23502 (N_23502,N_16328,N_19360);
xor U23503 (N_23503,N_19879,N_15824);
and U23504 (N_23504,N_18090,N_17820);
or U23505 (N_23505,N_16146,N_15296);
nand U23506 (N_23506,N_16134,N_16516);
xor U23507 (N_23507,N_17998,N_17403);
xnor U23508 (N_23508,N_19406,N_18320);
nor U23509 (N_23509,N_16884,N_18786);
and U23510 (N_23510,N_19501,N_17061);
xor U23511 (N_23511,N_17317,N_15424);
nand U23512 (N_23512,N_15413,N_15690);
nor U23513 (N_23513,N_17003,N_19242);
or U23514 (N_23514,N_18160,N_15185);
nor U23515 (N_23515,N_15597,N_19386);
xnor U23516 (N_23516,N_19830,N_16026);
or U23517 (N_23517,N_18271,N_18044);
xor U23518 (N_23518,N_15681,N_15614);
nand U23519 (N_23519,N_16375,N_17796);
nand U23520 (N_23520,N_19323,N_15164);
nand U23521 (N_23521,N_19515,N_18669);
xnor U23522 (N_23522,N_16645,N_15588);
nor U23523 (N_23523,N_18113,N_15147);
xor U23524 (N_23524,N_19212,N_16199);
or U23525 (N_23525,N_18630,N_19163);
or U23526 (N_23526,N_16841,N_17603);
nand U23527 (N_23527,N_17205,N_18664);
nand U23528 (N_23528,N_17581,N_17505);
nor U23529 (N_23529,N_16644,N_15165);
nand U23530 (N_23530,N_17465,N_17605);
nor U23531 (N_23531,N_19029,N_17622);
and U23532 (N_23532,N_19174,N_15379);
and U23533 (N_23533,N_18167,N_15359);
xnor U23534 (N_23534,N_18100,N_16170);
xnor U23535 (N_23535,N_18436,N_15548);
and U23536 (N_23536,N_18316,N_17081);
xor U23537 (N_23537,N_18723,N_16508);
nand U23538 (N_23538,N_19939,N_16126);
xor U23539 (N_23539,N_15878,N_18190);
nand U23540 (N_23540,N_16233,N_16000);
nor U23541 (N_23541,N_16642,N_19245);
nor U23542 (N_23542,N_16119,N_15347);
xnor U23543 (N_23543,N_15003,N_15185);
nand U23544 (N_23544,N_17036,N_15517);
nand U23545 (N_23545,N_19476,N_16403);
xnor U23546 (N_23546,N_19184,N_17863);
xor U23547 (N_23547,N_18816,N_15149);
nor U23548 (N_23548,N_15019,N_16679);
xor U23549 (N_23549,N_15943,N_17450);
or U23550 (N_23550,N_17389,N_18313);
nand U23551 (N_23551,N_19586,N_18305);
nor U23552 (N_23552,N_16447,N_15659);
or U23553 (N_23553,N_18575,N_15307);
xnor U23554 (N_23554,N_18931,N_19748);
and U23555 (N_23555,N_15999,N_18688);
and U23556 (N_23556,N_15553,N_15835);
or U23557 (N_23557,N_19712,N_15809);
nand U23558 (N_23558,N_19158,N_18555);
and U23559 (N_23559,N_17939,N_19939);
nor U23560 (N_23560,N_15937,N_16411);
and U23561 (N_23561,N_16779,N_16883);
nand U23562 (N_23562,N_17266,N_19987);
xor U23563 (N_23563,N_18655,N_16709);
xor U23564 (N_23564,N_16835,N_16580);
or U23565 (N_23565,N_15178,N_17336);
or U23566 (N_23566,N_15043,N_16898);
or U23567 (N_23567,N_18734,N_16041);
xor U23568 (N_23568,N_15878,N_19466);
nand U23569 (N_23569,N_17985,N_18385);
or U23570 (N_23570,N_15145,N_19783);
xor U23571 (N_23571,N_16702,N_19718);
and U23572 (N_23572,N_19910,N_17907);
and U23573 (N_23573,N_19625,N_19603);
nand U23574 (N_23574,N_18348,N_17100);
nand U23575 (N_23575,N_19939,N_15936);
nand U23576 (N_23576,N_15112,N_16114);
and U23577 (N_23577,N_16669,N_18708);
xnor U23578 (N_23578,N_17528,N_16423);
and U23579 (N_23579,N_18669,N_17597);
nand U23580 (N_23580,N_19845,N_16883);
xnor U23581 (N_23581,N_18775,N_18404);
xor U23582 (N_23582,N_15672,N_18339);
and U23583 (N_23583,N_18238,N_19561);
and U23584 (N_23584,N_16349,N_17874);
nand U23585 (N_23585,N_18480,N_18752);
nor U23586 (N_23586,N_19457,N_18109);
nand U23587 (N_23587,N_15193,N_18272);
or U23588 (N_23588,N_19415,N_19966);
nand U23589 (N_23589,N_19366,N_16954);
nand U23590 (N_23590,N_15801,N_16924);
nor U23591 (N_23591,N_17849,N_16787);
nor U23592 (N_23592,N_19068,N_16806);
and U23593 (N_23593,N_19544,N_19201);
nor U23594 (N_23594,N_16716,N_19759);
or U23595 (N_23595,N_16268,N_15031);
nor U23596 (N_23596,N_18800,N_15803);
xnor U23597 (N_23597,N_16703,N_16425);
nor U23598 (N_23598,N_17300,N_15638);
nor U23599 (N_23599,N_19609,N_18388);
nand U23600 (N_23600,N_16387,N_16347);
nor U23601 (N_23601,N_17131,N_19065);
or U23602 (N_23602,N_15292,N_16145);
nand U23603 (N_23603,N_18331,N_19787);
nand U23604 (N_23604,N_15404,N_16681);
nor U23605 (N_23605,N_17415,N_17040);
nor U23606 (N_23606,N_19717,N_18409);
xnor U23607 (N_23607,N_18763,N_15514);
or U23608 (N_23608,N_15723,N_15142);
and U23609 (N_23609,N_19743,N_15137);
and U23610 (N_23610,N_18593,N_18841);
xor U23611 (N_23611,N_19287,N_19254);
and U23612 (N_23612,N_16326,N_15753);
nand U23613 (N_23613,N_15080,N_16030);
nand U23614 (N_23614,N_15614,N_15281);
or U23615 (N_23615,N_17343,N_19728);
nand U23616 (N_23616,N_18466,N_17453);
nor U23617 (N_23617,N_18514,N_15815);
and U23618 (N_23618,N_19588,N_15743);
nor U23619 (N_23619,N_16551,N_15672);
nor U23620 (N_23620,N_18250,N_15296);
nor U23621 (N_23621,N_17019,N_18111);
nand U23622 (N_23622,N_16057,N_16229);
nand U23623 (N_23623,N_16303,N_19417);
and U23624 (N_23624,N_17115,N_15256);
nand U23625 (N_23625,N_15840,N_17278);
nor U23626 (N_23626,N_17043,N_18002);
nor U23627 (N_23627,N_18818,N_16336);
and U23628 (N_23628,N_17765,N_15134);
or U23629 (N_23629,N_15246,N_15019);
xor U23630 (N_23630,N_15832,N_19990);
or U23631 (N_23631,N_16177,N_18983);
and U23632 (N_23632,N_19800,N_17653);
xor U23633 (N_23633,N_18311,N_17478);
and U23634 (N_23634,N_19456,N_15708);
nor U23635 (N_23635,N_15029,N_15001);
nor U23636 (N_23636,N_17479,N_18404);
nand U23637 (N_23637,N_16749,N_15560);
or U23638 (N_23638,N_15305,N_15969);
nand U23639 (N_23639,N_19399,N_18289);
xnor U23640 (N_23640,N_16728,N_16532);
nand U23641 (N_23641,N_17973,N_15656);
and U23642 (N_23642,N_15594,N_17600);
nor U23643 (N_23643,N_18194,N_18391);
or U23644 (N_23644,N_18428,N_17226);
nand U23645 (N_23645,N_15272,N_18037);
xor U23646 (N_23646,N_16767,N_19834);
and U23647 (N_23647,N_19600,N_19010);
and U23648 (N_23648,N_15127,N_19570);
xnor U23649 (N_23649,N_18418,N_16050);
nor U23650 (N_23650,N_16879,N_16355);
nand U23651 (N_23651,N_15441,N_15408);
or U23652 (N_23652,N_15958,N_17916);
xnor U23653 (N_23653,N_17838,N_19908);
xor U23654 (N_23654,N_15463,N_19473);
or U23655 (N_23655,N_19877,N_15288);
nand U23656 (N_23656,N_19448,N_19950);
xnor U23657 (N_23657,N_17291,N_18439);
and U23658 (N_23658,N_19583,N_17539);
xor U23659 (N_23659,N_17807,N_16218);
and U23660 (N_23660,N_16530,N_17439);
nand U23661 (N_23661,N_16724,N_19353);
or U23662 (N_23662,N_15605,N_19604);
or U23663 (N_23663,N_15844,N_17422);
nor U23664 (N_23664,N_19161,N_16276);
xor U23665 (N_23665,N_19469,N_16103);
xor U23666 (N_23666,N_16090,N_17559);
nand U23667 (N_23667,N_15709,N_16085);
xor U23668 (N_23668,N_19753,N_15095);
nand U23669 (N_23669,N_16556,N_15435);
nor U23670 (N_23670,N_18490,N_18666);
nand U23671 (N_23671,N_19571,N_18823);
or U23672 (N_23672,N_15901,N_17725);
nand U23673 (N_23673,N_17474,N_16606);
and U23674 (N_23674,N_19445,N_18850);
xor U23675 (N_23675,N_16788,N_16015);
nand U23676 (N_23676,N_18361,N_19341);
or U23677 (N_23677,N_19176,N_18439);
xnor U23678 (N_23678,N_15715,N_17637);
and U23679 (N_23679,N_15051,N_19042);
nand U23680 (N_23680,N_17776,N_15082);
and U23681 (N_23681,N_18970,N_16459);
xor U23682 (N_23682,N_17145,N_16923);
nand U23683 (N_23683,N_17929,N_16822);
xnor U23684 (N_23684,N_18132,N_16085);
or U23685 (N_23685,N_19194,N_17888);
nand U23686 (N_23686,N_19297,N_16597);
nand U23687 (N_23687,N_15462,N_15954);
nor U23688 (N_23688,N_18242,N_18419);
or U23689 (N_23689,N_18587,N_16406);
or U23690 (N_23690,N_18567,N_17742);
nor U23691 (N_23691,N_15923,N_19689);
and U23692 (N_23692,N_18359,N_16453);
nand U23693 (N_23693,N_16059,N_19175);
or U23694 (N_23694,N_16560,N_17336);
xor U23695 (N_23695,N_15714,N_15303);
xnor U23696 (N_23696,N_18790,N_16904);
nand U23697 (N_23697,N_16753,N_17008);
xnor U23698 (N_23698,N_17011,N_16277);
and U23699 (N_23699,N_18138,N_17040);
nor U23700 (N_23700,N_16237,N_15262);
nand U23701 (N_23701,N_18157,N_15450);
nand U23702 (N_23702,N_19085,N_16182);
or U23703 (N_23703,N_16616,N_16837);
nand U23704 (N_23704,N_16893,N_16091);
nor U23705 (N_23705,N_15205,N_18733);
xnor U23706 (N_23706,N_16038,N_15895);
and U23707 (N_23707,N_15665,N_15544);
or U23708 (N_23708,N_18690,N_18108);
and U23709 (N_23709,N_18700,N_16188);
nand U23710 (N_23710,N_17659,N_17656);
nor U23711 (N_23711,N_15094,N_17258);
nor U23712 (N_23712,N_18293,N_17246);
and U23713 (N_23713,N_19995,N_15580);
nand U23714 (N_23714,N_16200,N_18025);
xor U23715 (N_23715,N_18141,N_17251);
and U23716 (N_23716,N_16888,N_15797);
or U23717 (N_23717,N_15349,N_17420);
or U23718 (N_23718,N_16304,N_15074);
nand U23719 (N_23719,N_17224,N_18496);
nand U23720 (N_23720,N_19333,N_16167);
and U23721 (N_23721,N_19456,N_17363);
xnor U23722 (N_23722,N_18247,N_19624);
nand U23723 (N_23723,N_15274,N_17619);
xor U23724 (N_23724,N_19222,N_19267);
and U23725 (N_23725,N_19491,N_15803);
nand U23726 (N_23726,N_18834,N_17318);
and U23727 (N_23727,N_16896,N_15173);
xor U23728 (N_23728,N_16138,N_19582);
and U23729 (N_23729,N_15926,N_19662);
or U23730 (N_23730,N_15966,N_18165);
and U23731 (N_23731,N_19857,N_19736);
nor U23732 (N_23732,N_15095,N_17054);
nor U23733 (N_23733,N_16927,N_18366);
or U23734 (N_23734,N_16883,N_17750);
or U23735 (N_23735,N_19646,N_16755);
or U23736 (N_23736,N_19186,N_15535);
xnor U23737 (N_23737,N_19723,N_16881);
xnor U23738 (N_23738,N_17915,N_15273);
nand U23739 (N_23739,N_16805,N_18320);
or U23740 (N_23740,N_17158,N_19303);
nand U23741 (N_23741,N_19268,N_15021);
nor U23742 (N_23742,N_17736,N_16027);
and U23743 (N_23743,N_16780,N_19195);
xnor U23744 (N_23744,N_19554,N_16168);
and U23745 (N_23745,N_16622,N_16163);
nand U23746 (N_23746,N_15557,N_18675);
xor U23747 (N_23747,N_17288,N_15697);
nand U23748 (N_23748,N_18718,N_19323);
and U23749 (N_23749,N_17635,N_16334);
or U23750 (N_23750,N_18468,N_16068);
nand U23751 (N_23751,N_15020,N_17763);
and U23752 (N_23752,N_17009,N_15494);
and U23753 (N_23753,N_17932,N_17068);
xor U23754 (N_23754,N_15585,N_15647);
nor U23755 (N_23755,N_19820,N_18049);
xnor U23756 (N_23756,N_16410,N_19219);
xor U23757 (N_23757,N_17655,N_15948);
xor U23758 (N_23758,N_16334,N_18997);
xor U23759 (N_23759,N_15912,N_16460);
xor U23760 (N_23760,N_15131,N_19206);
nor U23761 (N_23761,N_15228,N_16075);
nor U23762 (N_23762,N_16972,N_15146);
and U23763 (N_23763,N_18147,N_15164);
xor U23764 (N_23764,N_19965,N_16854);
or U23765 (N_23765,N_16894,N_19888);
xnor U23766 (N_23766,N_16392,N_16833);
nor U23767 (N_23767,N_19678,N_15472);
xor U23768 (N_23768,N_19952,N_17407);
and U23769 (N_23769,N_16602,N_18528);
xor U23770 (N_23770,N_19768,N_18131);
or U23771 (N_23771,N_17329,N_18605);
xor U23772 (N_23772,N_18675,N_17064);
or U23773 (N_23773,N_18622,N_18578);
nand U23774 (N_23774,N_18360,N_18184);
nand U23775 (N_23775,N_15277,N_16215);
xor U23776 (N_23776,N_17757,N_15198);
and U23777 (N_23777,N_15737,N_18425);
nand U23778 (N_23778,N_15566,N_15204);
and U23779 (N_23779,N_19131,N_18564);
and U23780 (N_23780,N_15952,N_18795);
nand U23781 (N_23781,N_17868,N_16947);
and U23782 (N_23782,N_19511,N_17322);
nor U23783 (N_23783,N_17568,N_19357);
nor U23784 (N_23784,N_19766,N_18580);
and U23785 (N_23785,N_16962,N_18425);
xnor U23786 (N_23786,N_19239,N_15856);
and U23787 (N_23787,N_18420,N_19125);
or U23788 (N_23788,N_19320,N_18958);
or U23789 (N_23789,N_16702,N_15561);
nor U23790 (N_23790,N_19335,N_15841);
nand U23791 (N_23791,N_17700,N_16649);
nor U23792 (N_23792,N_19851,N_19806);
and U23793 (N_23793,N_17557,N_19164);
and U23794 (N_23794,N_16419,N_18977);
or U23795 (N_23795,N_15975,N_17652);
and U23796 (N_23796,N_15695,N_17319);
nor U23797 (N_23797,N_19166,N_17077);
or U23798 (N_23798,N_19758,N_16903);
nor U23799 (N_23799,N_16333,N_18322);
nor U23800 (N_23800,N_15027,N_18231);
nand U23801 (N_23801,N_17380,N_18436);
nand U23802 (N_23802,N_16314,N_17280);
xnor U23803 (N_23803,N_15884,N_18084);
nor U23804 (N_23804,N_16610,N_19149);
nor U23805 (N_23805,N_17441,N_15528);
or U23806 (N_23806,N_18997,N_17238);
xor U23807 (N_23807,N_17528,N_18615);
and U23808 (N_23808,N_17909,N_16275);
xnor U23809 (N_23809,N_18633,N_18629);
nor U23810 (N_23810,N_16382,N_19544);
xnor U23811 (N_23811,N_18548,N_17997);
or U23812 (N_23812,N_15693,N_19220);
xnor U23813 (N_23813,N_16755,N_15779);
nor U23814 (N_23814,N_18132,N_17996);
and U23815 (N_23815,N_15476,N_16436);
or U23816 (N_23816,N_19132,N_15178);
xnor U23817 (N_23817,N_16498,N_15059);
and U23818 (N_23818,N_15339,N_16283);
nor U23819 (N_23819,N_15912,N_15259);
nor U23820 (N_23820,N_16182,N_18595);
xor U23821 (N_23821,N_19121,N_19326);
nand U23822 (N_23822,N_19599,N_16128);
xnor U23823 (N_23823,N_15944,N_19546);
xor U23824 (N_23824,N_15019,N_18459);
nand U23825 (N_23825,N_19482,N_15055);
or U23826 (N_23826,N_17033,N_17633);
xnor U23827 (N_23827,N_19476,N_17418);
xor U23828 (N_23828,N_17138,N_15292);
nand U23829 (N_23829,N_15698,N_16284);
and U23830 (N_23830,N_18784,N_16572);
or U23831 (N_23831,N_18084,N_16333);
xnor U23832 (N_23832,N_18525,N_15390);
xor U23833 (N_23833,N_15193,N_17652);
or U23834 (N_23834,N_19492,N_18230);
nor U23835 (N_23835,N_16000,N_17052);
and U23836 (N_23836,N_17143,N_16867);
xor U23837 (N_23837,N_18314,N_18073);
or U23838 (N_23838,N_19830,N_17127);
nor U23839 (N_23839,N_15976,N_15595);
nand U23840 (N_23840,N_15513,N_19664);
nand U23841 (N_23841,N_18113,N_19560);
or U23842 (N_23842,N_18582,N_15971);
or U23843 (N_23843,N_16909,N_15211);
and U23844 (N_23844,N_18505,N_18305);
nand U23845 (N_23845,N_17023,N_16561);
nor U23846 (N_23846,N_18286,N_16870);
nor U23847 (N_23847,N_16778,N_18223);
nand U23848 (N_23848,N_15217,N_19758);
xor U23849 (N_23849,N_16931,N_15804);
nand U23850 (N_23850,N_17910,N_18257);
nand U23851 (N_23851,N_15613,N_16739);
and U23852 (N_23852,N_16781,N_18647);
xor U23853 (N_23853,N_16056,N_16927);
nor U23854 (N_23854,N_16346,N_15327);
or U23855 (N_23855,N_17431,N_15073);
or U23856 (N_23856,N_17291,N_17246);
nor U23857 (N_23857,N_19987,N_19682);
or U23858 (N_23858,N_18074,N_19911);
nor U23859 (N_23859,N_19508,N_15208);
and U23860 (N_23860,N_19363,N_17182);
nor U23861 (N_23861,N_17915,N_16812);
xnor U23862 (N_23862,N_17281,N_15435);
and U23863 (N_23863,N_15980,N_17400);
nor U23864 (N_23864,N_19949,N_16947);
nor U23865 (N_23865,N_16515,N_16070);
xnor U23866 (N_23866,N_17514,N_18183);
xor U23867 (N_23867,N_18830,N_17047);
xor U23868 (N_23868,N_18032,N_19236);
nand U23869 (N_23869,N_15191,N_18210);
nand U23870 (N_23870,N_19857,N_18468);
nor U23871 (N_23871,N_17180,N_16366);
or U23872 (N_23872,N_17538,N_15297);
and U23873 (N_23873,N_17753,N_18070);
nand U23874 (N_23874,N_17553,N_17617);
nand U23875 (N_23875,N_16042,N_18759);
and U23876 (N_23876,N_18276,N_15713);
nand U23877 (N_23877,N_19145,N_19256);
or U23878 (N_23878,N_15207,N_19819);
or U23879 (N_23879,N_18941,N_17123);
nor U23880 (N_23880,N_15339,N_19358);
and U23881 (N_23881,N_16085,N_16288);
or U23882 (N_23882,N_19583,N_16241);
and U23883 (N_23883,N_16768,N_15455);
nand U23884 (N_23884,N_19152,N_17832);
xor U23885 (N_23885,N_17053,N_16158);
nand U23886 (N_23886,N_18905,N_17088);
nand U23887 (N_23887,N_17900,N_19431);
nor U23888 (N_23888,N_18275,N_18130);
xnor U23889 (N_23889,N_15972,N_19222);
nor U23890 (N_23890,N_16620,N_19213);
nor U23891 (N_23891,N_16886,N_19267);
nand U23892 (N_23892,N_17490,N_17253);
nor U23893 (N_23893,N_18587,N_19297);
nand U23894 (N_23894,N_18924,N_16688);
nor U23895 (N_23895,N_17783,N_16094);
and U23896 (N_23896,N_18070,N_15384);
or U23897 (N_23897,N_16250,N_15385);
nor U23898 (N_23898,N_15436,N_17410);
xnor U23899 (N_23899,N_17628,N_19553);
nor U23900 (N_23900,N_18798,N_19792);
or U23901 (N_23901,N_16956,N_16047);
nor U23902 (N_23902,N_15517,N_17785);
nor U23903 (N_23903,N_18474,N_18419);
nor U23904 (N_23904,N_17010,N_17868);
nor U23905 (N_23905,N_17691,N_18207);
and U23906 (N_23906,N_17731,N_16952);
nand U23907 (N_23907,N_19265,N_19790);
nand U23908 (N_23908,N_15642,N_16955);
and U23909 (N_23909,N_15860,N_15373);
or U23910 (N_23910,N_16652,N_19303);
nor U23911 (N_23911,N_15286,N_19760);
and U23912 (N_23912,N_17586,N_19553);
or U23913 (N_23913,N_16727,N_15930);
xnor U23914 (N_23914,N_16016,N_18384);
xnor U23915 (N_23915,N_17200,N_17313);
and U23916 (N_23916,N_19412,N_19778);
nor U23917 (N_23917,N_17268,N_15897);
nor U23918 (N_23918,N_16682,N_18446);
or U23919 (N_23919,N_15810,N_19967);
nor U23920 (N_23920,N_17333,N_19727);
nor U23921 (N_23921,N_18629,N_19283);
and U23922 (N_23922,N_17489,N_16623);
and U23923 (N_23923,N_15788,N_15607);
or U23924 (N_23924,N_15184,N_17657);
or U23925 (N_23925,N_17823,N_16421);
xnor U23926 (N_23926,N_15231,N_17678);
or U23927 (N_23927,N_19484,N_16423);
nor U23928 (N_23928,N_18414,N_17922);
xor U23929 (N_23929,N_18685,N_19034);
and U23930 (N_23930,N_19199,N_16545);
and U23931 (N_23931,N_18879,N_19482);
and U23932 (N_23932,N_19762,N_15754);
nor U23933 (N_23933,N_19551,N_18920);
nand U23934 (N_23934,N_19198,N_17190);
or U23935 (N_23935,N_18797,N_16140);
xor U23936 (N_23936,N_17481,N_16879);
xor U23937 (N_23937,N_17934,N_15409);
nand U23938 (N_23938,N_17106,N_15250);
nand U23939 (N_23939,N_16241,N_16473);
or U23940 (N_23940,N_16606,N_19106);
or U23941 (N_23941,N_19978,N_19991);
or U23942 (N_23942,N_19711,N_17366);
nand U23943 (N_23943,N_16471,N_18618);
xor U23944 (N_23944,N_18237,N_16697);
nor U23945 (N_23945,N_18151,N_16008);
nand U23946 (N_23946,N_18084,N_18104);
and U23947 (N_23947,N_17686,N_15374);
and U23948 (N_23948,N_18320,N_15763);
and U23949 (N_23949,N_16009,N_19072);
nor U23950 (N_23950,N_19426,N_16729);
or U23951 (N_23951,N_16477,N_18377);
nand U23952 (N_23952,N_15905,N_16979);
and U23953 (N_23953,N_18290,N_16676);
xor U23954 (N_23954,N_17607,N_16258);
xor U23955 (N_23955,N_19380,N_19480);
nand U23956 (N_23956,N_17137,N_16723);
or U23957 (N_23957,N_15094,N_19331);
and U23958 (N_23958,N_16188,N_16370);
and U23959 (N_23959,N_16004,N_16647);
nand U23960 (N_23960,N_17121,N_15672);
xnor U23961 (N_23961,N_19166,N_18087);
xnor U23962 (N_23962,N_17406,N_18307);
nor U23963 (N_23963,N_16222,N_15765);
xnor U23964 (N_23964,N_16532,N_19917);
xnor U23965 (N_23965,N_18998,N_16285);
or U23966 (N_23966,N_16854,N_15795);
and U23967 (N_23967,N_16253,N_16703);
xor U23968 (N_23968,N_17924,N_17319);
nor U23969 (N_23969,N_17591,N_15753);
nand U23970 (N_23970,N_15005,N_18459);
xor U23971 (N_23971,N_19050,N_15029);
and U23972 (N_23972,N_15990,N_18296);
and U23973 (N_23973,N_19866,N_18398);
or U23974 (N_23974,N_17120,N_15135);
xor U23975 (N_23975,N_17744,N_16831);
nor U23976 (N_23976,N_17987,N_15903);
xor U23977 (N_23977,N_18605,N_16958);
or U23978 (N_23978,N_18384,N_19234);
nand U23979 (N_23979,N_15374,N_15737);
nor U23980 (N_23980,N_16290,N_17837);
and U23981 (N_23981,N_15162,N_19807);
xor U23982 (N_23982,N_19062,N_15900);
or U23983 (N_23983,N_19264,N_17950);
and U23984 (N_23984,N_18249,N_18337);
nand U23985 (N_23985,N_18710,N_17472);
and U23986 (N_23986,N_19419,N_16574);
or U23987 (N_23987,N_15365,N_19886);
nand U23988 (N_23988,N_19894,N_16891);
and U23989 (N_23989,N_17249,N_18547);
and U23990 (N_23990,N_15959,N_18316);
and U23991 (N_23991,N_17617,N_19113);
or U23992 (N_23992,N_18264,N_19002);
xor U23993 (N_23993,N_18802,N_19878);
or U23994 (N_23994,N_18371,N_15426);
xnor U23995 (N_23995,N_18399,N_17030);
and U23996 (N_23996,N_16738,N_15811);
xnor U23997 (N_23997,N_16445,N_16416);
xor U23998 (N_23998,N_19823,N_19503);
and U23999 (N_23999,N_15418,N_19139);
and U24000 (N_24000,N_15975,N_16421);
nand U24001 (N_24001,N_19322,N_18848);
or U24002 (N_24002,N_17379,N_19387);
nor U24003 (N_24003,N_17957,N_15792);
nor U24004 (N_24004,N_18868,N_16587);
and U24005 (N_24005,N_18068,N_18534);
or U24006 (N_24006,N_16402,N_16373);
or U24007 (N_24007,N_16608,N_18503);
xnor U24008 (N_24008,N_18437,N_19739);
xor U24009 (N_24009,N_18454,N_15334);
nor U24010 (N_24010,N_17232,N_17934);
and U24011 (N_24011,N_19105,N_18986);
nor U24012 (N_24012,N_16073,N_17622);
xor U24013 (N_24013,N_16521,N_16091);
nor U24014 (N_24014,N_16352,N_17569);
nor U24015 (N_24015,N_17640,N_16753);
and U24016 (N_24016,N_19210,N_19305);
or U24017 (N_24017,N_16625,N_15001);
nor U24018 (N_24018,N_16027,N_17947);
and U24019 (N_24019,N_16462,N_19731);
or U24020 (N_24020,N_19708,N_16653);
and U24021 (N_24021,N_19898,N_17745);
xor U24022 (N_24022,N_16270,N_15496);
nor U24023 (N_24023,N_18398,N_16091);
xor U24024 (N_24024,N_17983,N_19916);
nand U24025 (N_24025,N_16961,N_18514);
nand U24026 (N_24026,N_17618,N_15469);
and U24027 (N_24027,N_19531,N_17165);
xor U24028 (N_24028,N_16525,N_19431);
and U24029 (N_24029,N_19291,N_19872);
or U24030 (N_24030,N_16382,N_17149);
xnor U24031 (N_24031,N_18726,N_15126);
and U24032 (N_24032,N_15024,N_19112);
nor U24033 (N_24033,N_15276,N_16222);
and U24034 (N_24034,N_18726,N_18283);
xor U24035 (N_24035,N_16567,N_17663);
nand U24036 (N_24036,N_15520,N_17741);
xor U24037 (N_24037,N_18633,N_15720);
or U24038 (N_24038,N_18963,N_19311);
or U24039 (N_24039,N_18461,N_17817);
and U24040 (N_24040,N_19294,N_18075);
or U24041 (N_24041,N_18300,N_16458);
xnor U24042 (N_24042,N_19152,N_18502);
nand U24043 (N_24043,N_17698,N_19049);
or U24044 (N_24044,N_19117,N_15291);
nor U24045 (N_24045,N_18826,N_15157);
and U24046 (N_24046,N_15119,N_15749);
or U24047 (N_24047,N_18656,N_18609);
and U24048 (N_24048,N_17660,N_16393);
xnor U24049 (N_24049,N_19692,N_16034);
nand U24050 (N_24050,N_16656,N_19621);
nand U24051 (N_24051,N_19712,N_17365);
and U24052 (N_24052,N_18115,N_18990);
nor U24053 (N_24053,N_18169,N_19154);
xnor U24054 (N_24054,N_19571,N_17841);
and U24055 (N_24055,N_16573,N_19416);
nand U24056 (N_24056,N_18971,N_19371);
and U24057 (N_24057,N_15686,N_19842);
nand U24058 (N_24058,N_16209,N_16102);
and U24059 (N_24059,N_19680,N_19207);
nor U24060 (N_24060,N_19858,N_16170);
or U24061 (N_24061,N_16720,N_15819);
and U24062 (N_24062,N_18949,N_16549);
nand U24063 (N_24063,N_17574,N_17165);
nand U24064 (N_24064,N_15643,N_18133);
nand U24065 (N_24065,N_19061,N_18116);
and U24066 (N_24066,N_17610,N_19452);
and U24067 (N_24067,N_16860,N_16039);
nand U24068 (N_24068,N_18267,N_18634);
xnor U24069 (N_24069,N_18583,N_16437);
xnor U24070 (N_24070,N_17898,N_19399);
and U24071 (N_24071,N_17905,N_19395);
or U24072 (N_24072,N_18208,N_15332);
xor U24073 (N_24073,N_15189,N_19551);
and U24074 (N_24074,N_15317,N_15856);
nand U24075 (N_24075,N_16515,N_19411);
nor U24076 (N_24076,N_19894,N_17191);
nand U24077 (N_24077,N_19345,N_17197);
nand U24078 (N_24078,N_15789,N_16005);
xnor U24079 (N_24079,N_17314,N_19223);
nand U24080 (N_24080,N_16706,N_17169);
nand U24081 (N_24081,N_19276,N_19457);
nand U24082 (N_24082,N_19503,N_19373);
xnor U24083 (N_24083,N_17431,N_17589);
xor U24084 (N_24084,N_19837,N_19392);
nor U24085 (N_24085,N_17138,N_15313);
and U24086 (N_24086,N_18215,N_17982);
xor U24087 (N_24087,N_16430,N_15401);
nor U24088 (N_24088,N_16135,N_16478);
or U24089 (N_24089,N_18564,N_16987);
or U24090 (N_24090,N_18202,N_19000);
nor U24091 (N_24091,N_19893,N_16997);
and U24092 (N_24092,N_15225,N_19777);
nand U24093 (N_24093,N_15114,N_15870);
nand U24094 (N_24094,N_17316,N_17202);
or U24095 (N_24095,N_15069,N_18400);
xor U24096 (N_24096,N_16657,N_19595);
or U24097 (N_24097,N_16441,N_16482);
nand U24098 (N_24098,N_17907,N_15075);
nor U24099 (N_24099,N_18666,N_19709);
and U24100 (N_24100,N_18142,N_16315);
nor U24101 (N_24101,N_19955,N_19868);
nor U24102 (N_24102,N_19104,N_19759);
or U24103 (N_24103,N_18035,N_15766);
or U24104 (N_24104,N_17796,N_16766);
or U24105 (N_24105,N_16447,N_18259);
xnor U24106 (N_24106,N_18427,N_17313);
and U24107 (N_24107,N_16344,N_18253);
and U24108 (N_24108,N_19559,N_17143);
nor U24109 (N_24109,N_18619,N_16433);
and U24110 (N_24110,N_15257,N_18291);
xnor U24111 (N_24111,N_16176,N_18786);
or U24112 (N_24112,N_18380,N_15310);
and U24113 (N_24113,N_15958,N_16624);
or U24114 (N_24114,N_16723,N_15195);
nand U24115 (N_24115,N_19204,N_17093);
nand U24116 (N_24116,N_16599,N_15902);
nand U24117 (N_24117,N_18931,N_16807);
or U24118 (N_24118,N_17633,N_16309);
and U24119 (N_24119,N_17822,N_17533);
nor U24120 (N_24120,N_19799,N_19957);
nand U24121 (N_24121,N_18020,N_18763);
nor U24122 (N_24122,N_19559,N_19365);
xnor U24123 (N_24123,N_15608,N_15993);
and U24124 (N_24124,N_16514,N_19729);
and U24125 (N_24125,N_15131,N_18329);
nor U24126 (N_24126,N_19140,N_16274);
nor U24127 (N_24127,N_17606,N_16537);
nand U24128 (N_24128,N_18135,N_15228);
and U24129 (N_24129,N_19668,N_15888);
and U24130 (N_24130,N_16013,N_16862);
and U24131 (N_24131,N_19118,N_16201);
nand U24132 (N_24132,N_16524,N_17429);
or U24133 (N_24133,N_19828,N_18545);
xor U24134 (N_24134,N_19445,N_15329);
or U24135 (N_24135,N_19034,N_18767);
and U24136 (N_24136,N_16450,N_15247);
nor U24137 (N_24137,N_17965,N_16072);
or U24138 (N_24138,N_19025,N_16807);
or U24139 (N_24139,N_18497,N_15154);
xnor U24140 (N_24140,N_17936,N_18036);
and U24141 (N_24141,N_15341,N_15622);
nor U24142 (N_24142,N_16751,N_19114);
or U24143 (N_24143,N_17334,N_17015);
xor U24144 (N_24144,N_15326,N_17311);
nor U24145 (N_24145,N_16496,N_16426);
or U24146 (N_24146,N_17715,N_16427);
and U24147 (N_24147,N_15933,N_16480);
and U24148 (N_24148,N_15910,N_16325);
or U24149 (N_24149,N_18882,N_15776);
and U24150 (N_24150,N_19221,N_19490);
nor U24151 (N_24151,N_17541,N_15674);
or U24152 (N_24152,N_17359,N_16076);
or U24153 (N_24153,N_18642,N_16069);
and U24154 (N_24154,N_18548,N_15262);
nand U24155 (N_24155,N_16451,N_18354);
and U24156 (N_24156,N_16483,N_18390);
and U24157 (N_24157,N_19320,N_19022);
and U24158 (N_24158,N_17609,N_16837);
nand U24159 (N_24159,N_17916,N_15358);
nor U24160 (N_24160,N_17948,N_17597);
or U24161 (N_24161,N_15580,N_15294);
and U24162 (N_24162,N_19657,N_16914);
nor U24163 (N_24163,N_15121,N_15485);
nor U24164 (N_24164,N_19105,N_16797);
or U24165 (N_24165,N_19082,N_17589);
xor U24166 (N_24166,N_16778,N_18128);
xor U24167 (N_24167,N_18669,N_15090);
nand U24168 (N_24168,N_19637,N_15304);
nor U24169 (N_24169,N_16896,N_15103);
nor U24170 (N_24170,N_18950,N_18112);
nand U24171 (N_24171,N_19095,N_17094);
nand U24172 (N_24172,N_16221,N_19956);
and U24173 (N_24173,N_18100,N_17022);
nor U24174 (N_24174,N_19337,N_19363);
xor U24175 (N_24175,N_18367,N_19849);
or U24176 (N_24176,N_17129,N_16185);
nand U24177 (N_24177,N_17476,N_16824);
xor U24178 (N_24178,N_18365,N_16727);
nand U24179 (N_24179,N_15002,N_19090);
xnor U24180 (N_24180,N_18997,N_15697);
nand U24181 (N_24181,N_19359,N_15999);
nand U24182 (N_24182,N_16164,N_16387);
xor U24183 (N_24183,N_15739,N_16542);
nand U24184 (N_24184,N_15737,N_17744);
xnor U24185 (N_24185,N_19609,N_16368);
nand U24186 (N_24186,N_15066,N_15252);
nand U24187 (N_24187,N_17530,N_16919);
nor U24188 (N_24188,N_15130,N_17331);
and U24189 (N_24189,N_18575,N_15184);
nand U24190 (N_24190,N_19318,N_18140);
nor U24191 (N_24191,N_19777,N_15789);
or U24192 (N_24192,N_18960,N_16216);
and U24193 (N_24193,N_17351,N_15283);
and U24194 (N_24194,N_16802,N_15253);
nor U24195 (N_24195,N_16732,N_19103);
nor U24196 (N_24196,N_17698,N_17953);
and U24197 (N_24197,N_17491,N_17646);
nand U24198 (N_24198,N_16925,N_17583);
or U24199 (N_24199,N_15990,N_19689);
or U24200 (N_24200,N_17549,N_19969);
and U24201 (N_24201,N_18673,N_16881);
nor U24202 (N_24202,N_16380,N_16693);
and U24203 (N_24203,N_15187,N_18732);
or U24204 (N_24204,N_18158,N_17964);
xor U24205 (N_24205,N_18569,N_17238);
and U24206 (N_24206,N_19918,N_16746);
nor U24207 (N_24207,N_16179,N_17058);
nor U24208 (N_24208,N_15708,N_19489);
and U24209 (N_24209,N_15982,N_15421);
and U24210 (N_24210,N_15606,N_15536);
and U24211 (N_24211,N_19078,N_17151);
and U24212 (N_24212,N_15038,N_19917);
and U24213 (N_24213,N_16558,N_16461);
or U24214 (N_24214,N_18161,N_16251);
xnor U24215 (N_24215,N_18549,N_19314);
or U24216 (N_24216,N_15245,N_17397);
or U24217 (N_24217,N_15526,N_15798);
nand U24218 (N_24218,N_17523,N_15310);
xor U24219 (N_24219,N_19704,N_18756);
nor U24220 (N_24220,N_16752,N_17327);
or U24221 (N_24221,N_19973,N_15686);
nor U24222 (N_24222,N_17279,N_19803);
xor U24223 (N_24223,N_15850,N_18912);
xnor U24224 (N_24224,N_15139,N_17317);
or U24225 (N_24225,N_19726,N_19272);
xnor U24226 (N_24226,N_15066,N_19517);
xnor U24227 (N_24227,N_18997,N_18674);
nand U24228 (N_24228,N_15602,N_15019);
xnor U24229 (N_24229,N_17919,N_16255);
and U24230 (N_24230,N_15915,N_18512);
nand U24231 (N_24231,N_19268,N_17939);
and U24232 (N_24232,N_15572,N_17939);
or U24233 (N_24233,N_18856,N_15233);
xnor U24234 (N_24234,N_18329,N_19407);
nor U24235 (N_24235,N_15081,N_16185);
nor U24236 (N_24236,N_18660,N_16844);
nor U24237 (N_24237,N_17318,N_17316);
xor U24238 (N_24238,N_19538,N_16382);
xor U24239 (N_24239,N_16466,N_16598);
or U24240 (N_24240,N_19215,N_15008);
nand U24241 (N_24241,N_17789,N_17099);
xor U24242 (N_24242,N_19173,N_19644);
nand U24243 (N_24243,N_18707,N_18037);
and U24244 (N_24244,N_16744,N_17445);
or U24245 (N_24245,N_18690,N_19828);
nand U24246 (N_24246,N_16892,N_17490);
and U24247 (N_24247,N_16522,N_15612);
or U24248 (N_24248,N_15436,N_17902);
or U24249 (N_24249,N_17364,N_15376);
and U24250 (N_24250,N_18782,N_16308);
or U24251 (N_24251,N_18462,N_17503);
or U24252 (N_24252,N_19935,N_16285);
xnor U24253 (N_24253,N_19691,N_19020);
and U24254 (N_24254,N_15554,N_16192);
xor U24255 (N_24255,N_17783,N_19844);
xor U24256 (N_24256,N_16859,N_16329);
nor U24257 (N_24257,N_15659,N_18082);
and U24258 (N_24258,N_17974,N_19465);
nor U24259 (N_24259,N_15719,N_15804);
nand U24260 (N_24260,N_17545,N_19003);
nor U24261 (N_24261,N_16399,N_16613);
nand U24262 (N_24262,N_16591,N_19621);
xnor U24263 (N_24263,N_17967,N_17389);
xor U24264 (N_24264,N_16126,N_17526);
xor U24265 (N_24265,N_16570,N_19757);
xor U24266 (N_24266,N_16094,N_18807);
nand U24267 (N_24267,N_15702,N_17918);
xnor U24268 (N_24268,N_15086,N_16484);
xor U24269 (N_24269,N_16331,N_17171);
or U24270 (N_24270,N_15674,N_16744);
and U24271 (N_24271,N_18666,N_17762);
nor U24272 (N_24272,N_19668,N_17848);
or U24273 (N_24273,N_15237,N_16031);
and U24274 (N_24274,N_16687,N_17287);
or U24275 (N_24275,N_15739,N_18743);
xnor U24276 (N_24276,N_19881,N_15908);
xor U24277 (N_24277,N_17692,N_16407);
xor U24278 (N_24278,N_19552,N_19360);
or U24279 (N_24279,N_15626,N_16008);
or U24280 (N_24280,N_19712,N_17506);
or U24281 (N_24281,N_18302,N_19147);
or U24282 (N_24282,N_15566,N_19110);
or U24283 (N_24283,N_19092,N_16587);
nand U24284 (N_24284,N_15059,N_17381);
or U24285 (N_24285,N_15536,N_18665);
or U24286 (N_24286,N_15059,N_15902);
and U24287 (N_24287,N_18361,N_15184);
nor U24288 (N_24288,N_16904,N_16040);
or U24289 (N_24289,N_18939,N_19555);
xnor U24290 (N_24290,N_19091,N_15986);
and U24291 (N_24291,N_15167,N_15776);
nand U24292 (N_24292,N_17780,N_17993);
nand U24293 (N_24293,N_19854,N_17027);
and U24294 (N_24294,N_16766,N_17099);
nor U24295 (N_24295,N_19619,N_16009);
nand U24296 (N_24296,N_16994,N_19942);
and U24297 (N_24297,N_15159,N_16271);
or U24298 (N_24298,N_18522,N_17477);
or U24299 (N_24299,N_19658,N_15141);
nand U24300 (N_24300,N_15007,N_17010);
xnor U24301 (N_24301,N_17715,N_18545);
nor U24302 (N_24302,N_18454,N_17267);
xnor U24303 (N_24303,N_19095,N_18616);
or U24304 (N_24304,N_18981,N_17169);
xnor U24305 (N_24305,N_16373,N_17500);
nor U24306 (N_24306,N_16706,N_15969);
and U24307 (N_24307,N_15522,N_17511);
xnor U24308 (N_24308,N_15193,N_17730);
or U24309 (N_24309,N_15397,N_15253);
xor U24310 (N_24310,N_15528,N_15415);
xnor U24311 (N_24311,N_15181,N_19626);
xnor U24312 (N_24312,N_15863,N_16270);
nor U24313 (N_24313,N_16315,N_17011);
and U24314 (N_24314,N_18629,N_15410);
or U24315 (N_24315,N_19277,N_17634);
nand U24316 (N_24316,N_16876,N_18918);
xor U24317 (N_24317,N_19815,N_19701);
nand U24318 (N_24318,N_15447,N_16449);
nand U24319 (N_24319,N_15686,N_19016);
nor U24320 (N_24320,N_19869,N_18440);
nor U24321 (N_24321,N_15104,N_19401);
nor U24322 (N_24322,N_15044,N_19905);
or U24323 (N_24323,N_15099,N_16922);
and U24324 (N_24324,N_15309,N_15737);
nand U24325 (N_24325,N_18772,N_16848);
xor U24326 (N_24326,N_19243,N_18941);
nand U24327 (N_24327,N_15637,N_17919);
nand U24328 (N_24328,N_16785,N_18747);
xnor U24329 (N_24329,N_19372,N_19949);
nor U24330 (N_24330,N_19314,N_15795);
xor U24331 (N_24331,N_18099,N_19915);
or U24332 (N_24332,N_16301,N_19690);
xnor U24333 (N_24333,N_18444,N_15246);
nand U24334 (N_24334,N_17718,N_15147);
or U24335 (N_24335,N_15068,N_16639);
or U24336 (N_24336,N_17284,N_15170);
and U24337 (N_24337,N_19495,N_18637);
or U24338 (N_24338,N_18285,N_19144);
and U24339 (N_24339,N_16748,N_15485);
nor U24340 (N_24340,N_19976,N_16854);
and U24341 (N_24341,N_17375,N_15890);
and U24342 (N_24342,N_16281,N_15139);
and U24343 (N_24343,N_19964,N_19150);
or U24344 (N_24344,N_18638,N_17192);
and U24345 (N_24345,N_17485,N_15366);
or U24346 (N_24346,N_16864,N_19351);
nand U24347 (N_24347,N_15107,N_19476);
nor U24348 (N_24348,N_18285,N_16390);
xor U24349 (N_24349,N_19163,N_18743);
and U24350 (N_24350,N_18867,N_15797);
and U24351 (N_24351,N_17053,N_19470);
or U24352 (N_24352,N_19080,N_19224);
or U24353 (N_24353,N_17485,N_19416);
nor U24354 (N_24354,N_17998,N_16645);
nand U24355 (N_24355,N_19100,N_18915);
nand U24356 (N_24356,N_18493,N_17699);
and U24357 (N_24357,N_19844,N_15400);
nand U24358 (N_24358,N_15046,N_17922);
or U24359 (N_24359,N_19677,N_16621);
nor U24360 (N_24360,N_16082,N_19630);
xnor U24361 (N_24361,N_16478,N_18149);
nor U24362 (N_24362,N_19722,N_17481);
and U24363 (N_24363,N_16657,N_18782);
and U24364 (N_24364,N_15386,N_18984);
and U24365 (N_24365,N_15457,N_15356);
and U24366 (N_24366,N_18647,N_17496);
or U24367 (N_24367,N_17528,N_17742);
or U24368 (N_24368,N_19199,N_16735);
and U24369 (N_24369,N_19795,N_17943);
nand U24370 (N_24370,N_17152,N_19609);
or U24371 (N_24371,N_15210,N_15234);
nor U24372 (N_24372,N_18463,N_19358);
xor U24373 (N_24373,N_18911,N_18408);
and U24374 (N_24374,N_19633,N_17049);
nor U24375 (N_24375,N_19216,N_15518);
xor U24376 (N_24376,N_15837,N_15084);
xnor U24377 (N_24377,N_18910,N_15316);
nor U24378 (N_24378,N_19143,N_18557);
and U24379 (N_24379,N_15561,N_16491);
xnor U24380 (N_24380,N_17760,N_15519);
nand U24381 (N_24381,N_15689,N_16564);
or U24382 (N_24382,N_16097,N_16415);
nand U24383 (N_24383,N_18820,N_16929);
or U24384 (N_24384,N_18485,N_19094);
xnor U24385 (N_24385,N_19159,N_19410);
xnor U24386 (N_24386,N_18080,N_19578);
xor U24387 (N_24387,N_18583,N_18507);
nand U24388 (N_24388,N_16156,N_15743);
nand U24389 (N_24389,N_19476,N_18584);
or U24390 (N_24390,N_17902,N_15636);
nor U24391 (N_24391,N_17643,N_17589);
or U24392 (N_24392,N_17102,N_18662);
or U24393 (N_24393,N_19378,N_15169);
or U24394 (N_24394,N_15234,N_18585);
nor U24395 (N_24395,N_16152,N_19216);
xor U24396 (N_24396,N_18370,N_19141);
xor U24397 (N_24397,N_18646,N_18466);
xor U24398 (N_24398,N_18740,N_17787);
or U24399 (N_24399,N_15789,N_15708);
and U24400 (N_24400,N_19763,N_16738);
or U24401 (N_24401,N_17139,N_18911);
nor U24402 (N_24402,N_18225,N_17826);
nor U24403 (N_24403,N_18667,N_17257);
nor U24404 (N_24404,N_17000,N_16452);
nor U24405 (N_24405,N_19680,N_17591);
nor U24406 (N_24406,N_15935,N_18360);
xnor U24407 (N_24407,N_16732,N_19190);
nand U24408 (N_24408,N_19086,N_15288);
nand U24409 (N_24409,N_16006,N_18699);
nor U24410 (N_24410,N_18548,N_19941);
and U24411 (N_24411,N_19591,N_15568);
nor U24412 (N_24412,N_19606,N_17809);
nor U24413 (N_24413,N_15609,N_17157);
nand U24414 (N_24414,N_17141,N_15537);
and U24415 (N_24415,N_17036,N_18268);
and U24416 (N_24416,N_17597,N_15640);
or U24417 (N_24417,N_18690,N_17333);
nor U24418 (N_24418,N_15962,N_19427);
xor U24419 (N_24419,N_17257,N_18004);
nand U24420 (N_24420,N_17974,N_19404);
and U24421 (N_24421,N_17507,N_19797);
xor U24422 (N_24422,N_19214,N_17408);
xnor U24423 (N_24423,N_19615,N_15007);
xor U24424 (N_24424,N_18126,N_16830);
nor U24425 (N_24425,N_18337,N_17385);
or U24426 (N_24426,N_15670,N_17611);
nand U24427 (N_24427,N_16280,N_17917);
xnor U24428 (N_24428,N_18244,N_16127);
or U24429 (N_24429,N_17866,N_19721);
nor U24430 (N_24430,N_19175,N_16596);
xnor U24431 (N_24431,N_17286,N_16598);
nor U24432 (N_24432,N_15064,N_15841);
xor U24433 (N_24433,N_18765,N_18139);
and U24434 (N_24434,N_19075,N_16204);
or U24435 (N_24435,N_18252,N_17445);
nand U24436 (N_24436,N_19405,N_16103);
nor U24437 (N_24437,N_18169,N_16597);
or U24438 (N_24438,N_19493,N_19525);
and U24439 (N_24439,N_16833,N_16115);
and U24440 (N_24440,N_18728,N_19067);
nand U24441 (N_24441,N_16852,N_18501);
or U24442 (N_24442,N_19665,N_15193);
xor U24443 (N_24443,N_19283,N_16344);
xor U24444 (N_24444,N_18542,N_15530);
or U24445 (N_24445,N_16012,N_18292);
or U24446 (N_24446,N_17925,N_18604);
xor U24447 (N_24447,N_19063,N_16161);
nor U24448 (N_24448,N_19023,N_18729);
xor U24449 (N_24449,N_16043,N_19290);
nor U24450 (N_24450,N_18221,N_17812);
or U24451 (N_24451,N_18607,N_16607);
xor U24452 (N_24452,N_19806,N_17186);
or U24453 (N_24453,N_19276,N_15845);
or U24454 (N_24454,N_19378,N_15080);
nor U24455 (N_24455,N_15744,N_17772);
and U24456 (N_24456,N_17873,N_17735);
xnor U24457 (N_24457,N_15190,N_18621);
nand U24458 (N_24458,N_19874,N_19805);
nand U24459 (N_24459,N_18171,N_17030);
xnor U24460 (N_24460,N_16518,N_18102);
xnor U24461 (N_24461,N_19408,N_17336);
nand U24462 (N_24462,N_15118,N_16940);
xnor U24463 (N_24463,N_16151,N_15216);
nor U24464 (N_24464,N_16989,N_16592);
nor U24465 (N_24465,N_15719,N_16300);
nor U24466 (N_24466,N_16337,N_16683);
nand U24467 (N_24467,N_15467,N_15704);
xor U24468 (N_24468,N_18105,N_16529);
or U24469 (N_24469,N_16011,N_15857);
or U24470 (N_24470,N_16054,N_19388);
xnor U24471 (N_24471,N_15508,N_17075);
nand U24472 (N_24472,N_17776,N_17358);
nand U24473 (N_24473,N_19598,N_19928);
and U24474 (N_24474,N_19101,N_17363);
nor U24475 (N_24475,N_16236,N_15268);
nand U24476 (N_24476,N_18238,N_17688);
and U24477 (N_24477,N_17324,N_15139);
or U24478 (N_24478,N_17138,N_15956);
nand U24479 (N_24479,N_18464,N_18977);
xor U24480 (N_24480,N_17034,N_17961);
and U24481 (N_24481,N_19381,N_15554);
nand U24482 (N_24482,N_17721,N_18949);
nor U24483 (N_24483,N_16296,N_18391);
or U24484 (N_24484,N_19090,N_16392);
nor U24485 (N_24485,N_19914,N_19985);
xor U24486 (N_24486,N_15758,N_16803);
xor U24487 (N_24487,N_19136,N_15877);
and U24488 (N_24488,N_18858,N_19172);
nor U24489 (N_24489,N_19151,N_17340);
nor U24490 (N_24490,N_15456,N_15998);
and U24491 (N_24491,N_17601,N_18087);
nor U24492 (N_24492,N_18530,N_18804);
nand U24493 (N_24493,N_18366,N_15697);
nand U24494 (N_24494,N_17413,N_19720);
nor U24495 (N_24495,N_17502,N_19934);
xor U24496 (N_24496,N_16646,N_15051);
xnor U24497 (N_24497,N_18430,N_15675);
nor U24498 (N_24498,N_17908,N_15675);
or U24499 (N_24499,N_19845,N_18184);
xnor U24500 (N_24500,N_16769,N_18412);
or U24501 (N_24501,N_19809,N_15824);
or U24502 (N_24502,N_19495,N_17406);
and U24503 (N_24503,N_19631,N_17177);
xor U24504 (N_24504,N_17295,N_17017);
or U24505 (N_24505,N_17258,N_17369);
nand U24506 (N_24506,N_15729,N_16016);
nand U24507 (N_24507,N_16153,N_16654);
and U24508 (N_24508,N_18609,N_17567);
and U24509 (N_24509,N_17202,N_16538);
or U24510 (N_24510,N_16317,N_16273);
and U24511 (N_24511,N_15590,N_15227);
and U24512 (N_24512,N_18141,N_19083);
nand U24513 (N_24513,N_16910,N_17972);
nor U24514 (N_24514,N_19449,N_17073);
xnor U24515 (N_24515,N_18271,N_15004);
xnor U24516 (N_24516,N_19166,N_18036);
or U24517 (N_24517,N_16638,N_18747);
xnor U24518 (N_24518,N_18850,N_15078);
xor U24519 (N_24519,N_18874,N_16096);
xor U24520 (N_24520,N_15160,N_19818);
nor U24521 (N_24521,N_15398,N_18326);
nand U24522 (N_24522,N_15655,N_17857);
and U24523 (N_24523,N_16967,N_18105);
or U24524 (N_24524,N_17381,N_16977);
and U24525 (N_24525,N_15969,N_17267);
nand U24526 (N_24526,N_18365,N_17302);
xnor U24527 (N_24527,N_15059,N_18226);
nor U24528 (N_24528,N_17379,N_16276);
nor U24529 (N_24529,N_17416,N_16468);
nand U24530 (N_24530,N_19482,N_19130);
nand U24531 (N_24531,N_17686,N_15655);
and U24532 (N_24532,N_16221,N_17176);
or U24533 (N_24533,N_16475,N_19477);
nor U24534 (N_24534,N_19853,N_15378);
xor U24535 (N_24535,N_18874,N_16033);
and U24536 (N_24536,N_16430,N_19902);
xor U24537 (N_24537,N_19228,N_17530);
or U24538 (N_24538,N_18296,N_16255);
nand U24539 (N_24539,N_17846,N_15791);
xor U24540 (N_24540,N_17926,N_18148);
nand U24541 (N_24541,N_18230,N_18904);
nor U24542 (N_24542,N_18575,N_15047);
nor U24543 (N_24543,N_19926,N_19094);
xnor U24544 (N_24544,N_17626,N_15339);
nand U24545 (N_24545,N_18873,N_18004);
nand U24546 (N_24546,N_15348,N_15163);
xnor U24547 (N_24547,N_17881,N_19888);
nor U24548 (N_24548,N_15658,N_16099);
and U24549 (N_24549,N_15542,N_17343);
nand U24550 (N_24550,N_15504,N_18532);
or U24551 (N_24551,N_17479,N_16040);
nor U24552 (N_24552,N_19817,N_15097);
and U24553 (N_24553,N_17132,N_18251);
nand U24554 (N_24554,N_17023,N_19510);
nand U24555 (N_24555,N_18918,N_15486);
or U24556 (N_24556,N_16415,N_17005);
xnor U24557 (N_24557,N_19621,N_17579);
xnor U24558 (N_24558,N_16311,N_15544);
nor U24559 (N_24559,N_17202,N_19729);
and U24560 (N_24560,N_15048,N_15303);
xnor U24561 (N_24561,N_18011,N_17230);
or U24562 (N_24562,N_16169,N_19798);
nor U24563 (N_24563,N_15695,N_16187);
nand U24564 (N_24564,N_19891,N_15766);
or U24565 (N_24565,N_18520,N_16896);
nor U24566 (N_24566,N_19280,N_16011);
xor U24567 (N_24567,N_17094,N_19408);
xor U24568 (N_24568,N_16000,N_15149);
nor U24569 (N_24569,N_18017,N_18992);
nand U24570 (N_24570,N_18251,N_16182);
or U24571 (N_24571,N_17465,N_18949);
nand U24572 (N_24572,N_18944,N_19909);
nor U24573 (N_24573,N_18815,N_17437);
nand U24574 (N_24574,N_18611,N_15589);
xor U24575 (N_24575,N_16203,N_17875);
nor U24576 (N_24576,N_19697,N_16092);
nor U24577 (N_24577,N_17486,N_19197);
nand U24578 (N_24578,N_15785,N_19929);
and U24579 (N_24579,N_16550,N_18435);
xnor U24580 (N_24580,N_19510,N_18167);
and U24581 (N_24581,N_19266,N_15841);
xor U24582 (N_24582,N_17649,N_15002);
or U24583 (N_24583,N_19653,N_19236);
and U24584 (N_24584,N_19191,N_17049);
or U24585 (N_24585,N_19112,N_17681);
or U24586 (N_24586,N_18594,N_17495);
nor U24587 (N_24587,N_16145,N_15398);
and U24588 (N_24588,N_19702,N_16543);
or U24589 (N_24589,N_19392,N_19640);
nor U24590 (N_24590,N_16984,N_18588);
nand U24591 (N_24591,N_18918,N_19172);
xnor U24592 (N_24592,N_17877,N_15603);
nor U24593 (N_24593,N_17584,N_19794);
or U24594 (N_24594,N_17851,N_16766);
nor U24595 (N_24595,N_19677,N_17411);
or U24596 (N_24596,N_19137,N_16618);
xnor U24597 (N_24597,N_16597,N_15915);
xnor U24598 (N_24598,N_18614,N_16818);
nor U24599 (N_24599,N_16866,N_18749);
nor U24600 (N_24600,N_19838,N_16263);
nand U24601 (N_24601,N_15832,N_15067);
xnor U24602 (N_24602,N_16033,N_16242);
nor U24603 (N_24603,N_19186,N_19865);
xnor U24604 (N_24604,N_19845,N_15204);
or U24605 (N_24605,N_19991,N_16051);
nand U24606 (N_24606,N_17060,N_18807);
or U24607 (N_24607,N_19395,N_19786);
nor U24608 (N_24608,N_16483,N_15053);
or U24609 (N_24609,N_16996,N_15869);
nor U24610 (N_24610,N_19087,N_19458);
nand U24611 (N_24611,N_16824,N_17624);
or U24612 (N_24612,N_15462,N_17962);
nand U24613 (N_24613,N_15840,N_17344);
xnor U24614 (N_24614,N_15805,N_17413);
xor U24615 (N_24615,N_15589,N_18225);
xor U24616 (N_24616,N_15754,N_18461);
and U24617 (N_24617,N_16847,N_16473);
xor U24618 (N_24618,N_16868,N_19731);
nor U24619 (N_24619,N_15532,N_18956);
nor U24620 (N_24620,N_17081,N_17226);
or U24621 (N_24621,N_17749,N_15503);
nor U24622 (N_24622,N_16603,N_15330);
nor U24623 (N_24623,N_16971,N_19631);
nor U24624 (N_24624,N_17204,N_15206);
and U24625 (N_24625,N_16372,N_15339);
and U24626 (N_24626,N_19755,N_17320);
and U24627 (N_24627,N_19112,N_19097);
nand U24628 (N_24628,N_15770,N_19410);
nand U24629 (N_24629,N_15531,N_19910);
or U24630 (N_24630,N_17263,N_15442);
nor U24631 (N_24631,N_17723,N_16984);
nand U24632 (N_24632,N_15489,N_18557);
or U24633 (N_24633,N_18504,N_16820);
or U24634 (N_24634,N_17644,N_18181);
and U24635 (N_24635,N_18756,N_16627);
and U24636 (N_24636,N_16605,N_15671);
xor U24637 (N_24637,N_15930,N_19256);
and U24638 (N_24638,N_17280,N_18738);
nor U24639 (N_24639,N_19772,N_18772);
xnor U24640 (N_24640,N_19997,N_16255);
or U24641 (N_24641,N_19626,N_16705);
xor U24642 (N_24642,N_16832,N_16175);
xnor U24643 (N_24643,N_18082,N_15774);
nand U24644 (N_24644,N_19281,N_19185);
or U24645 (N_24645,N_15839,N_16930);
xor U24646 (N_24646,N_17430,N_16173);
and U24647 (N_24647,N_18247,N_18417);
xnor U24648 (N_24648,N_19104,N_19830);
xnor U24649 (N_24649,N_15331,N_17768);
xor U24650 (N_24650,N_19327,N_15904);
or U24651 (N_24651,N_16820,N_15196);
nor U24652 (N_24652,N_19882,N_19527);
or U24653 (N_24653,N_15449,N_16280);
or U24654 (N_24654,N_15142,N_15380);
and U24655 (N_24655,N_16267,N_17906);
and U24656 (N_24656,N_19215,N_15227);
nand U24657 (N_24657,N_15248,N_16080);
or U24658 (N_24658,N_15273,N_19686);
xnor U24659 (N_24659,N_17602,N_16486);
and U24660 (N_24660,N_15024,N_15740);
and U24661 (N_24661,N_15408,N_17315);
nor U24662 (N_24662,N_15762,N_18325);
nand U24663 (N_24663,N_17691,N_15961);
or U24664 (N_24664,N_18589,N_17208);
or U24665 (N_24665,N_15176,N_17763);
or U24666 (N_24666,N_19238,N_19854);
nor U24667 (N_24667,N_19239,N_18426);
xor U24668 (N_24668,N_18280,N_18185);
nor U24669 (N_24669,N_15503,N_17009);
or U24670 (N_24670,N_19102,N_17176);
nor U24671 (N_24671,N_15868,N_15458);
nor U24672 (N_24672,N_18431,N_19298);
xor U24673 (N_24673,N_16425,N_17283);
or U24674 (N_24674,N_17592,N_16195);
xor U24675 (N_24675,N_17593,N_19784);
and U24676 (N_24676,N_19501,N_17889);
nor U24677 (N_24677,N_15365,N_18745);
xor U24678 (N_24678,N_16047,N_18341);
nor U24679 (N_24679,N_19533,N_16578);
nand U24680 (N_24680,N_19967,N_17973);
nand U24681 (N_24681,N_19520,N_17576);
nor U24682 (N_24682,N_19143,N_16141);
or U24683 (N_24683,N_17059,N_19128);
xnor U24684 (N_24684,N_17522,N_15017);
xnor U24685 (N_24685,N_16841,N_15038);
xnor U24686 (N_24686,N_18984,N_15303);
or U24687 (N_24687,N_18742,N_19087);
or U24688 (N_24688,N_18593,N_16684);
xnor U24689 (N_24689,N_15080,N_19674);
xnor U24690 (N_24690,N_17361,N_16676);
nor U24691 (N_24691,N_17505,N_15895);
nor U24692 (N_24692,N_17271,N_16953);
or U24693 (N_24693,N_16492,N_15182);
nor U24694 (N_24694,N_15757,N_18907);
nand U24695 (N_24695,N_19130,N_19322);
nor U24696 (N_24696,N_19334,N_16246);
and U24697 (N_24697,N_18973,N_17431);
nor U24698 (N_24698,N_16410,N_15515);
xor U24699 (N_24699,N_17692,N_18924);
or U24700 (N_24700,N_19684,N_16267);
and U24701 (N_24701,N_19740,N_17062);
xor U24702 (N_24702,N_17148,N_17874);
or U24703 (N_24703,N_19446,N_18445);
nand U24704 (N_24704,N_16467,N_16709);
nor U24705 (N_24705,N_19093,N_16384);
nor U24706 (N_24706,N_19776,N_18240);
xor U24707 (N_24707,N_16208,N_18648);
nor U24708 (N_24708,N_18716,N_19687);
nand U24709 (N_24709,N_16574,N_15689);
or U24710 (N_24710,N_17091,N_15266);
and U24711 (N_24711,N_15428,N_17437);
nand U24712 (N_24712,N_18865,N_15216);
or U24713 (N_24713,N_19653,N_15676);
or U24714 (N_24714,N_19446,N_17113);
and U24715 (N_24715,N_19655,N_17690);
nor U24716 (N_24716,N_17785,N_18031);
nor U24717 (N_24717,N_17369,N_17051);
or U24718 (N_24718,N_18539,N_16821);
nor U24719 (N_24719,N_18350,N_15394);
and U24720 (N_24720,N_15841,N_16589);
xnor U24721 (N_24721,N_18154,N_17513);
or U24722 (N_24722,N_15103,N_16837);
and U24723 (N_24723,N_16186,N_17053);
nor U24724 (N_24724,N_16505,N_17053);
nor U24725 (N_24725,N_17771,N_17628);
or U24726 (N_24726,N_18885,N_15304);
nand U24727 (N_24727,N_15041,N_16327);
xor U24728 (N_24728,N_17372,N_16161);
nor U24729 (N_24729,N_18793,N_19084);
nand U24730 (N_24730,N_17087,N_15338);
xor U24731 (N_24731,N_18635,N_15016);
and U24732 (N_24732,N_18718,N_17508);
or U24733 (N_24733,N_15452,N_19532);
and U24734 (N_24734,N_15640,N_17126);
nand U24735 (N_24735,N_17058,N_16684);
xnor U24736 (N_24736,N_19618,N_19491);
or U24737 (N_24737,N_16900,N_15263);
and U24738 (N_24738,N_15502,N_15769);
nor U24739 (N_24739,N_16890,N_16995);
or U24740 (N_24740,N_15180,N_15454);
nand U24741 (N_24741,N_17697,N_18556);
and U24742 (N_24742,N_18876,N_18836);
xor U24743 (N_24743,N_17957,N_15555);
and U24744 (N_24744,N_15927,N_18831);
nor U24745 (N_24745,N_15742,N_18672);
and U24746 (N_24746,N_18913,N_18315);
and U24747 (N_24747,N_19149,N_18381);
or U24748 (N_24748,N_17266,N_16882);
nor U24749 (N_24749,N_19818,N_17229);
xor U24750 (N_24750,N_16950,N_19878);
or U24751 (N_24751,N_17276,N_19784);
nand U24752 (N_24752,N_16856,N_15993);
nor U24753 (N_24753,N_15239,N_17675);
xnor U24754 (N_24754,N_16035,N_16975);
xor U24755 (N_24755,N_17072,N_15739);
and U24756 (N_24756,N_19882,N_18162);
and U24757 (N_24757,N_18283,N_18973);
and U24758 (N_24758,N_19968,N_18364);
or U24759 (N_24759,N_15177,N_16663);
nor U24760 (N_24760,N_18775,N_18655);
nor U24761 (N_24761,N_17413,N_17479);
xor U24762 (N_24762,N_16496,N_15071);
nand U24763 (N_24763,N_19996,N_15119);
or U24764 (N_24764,N_19596,N_18690);
nand U24765 (N_24765,N_15680,N_16896);
and U24766 (N_24766,N_15609,N_17209);
nor U24767 (N_24767,N_17196,N_16437);
nand U24768 (N_24768,N_15911,N_19671);
nand U24769 (N_24769,N_15217,N_17374);
or U24770 (N_24770,N_18613,N_15023);
or U24771 (N_24771,N_18671,N_16472);
nor U24772 (N_24772,N_16846,N_15440);
xor U24773 (N_24773,N_18621,N_18085);
xnor U24774 (N_24774,N_15390,N_16369);
xnor U24775 (N_24775,N_16647,N_16063);
and U24776 (N_24776,N_19450,N_18526);
and U24777 (N_24777,N_19300,N_19175);
and U24778 (N_24778,N_17495,N_19321);
nand U24779 (N_24779,N_16556,N_18362);
nor U24780 (N_24780,N_18335,N_16887);
xnor U24781 (N_24781,N_19355,N_18503);
nor U24782 (N_24782,N_19200,N_19876);
or U24783 (N_24783,N_16937,N_15097);
or U24784 (N_24784,N_18781,N_16775);
xor U24785 (N_24785,N_18267,N_15979);
nand U24786 (N_24786,N_16942,N_16725);
nor U24787 (N_24787,N_18055,N_18088);
nor U24788 (N_24788,N_15162,N_17243);
xnor U24789 (N_24789,N_18234,N_17785);
xnor U24790 (N_24790,N_16769,N_15368);
nand U24791 (N_24791,N_19691,N_17664);
nand U24792 (N_24792,N_19230,N_18896);
nor U24793 (N_24793,N_18062,N_16677);
xor U24794 (N_24794,N_18721,N_18890);
nand U24795 (N_24795,N_18234,N_15053);
or U24796 (N_24796,N_19724,N_19839);
nor U24797 (N_24797,N_19006,N_15468);
xnor U24798 (N_24798,N_16334,N_18876);
nor U24799 (N_24799,N_15204,N_16726);
xor U24800 (N_24800,N_18863,N_19445);
nand U24801 (N_24801,N_17390,N_17208);
nor U24802 (N_24802,N_15929,N_17225);
and U24803 (N_24803,N_16273,N_18541);
nand U24804 (N_24804,N_18780,N_16264);
nor U24805 (N_24805,N_19300,N_18461);
or U24806 (N_24806,N_18486,N_19956);
xor U24807 (N_24807,N_18251,N_17537);
and U24808 (N_24808,N_16994,N_15890);
nand U24809 (N_24809,N_15633,N_16807);
or U24810 (N_24810,N_17773,N_17316);
and U24811 (N_24811,N_19877,N_17811);
and U24812 (N_24812,N_16680,N_18951);
nor U24813 (N_24813,N_19840,N_17163);
xnor U24814 (N_24814,N_16029,N_19407);
and U24815 (N_24815,N_15700,N_18876);
or U24816 (N_24816,N_15591,N_19127);
nand U24817 (N_24817,N_18921,N_19482);
and U24818 (N_24818,N_15174,N_17322);
or U24819 (N_24819,N_17560,N_15016);
xnor U24820 (N_24820,N_19209,N_18747);
nand U24821 (N_24821,N_16494,N_16760);
or U24822 (N_24822,N_18097,N_17381);
nand U24823 (N_24823,N_15309,N_19750);
or U24824 (N_24824,N_18330,N_17534);
nor U24825 (N_24825,N_16657,N_19733);
and U24826 (N_24826,N_18463,N_15357);
xnor U24827 (N_24827,N_15100,N_19707);
and U24828 (N_24828,N_15781,N_15415);
xnor U24829 (N_24829,N_19148,N_18528);
nand U24830 (N_24830,N_18045,N_17607);
and U24831 (N_24831,N_17729,N_15949);
xor U24832 (N_24832,N_16559,N_16595);
xor U24833 (N_24833,N_18973,N_16037);
and U24834 (N_24834,N_17757,N_15874);
or U24835 (N_24835,N_18158,N_15111);
nand U24836 (N_24836,N_15705,N_17983);
nand U24837 (N_24837,N_16226,N_16303);
xnor U24838 (N_24838,N_18542,N_15578);
or U24839 (N_24839,N_16556,N_18497);
nor U24840 (N_24840,N_17906,N_18461);
nand U24841 (N_24841,N_16827,N_17967);
and U24842 (N_24842,N_16859,N_15559);
xor U24843 (N_24843,N_15389,N_16101);
or U24844 (N_24844,N_16313,N_16897);
and U24845 (N_24845,N_15342,N_18746);
xnor U24846 (N_24846,N_17117,N_19290);
nand U24847 (N_24847,N_17492,N_16882);
nand U24848 (N_24848,N_18081,N_18946);
or U24849 (N_24849,N_16784,N_16918);
and U24850 (N_24850,N_18428,N_16558);
and U24851 (N_24851,N_18237,N_17128);
xnor U24852 (N_24852,N_17240,N_15663);
nor U24853 (N_24853,N_17455,N_18946);
nand U24854 (N_24854,N_15594,N_19962);
or U24855 (N_24855,N_18665,N_16949);
and U24856 (N_24856,N_17778,N_17528);
or U24857 (N_24857,N_17077,N_19248);
xnor U24858 (N_24858,N_17850,N_17610);
and U24859 (N_24859,N_16498,N_16348);
or U24860 (N_24860,N_16932,N_19772);
nand U24861 (N_24861,N_17096,N_18813);
or U24862 (N_24862,N_18342,N_16523);
xnor U24863 (N_24863,N_17103,N_19908);
xnor U24864 (N_24864,N_19585,N_17698);
and U24865 (N_24865,N_18831,N_15214);
xnor U24866 (N_24866,N_16874,N_16911);
and U24867 (N_24867,N_16203,N_15669);
and U24868 (N_24868,N_16965,N_18477);
nor U24869 (N_24869,N_15707,N_15865);
or U24870 (N_24870,N_17623,N_15863);
or U24871 (N_24871,N_19565,N_17471);
nor U24872 (N_24872,N_15369,N_16859);
or U24873 (N_24873,N_19813,N_15971);
xnor U24874 (N_24874,N_17239,N_17790);
nand U24875 (N_24875,N_15054,N_18136);
or U24876 (N_24876,N_17163,N_19449);
and U24877 (N_24877,N_18876,N_18067);
nor U24878 (N_24878,N_15864,N_15701);
xor U24879 (N_24879,N_18966,N_17237);
nor U24880 (N_24880,N_15847,N_17885);
or U24881 (N_24881,N_18877,N_17436);
xnor U24882 (N_24882,N_15921,N_15991);
or U24883 (N_24883,N_19975,N_16955);
xor U24884 (N_24884,N_16370,N_15902);
and U24885 (N_24885,N_19402,N_18867);
nor U24886 (N_24886,N_15332,N_15383);
nand U24887 (N_24887,N_18691,N_18897);
and U24888 (N_24888,N_15988,N_19538);
xnor U24889 (N_24889,N_19934,N_18859);
nor U24890 (N_24890,N_18892,N_17124);
and U24891 (N_24891,N_17599,N_15998);
and U24892 (N_24892,N_17287,N_16349);
xnor U24893 (N_24893,N_15487,N_18056);
or U24894 (N_24894,N_15495,N_19801);
nor U24895 (N_24895,N_16188,N_15774);
nor U24896 (N_24896,N_19227,N_18108);
or U24897 (N_24897,N_19183,N_15480);
and U24898 (N_24898,N_16960,N_15605);
and U24899 (N_24899,N_16267,N_18508);
and U24900 (N_24900,N_15871,N_18049);
xnor U24901 (N_24901,N_15008,N_17720);
xor U24902 (N_24902,N_18981,N_19194);
xor U24903 (N_24903,N_18392,N_16977);
nor U24904 (N_24904,N_19192,N_18785);
xor U24905 (N_24905,N_15054,N_16362);
and U24906 (N_24906,N_15611,N_16970);
nor U24907 (N_24907,N_19890,N_15206);
and U24908 (N_24908,N_16935,N_18110);
xor U24909 (N_24909,N_15352,N_19379);
or U24910 (N_24910,N_16060,N_15849);
nor U24911 (N_24911,N_18032,N_17521);
or U24912 (N_24912,N_18103,N_15036);
or U24913 (N_24913,N_15781,N_17913);
nand U24914 (N_24914,N_15282,N_17068);
nor U24915 (N_24915,N_19442,N_18083);
nand U24916 (N_24916,N_17953,N_19735);
and U24917 (N_24917,N_19410,N_15068);
nor U24918 (N_24918,N_17223,N_15337);
and U24919 (N_24919,N_16333,N_16021);
nor U24920 (N_24920,N_18086,N_16820);
xnor U24921 (N_24921,N_17897,N_17458);
and U24922 (N_24922,N_16458,N_16469);
nand U24923 (N_24923,N_19368,N_19978);
xnor U24924 (N_24924,N_17379,N_17407);
nor U24925 (N_24925,N_19658,N_15721);
or U24926 (N_24926,N_17242,N_16291);
nand U24927 (N_24927,N_17429,N_17431);
or U24928 (N_24928,N_17459,N_15537);
xor U24929 (N_24929,N_16036,N_16729);
nand U24930 (N_24930,N_19984,N_18023);
nor U24931 (N_24931,N_19801,N_19073);
and U24932 (N_24932,N_18456,N_18372);
nor U24933 (N_24933,N_15084,N_18603);
nand U24934 (N_24934,N_16653,N_17442);
or U24935 (N_24935,N_16076,N_15052);
xor U24936 (N_24936,N_17688,N_19040);
xnor U24937 (N_24937,N_18398,N_17227);
or U24938 (N_24938,N_15441,N_15927);
or U24939 (N_24939,N_16625,N_19475);
nand U24940 (N_24940,N_17839,N_19200);
nor U24941 (N_24941,N_19573,N_15936);
and U24942 (N_24942,N_16127,N_15616);
and U24943 (N_24943,N_16330,N_19347);
and U24944 (N_24944,N_18019,N_16678);
xor U24945 (N_24945,N_15481,N_15368);
xnor U24946 (N_24946,N_18624,N_15290);
and U24947 (N_24947,N_18935,N_19875);
nor U24948 (N_24948,N_18639,N_16660);
or U24949 (N_24949,N_17623,N_17755);
xnor U24950 (N_24950,N_16511,N_18515);
nor U24951 (N_24951,N_19539,N_19651);
nor U24952 (N_24952,N_19304,N_18916);
xor U24953 (N_24953,N_17674,N_17762);
and U24954 (N_24954,N_18121,N_15479);
nand U24955 (N_24955,N_19564,N_18780);
nand U24956 (N_24956,N_19789,N_17305);
nand U24957 (N_24957,N_15718,N_16877);
and U24958 (N_24958,N_19985,N_19804);
and U24959 (N_24959,N_15242,N_16172);
xor U24960 (N_24960,N_15336,N_15803);
nand U24961 (N_24961,N_19161,N_15681);
and U24962 (N_24962,N_17500,N_18392);
or U24963 (N_24963,N_16850,N_15967);
xor U24964 (N_24964,N_15270,N_16465);
nor U24965 (N_24965,N_18939,N_18866);
and U24966 (N_24966,N_18461,N_18736);
nand U24967 (N_24967,N_16283,N_19645);
xnor U24968 (N_24968,N_18607,N_15734);
nor U24969 (N_24969,N_18356,N_17451);
or U24970 (N_24970,N_16992,N_16086);
and U24971 (N_24971,N_17676,N_18771);
or U24972 (N_24972,N_17590,N_16072);
and U24973 (N_24973,N_18172,N_16731);
xor U24974 (N_24974,N_19309,N_18050);
nor U24975 (N_24975,N_15671,N_19026);
and U24976 (N_24976,N_17621,N_18824);
nor U24977 (N_24977,N_18218,N_18401);
and U24978 (N_24978,N_16573,N_17188);
xnor U24979 (N_24979,N_16718,N_19578);
xor U24980 (N_24980,N_15744,N_17061);
or U24981 (N_24981,N_16741,N_19474);
nor U24982 (N_24982,N_18587,N_18656);
or U24983 (N_24983,N_18690,N_16015);
xor U24984 (N_24984,N_19822,N_15978);
xnor U24985 (N_24985,N_19690,N_17542);
and U24986 (N_24986,N_17961,N_19823);
nand U24987 (N_24987,N_16077,N_17653);
nand U24988 (N_24988,N_19568,N_18915);
and U24989 (N_24989,N_15371,N_18717);
nand U24990 (N_24990,N_16117,N_18560);
and U24991 (N_24991,N_15795,N_15558);
nor U24992 (N_24992,N_19618,N_18803);
or U24993 (N_24993,N_18006,N_17250);
and U24994 (N_24994,N_18048,N_19932);
nand U24995 (N_24995,N_19225,N_19323);
xnor U24996 (N_24996,N_15349,N_17944);
nor U24997 (N_24997,N_19694,N_17808);
xnor U24998 (N_24998,N_17827,N_19995);
or U24999 (N_24999,N_18683,N_19510);
and U25000 (N_25000,N_24985,N_24816);
and U25001 (N_25001,N_23748,N_23631);
nor U25002 (N_25002,N_20321,N_22729);
xnor U25003 (N_25003,N_22973,N_24505);
nand U25004 (N_25004,N_24690,N_22850);
nand U25005 (N_25005,N_23227,N_21470);
nand U25006 (N_25006,N_23970,N_21310);
and U25007 (N_25007,N_24819,N_24008);
nor U25008 (N_25008,N_20336,N_21489);
nor U25009 (N_25009,N_24097,N_21085);
and U25010 (N_25010,N_20348,N_22263);
nand U25011 (N_25011,N_20258,N_20666);
nor U25012 (N_25012,N_24462,N_22976);
nor U25013 (N_25013,N_22943,N_21645);
or U25014 (N_25014,N_20057,N_24770);
or U25015 (N_25015,N_21833,N_24026);
and U25016 (N_25016,N_21118,N_24879);
and U25017 (N_25017,N_20520,N_23729);
nor U25018 (N_25018,N_23542,N_22359);
nor U25019 (N_25019,N_20072,N_21854);
nor U25020 (N_25020,N_24253,N_22388);
or U25021 (N_25021,N_20964,N_21652);
and U25022 (N_25022,N_22327,N_20312);
or U25023 (N_25023,N_24906,N_23098);
xor U25024 (N_25024,N_22269,N_20712);
nor U25025 (N_25025,N_21122,N_20539);
or U25026 (N_25026,N_20077,N_21597);
nand U25027 (N_25027,N_20836,N_24521);
xor U25028 (N_25028,N_21098,N_20103);
nand U25029 (N_25029,N_23440,N_20904);
and U25030 (N_25030,N_22339,N_24749);
xnor U25031 (N_25031,N_21314,N_21982);
xnor U25032 (N_25032,N_24017,N_24844);
or U25033 (N_25033,N_20415,N_20105);
nand U25034 (N_25034,N_20531,N_20014);
and U25035 (N_25035,N_24832,N_24109);
nand U25036 (N_25036,N_23708,N_23630);
and U25037 (N_25037,N_21447,N_22271);
nand U25038 (N_25038,N_22362,N_20365);
nand U25039 (N_25039,N_23129,N_23859);
nand U25040 (N_25040,N_24110,N_21491);
nor U25041 (N_25041,N_23716,N_20062);
nand U25042 (N_25042,N_22354,N_20085);
nor U25043 (N_25043,N_24227,N_23459);
and U25044 (N_25044,N_21146,N_20752);
and U25045 (N_25045,N_22533,N_21378);
nand U25046 (N_25046,N_21550,N_20182);
xnor U25047 (N_25047,N_24432,N_24422);
and U25048 (N_25048,N_23948,N_21772);
xor U25049 (N_25049,N_22617,N_23502);
nor U25050 (N_25050,N_22484,N_20601);
or U25051 (N_25051,N_20777,N_20392);
and U25052 (N_25052,N_23993,N_22952);
and U25053 (N_25053,N_23787,N_24986);
and U25054 (N_25054,N_23928,N_21835);
nand U25055 (N_25055,N_22471,N_23485);
or U25056 (N_25056,N_21104,N_23964);
or U25057 (N_25057,N_21192,N_22261);
or U25058 (N_25058,N_22136,N_22657);
nor U25059 (N_25059,N_22485,N_23403);
and U25060 (N_25060,N_24914,N_20656);
nor U25061 (N_25061,N_23963,N_22308);
nor U25062 (N_25062,N_20221,N_23126);
and U25063 (N_25063,N_24936,N_22955);
nand U25064 (N_25064,N_21025,N_20892);
nand U25065 (N_25065,N_22857,N_22515);
or U25066 (N_25066,N_24774,N_22065);
or U25067 (N_25067,N_20242,N_20687);
nand U25068 (N_25068,N_24766,N_20146);
nand U25069 (N_25069,N_23395,N_24988);
xor U25070 (N_25070,N_22145,N_20201);
nor U25071 (N_25071,N_21700,N_23333);
or U25072 (N_25072,N_22814,N_23592);
and U25073 (N_25073,N_21404,N_24741);
and U25074 (N_25074,N_23105,N_22512);
and U25075 (N_25075,N_24778,N_22006);
nand U25076 (N_25076,N_20208,N_20993);
or U25077 (N_25077,N_21548,N_24417);
or U25078 (N_25078,N_20556,N_24689);
nor U25079 (N_25079,N_23558,N_23419);
xor U25080 (N_25080,N_22525,N_23524);
and U25081 (N_25081,N_24859,N_22299);
nor U25082 (N_25082,N_24365,N_20330);
nand U25083 (N_25083,N_24238,N_24686);
and U25084 (N_25084,N_20311,N_24871);
nand U25085 (N_25085,N_22808,N_22004);
and U25086 (N_25086,N_20517,N_20740);
and U25087 (N_25087,N_23140,N_22390);
xnor U25088 (N_25088,N_23275,N_24501);
or U25089 (N_25089,N_20518,N_20716);
nand U25090 (N_25090,N_23173,N_24272);
xnor U25091 (N_25091,N_20549,N_24362);
and U25092 (N_25092,N_22750,N_20200);
nor U25093 (N_25093,N_23297,N_22555);
nand U25094 (N_25094,N_22612,N_22405);
or U25095 (N_25095,N_24033,N_23516);
nand U25096 (N_25096,N_24918,N_20481);
nand U25097 (N_25097,N_24642,N_22895);
nand U25098 (N_25098,N_23842,N_24604);
or U25099 (N_25099,N_20043,N_22904);
nand U25100 (N_25100,N_23888,N_24948);
and U25101 (N_25101,N_24546,N_21091);
and U25102 (N_25102,N_24554,N_20009);
nor U25103 (N_25103,N_21893,N_24301);
or U25104 (N_25104,N_22276,N_23474);
nor U25105 (N_25105,N_24153,N_24876);
nand U25106 (N_25106,N_21620,N_21115);
nand U25107 (N_25107,N_21871,N_21302);
xor U25108 (N_25108,N_21913,N_24128);
or U25109 (N_25109,N_20135,N_20432);
nand U25110 (N_25110,N_24565,N_22012);
nand U25111 (N_25111,N_23322,N_24754);
and U25112 (N_25112,N_23118,N_22113);
xnor U25113 (N_25113,N_20960,N_24015);
xor U25114 (N_25114,N_24336,N_23903);
or U25115 (N_25115,N_21441,N_21509);
and U25116 (N_25116,N_24675,N_24477);
xor U25117 (N_25117,N_20835,N_21094);
nor U25118 (N_25118,N_21594,N_24573);
nor U25119 (N_25119,N_23229,N_22459);
xor U25120 (N_25120,N_24898,N_22165);
xnor U25121 (N_25121,N_24994,N_22310);
or U25122 (N_25122,N_24930,N_20820);
nand U25123 (N_25123,N_21572,N_20143);
nand U25124 (N_25124,N_23498,N_22461);
and U25125 (N_25125,N_20529,N_20924);
or U25126 (N_25126,N_23804,N_21939);
nor U25127 (N_25127,N_21328,N_20231);
nand U25128 (N_25128,N_23201,N_23839);
nand U25129 (N_25129,N_20025,N_22081);
xnor U25130 (N_25130,N_21464,N_23441);
xnor U25131 (N_25131,N_20262,N_22279);
nor U25132 (N_25132,N_24562,N_21512);
or U25133 (N_25133,N_20339,N_21945);
nor U25134 (N_25134,N_21420,N_20660);
nand U25135 (N_25135,N_20535,N_21671);
or U25136 (N_25136,N_22789,N_24959);
or U25137 (N_25137,N_21380,N_22598);
nand U25138 (N_25138,N_20615,N_20706);
nor U25139 (N_25139,N_23230,N_21087);
nand U25140 (N_25140,N_24455,N_20466);
nand U25141 (N_25141,N_23503,N_20923);
xnor U25142 (N_25142,N_24529,N_21475);
and U25143 (N_25143,N_20408,N_20310);
and U25144 (N_25144,N_23973,N_23810);
xor U25145 (N_25145,N_24831,N_23952);
nor U25146 (N_25146,N_20910,N_22409);
or U25147 (N_25147,N_21851,N_24144);
and U25148 (N_25148,N_21775,N_20497);
nand U25149 (N_25149,N_21354,N_23185);
or U25150 (N_25150,N_21458,N_21413);
nand U25151 (N_25151,N_20824,N_21804);
and U25152 (N_25152,N_24108,N_22051);
and U25153 (N_25153,N_22511,N_22643);
or U25154 (N_25154,N_20436,N_22882);
xor U25155 (N_25155,N_21181,N_21957);
or U25156 (N_25156,N_20176,N_22684);
xnor U25157 (N_25157,N_21587,N_21824);
or U25158 (N_25158,N_21865,N_21735);
xnor U25159 (N_25159,N_21051,N_22840);
and U25160 (N_25160,N_24345,N_24276);
nor U25161 (N_25161,N_21030,N_21435);
nor U25162 (N_25162,N_22671,N_24273);
nor U25163 (N_25163,N_24240,N_20915);
and U25164 (N_25164,N_24528,N_20902);
nand U25165 (N_25165,N_21558,N_21371);
nand U25166 (N_25166,N_23217,N_20796);
xor U25167 (N_25167,N_22947,N_21717);
nor U25168 (N_25168,N_22000,N_24897);
xnor U25169 (N_25169,N_23056,N_21480);
nand U25170 (N_25170,N_20050,N_24192);
or U25171 (N_25171,N_21336,N_23020);
xnor U25172 (N_25172,N_20872,N_21954);
xor U25173 (N_25173,N_24349,N_23417);
and U25174 (N_25174,N_23966,N_22008);
or U25175 (N_25175,N_20477,N_21638);
nor U25176 (N_25176,N_21670,N_22198);
nor U25177 (N_25177,N_23041,N_22188);
nand U25178 (N_25178,N_20921,N_22727);
or U25179 (N_25179,N_21061,N_22394);
xor U25180 (N_25180,N_24834,N_22924);
nor U25181 (N_25181,N_24630,N_24090);
and U25182 (N_25182,N_23747,N_21100);
or U25183 (N_25183,N_21204,N_20111);
and U25184 (N_25184,N_24025,N_24550);
or U25185 (N_25185,N_20770,N_22007);
and U25186 (N_25186,N_21217,N_22697);
or U25187 (N_25187,N_23366,N_24408);
xor U25188 (N_25188,N_21516,N_23865);
nand U25189 (N_25189,N_22427,N_23458);
nor U25190 (N_25190,N_20616,N_22067);
or U25191 (N_25191,N_24329,N_21171);
or U25192 (N_25192,N_24862,N_24924);
xor U25193 (N_25193,N_22756,N_22175);
nor U25194 (N_25194,N_24137,N_24639);
or U25195 (N_25195,N_21578,N_24036);
xnor U25196 (N_25196,N_24631,N_20744);
xnor U25197 (N_25197,N_21968,N_21964);
nor U25198 (N_25198,N_21860,N_21570);
nor U25199 (N_25199,N_20426,N_22798);
nand U25200 (N_25200,N_23734,N_24139);
and U25201 (N_25201,N_22606,N_21052);
and U25202 (N_25202,N_22329,N_24698);
xor U25203 (N_25203,N_20949,N_20070);
nand U25204 (N_25204,N_21333,N_20459);
nor U25205 (N_25205,N_24552,N_22738);
and U25206 (N_25206,N_21451,N_21669);
xor U25207 (N_25207,N_21569,N_24467);
or U25208 (N_25208,N_20505,N_21478);
or U25209 (N_25209,N_22181,N_21842);
nand U25210 (N_25210,N_22824,N_21600);
nand U25211 (N_25211,N_21285,N_21011);
xor U25212 (N_25212,N_22849,N_22040);
xor U25213 (N_25213,N_22066,N_21158);
or U25214 (N_25214,N_23142,N_20044);
and U25215 (N_25215,N_23713,N_24045);
nor U25216 (N_25216,N_20418,N_20906);
nor U25217 (N_25217,N_21015,N_24743);
nand U25218 (N_25218,N_21143,N_24849);
nor U25219 (N_25219,N_20711,N_20975);
or U25220 (N_25220,N_20457,N_23326);
or U25221 (N_25221,N_24629,N_22831);
xnor U25222 (N_25222,N_22477,N_20771);
and U25223 (N_25223,N_21004,N_22349);
xnor U25224 (N_25224,N_22043,N_23397);
or U25225 (N_25225,N_22975,N_20598);
xnor U25226 (N_25226,N_21872,N_22422);
nor U25227 (N_25227,N_20296,N_23742);
nor U25228 (N_25228,N_21107,N_24224);
nand U25229 (N_25229,N_24549,N_22472);
nand U25230 (N_25230,N_22642,N_24157);
and U25231 (N_25231,N_22543,N_24474);
xor U25232 (N_25232,N_22335,N_22694);
xor U25233 (N_25233,N_22868,N_20259);
xnor U25234 (N_25234,N_20470,N_23306);
or U25235 (N_25235,N_21236,N_20186);
nor U25236 (N_25236,N_21844,N_22383);
nor U25237 (N_25237,N_20414,N_23323);
and U25238 (N_25238,N_23702,N_24995);
xnor U25239 (N_25239,N_22576,N_22295);
xor U25240 (N_25240,N_21729,N_21921);
nand U25241 (N_25241,N_20343,N_20506);
nand U25242 (N_25242,N_23514,N_22412);
xor U25243 (N_25243,N_24018,N_22781);
nor U25244 (N_25244,N_22408,N_22954);
xor U25245 (N_25245,N_24006,N_20073);
nor U25246 (N_25246,N_22011,N_20484);
or U25247 (N_25247,N_20156,N_20594);
xnor U25248 (N_25248,N_22297,N_22410);
nand U25249 (N_25249,N_24804,N_23840);
xnor U25250 (N_25250,N_22579,N_21581);
xor U25251 (N_25251,N_23589,N_20357);
and U25252 (N_25252,N_23621,N_23219);
xnor U25253 (N_25253,N_22149,N_23953);
or U25254 (N_25254,N_23469,N_24797);
or U25255 (N_25255,N_24368,N_22714);
nor U25256 (N_25256,N_20691,N_23145);
and U25257 (N_25257,N_24829,N_21226);
nand U25258 (N_25258,N_20188,N_21714);
or U25259 (N_25259,N_23990,N_20468);
nand U25260 (N_25260,N_20736,N_22233);
and U25261 (N_25261,N_20049,N_24933);
xnor U25262 (N_25262,N_23018,N_23940);
and U25263 (N_25263,N_20213,N_20507);
xor U25264 (N_25264,N_24634,N_20575);
and U25265 (N_25265,N_23452,N_22507);
nand U25266 (N_25266,N_23282,N_20404);
nand U25267 (N_25267,N_22280,N_21116);
nand U25268 (N_25268,N_22888,N_22420);
nor U25269 (N_25269,N_21223,N_23921);
and U25270 (N_25270,N_24100,N_24817);
nand U25271 (N_25271,N_24316,N_24334);
nand U25272 (N_25272,N_22722,N_22298);
or U25273 (N_25273,N_21154,N_23036);
and U25274 (N_25274,N_23980,N_24013);
or U25275 (N_25275,N_22561,N_23535);
or U25276 (N_25276,N_20688,N_24023);
nand U25277 (N_25277,N_21395,N_21666);
or U25278 (N_25278,N_23208,N_23468);
and U25279 (N_25279,N_22518,N_24092);
nor U25280 (N_25280,N_20021,N_23189);
nor U25281 (N_25281,N_23360,N_24074);
nand U25282 (N_25282,N_23232,N_20672);
nand U25283 (N_25283,N_22775,N_20197);
and U25284 (N_25284,N_22964,N_22192);
and U25285 (N_25285,N_21267,N_22361);
and U25286 (N_25286,N_21180,N_23316);
xor U25287 (N_25287,N_22226,N_23566);
or U25288 (N_25288,N_21047,N_23753);
nand U25289 (N_25289,N_23159,N_23603);
or U25290 (N_25290,N_24626,N_23342);
or U25291 (N_25291,N_22128,N_24676);
nor U25292 (N_25292,N_22711,N_23773);
nor U25293 (N_25293,N_23269,N_22933);
xor U25294 (N_25294,N_21448,N_24027);
xor U25295 (N_25295,N_20115,N_24458);
nand U25296 (N_25296,N_21561,N_21280);
xnor U25297 (N_25297,N_24793,N_20985);
nand U25298 (N_25298,N_20780,N_24715);
nand U25299 (N_25299,N_22971,N_20852);
nor U25300 (N_25300,N_20374,N_20552);
nand U25301 (N_25301,N_23837,N_24535);
nor U25302 (N_25302,N_23162,N_20126);
nand U25303 (N_25303,N_24395,N_24448);
or U25304 (N_25304,N_20381,N_24009);
and U25305 (N_25305,N_23934,N_23075);
and U25306 (N_25306,N_21625,N_20088);
nor U25307 (N_25307,N_24579,N_22013);
or U25308 (N_25308,N_21461,N_22632);
xor U25309 (N_25309,N_21609,N_20557);
nor U25310 (N_25310,N_20205,N_22475);
and U25311 (N_25311,N_21126,N_23685);
or U25312 (N_25312,N_23423,N_23594);
or U25313 (N_25313,N_20589,N_24730);
or U25314 (N_25314,N_24940,N_23493);
and U25315 (N_25315,N_20763,N_21276);
and U25316 (N_25316,N_21861,N_23299);
or U25317 (N_25317,N_20095,N_20925);
and U25318 (N_25318,N_23668,N_22950);
or U25319 (N_25319,N_21039,N_20797);
xnor U25320 (N_25320,N_23038,N_24893);
or U25321 (N_25321,N_23760,N_24416);
and U25322 (N_25322,N_20075,N_20894);
nor U25323 (N_25323,N_21640,N_22870);
xor U25324 (N_25324,N_22122,N_21403);
or U25325 (N_25325,N_23660,N_23573);
nor U25326 (N_25326,N_21674,N_20652);
or U25327 (N_25327,N_21303,N_24719);
or U25328 (N_25328,N_23023,N_24711);
xor U25329 (N_25329,N_24439,N_23611);
xor U25330 (N_25330,N_23650,N_23280);
nor U25331 (N_25331,N_23207,N_21022);
or U25332 (N_25332,N_22830,N_24098);
nor U25333 (N_25333,N_24657,N_21383);
nor U25334 (N_25334,N_23119,N_21330);
nand U25335 (N_25335,N_22197,N_24801);
nand U25336 (N_25336,N_21618,N_23571);
nor U25337 (N_25337,N_21396,N_20503);
nand U25338 (N_25338,N_24902,N_23051);
nor U25339 (N_25339,N_21787,N_24520);
or U25340 (N_25340,N_20022,N_21456);
and U25341 (N_25341,N_22935,N_22473);
or U25342 (N_25342,N_22776,N_24409);
nor U25343 (N_25343,N_21334,N_20192);
or U25344 (N_25344,N_24468,N_21651);
xor U25345 (N_25345,N_24245,N_21928);
nand U25346 (N_25346,N_20756,N_22658);
and U25347 (N_25347,N_21562,N_24075);
nor U25348 (N_25348,N_24830,N_21849);
nand U25349 (N_25349,N_23026,N_24523);
nor U25350 (N_25350,N_22526,N_20927);
xnor U25351 (N_25351,N_23690,N_23301);
or U25352 (N_25352,N_20212,N_22024);
nor U25353 (N_25353,N_21631,N_22910);
nor U25354 (N_25354,N_21536,N_23532);
or U25355 (N_25355,N_20318,N_24476);
and U25356 (N_25356,N_20145,N_21757);
nand U25357 (N_25357,N_22490,N_23444);
xnor U25358 (N_25358,N_20370,N_20167);
or U25359 (N_25359,N_20634,N_24358);
xor U25360 (N_25360,N_21024,N_21504);
nand U25361 (N_25361,N_21782,N_21771);
or U25362 (N_25362,N_20138,N_20846);
and U25363 (N_25363,N_23749,N_20319);
and U25364 (N_25364,N_24185,N_21457);
or U25365 (N_25365,N_22590,N_21227);
nor U25366 (N_25366,N_21324,N_20401);
and U25367 (N_25367,N_20513,N_22562);
or U25368 (N_25368,N_20413,N_23587);
xor U25369 (N_25369,N_24263,N_21364);
and U25370 (N_25370,N_22099,N_24612);
nor U25371 (N_25371,N_23698,N_24732);
xor U25372 (N_25372,N_23769,N_24480);
and U25373 (N_25373,N_24919,N_22681);
xor U25374 (N_25374,N_23143,N_22676);
and U25375 (N_25375,N_24663,N_23347);
and U25376 (N_25376,N_21372,N_22324);
nor U25377 (N_25377,N_22832,N_21783);
or U25378 (N_25378,N_24172,N_21831);
nand U25379 (N_25379,N_22692,N_21273);
nand U25380 (N_25380,N_20019,N_22730);
xor U25381 (N_25381,N_21230,N_23941);
nand U25382 (N_25382,N_23955,N_20766);
and U25383 (N_25383,N_20117,N_21485);
or U25384 (N_25384,N_20538,N_24839);
and U25385 (N_25385,N_20362,N_22033);
nand U25386 (N_25386,N_22417,N_22185);
nand U25387 (N_25387,N_21994,N_20499);
nand U25388 (N_25388,N_22186,N_21539);
and U25389 (N_25389,N_21883,N_24709);
xnor U25390 (N_25390,N_24099,N_24522);
xor U25391 (N_25391,N_23949,N_20196);
or U25392 (N_25392,N_24542,N_23596);
and U25393 (N_25393,N_24035,N_23309);
and U25394 (N_25394,N_22183,N_21710);
or U25395 (N_25395,N_20651,N_21978);
or U25396 (N_25396,N_22682,N_20764);
xor U25397 (N_25397,N_23178,N_21727);
nand U25398 (N_25398,N_21773,N_21863);
xnor U25399 (N_25399,N_20092,N_20467);
nor U25400 (N_25400,N_20074,N_23035);
or U25401 (N_25401,N_21028,N_24916);
xnor U25402 (N_25402,N_20920,N_23580);
nand U25403 (N_25403,N_23362,N_23745);
xnor U25404 (N_25404,N_21744,N_22760);
xor U25405 (N_25405,N_21760,N_24174);
nor U25406 (N_25406,N_22281,N_22645);
nor U25407 (N_25407,N_20291,N_20372);
xnor U25408 (N_25408,N_22646,N_23058);
nor U25409 (N_25409,N_23268,N_23103);
or U25410 (N_25410,N_20178,N_22104);
xnor U25411 (N_25411,N_24383,N_21275);
and U25412 (N_25412,N_23860,N_23238);
or U25413 (N_25413,N_21626,N_24255);
xor U25414 (N_25414,N_23557,N_24122);
nor U25415 (N_25415,N_21277,N_23202);
and U25416 (N_25416,N_21668,N_22647);
and U25417 (N_25417,N_24003,N_20034);
or U25418 (N_25418,N_24581,N_23539);
nor U25419 (N_25419,N_21960,N_21915);
or U25420 (N_25420,N_20784,N_20772);
and U25421 (N_25421,N_24519,N_21345);
or U25422 (N_25422,N_24087,N_22196);
xnor U25423 (N_25423,N_22106,N_23291);
nand U25424 (N_25424,N_24688,N_20303);
and U25425 (N_25425,N_22190,N_20534);
xnor U25426 (N_25426,N_23572,N_24105);
and U25427 (N_25427,N_23007,N_21393);
or U25428 (N_25428,N_22450,N_21429);
or U25429 (N_25429,N_22670,N_24925);
nand U25430 (N_25430,N_20700,N_24430);
nor U25431 (N_25431,N_23287,N_23180);
or U25432 (N_25432,N_20136,N_20982);
or U25433 (N_25433,N_22531,N_24670);
xnor U25434 (N_25434,N_20287,N_20775);
or U25435 (N_25435,N_21822,N_20787);
nand U25436 (N_25436,N_23544,N_20645);
nor U25437 (N_25437,N_20174,N_21397);
nor U25438 (N_25438,N_23707,N_23272);
and U25439 (N_25439,N_20653,N_21808);
nor U25440 (N_25440,N_24725,N_22628);
nand U25441 (N_25441,N_22002,N_21832);
or U25442 (N_25442,N_21595,N_23063);
or U25443 (N_25443,N_24116,N_20859);
and U25444 (N_25444,N_20495,N_24216);
and U25445 (N_25445,N_24660,N_21980);
xnor U25446 (N_25446,N_21552,N_22063);
and U25447 (N_25447,N_23700,N_22983);
nor U25448 (N_25448,N_22791,N_22132);
or U25449 (N_25449,N_23388,N_24168);
or U25450 (N_25450,N_21242,N_21013);
and U25451 (N_25451,N_23199,N_23121);
or U25452 (N_25452,N_22965,N_22080);
nand U25453 (N_25453,N_22238,N_21411);
xor U25454 (N_25454,N_22786,N_24824);
or U25455 (N_25455,N_22497,N_22918);
nor U25456 (N_25456,N_22594,N_23826);
or U25457 (N_25457,N_21763,N_21696);
xnor U25458 (N_25458,N_24364,N_21002);
nand U25459 (N_25459,N_23615,N_20790);
or U25460 (N_25460,N_23310,N_20301);
nand U25461 (N_25461,N_24215,N_24576);
nor U25462 (N_25462,N_22701,N_23848);
or U25463 (N_25463,N_21747,N_23847);
and U25464 (N_25464,N_24762,N_21912);
nor U25465 (N_25465,N_24206,N_24979);
and U25466 (N_25466,N_20568,N_20055);
xnor U25467 (N_25467,N_22746,N_20860);
and U25468 (N_25468,N_23661,N_24805);
and U25469 (N_25469,N_21066,N_23314);
nor U25470 (N_25470,N_20685,N_24314);
nor U25471 (N_25471,N_20154,N_21499);
or U25472 (N_25472,N_21291,N_21507);
nor U25473 (N_25473,N_20584,N_22350);
xnor U25474 (N_25474,N_21848,N_20704);
nand U25475 (N_25475,N_20363,N_20458);
nor U25476 (N_25476,N_20001,N_20328);
xor U25477 (N_25477,N_23355,N_22005);
nand U25478 (N_25478,N_20675,N_24126);
nand U25479 (N_25479,N_23182,N_24784);
nor U25480 (N_25480,N_21962,N_23656);
or U25481 (N_25481,N_20795,N_22580);
nor U25482 (N_25482,N_24848,N_21218);
xor U25483 (N_25483,N_20637,N_24303);
or U25484 (N_25484,N_21999,N_20107);
xor U25485 (N_25485,N_21564,N_20958);
xnor U25486 (N_25486,N_23538,N_20079);
nand U25487 (N_25487,N_21391,N_23914);
and U25488 (N_25488,N_23273,N_20185);
or U25489 (N_25489,N_22082,N_20373);
nand U25490 (N_25490,N_24894,N_23002);
xor U25491 (N_25491,N_24393,N_24435);
or U25492 (N_25492,N_21575,N_21781);
nand U25493 (N_25493,N_20173,N_22721);
nor U25494 (N_25494,N_22219,N_21077);
and U25495 (N_25495,N_24052,N_24896);
nand U25496 (N_25496,N_20276,N_24293);
and U25497 (N_25497,N_23500,N_22650);
nor U25498 (N_25498,N_21813,N_20851);
nand U25499 (N_25499,N_23482,N_23869);
and U25500 (N_25500,N_20988,N_23739);
nor U25501 (N_25501,N_22680,N_20638);
nand U25502 (N_25502,N_20669,N_24912);
nor U25503 (N_25503,N_24078,N_21138);
and U25504 (N_25504,N_20883,N_23165);
or U25505 (N_25505,N_20140,N_24019);
or U25506 (N_25506,N_23728,N_20035);
nor U25507 (N_25507,N_22847,N_23696);
nand U25508 (N_25508,N_22074,N_23256);
or U25509 (N_25509,N_21349,N_24187);
nor U25510 (N_25510,N_23732,N_23641);
xnor U25511 (N_25511,N_23876,N_21102);
nand U25512 (N_25512,N_21418,N_22946);
nor U25513 (N_25513,N_22211,N_21565);
nand U25514 (N_25514,N_24742,N_23427);
nor U25515 (N_25515,N_21955,N_21282);
and U25516 (N_25516,N_24755,N_21257);
and U25517 (N_25517,N_22131,N_24645);
nand U25518 (N_25518,N_22959,N_23833);
xnor U25519 (N_25519,N_21058,N_24737);
and U25520 (N_25520,N_24788,N_21086);
and U25521 (N_25521,N_20800,N_22057);
nand U25522 (N_25522,N_24471,N_21071);
or U25523 (N_25523,N_22352,N_23146);
and U25524 (N_25524,N_23400,N_22793);
nand U25525 (N_25525,N_22030,N_22618);
xnor U25526 (N_25526,N_24152,N_24888);
or U25527 (N_25527,N_24591,N_23890);
nor U25528 (N_25528,N_22817,N_20108);
xnor U25529 (N_25529,N_22483,N_22139);
or U25530 (N_25530,N_21286,N_20697);
and U25531 (N_25531,N_20733,N_23751);
xnor U25532 (N_25532,N_21164,N_22720);
xor U25533 (N_25533,N_20302,N_21501);
xnor U25534 (N_25534,N_23779,N_21069);
or U25535 (N_25535,N_22332,N_23923);
nor U25536 (N_25536,N_24736,N_24038);
or U25537 (N_25537,N_24753,N_20957);
nand U25538 (N_25538,N_22581,N_24632);
xnor U25539 (N_25539,N_20453,N_24096);
nand U25540 (N_25540,N_20662,N_23861);
xnor U25541 (N_25541,N_22920,N_23722);
or U25542 (N_25542,N_20994,N_24509);
nand U25543 (N_25543,N_20183,N_24989);
nor U25544 (N_25544,N_24489,N_21460);
or U25545 (N_25545,N_22768,N_21571);
nor U25546 (N_25546,N_23244,N_22818);
xor U25547 (N_25547,N_24195,N_22559);
nor U25548 (N_25548,N_21937,N_20322);
and U25549 (N_25549,N_24107,N_20273);
nand U25550 (N_25550,N_23014,N_23149);
or U25551 (N_25551,N_23251,N_23470);
nor U25552 (N_25552,N_20046,N_20332);
xor U25553 (N_25553,N_20006,N_21119);
xnor U25554 (N_25554,N_23726,N_21377);
or U25555 (N_25555,N_20485,N_21802);
xnor U25556 (N_25556,N_23339,N_24502);
and U25557 (N_25557,N_23561,N_24007);
nor U25558 (N_25558,N_23899,N_24648);
or U25559 (N_25559,N_22460,N_22262);
and U25560 (N_25560,N_21741,N_23065);
or U25561 (N_25561,N_20720,N_22338);
xnor U25562 (N_25562,N_20283,N_20665);
and U25563 (N_25563,N_21716,N_22479);
or U25564 (N_25564,N_21614,N_20405);
nand U25565 (N_25565,N_21199,N_24853);
or U25566 (N_25566,N_24511,N_20550);
nor U25567 (N_25567,N_21549,N_20471);
nor U25568 (N_25568,N_21161,N_21067);
nand U25569 (N_25569,N_20290,N_24957);
xnor U25570 (N_25570,N_20000,N_20583);
xnor U25571 (N_25571,N_24366,N_24059);
or U25572 (N_25572,N_23563,N_23478);
and U25573 (N_25573,N_21560,N_21970);
nor U25574 (N_25574,N_24398,N_21637);
nor U25575 (N_25575,N_22799,N_21701);
and U25576 (N_25576,N_24264,N_20109);
xor U25577 (N_25577,N_23693,N_21021);
nor U25578 (N_25578,N_24729,N_23962);
nand U25579 (N_25579,N_22230,N_24566);
nor U25580 (N_25580,N_23016,N_24296);
and U25581 (N_25581,N_24929,N_22908);
xnor U25582 (N_25582,N_24548,N_22740);
xnor U25583 (N_25583,N_22463,N_22529);
or U25584 (N_25584,N_22995,N_21916);
or U25585 (N_25585,N_24179,N_24262);
xor U25586 (N_25586,N_24993,N_23652);
nand U25587 (N_25587,N_23593,N_24647);
or U25588 (N_25588,N_21177,N_24400);
or U25589 (N_25589,N_24852,N_22302);
nor U25590 (N_25590,N_23341,N_24637);
nand U25591 (N_25591,N_21121,N_20344);
nor U25592 (N_25592,N_24029,N_20162);
nand U25593 (N_25593,N_22755,N_22687);
or U25594 (N_25594,N_22377,N_20963);
nand U25595 (N_25595,N_20602,N_20225);
xnor U25596 (N_25596,N_23640,N_24710);
and U25597 (N_25597,N_23796,N_21208);
xor U25598 (N_25598,N_23492,N_22540);
or U25599 (N_25599,N_20220,N_22506);
nand U25600 (N_25600,N_24682,N_23546);
nand U25601 (N_25601,N_23374,N_24378);
nor U25602 (N_25602,N_21694,N_22856);
or U25603 (N_25603,N_20391,N_22214);
nand U25604 (N_25604,N_20422,N_22800);
or U25605 (N_25605,N_24492,N_22842);
nor U25606 (N_25606,N_21482,N_20359);
and U25607 (N_25607,N_23132,N_22103);
or U25608 (N_25608,N_22528,N_20661);
xnor U25609 (N_25609,N_23536,N_23951);
or U25610 (N_25610,N_23084,N_21984);
nor U25611 (N_25611,N_22382,N_23910);
and U25612 (N_25612,N_23520,N_22256);
nand U25613 (N_25613,N_20970,N_23116);
xor U25614 (N_25614,N_21135,N_21720);
and U25615 (N_25615,N_22916,N_21784);
or U25616 (N_25616,N_21707,N_23073);
or U25617 (N_25617,N_24712,N_20051);
or U25618 (N_25618,N_21184,N_21083);
nand U25619 (N_25619,N_20801,N_21417);
nand U25620 (N_25620,N_21350,N_22605);
or U25621 (N_25621,N_23069,N_20184);
nand U25622 (N_25622,N_20996,N_22980);
xnor U25623 (N_25623,N_22366,N_20443);
and U25624 (N_25624,N_22387,N_20781);
and U25625 (N_25625,N_24799,N_20715);
xnor U25626 (N_25626,N_22428,N_23961);
xor U25627 (N_25627,N_23401,N_23584);
nand U25628 (N_25628,N_22117,N_23515);
and U25629 (N_25629,N_20171,N_23827);
nand U25630 (N_25630,N_24703,N_22593);
nand U25631 (N_25631,N_21279,N_20916);
or U25632 (N_25632,N_23177,N_24790);
xnor U25633 (N_25633,N_22630,N_20351);
xor U25634 (N_25634,N_22121,N_23612);
or U25635 (N_25635,N_22801,N_21385);
or U25636 (N_25636,N_24789,N_20636);
nor U25637 (N_25637,N_23186,N_20515);
nand U25638 (N_25638,N_20918,N_22889);
nand U25639 (N_25639,N_20895,N_20746);
nor U25640 (N_25640,N_22530,N_22498);
nor U25641 (N_25641,N_23771,N_20010);
or U25642 (N_25642,N_21449,N_23813);
nor U25643 (N_25643,N_24807,N_22474);
and U25644 (N_25644,N_20750,N_23724);
xor U25645 (N_25645,N_21546,N_22848);
and U25646 (N_25646,N_24761,N_21780);
nor U25647 (N_25647,N_21081,N_23846);
nor U25648 (N_25648,N_23215,N_24706);
nand U25649 (N_25649,N_20340,N_24384);
nand U25650 (N_25650,N_21524,N_23398);
and U25651 (N_25651,N_20850,N_20395);
nand U25652 (N_25652,N_20757,N_23528);
or U25653 (N_25653,N_24623,N_20350);
nor U25654 (N_25654,N_20832,N_23336);
nand U25655 (N_25655,N_23442,N_21231);
and U25656 (N_25656,N_23279,N_20622);
and U25657 (N_25657,N_24080,N_23099);
or U25658 (N_25658,N_23370,N_20773);
xnor U25659 (N_25659,N_23936,N_23908);
and U25660 (N_25660,N_24935,N_20224);
xor U25661 (N_25661,N_23644,N_22379);
xor U25662 (N_25662,N_24030,N_24084);
and U25663 (N_25663,N_23190,N_23554);
and U25664 (N_25664,N_22690,N_23350);
nand U25665 (N_25665,N_24903,N_23088);
or U25666 (N_25666,N_23675,N_22255);
and U25667 (N_25667,N_24845,N_22931);
or U25668 (N_25668,N_22252,N_20246);
and U25669 (N_25669,N_23808,N_24757);
and U25670 (N_25670,N_24203,N_21777);
nand U25671 (N_25671,N_22820,N_21238);
nor U25672 (N_25672,N_24747,N_24800);
or U25673 (N_25673,N_21440,N_24024);
xor U25674 (N_25674,N_23534,N_23243);
and U25675 (N_25675,N_21342,N_21405);
or U25676 (N_25676,N_22331,N_23986);
xnor U25677 (N_25677,N_20255,N_22909);
nor U25678 (N_25678,N_21148,N_24498);
nand U25679 (N_25679,N_23704,N_23809);
and U25680 (N_25680,N_21870,N_22871);
nand U25681 (N_25681,N_23591,N_24716);
nor U25682 (N_25682,N_22055,N_24700);
nor U25683 (N_25683,N_21487,N_22782);
xnor U25684 (N_25684,N_23559,N_22536);
nand U25685 (N_25685,N_22129,N_24782);
and U25686 (N_25686,N_24618,N_24889);
nor U25687 (N_25687,N_20110,N_21910);
nand U25688 (N_25688,N_22270,N_21559);
xnor U25689 (N_25689,N_23172,N_23331);
nor U25690 (N_25690,N_21497,N_21965);
or U25691 (N_25691,N_23586,N_21374);
nor U25692 (N_25692,N_20947,N_20123);
and U25693 (N_25693,N_23319,N_23409);
or U25694 (N_25694,N_23107,N_21297);
xor U25695 (N_25695,N_24242,N_24699);
nor U25696 (N_25696,N_22990,N_21312);
nand U25697 (N_25697,N_24680,N_24543);
nand U25698 (N_25698,N_21348,N_20912);
nand U25699 (N_25699,N_24181,N_24978);
nand U25700 (N_25700,N_23582,N_22232);
or U25701 (N_25701,N_21523,N_22247);
and U25702 (N_25702,N_20649,N_23606);
or U25703 (N_25703,N_24544,N_21419);
nor U25704 (N_25704,N_22553,N_21554);
nand U25705 (N_25705,N_21185,N_20768);
nor U25706 (N_25706,N_20402,N_23226);
nor U25707 (N_25707,N_23673,N_22449);
nand U25708 (N_25708,N_24526,N_22019);
or U25709 (N_25709,N_21615,N_24597);
nor U25710 (N_25710,N_21719,N_24425);
or U25711 (N_25711,N_21167,N_20037);
nor U25712 (N_25712,N_23947,N_20628);
nor U25713 (N_25713,N_23368,N_22930);
nand U25714 (N_25714,N_23560,N_21062);
xnor U25715 (N_25715,N_20931,N_21465);
or U25716 (N_25716,N_21245,N_21768);
xor U25717 (N_25717,N_21237,N_20323);
and U25718 (N_25718,N_20437,N_21917);
nand U25719 (N_25719,N_24000,N_22141);
nand U25720 (N_25720,N_20609,N_22615);
nand U25721 (N_25721,N_21517,N_20717);
and U25722 (N_25722,N_20081,N_24191);
nand U25723 (N_25723,N_23883,N_24198);
or U25724 (N_25724,N_24945,N_24731);
nand U25725 (N_25725,N_22926,N_21909);
nor U25726 (N_25726,N_21519,N_24136);
nand U25727 (N_25727,N_23526,N_24178);
xor U25728 (N_25728,N_22733,N_24704);
and U25729 (N_25729,N_20705,N_22493);
nor U25730 (N_25730,N_23377,N_23393);
and U25731 (N_25731,N_23475,N_21304);
nor U25732 (N_25732,N_21454,N_24487);
or U25733 (N_25733,N_20792,N_22250);
and U25734 (N_25734,N_24091,N_22003);
xor U25735 (N_25735,N_24792,N_21672);
and U25736 (N_25736,N_21174,N_22061);
nand U25737 (N_25737,N_20762,N_22763);
nor U25738 (N_25738,N_24850,N_20874);
and U25739 (N_25739,N_20100,N_20681);
xor U25740 (N_25740,N_20953,N_24083);
xor U25741 (N_25741,N_24661,N_22996);
and U25742 (N_25742,N_22077,N_20579);
and U25743 (N_25743,N_20839,N_21568);
nand U25744 (N_25744,N_24291,N_22899);
and U25745 (N_25745,N_22874,N_21031);
xor U25746 (N_25746,N_22431,N_24440);
and U25747 (N_25747,N_21991,N_23692);
or U25748 (N_25748,N_23674,N_20040);
nand U25749 (N_25749,N_22879,N_21496);
nor U25750 (N_25750,N_23944,N_23312);
and U25751 (N_25751,N_22014,N_24382);
or U25752 (N_25752,N_21020,N_20991);
nand U25753 (N_25753,N_22578,N_22853);
and U25754 (N_25754,N_23857,N_23439);
and U25755 (N_25755,N_23138,N_20120);
and U25756 (N_25756,N_23196,N_24210);
nand U25757 (N_25757,N_20939,N_22863);
nor U25758 (N_25758,N_21446,N_23505);
xnor U25759 (N_25759,N_21702,N_21953);
xnor U25760 (N_25760,N_21209,N_21769);
and U25761 (N_25761,N_20545,N_23104);
nand U25762 (N_25762,N_21123,N_22591);
or U25763 (N_25763,N_24407,N_23170);
xor U25764 (N_25764,N_22978,N_24387);
and U25765 (N_25765,N_20644,N_20412);
and U25766 (N_25766,N_24609,N_23487);
nand U25767 (N_25767,N_23153,N_24694);
or U25768 (N_25768,N_22906,N_23009);
nor U25769 (N_25769,N_22859,N_21879);
xor U25770 (N_25770,N_22370,N_23415);
nor U25771 (N_25771,N_24857,N_20713);
nand U25772 (N_25772,N_21467,N_23298);
nor U25773 (N_25773,N_23977,N_23183);
nor U25774 (N_25774,N_21251,N_24346);
or U25775 (N_25775,N_22881,N_23443);
nand U25776 (N_25776,N_24514,N_23531);
and U25777 (N_25777,N_23025,N_22415);
or U25778 (N_25778,N_21837,N_23017);
nor U25779 (N_25779,N_24678,N_21406);
and U25780 (N_25780,N_23262,N_22378);
or U25781 (N_25781,N_20587,N_20309);
and U25782 (N_25782,N_23996,N_22114);
and U25783 (N_25783,N_20540,N_23290);
or U25784 (N_25784,N_24787,N_21322);
xnor U25785 (N_25785,N_20494,N_20782);
or U25786 (N_25786,N_24449,N_24201);
nor U25787 (N_25787,N_21425,N_23288);
nor U25788 (N_25788,N_23583,N_22753);
nand U25789 (N_25789,N_23886,N_20596);
and U25790 (N_25790,N_21792,N_22735);
or U25791 (N_25791,N_23844,N_22195);
and U25792 (N_25792,N_22440,N_22981);
nand U25793 (N_25793,N_21409,N_20371);
nand U25794 (N_25794,N_22333,N_23551);
nand U25795 (N_25795,N_21045,N_23246);
or U25796 (N_25796,N_23922,N_21724);
and U25797 (N_25797,N_23689,N_23825);
or U25798 (N_25798,N_23897,N_21754);
and U25799 (N_25799,N_24956,N_22500);
and U25800 (N_25800,N_22451,N_24810);
nand U25801 (N_25801,N_21547,N_21765);
xor U25802 (N_25802,N_22601,N_23117);
or U25803 (N_25803,N_20728,N_21911);
or U25804 (N_25804,N_24607,N_24939);
and U25805 (N_25805,N_22444,N_22663);
xnor U25806 (N_25806,N_23463,N_23609);
nand U25807 (N_25807,N_23547,N_23048);
nand U25808 (N_25808,N_20938,N_20450);
nor U25809 (N_25809,N_24911,N_20133);
or U25810 (N_25810,N_20274,N_21188);
nor U25811 (N_25811,N_24765,N_20346);
nand U25812 (N_25812,N_20089,N_21427);
nor U25813 (N_25813,N_20677,N_21555);
or U25814 (N_25814,N_24156,N_21576);
nand U25815 (N_25815,N_22396,N_20853);
nand U25816 (N_25816,N_23406,N_22901);
and U25817 (N_25817,N_22969,N_20737);
xor U25818 (N_25818,N_24332,N_24042);
xnor U25819 (N_25819,N_24578,N_24113);
and U25820 (N_25820,N_23864,N_24697);
nand U25821 (N_25821,N_24941,N_24828);
xnor U25822 (N_25822,N_20153,N_20543);
nor U25823 (N_25823,N_21819,N_21975);
or U25824 (N_25824,N_24367,N_20980);
xor U25825 (N_25825,N_21922,N_24837);
and U25826 (N_25826,N_21382,N_21514);
nand U25827 (N_25827,N_23029,N_23303);
nand U25828 (N_25828,N_20600,N_22796);
nor U25829 (N_25829,N_22940,N_23782);
xnor U25830 (N_25830,N_22659,N_21828);
and U25831 (N_25831,N_21283,N_21518);
and U25832 (N_25832,N_22678,N_23604);
nand U25833 (N_25833,N_24960,N_22696);
or U25834 (N_25834,N_24292,N_24189);
and U25835 (N_25835,N_21096,N_22430);
xnor U25836 (N_25836,N_22070,N_21387);
nor U25837 (N_25837,N_20553,N_24668);
and U25838 (N_25838,N_23144,N_22487);
nand U25839 (N_25839,N_24162,N_22679);
xnor U25840 (N_25840,N_22244,N_22135);
or U25841 (N_25841,N_24010,N_20433);
xnor U25842 (N_25842,N_20141,N_22268);
nor U25843 (N_25843,N_24324,N_21657);
and U25844 (N_25844,N_21839,N_21840);
or U25845 (N_25845,N_21584,N_24048);
nor U25846 (N_25846,N_22858,N_23906);
xnor U25847 (N_25847,N_23338,N_24880);
nor U25848 (N_25848,N_23634,N_21018);
or U25849 (N_25849,N_20876,N_22836);
or U25850 (N_25850,N_23626,N_21914);
xor U25851 (N_25851,N_20118,N_20856);
or U25852 (N_25852,N_20827,N_24602);
nand U25853 (N_25853,N_22737,N_21627);
or U25854 (N_25854,N_21850,N_22838);
and U25855 (N_25855,N_20347,N_23192);
nor U25856 (N_25856,N_22342,N_21182);
nor U25857 (N_25857,N_22434,N_20558);
xor U25858 (N_25858,N_21619,N_21924);
or U25859 (N_25859,N_21538,N_20621);
nor U25860 (N_25860,N_21006,N_21567);
or U25861 (N_25861,N_21438,N_24551);
or U25862 (N_25862,N_20703,N_21139);
or U25863 (N_25863,N_20462,N_21761);
or U25864 (N_25864,N_24300,N_23079);
or U25865 (N_25865,N_21942,N_21084);
xnor U25866 (N_25866,N_22648,N_24763);
and U25867 (N_25867,N_24134,N_21337);
and U25868 (N_25868,N_20863,N_23094);
nand U25869 (N_25869,N_21007,N_21739);
nand U25870 (N_25870,N_20606,N_21253);
nor U25871 (N_25871,N_21414,N_21114);
nor U25872 (N_25872,N_21825,N_22649);
xnor U25873 (N_25873,N_20555,N_23357);
xor U25874 (N_25874,N_20397,N_20493);
nor U25875 (N_25875,N_24308,N_20592);
nand U25876 (N_25876,N_21239,N_21997);
xnor U25877 (N_25877,N_24369,N_21407);
or U25878 (N_25878,N_21325,N_24891);
nor U25879 (N_25879,N_22039,N_23293);
or U25880 (N_25880,N_20873,N_23590);
nor U25881 (N_25881,N_21463,N_22538);
and U25882 (N_25882,N_23096,N_24271);
nor U25883 (N_25883,N_22321,N_23576);
nand U25884 (N_25884,N_24721,N_24781);
or U25885 (N_25885,N_21178,N_23447);
xnor U25886 (N_25886,N_24041,N_23266);
or U25887 (N_25887,N_22569,N_20646);
nand U25888 (N_25888,N_24016,N_24305);
and U25889 (N_25889,N_21990,N_21943);
nor U25890 (N_25890,N_24465,N_24143);
and U25891 (N_25891,N_23943,N_21818);
xor U25892 (N_25892,N_24983,N_23828);
and U25893 (N_25893,N_23307,N_22010);
or U25894 (N_25894,N_23904,N_22446);
or U25895 (N_25895,N_23077,N_20643);
and U25896 (N_25896,N_24343,N_20678);
nand U25897 (N_25897,N_21168,N_24063);
xor U25898 (N_25898,N_23195,N_22300);
nor U25899 (N_25899,N_24907,N_22521);
and U25900 (N_25900,N_20094,N_24127);
and U25901 (N_25901,N_22695,N_20059);
and U25902 (N_25902,N_24555,N_23994);
nand U25903 (N_25903,N_20586,N_23617);
nor U25904 (N_25904,N_23794,N_20799);
nand U25905 (N_25905,N_22807,N_22231);
or U25906 (N_25906,N_23166,N_20048);
and U25907 (N_25907,N_22022,N_24286);
or U25908 (N_25908,N_22317,N_20565);
and U25909 (N_25909,N_20449,N_22774);
nor U25910 (N_25910,N_20445,N_23446);
nand U25911 (N_25911,N_24513,N_22948);
xnor U25912 (N_25912,N_22199,N_22058);
nand U25913 (N_25913,N_22386,N_20674);
and U25914 (N_25914,N_21525,N_24967);
or U25915 (N_25915,N_21579,N_22886);
nand U25916 (N_25916,N_21117,N_24188);
xor U25917 (N_25917,N_21155,N_22228);
nand U25918 (N_25918,N_21873,N_22177);
xnor U25919 (N_25919,N_22180,N_22880);
and U25920 (N_25920,N_22438,N_24600);
xnor U25921 (N_25921,N_23212,N_21057);
or U25922 (N_25922,N_24220,N_23733);
xnor U25923 (N_25923,N_22873,N_23757);
nor U25924 (N_25924,N_22194,N_24965);
nor U25925 (N_25925,N_21343,N_22570);
nor U25926 (N_25926,N_23250,N_20566);
nor U25927 (N_25927,N_24093,N_21926);
and U25928 (N_25928,N_23097,N_24841);
or U25929 (N_25929,N_23659,N_24846);
and U25930 (N_25930,N_20544,N_23379);
nor U25931 (N_25931,N_22810,N_24257);
and U25932 (N_25932,N_20268,N_21032);
xnor U25933 (N_25933,N_20990,N_23647);
or U25934 (N_25934,N_23570,N_20671);
and U25935 (N_25935,N_22574,N_22784);
and U25936 (N_25936,N_20315,N_23078);
and U25937 (N_25937,N_24486,N_23085);
or U25938 (N_25938,N_20843,N_21503);
xnor U25939 (N_25939,N_24081,N_20899);
xor U25940 (N_25940,N_21012,N_24184);
and U25941 (N_25941,N_23995,N_21814);
nand U25942 (N_25942,N_22147,N_23187);
nand U25943 (N_25943,N_20702,N_21288);
or U25944 (N_25944,N_20389,N_24072);
and U25945 (N_25945,N_24375,N_20033);
nand U25946 (N_25946,N_21522,N_23613);
and U25947 (N_25947,N_20919,N_20387);
xor U25948 (N_25948,N_21481,N_23954);
or U25949 (N_25949,N_22495,N_20683);
nand U25950 (N_25950,N_24149,N_23426);
nor U25951 (N_25951,N_22552,N_23664);
xor U25952 (N_25952,N_22411,N_22719);
or U25953 (N_25953,N_21712,N_22050);
xor U25954 (N_25954,N_22542,N_21290);
or U25955 (N_25955,N_21243,N_21845);
nand U25956 (N_25956,N_20004,N_23797);
or U25957 (N_25957,N_24691,N_21179);
nand U25958 (N_25958,N_20530,N_22257);
or U25959 (N_25959,N_24247,N_23090);
and U25960 (N_25960,N_21014,N_23414);
or U25961 (N_25961,N_22224,N_20611);
nor U25962 (N_25962,N_23161,N_20489);
nand U25963 (N_25963,N_24671,N_21203);
xor U25964 (N_25964,N_23386,N_24070);
xnor U25965 (N_25965,N_20619,N_22358);
or U25966 (N_25966,N_21080,N_23646);
and U25967 (N_25967,N_21610,N_21799);
and U25968 (N_25968,N_21269,N_24714);
xnor U25969 (N_25969,N_24723,N_21902);
nand U25970 (N_25970,N_20007,N_24794);
and U25971 (N_25971,N_24868,N_20647);
or U25972 (N_25972,N_20858,N_24679);
or U25973 (N_25973,N_21068,N_21875);
nor U25974 (N_25974,N_24260,N_22966);
nor U25975 (N_25975,N_20828,N_23450);
and U25976 (N_25976,N_22549,N_20692);
or U25977 (N_25977,N_22656,N_22982);
nand U25978 (N_25978,N_22089,N_24938);
or U25979 (N_25979,N_24085,N_21434);
nor U25980 (N_25980,N_21159,N_21630);
and U25981 (N_25981,N_21320,N_20366);
xnor U25982 (N_25982,N_24246,N_23909);
xnor U25983 (N_25983,N_20353,N_20429);
xnor U25984 (N_25984,N_23862,N_22809);
and U25985 (N_25985,N_20219,N_24297);
xor U25986 (N_25986,N_21241,N_21698);
xor U25987 (N_25987,N_24190,N_21577);
or U25988 (N_25988,N_23070,N_24649);
nor U25989 (N_25989,N_22042,N_20228);
or U25990 (N_25990,N_22708,N_23901);
xor U25991 (N_25991,N_21959,N_23933);
nand U25992 (N_25992,N_20427,N_24650);
nand U25993 (N_25993,N_23225,N_24567);
or U25994 (N_25994,N_24883,N_24777);
and U25995 (N_25995,N_23932,N_20066);
xor U25996 (N_25996,N_20388,N_23854);
or U25997 (N_25997,N_20253,N_21293);
xnor U25998 (N_25998,N_21370,N_22957);
or U25999 (N_25999,N_23408,N_20585);
xnor U26000 (N_26000,N_21796,N_22514);
or U26001 (N_26001,N_23224,N_20411);
and U26002 (N_26002,N_21023,N_22274);
and U26003 (N_26003,N_20934,N_23710);
and U26004 (N_26004,N_23711,N_22100);
and U26005 (N_26005,N_23812,N_22734);
and U26006 (N_26006,N_24032,N_21815);
xor U26007 (N_26007,N_20227,N_21821);
nor U26008 (N_26008,N_24044,N_21834);
xnor U26009 (N_26009,N_24508,N_24510);
nand U26010 (N_26010,N_23971,N_21738);
nor U26011 (N_26011,N_22968,N_22486);
xor U26012 (N_26012,N_22130,N_24669);
or U26013 (N_26013,N_24798,N_24067);
nor U26014 (N_26014,N_22445,N_21305);
xnor U26015 (N_26015,N_21459,N_23657);
nand U26016 (N_26016,N_22504,N_22872);
or U26017 (N_26017,N_21347,N_22739);
xor U26018 (N_26018,N_23130,N_24235);
and U26019 (N_26019,N_23239,N_20294);
xor U26020 (N_26020,N_22544,N_22016);
or U26021 (N_26021,N_21663,N_23655);
nand U26022 (N_26022,N_22137,N_21992);
nand U26023 (N_26023,N_22675,N_20831);
xor U26024 (N_26024,N_20900,N_23958);
nand U26025 (N_26025,N_23115,N_22047);
nand U26026 (N_26026,N_23815,N_24357);
and U26027 (N_26027,N_22375,N_24900);
nand U26028 (N_26028,N_24444,N_22347);
nor U26029 (N_26029,N_23548,N_20203);
nand U26030 (N_26030,N_24261,N_21214);
nor U26031 (N_26031,N_20533,N_20400);
xor U26032 (N_26032,N_22566,N_23488);
xnor U26033 (N_26033,N_23356,N_20382);
nor U26034 (N_26034,N_20289,N_21316);
nor U26035 (N_26035,N_24823,N_22264);
xnor U26036 (N_26036,N_23902,N_24972);
or U26037 (N_26037,N_20032,N_21206);
nand U26038 (N_26038,N_22289,N_23438);
and U26039 (N_26039,N_24347,N_21095);
and U26040 (N_26040,N_24479,N_21591);
nor U26041 (N_26041,N_21961,N_24955);
or U26042 (N_26042,N_21628,N_21996);
xnor U26043 (N_26043,N_21355,N_21746);
and U26044 (N_26044,N_23061,N_24667);
nand U26045 (N_26045,N_20071,N_21296);
or U26046 (N_26046,N_20524,N_23956);
nand U26047 (N_26047,N_24655,N_21859);
or U26048 (N_26048,N_23363,N_21946);
nand U26049 (N_26049,N_21294,N_24937);
xor U26050 (N_26050,N_22309,N_24931);
nor U26051 (N_26051,N_21207,N_21037);
or U26052 (N_26052,N_21059,N_22917);
nand U26053 (N_26053,N_24319,N_21453);
or U26054 (N_26054,N_24337,N_21075);
and U26055 (N_26055,N_21196,N_20245);
nand U26056 (N_26056,N_20588,N_20965);
and U26057 (N_26057,N_23200,N_21676);
nand U26058 (N_26058,N_21140,N_24811);
or U26059 (N_26059,N_24575,N_23687);
xnor U26060 (N_26060,N_22993,N_23816);
nand U26061 (N_26061,N_23030,N_24338);
and U26062 (N_26062,N_22079,N_23682);
or U26063 (N_26063,N_22085,N_21927);
and U26064 (N_26064,N_21346,N_20130);
or U26065 (N_26065,N_24076,N_21332);
and U26066 (N_26066,N_21498,N_24391);
nor U26067 (N_26067,N_20295,N_21827);
or U26068 (N_26068,N_21359,N_20879);
nor U26069 (N_26069,N_20512,N_24441);
nand U26070 (N_26070,N_20023,N_22187);
or U26071 (N_26071,N_23216,N_23555);
nand U26072 (N_26072,N_21019,N_21543);
or U26073 (N_26073,N_20206,N_24226);
and U26074 (N_26074,N_23154,N_21582);
nor U26075 (N_26075,N_24167,N_24616);
xnor U26076 (N_26076,N_22397,N_24808);
or U26077 (N_26077,N_22742,N_22637);
and U26078 (N_26078,N_22823,N_22153);
xor U26079 (N_26079,N_21169,N_21836);
nand U26080 (N_26080,N_22534,N_20266);
xnor U26081 (N_26081,N_24601,N_22367);
or U26082 (N_26082,N_22607,N_24946);
or U26083 (N_26083,N_20486,N_24118);
xnor U26084 (N_26084,N_21187,N_24976);
xor U26085 (N_26085,N_24208,N_23765);
and U26086 (N_26086,N_24371,N_24507);
nor U26087 (N_26087,N_24490,N_22035);
xnor U26088 (N_26088,N_22259,N_20017);
and U26089 (N_26089,N_21442,N_23569);
and U26090 (N_26090,N_22779,N_23998);
xor U26091 (N_26091,N_22728,N_21585);
or U26092 (N_26092,N_23052,N_21580);
xor U26093 (N_26093,N_24451,N_24769);
xnor U26094 (N_26094,N_24040,N_20461);
and U26095 (N_26095,N_20271,N_22015);
nand U26096 (N_26096,N_23479,N_21426);
nor U26097 (N_26097,N_22963,N_23625);
or U26098 (N_26098,N_23472,N_24536);
and U26099 (N_26099,N_23274,N_23550);
or U26100 (N_26100,N_21653,N_20871);
nor U26101 (N_26101,N_20695,N_22661);
xor U26102 (N_26102,N_21274,N_20569);
or U26103 (N_26103,N_24064,N_23168);
nand U26104 (N_26104,N_20137,N_21323);
xnor U26105 (N_26105,N_24856,N_22655);
nor U26106 (N_26106,N_24249,N_22273);
and U26107 (N_26107,N_21268,N_20933);
or U26108 (N_26108,N_22204,N_20243);
and U26109 (N_26109,N_22170,N_24658);
or U26110 (N_26110,N_23364,N_21553);
xor U26111 (N_26111,N_21935,N_20709);
and U26112 (N_26112,N_20577,N_23770);
and U26113 (N_26113,N_20378,N_22155);
nor U26114 (N_26114,N_24969,N_24539);
xor U26115 (N_26115,N_22766,N_22960);
nor U26116 (N_26116,N_21704,N_22845);
or U26117 (N_26117,N_24619,N_23382);
nor U26118 (N_26118,N_21175,N_20696);
nand U26119 (N_26119,N_20207,N_21726);
and U26120 (N_26120,N_20610,N_21679);
xor U26121 (N_26121,N_24237,N_23134);
nor U26122 (N_26122,N_20978,N_24344);
and U26123 (N_26123,N_20380,N_21730);
or U26124 (N_26124,N_22790,N_23719);
and U26125 (N_26125,N_20250,N_21642);
xnor U26126 (N_26126,N_21260,N_20364);
xnor U26127 (N_26127,N_21157,N_23752);
or U26128 (N_26128,N_23343,N_22866);
xnor U26129 (N_26129,N_23777,N_20502);
xor U26130 (N_26130,N_23654,N_22551);
xor U26131 (N_26131,N_22653,N_22869);
or U26132 (N_26132,N_22805,N_22462);
xnor U26133 (N_26133,N_23871,N_22116);
xor U26134 (N_26134,N_22956,N_20193);
and U26135 (N_26135,N_20812,N_21351);
xnor U26136 (N_26136,N_23518,N_22877);
nand U26137 (N_26137,N_22118,N_24750);
and U26138 (N_26138,N_22161,N_20952);
and U26139 (N_26139,N_22403,N_21983);
nand U26140 (N_26140,N_23565,N_23220);
nand U26141 (N_26141,N_24611,N_21801);
or U26142 (N_26142,N_24553,N_22164);
and U26143 (N_26143,N_23568,N_22158);
and U26144 (N_26144,N_23321,N_23380);
nor U26145 (N_26145,N_20932,N_20134);
or U26146 (N_26146,N_21313,N_21857);
nand U26147 (N_26147,N_20263,N_23437);
or U26148 (N_26148,N_21353,N_20435);
nor U26149 (N_26149,N_21142,N_20818);
and U26150 (N_26150,N_22686,N_24734);
and U26151 (N_26151,N_23141,N_21588);
and U26152 (N_26152,N_20854,N_24867);
or U26153 (N_26153,N_23418,N_24225);
and U26154 (N_26154,N_21149,N_22898);
xor U26155 (N_26155,N_22929,N_22625);
and U26156 (N_26156,N_20891,N_22762);
xnor U26157 (N_26157,N_22029,N_21958);
xnor U26158 (N_26158,N_24289,N_20053);
xor U26159 (N_26159,N_24146,N_20327);
nand U26160 (N_26160,N_21551,N_24450);
nor U26161 (N_26161,N_21368,N_20217);
nand U26162 (N_26162,N_20805,N_20979);
nor U26163 (N_26163,N_21265,N_21838);
or U26164 (N_26164,N_22095,N_23037);
or U26165 (N_26165,N_24342,N_24061);
and U26166 (N_26166,N_21373,N_24302);
and U26167 (N_26167,N_24659,N_22994);
nand U26168 (N_26168,N_20265,N_21762);
nand U26169 (N_26169,N_24643,N_21375);
and U26170 (N_26170,N_23881,N_23629);
nand U26171 (N_26171,N_20626,N_24313);
nor U26172 (N_26172,N_20885,N_24635);
or U26173 (N_26173,N_24424,N_21254);
or U26174 (N_26174,N_22860,N_24133);
nor U26175 (N_26175,N_22568,N_24278);
nor U26176 (N_26176,N_22611,N_21363);
or U26177 (N_26177,N_21731,N_23889);
and U26178 (N_26178,N_24651,N_21737);
and U26179 (N_26179,N_23054,N_22307);
and U26180 (N_26180,N_21686,N_23013);
nand U26181 (N_26181,N_20159,N_20522);
nor U26182 (N_26182,N_22811,N_21690);
or U26183 (N_26183,N_24125,N_24318);
nor U26184 (N_26184,N_24890,N_22478);
or U26185 (N_26185,N_24997,N_20124);
xnor U26186 (N_26186,N_22221,N_23984);
or U26187 (N_26187,N_23721,N_22777);
xnor U26188 (N_26188,N_23931,N_20999);
or U26189 (N_26189,N_24095,N_21891);
nor U26190 (N_26190,N_21682,N_23703);
and U26191 (N_26191,N_22691,N_24028);
nor U26192 (N_26192,N_23292,N_23924);
and U26193 (N_26193,N_22595,N_20488);
and U26194 (N_26194,N_21246,N_20560);
nand U26195 (N_26195,N_24744,N_20064);
nor U26196 (N_26196,N_22245,N_21592);
nor U26197 (N_26197,N_21001,N_20166);
xor U26198 (N_26198,N_20861,N_24470);
and U26199 (N_26199,N_21649,N_21948);
xor U26200 (N_26200,N_21973,N_22839);
nor U26201 (N_26201,N_24717,N_20580);
and U26202 (N_26202,N_20390,N_24855);
or U26203 (N_26203,N_23081,N_22441);
xnor U26204 (N_26204,N_23972,N_22110);
nand U26205 (N_26205,N_21278,N_22093);
xnor U26206 (N_26206,N_23762,N_22945);
nand U26207 (N_26207,N_24835,N_22169);
and U26208 (N_26208,N_21566,N_20170);
and U26209 (N_26209,N_22215,N_23223);
xor U26210 (N_26210,N_22915,N_24534);
or U26211 (N_26211,N_24910,N_21125);
xor U26212 (N_26212,N_21732,N_22748);
and U26213 (N_26213,N_23236,N_23818);
xnor U26214 (N_26214,N_20971,N_21803);
and U26215 (N_26215,N_20355,N_21366);
nand U26216 (N_26216,N_20969,N_23601);
xor U26217 (N_26217,N_20406,N_22173);
nor U26218 (N_26218,N_23793,N_21874);
nor U26219 (N_26219,N_24656,N_20604);
nand U26220 (N_26220,N_22723,N_20973);
nand U26221 (N_26221,N_22876,N_20956);
nand U26222 (N_26222,N_22146,N_21437);
nand U26223 (N_26223,N_23112,N_22112);
and U26224 (N_26224,N_24411,N_23767);
or U26225 (N_26225,N_23510,N_20595);
or U26226 (N_26226,N_21736,N_24662);
nor U26227 (N_26227,N_20834,N_24556);
xnor U26228 (N_26228,N_22059,N_21635);
and U26229 (N_26229,N_24860,N_20618);
nor U26230 (N_26230,N_22119,N_21394);
xor U26231 (N_26231,N_23527,N_22303);
or U26232 (N_26232,N_23193,N_21778);
nor U26233 (N_26233,N_24702,N_20444);
nor U26234 (N_26234,N_20693,N_21703);
xor U26235 (N_26235,N_22535,N_20803);
nand U26236 (N_26236,N_20721,N_23519);
nand U26237 (N_26237,N_21947,N_24785);
or U26238 (N_26238,N_24958,N_20305);
and U26239 (N_26239,N_22282,N_21574);
or U26240 (N_26240,N_22171,N_20676);
or U26241 (N_26241,N_20226,N_20527);
xor U26242 (N_26242,N_20264,N_20730);
nor U26243 (N_26243,N_23530,N_22071);
nor U26244 (N_26244,N_24205,N_24527);
or U26245 (N_26245,N_20808,N_23158);
or U26246 (N_26246,N_20838,N_22319);
nand U26247 (N_26247,N_22229,N_22509);
or U26248 (N_26248,N_22769,N_21190);
nor U26249 (N_26249,N_23853,N_21688);
or U26250 (N_26250,N_22638,N_22278);
and U26251 (N_26251,N_20020,N_21339);
and U26252 (N_26252,N_24973,N_21520);
xnor U26253 (N_26253,N_21728,N_22852);
nor U26254 (N_26254,N_24421,N_22563);
xnor U26255 (N_26255,N_24148,N_20778);
nor U26256 (N_26256,N_21812,N_22705);
nor U26257 (N_26257,N_23318,N_23525);
nor U26258 (N_26258,N_20884,N_21259);
nor U26259 (N_26259,N_23750,N_22812);
xnor U26260 (N_26260,N_24759,N_20099);
nor U26261 (N_26261,N_22044,N_22320);
nor U26262 (N_26262,N_23537,N_23822);
nand U26263 (N_26263,N_20442,N_20590);
nand U26264 (N_26264,N_23101,N_22108);
and U26265 (N_26265,N_20726,N_22020);
xor U26266 (N_26266,N_22702,N_20298);
nor U26267 (N_26267,N_23878,N_21431);
nor U26268 (N_26268,N_23125,N_24934);
nor U26269 (N_26269,N_23481,N_22556);
nor U26270 (N_26270,N_20877,N_23880);
nor U26271 (N_26271,N_20732,N_24231);
and U26272 (N_26272,N_23240,N_24359);
nor U26273 (N_26273,N_23723,N_24641);
nor U26274 (N_26274,N_23875,N_21706);
xor U26275 (N_26275,N_24713,N_23979);
or U26276 (N_26276,N_21219,N_21493);
and U26277 (N_26277,N_21141,N_22418);
nor U26278 (N_26278,N_21356,N_20076);
or U26279 (N_26279,N_22025,N_21432);
nor U26280 (N_26280,N_21428,N_24493);
nor U26281 (N_26281,N_24954,N_22603);
xor U26282 (N_26282,N_20496,N_22212);
or U26283 (N_26283,N_24460,N_23428);
nor U26284 (N_26284,N_20842,N_23047);
or U26285 (N_26285,N_24155,N_20331);
or U26286 (N_26286,N_21877,N_21632);
nor U26287 (N_26287,N_23706,N_24037);
and U26288 (N_26288,N_24497,N_21108);
and U26289 (N_26289,N_23595,N_22399);
nand U26290 (N_26290,N_23284,N_20204);
or U26291 (N_26291,N_22239,N_23819);
xnor U26292 (N_26292,N_20554,N_20559);
nor U26293 (N_26293,N_23845,N_23684);
nor U26294 (N_26294,N_20630,N_22290);
nand U26295 (N_26295,N_23445,N_20361);
and U26296 (N_26296,N_23113,N_20612);
and U26297 (N_26297,N_22704,N_24516);
xnor U26298 (N_26298,N_23420,N_21810);
xor U26299 (N_26299,N_21271,N_20654);
nand U26300 (N_26300,N_21469,N_20476);
or U26301 (N_26301,N_24399,N_23507);
and U26302 (N_26302,N_20984,N_22210);
and U26303 (N_26303,N_20655,N_23260);
xnor U26304 (N_26304,N_20868,N_23879);
xor U26305 (N_26305,N_22348,N_23000);
nor U26306 (N_26306,N_21415,N_22501);
xnor U26307 (N_26307,N_20917,N_20823);
nand U26308 (N_26308,N_22609,N_23628);
nor U26309 (N_26309,N_21381,N_20342);
nand U26310 (N_26310,N_24094,N_21675);
nor U26311 (N_26311,N_22524,N_23676);
nand U26312 (N_26312,N_20617,N_21134);
or U26313 (N_26313,N_24376,N_22034);
nand U26314 (N_26314,N_23545,N_23449);
nand U26315 (N_26315,N_23402,N_20235);
nor U26316 (N_26316,N_20825,N_23194);
and U26317 (N_26317,N_20013,N_20936);
xor U26318 (N_26318,N_21963,N_21846);
or U26319 (N_26319,N_23543,N_20091);
nor U26320 (N_26320,N_22517,N_24620);
or U26321 (N_26321,N_21923,N_21063);
nand U26322 (N_26322,N_20003,N_21317);
and U26323 (N_26323,N_20760,N_21392);
and U26324 (N_26324,N_21443,N_22896);
nand U26325 (N_26325,N_22709,N_21885);
xor U26326 (N_26326,N_20008,N_21573);
xnor U26327 (N_26327,N_20180,N_20620);
or U26328 (N_26328,N_24311,N_20026);
or U26329 (N_26329,N_22999,N_21264);
nor U26330 (N_26330,N_24114,N_22154);
xnor U26331 (N_26331,N_21112,N_24429);
or U26332 (N_26332,N_23597,N_21399);
or U26333 (N_26333,N_22741,N_23929);
or U26334 (N_26334,N_23863,N_21255);
xor U26335 (N_26335,N_24814,N_21315);
and U26336 (N_26336,N_24464,N_20735);
nand U26337 (N_26337,N_20761,N_24427);
or U26338 (N_26338,N_20943,N_21202);
nand U26339 (N_26339,N_23457,N_23982);
nor U26340 (N_26340,N_24039,N_21949);
nand U26341 (N_26341,N_22599,N_22949);
nand U26342 (N_26342,N_22788,N_23111);
or U26343 (N_26343,N_20116,N_21662);
nand U26344 (N_26344,N_22622,N_21073);
nand U26345 (N_26345,N_20215,N_20804);
xor U26346 (N_26346,N_22919,N_23658);
xnor U26347 (N_26347,N_23302,N_24980);
xnor U26348 (N_26348,N_20561,N_20624);
and U26349 (N_26349,N_22669,N_21709);
or U26350 (N_26350,N_20749,N_22677);
nand U26351 (N_26351,N_24065,N_24664);
nor U26352 (N_26352,N_23499,N_22890);
nor U26353 (N_26353,N_23404,N_21029);
or U26354 (N_26354,N_23755,N_20983);
and U26355 (N_26355,N_21750,N_24538);
and U26356 (N_26356,N_22897,N_24420);
or U26357 (N_26357,N_23841,N_23999);
or U26358 (N_26358,N_20080,N_22023);
and U26359 (N_26359,N_24652,N_24724);
nor U26360 (N_26360,N_21590,N_22364);
xor U26361 (N_26361,N_21633,N_24953);
or U26362 (N_26362,N_22571,N_24101);
and U26363 (N_26363,N_23513,N_24171);
or U26364 (N_26364,N_23605,N_20641);
and U26365 (N_26365,N_21940,N_21145);
and U26366 (N_26366,N_21369,N_23988);
or U26367 (N_26367,N_20038,N_22523);
xnor U26368 (N_26368,N_23169,N_24012);
nand U26369 (N_26369,N_24560,N_22351);
xnor U26370 (N_26370,N_23504,N_22583);
nand U26371 (N_26371,N_23093,N_22334);
and U26372 (N_26372,N_23789,N_20521);
or U26373 (N_26373,N_22157,N_23553);
or U26374 (N_26374,N_21044,N_21908);
or U26375 (N_26375,N_23066,N_20708);
xnor U26376 (N_26376,N_23870,N_20523);
nand U26377 (N_26377,N_21234,N_23004);
or U26378 (N_26378,N_21309,N_23462);
nand U26379 (N_26379,N_24213,N_20625);
nor U26380 (N_26380,N_23255,N_23836);
nor U26381 (N_26381,N_23156,N_23456);
nand U26382 (N_26382,N_22693,N_20152);
xor U26383 (N_26383,N_24496,N_23768);
or U26384 (N_26384,N_23378,N_20209);
nor U26385 (N_26385,N_22587,N_23050);
and U26386 (N_26386,N_21583,N_23686);
nor U26387 (N_26387,N_22608,N_24034);
nand U26388 (N_26388,N_24863,N_22266);
nand U26389 (N_26389,N_23188,N_20514);
nor U26390 (N_26390,N_23191,N_20490);
xor U26391 (N_26391,N_21205,N_20698);
nand U26392 (N_26392,N_23425,N_20015);
and U26393 (N_26393,N_22991,N_23868);
and U26394 (N_26394,N_21439,N_20360);
and U26395 (N_26395,N_24594,N_24854);
or U26396 (N_26396,N_24982,N_21862);
nand U26397 (N_26397,N_24826,N_23448);
nor U26398 (N_26398,N_21471,N_21697);
nand U26399 (N_26399,N_22813,N_21128);
and U26400 (N_26400,N_22987,N_22747);
or U26401 (N_26401,N_20104,N_20210);
nor U26402 (N_26402,N_23791,N_24558);
and U26403 (N_26403,N_21421,N_20567);
xnor U26404 (N_26404,N_24895,N_20011);
xnor U26405 (N_26405,N_24401,N_22688);
or U26406 (N_26406,N_22111,N_21820);
nor U26407 (N_26407,N_22986,N_23184);
or U26408 (N_26408,N_21193,N_22038);
xnor U26409 (N_26409,N_24772,N_22602);
xor U26410 (N_26410,N_24419,N_23059);
and U26411 (N_26411,N_21120,N_21466);
xnor U26412 (N_26412,N_23351,N_21462);
and U26413 (N_26413,N_20510,N_22560);
and U26414 (N_26414,N_23124,N_24244);
or U26415 (N_26415,N_21110,N_23946);
and U26416 (N_26416,N_24138,N_21436);
or U26417 (N_26417,N_23974,N_23392);
and U26418 (N_26418,N_20581,N_24111);
and U26419 (N_26419,N_20977,N_21064);
and U26420 (N_26420,N_23761,N_20491);
and U26421 (N_26421,N_22225,N_22794);
nor U26422 (N_26422,N_24728,N_23281);
or U26423 (N_26423,N_23435,N_22953);
and U26424 (N_26424,N_22745,N_23645);
and U26425 (N_26425,N_21232,N_24243);
and U26426 (N_26426,N_21897,N_24606);
nand U26427 (N_26427,N_21665,N_23663);
and U26428 (N_26428,N_21941,N_23466);
nand U26429 (N_26429,N_23850,N_21479);
and U26430 (N_26430,N_21751,N_21455);
or U26431 (N_26431,N_23349,N_24990);
nor U26432 (N_26432,N_20251,N_21250);
nand U26433 (N_26433,N_22754,N_20285);
xor U26434 (N_26434,N_22203,N_20686);
nand U26435 (N_26435,N_23477,N_20403);
nor U26436 (N_26436,N_24412,N_22710);
and U26437 (N_26437,N_23562,N_22304);
nor U26438 (N_26438,N_23480,N_24004);
nand U26439 (N_26439,N_24796,N_21931);
or U26440 (N_26440,N_24767,N_23679);
nor U26441 (N_26441,N_23471,N_20308);
or U26442 (N_26442,N_23669,N_20297);
or U26443 (N_26443,N_24776,N_23743);
nor U26444 (N_26444,N_22163,N_24541);
and U26445 (N_26445,N_22833,N_24131);
and U26446 (N_26446,N_24182,N_20187);
nand U26447 (N_26447,N_20169,N_21987);
nor U26448 (N_26448,N_24014,N_21636);
nor U26449 (N_26449,N_21042,N_21793);
nand U26450 (N_26450,N_20741,N_21176);
and U26451 (N_26451,N_23259,N_22254);
nor U26452 (N_26452,N_23824,N_21272);
or U26453 (N_26453,N_22699,N_22803);
nand U26454 (N_26454,N_20847,N_21888);
or U26455 (N_26455,N_22436,N_22209);
xor U26456 (N_26456,N_20260,N_20456);
and U26457 (N_26457,N_21607,N_20063);
nand U26458 (N_26458,N_21722,N_21887);
and U26459 (N_26459,N_20526,N_24252);
or U26460 (N_26460,N_22454,N_24815);
or U26461 (N_26461,N_23436,N_21008);
and U26462 (N_26462,N_21450,N_24595);
or U26463 (N_26463,N_22092,N_23454);
or U26464 (N_26464,N_23866,N_24843);
nand U26465 (N_26465,N_21506,N_23205);
xnor U26466 (N_26466,N_20500,N_20629);
and U26467 (N_26467,N_21211,N_24596);
or U26468 (N_26468,N_23867,N_24073);
and U26469 (N_26469,N_23872,N_22572);
and U26470 (N_26470,N_22201,N_22357);
xor U26471 (N_26471,N_20455,N_24653);
or U26472 (N_26472,N_20031,N_24333);
or U26473 (N_26473,N_24390,N_23076);
and U26474 (N_26474,N_22584,N_22731);
and U26475 (N_26475,N_22162,N_20195);
nor U26476 (N_26476,N_23800,N_22616);
or U26477 (N_26477,N_23600,N_22235);
nor U26478 (N_26478,N_20097,N_21490);
or U26479 (N_26479,N_24466,N_22176);
nand U26480 (N_26480,N_22761,N_23148);
nor U26481 (N_26481,N_23032,N_24173);
and U26482 (N_26482,N_24454,N_20532);
nand U26483 (N_26483,N_21742,N_24280);
and U26484 (N_26484,N_24827,N_20256);
and U26485 (N_26485,N_20528,N_24282);
and U26486 (N_26486,N_22330,N_21213);
nand U26487 (N_26487,N_20547,N_20889);
nor U26488 (N_26488,N_20793,N_23807);
nand U26489 (N_26489,N_23701,N_24571);
nand U26490 (N_26490,N_24636,N_24428);
xnor U26491 (N_26491,N_24218,N_22435);
nand U26492 (N_26492,N_24494,N_23311);
or U26493 (N_26493,N_23983,N_23080);
nand U26494 (N_26494,N_24614,N_21855);
nand U26495 (N_26495,N_21667,N_20922);
nand U26496 (N_26496,N_21596,N_23616);
and U26497 (N_26497,N_24380,N_20083);
xnor U26498 (N_26498,N_20487,N_22258);
or U26499 (N_26499,N_24211,N_21027);
nand U26500 (N_26500,N_23783,N_20002);
and U26501 (N_26501,N_20024,N_21856);
nand U26502 (N_26502,N_20670,N_23575);
nand U26503 (N_26503,N_20469,N_22577);
nor U26504 (N_26504,N_22385,N_23383);
nand U26505 (N_26505,N_20114,N_21774);
xor U26506 (N_26506,N_24312,N_24812);
or U26507 (N_26507,N_22843,N_22667);
nor U26508 (N_26508,N_22841,N_23976);
nor U26509 (N_26509,N_20181,N_23775);
and U26510 (N_26510,N_22951,N_20483);
nand U26511 (N_26511,N_21183,N_24317);
xor U26512 (N_26512,N_20269,N_24499);
nor U26513 (N_26513,N_22907,N_23128);
nor U26514 (N_26514,N_24991,N_24281);
nand U26515 (N_26515,N_20946,N_23564);
or U26516 (N_26516,N_20061,N_23422);
xnor U26517 (N_26517,N_24475,N_24350);
nand U26518 (N_26518,N_23648,N_20631);
or U26519 (N_26519,N_23830,N_21920);
nand U26520 (N_26520,N_22369,N_24758);
xnor U26521 (N_26521,N_21365,N_23817);
nor U26522 (N_26522,N_24592,N_22102);
nor U26523 (N_26523,N_24077,N_22227);
and U26524 (N_26524,N_21869,N_22001);
and U26525 (N_26525,N_23264,N_20734);
nand U26526 (N_26526,N_20767,N_21892);
nand U26527 (N_26527,N_22017,N_24269);
or U26528 (N_26528,N_22138,N_22780);
and U26529 (N_26529,N_21390,N_22056);
nand U26530 (N_26530,N_21152,N_21986);
xnor U26531 (N_26531,N_21641,N_20155);
xnor U26532 (N_26532,N_21295,N_22939);
xnor U26533 (N_26533,N_23127,N_20738);
xnor U26534 (N_26534,N_23670,N_24120);
xor U26535 (N_26535,N_20060,N_22567);
nor U26536 (N_26536,N_22944,N_23610);
nand U26537 (N_26537,N_22502,N_22481);
or U26538 (N_26538,N_22421,N_21261);
or U26539 (N_26539,N_20286,N_21424);
nor U26540 (N_26540,N_22673,N_21806);
nand U26541 (N_26541,N_24726,N_22582);
nand U26542 (N_26542,N_20648,N_20041);
nor U26543 (N_26543,N_24786,N_22220);
nor U26544 (N_26544,N_21106,N_22371);
or U26545 (N_26545,N_20157,N_20354);
xnor U26546 (N_26546,N_20275,N_24164);
or U26547 (N_26547,N_20867,N_24917);
nor U26548 (N_26548,N_20862,N_22336);
nor U26549 (N_26549,N_23574,N_24733);
nand U26550 (N_26550,N_21677,N_21089);
nor U26551 (N_26551,N_21056,N_24217);
nand U26552 (N_26552,N_23730,N_24875);
or U26553 (N_26553,N_20896,N_20106);
and U26554 (N_26554,N_21048,N_22905);
and U26555 (N_26555,N_22380,N_24086);
xor U26556 (N_26556,N_24878,N_24927);
nand U26557 (N_26557,N_20945,N_22216);
nand U26558 (N_26558,N_24199,N_21306);
xnor U26559 (N_26559,N_22992,N_23874);
nand U26560 (N_26560,N_21049,N_24330);
or U26561 (N_26561,N_20189,N_21321);
or U26562 (N_26562,N_20959,N_22970);
or U26563 (N_26563,N_21755,N_22565);
or U26564 (N_26564,N_23110,N_21540);
nor U26565 (N_26565,N_21650,N_23894);
xor U26566 (N_26566,N_21759,N_23823);
xnor U26567 (N_26567,N_22433,N_20765);
nand U26568 (N_26568,N_23330,N_22773);
and U26569 (N_26569,N_21137,N_24323);
nand U26570 (N_26570,N_21655,N_22037);
or U26571 (N_26571,N_22489,N_20955);
and U26572 (N_26572,N_24123,N_23917);
nor U26573 (N_26573,N_23131,N_21200);
nor U26574 (N_26574,N_21147,N_21795);
nand U26575 (N_26575,N_20866,N_23523);
or U26576 (N_26576,N_21235,N_24445);
nand U26577 (N_26577,N_22395,N_20087);
xor U26578 (N_26578,N_23043,N_24373);
and U26579 (N_26579,N_20054,N_20039);
or U26580 (N_26580,N_24672,N_21644);
and U26581 (N_26581,N_24176,N_22086);
xnor U26582 (N_26582,N_21040,N_23486);
xor U26583 (N_26583,N_20819,N_22835);
xnor U26584 (N_26584,N_22109,N_23034);
nand U26585 (N_26585,N_24154,N_21867);
xor U26586 (N_26586,N_24621,N_23925);
nand U26587 (N_26587,N_20509,N_22631);
nor U26588 (N_26588,N_24361,N_20045);
or U26589 (N_26589,N_22532,N_24605);
and U26590 (N_26590,N_24434,N_23337);
nand U26591 (N_26591,N_22828,N_23918);
and U26592 (N_26592,N_20383,N_21308);
xor U26593 (N_26593,N_20376,N_23699);
and U26594 (N_26594,N_21046,N_21899);
and U26595 (N_26595,N_24437,N_22815);
xor U26596 (N_26596,N_22049,N_21201);
or U26597 (N_26597,N_23667,N_20464);
nor U26598 (N_26598,N_21170,N_24984);
and U26599 (N_26599,N_21785,N_21603);
nor U26600 (N_26600,N_24887,N_20974);
or U26601 (N_26601,N_22312,N_23989);
nor U26602 (N_26602,N_21684,N_20998);
nor U26603 (N_26603,N_20901,N_22360);
xnor U26604 (N_26604,N_23494,N_21430);
or U26605 (N_26605,N_22482,N_20307);
or U26606 (N_26606,N_24140,N_23157);
xnor U26607 (N_26607,N_21617,N_20714);
nor U26608 (N_26608,N_23015,N_20480);
nor U26609 (N_26609,N_21689,N_24214);
nor U26610 (N_26610,N_24633,N_23885);
and U26611 (N_26611,N_23315,N_24327);
nor U26612 (N_26612,N_22825,N_20935);
and U26613 (N_26613,N_22189,N_24585);
and U26614 (N_26614,N_23027,N_20478);
xor U26615 (N_26615,N_21979,N_22887);
or U26616 (N_26616,N_21807,N_20247);
nand U26617 (N_26617,N_23957,N_22505);
and U26618 (N_26618,N_20972,N_22668);
xnor U26619 (N_26619,N_23967,N_21643);
or U26620 (N_26620,N_24638,N_23517);
and U26621 (N_26621,N_22374,N_20657);
and U26622 (N_26622,N_23766,N_23852);
and U26623 (N_26623,N_21852,N_24469);
xnor U26624 (N_26624,N_21950,N_21692);
nor U26625 (N_26625,N_23758,N_21065);
nand U26626 (N_26626,N_23992,N_24055);
nor U26627 (N_26627,N_23666,N_20234);
xnor U26628 (N_26628,N_21611,N_21623);
nand U26629 (N_26629,N_24414,N_24265);
xnor U26630 (N_26630,N_23203,N_21055);
or U26631 (N_26631,N_22759,N_22425);
or U26632 (N_26632,N_20632,N_24970);
nor U26633 (N_26633,N_21162,N_24877);
nor U26634 (N_26634,N_21889,N_23877);
and U26635 (N_26635,N_24915,N_23737);
nand U26636 (N_26636,N_23040,N_20603);
xor U26637 (N_26637,N_24500,N_24806);
nor U26638 (N_26638,N_24283,N_24589);
xnor U26639 (N_26639,N_21695,N_21009);
nor U26640 (N_26640,N_23919,N_21621);
or U26641 (N_26641,N_22545,N_23598);
or U26642 (N_26642,N_24899,N_21976);
xnor U26643 (N_26643,N_21513,N_23399);
nor U26644 (N_26644,N_20325,N_24241);
or U26645 (N_26645,N_23735,N_22837);
nor U26646 (N_26646,N_24254,N_20729);
and U26647 (N_26647,N_23490,N_24751);
or U26648 (N_26648,N_20338,N_23365);
and U26649 (N_26649,N_20742,N_22105);
nand U26650 (N_26650,N_21800,N_21882);
nand U26651 (N_26651,N_24426,N_22277);
xor U26652 (N_26652,N_23164,N_21494);
and U26653 (N_26653,N_21647,N_23150);
or U26654 (N_26654,N_24484,N_24971);
or U26655 (N_26655,N_22827,N_20420);
xnor U26656 (N_26656,N_20593,N_23756);
or U26657 (N_26657,N_24998,N_22031);
nor U26658 (N_26658,N_23320,N_24738);
and U26659 (N_26659,N_23945,N_24768);
nand U26660 (N_26660,N_22311,N_23795);
xor U26661 (N_26661,N_23802,N_20158);
and U26662 (N_26662,N_20798,N_21971);
or U26663 (N_26663,N_22546,N_22554);
nor U26664 (N_26664,N_22294,N_22564);
and U26665 (N_26665,N_22698,N_22260);
nand U26666 (N_26666,N_21683,N_20356);
nor U26667 (N_26667,N_22292,N_21988);
or U26668 (N_26668,N_23884,N_24069);
and U26669 (N_26669,N_23433,N_20029);
and U26670 (N_26670,N_24258,N_23432);
and U26671 (N_26671,N_23369,N_22787);
and U26672 (N_26672,N_22337,N_22340);
xor U26673 (N_26673,N_20028,N_20682);
or U26674 (N_26674,N_24615,N_22865);
nand U26675 (N_26675,N_23942,N_23067);
and U26676 (N_26676,N_22624,N_24540);
and U26677 (N_26677,N_22120,N_24256);
xnor U26678 (N_26678,N_21444,N_23618);
xor U26679 (N_26679,N_23579,N_24402);
xnor U26680 (N_26680,N_22316,N_23160);
or U26681 (N_26681,N_23759,N_24177);
nand U26682 (N_26682,N_24981,N_23907);
and U26683 (N_26683,N_21053,N_21533);
xnor U26684 (N_26684,N_23033,N_24228);
nor U26685 (N_26685,N_24150,N_21244);
xor U26686 (N_26686,N_21629,N_22962);
xnor U26687 (N_26687,N_24869,N_23248);
or U26688 (N_26688,N_24204,N_20511);
nor U26689 (N_26689,N_23567,N_24818);
or U26690 (N_26690,N_22275,N_20377);
nor U26691 (N_26691,N_22098,N_22344);
and U26692 (N_26692,N_20786,N_24161);
nand U26693 (N_26693,N_20913,N_22413);
and U26694 (N_26694,N_23006,N_24071);
or U26695 (N_26695,N_21521,N_24622);
xnor U26696 (N_26696,N_22988,N_22867);
and U26697 (N_26697,N_22287,N_20149);
nand U26698 (N_26698,N_23329,N_23060);
xnor U26699 (N_26699,N_24066,N_21132);
xnor U26700 (N_26700,N_21878,N_22416);
xnor U26701 (N_26701,N_22028,N_20725);
xor U26702 (N_26702,N_21224,N_22053);
xnor U26703 (N_26703,N_24320,N_24160);
and U26704 (N_26704,N_21981,N_21508);
nand U26705 (N_26705,N_22423,N_24298);
or U26706 (N_26706,N_24089,N_20914);
and U26707 (N_26707,N_22205,N_22107);
nor U26708 (N_26708,N_20430,N_20748);
xor U26709 (N_26709,N_20664,N_21035);
nor U26710 (N_26710,N_20434,N_22094);
nor U26711 (N_26711,N_23638,N_23221);
nor U26712 (N_26712,N_23373,N_21289);
nand U26713 (N_26713,N_22633,N_20052);
xor U26714 (N_26714,N_20179,N_24531);
xor U26715 (N_26715,N_24870,N_22243);
nor U26716 (N_26716,N_24001,N_23744);
nor U26717 (N_26717,N_22715,N_24756);
nor U26718 (N_26718,N_21422,N_23133);
or U26719 (N_26719,N_23602,N_22283);
and U26720 (N_26720,N_21160,N_23838);
xor U26721 (N_26721,N_21113,N_22151);
nand U26722 (N_26722,N_20755,N_23455);
xnor U26723 (N_26723,N_20281,N_23821);
nor U26724 (N_26724,N_22846,N_22496);
and U26725 (N_26725,N_20139,N_20326);
and U26726 (N_26726,N_23489,N_20829);
xnor U26727 (N_26727,N_24325,N_21884);
and U26728 (N_26728,N_21589,N_23892);
nor U26729 (N_26729,N_20701,N_20272);
xor U26730 (N_26730,N_21880,N_24005);
nand U26731 (N_26731,N_22864,N_21876);
nor U26732 (N_26732,N_20306,N_21989);
nand U26733 (N_26733,N_21492,N_24695);
nor U26734 (N_26734,N_20722,N_23253);
xor U26735 (N_26735,N_21791,N_23714);
nand U26736 (N_26736,N_21788,N_24142);
and U26737 (N_26737,N_22143,N_22291);
xnor U26738 (N_26738,N_22429,N_23938);
nor U26739 (N_26739,N_22627,N_21225);
xnor U26740 (N_26740,N_21195,N_21398);
nor U26741 (N_26741,N_22732,N_22652);
and U26742 (N_26742,N_20237,N_22997);
and U26743 (N_26743,N_21864,N_23927);
xnor U26744 (N_26744,N_24377,N_21331);
xnor U26745 (N_26745,N_24348,N_22503);
nor U26746 (N_26746,N_22458,N_24410);
and U26747 (N_26747,N_24608,N_22152);
and U26748 (N_26748,N_21256,N_23916);
and U26749 (N_26749,N_20352,N_21127);
and U26750 (N_26750,N_23135,N_22406);
xnor U26751 (N_26751,N_24613,N_24892);
or U26752 (N_26752,N_22174,N_22148);
and U26753 (N_26753,N_21078,N_24557);
xor U26754 (N_26754,N_22685,N_22467);
nand U26755 (N_26755,N_22200,N_23473);
or U26756 (N_26756,N_22834,N_22961);
or U26757 (N_26757,N_20880,N_23588);
nor U26758 (N_26758,N_22315,N_23556);
nor U26759 (N_26759,N_20042,N_21054);
xor U26760 (N_26760,N_24681,N_22703);
or U26761 (N_26761,N_23460,N_21233);
nand U26762 (N_26762,N_22639,N_20160);
xnor U26763 (N_26763,N_20398,N_20811);
xnor U26764 (N_26764,N_24250,N_23898);
nand U26765 (N_26765,N_21088,N_23843);
nand U26766 (N_26766,N_21766,N_20930);
nand U26767 (N_26767,N_22520,N_24147);
or U26768 (N_26768,N_24922,N_20270);
nand U26769 (N_26769,N_23814,N_20333);
nand U26770 (N_26770,N_21843,N_20214);
or U26771 (N_26771,N_20121,N_23832);
nor U26772 (N_26772,N_23533,N_22785);
and U26773 (N_26773,N_22251,N_24389);
or U26774 (N_26774,N_21537,N_20961);
and U26775 (N_26775,N_24413,N_20369);
nand U26776 (N_26776,N_21748,N_23277);
nand U26777 (N_26777,N_20473,N_24503);
and U26778 (N_26778,N_21932,N_24921);
xnor U26779 (N_26779,N_23285,N_21853);
nand U26780 (N_26780,N_24684,N_20633);
and U26781 (N_26781,N_23086,N_20349);
nand U26782 (N_26782,N_21659,N_23100);
or U26783 (N_26783,N_23412,N_22009);
nand U26784 (N_26784,N_21477,N_24752);
xor U26785 (N_26785,N_22223,N_21977);
xnor U26786 (N_26786,N_23411,N_24381);
nand U26787 (N_26787,N_22126,N_23511);
and U26788 (N_26788,N_24873,N_21673);
or U26789 (N_26789,N_21335,N_24472);
nor U26790 (N_26790,N_20086,N_23774);
and U26791 (N_26791,N_20386,N_24884);
or U26792 (N_26792,N_20542,N_21124);
nand U26793 (N_26793,N_22426,N_22133);
nor U26794 (N_26794,N_22323,N_24952);
nor U26795 (N_26795,N_22573,N_21386);
or U26796 (N_26796,N_21173,N_23637);
xnor U26797 (N_26797,N_24942,N_22783);
xnor U26798 (N_26798,N_24002,N_20942);
and U26799 (N_26799,N_21919,N_20463);
xor U26800 (N_26800,N_21612,N_20642);
and U26801 (N_26801,N_23975,N_23396);
nand U26802 (N_26802,N_22469,N_22891);
and U26803 (N_26803,N_24840,N_20148);
xor U26804 (N_26804,N_23010,N_20069);
and U26805 (N_26805,N_21966,N_24570);
nor U26806 (N_26806,N_24909,N_23413);
xnor U26807 (N_26807,N_20551,N_21318);
nand U26808 (N_26808,N_23174,N_22076);
xnor U26809 (N_26809,N_22589,N_21817);
or U26810 (N_26810,N_20425,N_20367);
nand U26811 (N_26811,N_22979,N_22368);
and U26812 (N_26812,N_20440,N_24284);
nor U26813 (N_26813,N_21532,N_23585);
and U26814 (N_26814,N_23978,N_20563);
nor U26815 (N_26815,N_24341,N_22363);
nand U26816 (N_26816,N_24079,N_22792);
nor U26817 (N_26817,N_22922,N_21017);
nor U26818 (N_26818,N_21131,N_23614);
nor U26819 (N_26819,N_21252,N_21416);
or U26820 (N_26820,N_22592,N_22166);
xnor U26821 (N_26821,N_22464,N_21886);
or U26822 (N_26822,N_22651,N_21338);
nand U26823 (N_26823,N_21529,N_23139);
nor U26824 (N_26824,N_20396,N_22134);
and U26825 (N_26825,N_20236,N_24833);
nor U26826 (N_26826,N_24901,N_22537);
or U26827 (N_26827,N_20252,N_23691);
and U26828 (N_26828,N_24908,N_22296);
nand U26829 (N_26829,N_22547,N_24740);
nor U26830 (N_26830,N_24603,N_24011);
xnor U26831 (N_26831,N_22934,N_24515);
or U26832 (N_26832,N_20751,N_20650);
nand U26833 (N_26833,N_23599,N_20791);
and U26834 (N_26834,N_22829,N_24060);
xnor U26835 (N_26835,N_20202,N_21823);
nand U26836 (N_26836,N_24268,N_23092);
or U26837 (N_26837,N_22510,N_23495);
and U26838 (N_26838,N_21510,N_22237);
nor U26839 (N_26839,N_23387,N_20826);
and U26840 (N_26840,N_21764,N_24951);
nor U26841 (N_26841,N_23270,N_22621);
or U26842 (N_26842,N_22447,N_21646);
nand U26843 (N_26843,N_21144,N_21725);
or U26844 (N_26844,N_23653,N_20058);
xor U26845 (N_26845,N_21634,N_22301);
or U26846 (N_26846,N_22343,N_24491);
xnor U26847 (N_26847,N_24166,N_24396);
and U26848 (N_26848,N_20292,N_24354);
nor U26849 (N_26849,N_20571,N_23678);
and U26850 (N_26850,N_20888,N_22644);
nor U26851 (N_26851,N_23044,N_21074);
or U26852 (N_26852,N_21360,N_20112);
or U26853 (N_26853,N_22539,N_20613);
and U26854 (N_26854,N_22558,N_24783);
or U26855 (N_26855,N_22246,N_20941);
nor U26856 (N_26856,N_22893,N_24773);
and U26857 (N_26857,N_24577,N_22193);
and U26858 (N_26858,N_21606,N_22640);
nand U26859 (N_26859,N_21993,N_22654);
nand U26860 (N_26860,N_23231,N_23228);
xnor U26861 (N_26861,N_23803,N_20909);
xor U26862 (N_26862,N_23736,N_24905);
nor U26863 (N_26863,N_20881,N_20142);
nand U26864 (N_26864,N_20562,N_21758);
nand U26865 (N_26865,N_21222,N_21060);
nand U26866 (N_26866,N_20131,N_23305);
nor U26867 (N_26867,N_21483,N_24453);
or U26868 (N_26868,N_22027,N_20951);
or U26869 (N_26869,N_20005,N_22202);
and U26870 (N_26870,N_22156,N_20779);
and U26871 (N_26871,N_21531,N_22140);
or U26872 (N_26872,N_23781,N_24780);
xor U26873 (N_26873,N_23167,N_20788);
xor U26874 (N_26874,N_24307,N_21708);
xnor U26875 (N_26875,N_20065,N_23831);
and U26876 (N_26876,N_23577,N_21000);
xor U26877 (N_26877,N_21900,N_20614);
xnor U26878 (N_26878,N_20098,N_24299);
and U26879 (N_26879,N_23788,N_20446);
xnor U26880 (N_26880,N_24202,N_20239);
and U26881 (N_26881,N_22207,N_24654);
nand U26882 (N_26882,N_20222,N_24739);
xor U26883 (N_26883,N_24720,N_22284);
nor U26884 (N_26884,N_20093,N_24949);
nand U26885 (N_26885,N_21557,N_20869);
and U26886 (N_26886,N_22765,N_21515);
xor U26887 (N_26887,N_23913,N_23697);
nor U26888 (N_26888,N_21408,N_20950);
nor U26889 (N_26889,N_20573,N_24212);
and U26890 (N_26890,N_20423,N_20822);
and U26891 (N_26891,N_21093,N_20190);
and U26892 (N_26892,N_24764,N_21535);
nor U26893 (N_26893,N_22045,N_20067);
or U26894 (N_26894,N_21586,N_23738);
and U26895 (N_26895,N_21452,N_23222);
nand U26896 (N_26896,N_21357,N_21906);
nor U26897 (N_26897,N_20399,N_20416);
or U26898 (N_26898,N_22770,N_21830);
and U26899 (N_26899,N_23267,N_22937);
or U26900 (N_26900,N_23772,N_22414);
or U26901 (N_26901,N_21685,N_20769);
nand U26902 (N_26902,N_24488,N_22150);
nor U26903 (N_26903,N_20783,N_22743);
xor U26904 (N_26904,N_20410,N_21258);
nand U26905 (N_26905,N_22234,N_21151);
and U26906 (N_26906,N_22069,N_22401);
xnor U26907 (N_26907,N_21952,N_23464);
nor U26908 (N_26908,N_22090,N_24881);
nor U26909 (N_26909,N_22432,N_21660);
and U26910 (N_26910,N_24559,N_20578);
nor U26911 (N_26911,N_24456,N_20409);
and U26912 (N_26912,N_23491,N_24722);
and U26913 (N_26913,N_20981,N_24267);
nand U26914 (N_26914,N_22707,N_22984);
or U26915 (N_26915,N_21082,N_23405);
nor U26916 (N_26916,N_21951,N_22516);
and U26917 (N_26917,N_21401,N_20546);
xnor U26918 (N_26918,N_20680,N_24406);
or U26919 (N_26919,N_24545,N_23012);
nand U26920 (N_26920,N_21680,N_22641);
xor U26921 (N_26921,N_24058,N_22096);
or U26922 (N_26922,N_24795,N_22744);
xor U26923 (N_26923,N_21967,N_23778);
or U26924 (N_26924,N_21745,N_21165);
xnor U26925 (N_26925,N_22894,N_24233);
or U26926 (N_26926,N_24452,N_23181);
nor U26927 (N_26927,N_20194,N_22442);
nand U26928 (N_26928,N_23087,N_20802);
and U26929 (N_26929,N_21601,N_24974);
xor U26930 (N_26930,N_22322,N_24141);
and U26931 (N_26931,N_21936,N_21412);
xnor U26932 (N_26932,N_21361,N_23608);
and U26933 (N_26933,N_23286,N_23801);
and U26934 (N_26934,N_23344,N_23042);
nor U26935 (N_26935,N_22527,N_20605);
and U26936 (N_26936,N_21389,N_21938);
xnor U26937 (N_26937,N_23451,N_24599);
nand U26938 (N_26938,N_21344,N_22041);
nor U26939 (N_26939,N_20719,N_23001);
nor U26940 (N_26940,N_23636,N_23102);
and U26941 (N_26941,N_22439,N_22078);
xnor U26942 (N_26942,N_24872,N_20570);
nor U26943 (N_26943,N_22087,N_22491);
xnor U26944 (N_26944,N_24386,N_24809);
nand U26945 (N_26945,N_21410,N_23348);
or U26946 (N_26946,N_20223,N_24170);
nor U26947 (N_26947,N_22854,N_24987);
nand U26948 (N_26948,N_22613,N_23072);
and U26949 (N_26949,N_23643,N_21756);
nor U26950 (N_26950,N_21034,N_20673);
and U26951 (N_26951,N_24112,N_20870);
and U26952 (N_26952,N_21172,N_20882);
nand U26953 (N_26953,N_23725,N_24279);
or U26954 (N_26954,N_24223,N_23501);
nor U26955 (N_26955,N_22054,N_23712);
and U26956 (N_26956,N_23950,N_24858);
nand U26957 (N_26957,N_24885,N_24169);
or U26958 (N_26958,N_22068,N_23552);
nor U26959 (N_26959,N_23741,N_20659);
or U26960 (N_26960,N_20724,N_24825);
xor U26961 (N_26961,N_23483,N_24236);
xnor U26962 (N_26962,N_23720,N_24598);
nor U26963 (N_26963,N_22384,N_20113);
nand U26964 (N_26964,N_21995,N_24197);
nand U26965 (N_26965,N_22597,N_23416);
nor U26966 (N_26966,N_24483,N_21678);
or U26967 (N_26967,N_22989,N_23911);
nand U26968 (N_26968,N_22046,N_20199);
and U26969 (N_26969,N_20710,N_23935);
nand U26970 (N_26970,N_24820,N_22548);
and U26971 (N_26971,N_22914,N_22470);
or U26972 (N_26972,N_24674,N_24836);
nor U26973 (N_26973,N_24813,N_20475);
or U26974 (N_26974,N_22457,N_23677);
xnor U26975 (N_26975,N_21092,N_23294);
xor U26976 (N_26976,N_21809,N_21654);
and U26977 (N_26977,N_23926,N_22855);
nand U26978 (N_26978,N_22575,N_20997);
nor U26979 (N_26979,N_24996,N_22492);
xor U26980 (N_26980,N_23271,N_23991);
xor U26981 (N_26981,N_23541,N_22305);
and U26982 (N_26982,N_22456,N_23019);
nor U26983 (N_26983,N_23855,N_21090);
xnor U26984 (N_26984,N_24574,N_23453);
or U26985 (N_26985,N_22797,N_23705);
nor U26986 (N_26986,N_20078,N_24062);
and U26987 (N_26987,N_20815,N_21998);
and U26988 (N_26988,N_22448,N_24290);
nand U26989 (N_26989,N_20278,N_23731);
and U26990 (N_26990,N_21895,N_24322);
or U26991 (N_26991,N_24442,N_20937);
nor U26992 (N_26992,N_20101,N_23790);
xor U26993 (N_26993,N_24457,N_22326);
nand U26994 (N_26994,N_22167,N_24266);
or U26995 (N_26995,N_20337,N_20816);
and U26996 (N_26996,N_24295,N_22903);
xor U26997 (N_26997,N_22662,N_20774);
xor U26998 (N_26998,N_21026,N_23237);
xor U26999 (N_26999,N_23799,N_20627);
xnor U27000 (N_27000,N_24727,N_23082);
nand U27001 (N_27001,N_21472,N_22179);
nor U27002 (N_27002,N_20807,N_22932);
or U27003 (N_27003,N_24443,N_22088);
nor U27004 (N_27004,N_23786,N_22265);
nand U27005 (N_27005,N_21903,N_21545);
nand U27006 (N_27006,N_24861,N_24423);
nor U27007 (N_27007,N_23987,N_24135);
nor U27008 (N_27008,N_23887,N_24803);
nor U27009 (N_27009,N_22757,N_22751);
or U27010 (N_27010,N_24288,N_23811);
nand U27011 (N_27011,N_24718,N_22660);
nor U27012 (N_27012,N_20640,N_20679);
xnor U27013 (N_27013,N_21956,N_22634);
and U27014 (N_27014,N_20875,N_22900);
nand U27015 (N_27015,N_23361,N_21894);
nor U27016 (N_27016,N_22443,N_23340);
nand U27017 (N_27017,N_21790,N_22286);
xnor U27018 (N_27018,N_23642,N_22878);
and U27019 (N_27019,N_22875,N_24326);
or U27020 (N_27020,N_21816,N_20658);
and U27021 (N_27021,N_22453,N_23937);
nor U27022 (N_27022,N_24842,N_24103);
and U27023 (N_27023,N_24708,N_22144);
nand U27024 (N_27024,N_21944,N_24610);
xnor U27025 (N_27025,N_23512,N_23258);
or U27026 (N_27026,N_22862,N_21240);
xnor U27027 (N_27027,N_24944,N_22021);
nand U27028 (N_27028,N_22689,N_20898);
nor U27029 (N_27029,N_21299,N_21904);
xor U27030 (N_27030,N_23915,N_23206);
nor U27031 (N_27031,N_22522,N_23912);
nor U27032 (N_27032,N_20334,N_20175);
and U27033 (N_27033,N_21326,N_23968);
nand U27034 (N_27034,N_21797,N_20282);
nand U27035 (N_27035,N_23960,N_22488);
xnor U27036 (N_27036,N_20707,N_22716);
nor U27037 (N_27037,N_23476,N_22249);
or U27038 (N_27038,N_22437,N_21776);
nor U27039 (N_27039,N_20447,N_24683);
or U27040 (N_27040,N_24568,N_21281);
nor U27041 (N_27041,N_23039,N_21248);
nor U27042 (N_27042,N_23375,N_22802);
and U27043 (N_27043,N_22923,N_21166);
and U27044 (N_27044,N_24473,N_24866);
nor U27045 (N_27045,N_22452,N_23068);
nor U27046 (N_27046,N_22550,N_20574);
nand U27047 (N_27047,N_24530,N_21210);
or U27048 (N_27048,N_24696,N_23969);
nor U27049 (N_27049,N_23985,N_22341);
and U27050 (N_27050,N_24932,N_22541);
or U27051 (N_27051,N_22499,N_20431);
nor U27052 (N_27052,N_20845,N_23549);
and U27053 (N_27053,N_21767,N_24802);
or U27054 (N_27054,N_23317,N_22217);
xor U27055 (N_27055,N_21544,N_23114);
nand U27056 (N_27056,N_20299,N_20211);
nor U27057 (N_27057,N_24461,N_20424);
xor U27058 (N_27058,N_21041,N_21930);
nor U27059 (N_27059,N_24339,N_21789);
and U27060 (N_27060,N_21010,N_22664);
xor U27061 (N_27061,N_22619,N_24874);
and U27062 (N_27062,N_20944,N_20012);
nand U27063 (N_27063,N_21934,N_23346);
or U27064 (N_27064,N_20926,N_24207);
and U27065 (N_27065,N_20096,N_22402);
and U27066 (N_27066,N_20284,N_22758);
nor U27067 (N_27067,N_24735,N_20277);
nor U27068 (N_27068,N_24588,N_21400);
nor U27069 (N_27069,N_20830,N_24438);
xor U27070 (N_27070,N_21500,N_21779);
nand U27071 (N_27071,N_23296,N_24963);
xnor U27072 (N_27072,N_20986,N_22400);
or U27073 (N_27073,N_23022,N_23045);
nand U27074 (N_27074,N_24966,N_20817);
and U27075 (N_27075,N_24117,N_22911);
nor U27076 (N_27076,N_24923,N_21898);
or U27077 (N_27077,N_22242,N_21229);
and U27078 (N_27078,N_20668,N_23681);
and U27079 (N_27079,N_21734,N_20903);
or U27080 (N_27080,N_22392,N_22972);
nor U27081 (N_27081,N_22494,N_20855);
nor U27082 (N_27082,N_24379,N_23798);
nand U27083 (N_27083,N_21743,N_24370);
xnor U27084 (N_27084,N_24587,N_20501);
or U27085 (N_27085,N_23123,N_20460);
nor U27086 (N_27086,N_24524,N_20667);
nand U27087 (N_27087,N_21133,N_22892);
and U27088 (N_27088,N_20375,N_22819);
nand U27089 (N_27089,N_21896,N_22985);
xor U27090 (N_27090,N_20439,N_21262);
or U27091 (N_27091,N_20150,N_22272);
nor U27092 (N_27092,N_23353,N_20537);
or U27093 (N_27093,N_23633,N_23540);
or U27094 (N_27094,N_20849,N_20317);
or U27095 (N_27095,N_21476,N_23776);
nor U27096 (N_27096,N_22356,N_24821);
and U27097 (N_27097,N_22826,N_24335);
nand U27098 (N_27098,N_21699,N_23820);
or U27099 (N_27099,N_23249,N_23784);
nand U27100 (N_27100,N_20690,N_24229);
or U27101 (N_27101,N_22938,N_20241);
or U27102 (N_27102,N_22115,N_21608);
nand U27103 (N_27103,N_21502,N_24865);
xor U27104 (N_27104,N_23849,N_20102);
nor U27105 (N_27105,N_22206,N_20232);
xnor U27106 (N_27106,N_23858,N_23354);
nor U27107 (N_27107,N_20597,N_23467);
nor U27108 (N_27108,N_21713,N_23214);
xor U27109 (N_27109,N_24512,N_20047);
and U27110 (N_27110,N_20948,N_23434);
and U27111 (N_27111,N_23662,N_21005);
or U27112 (N_27112,N_24270,N_24355);
or U27113 (N_27113,N_24525,N_24582);
and U27114 (N_27114,N_21263,N_23359);
xnor U27115 (N_27115,N_23147,N_23805);
or U27116 (N_27116,N_21604,N_22060);
xor U27117 (N_27117,N_24640,N_23421);
and U27118 (N_27118,N_21486,N_21003);
xnor U27119 (N_27119,N_20789,N_23389);
xor U27120 (N_27120,N_21103,N_20068);
xor U27121 (N_27121,N_20316,N_24403);
and U27122 (N_27122,N_21043,N_22586);
or U27123 (N_27123,N_20238,N_22365);
xnor U27124 (N_27124,N_24745,N_22861);
nand U27125 (N_27125,N_22725,N_24482);
and U27126 (N_27126,N_24463,N_24385);
xnor U27127 (N_27127,N_20718,N_22236);
nand U27128 (N_27128,N_24775,N_22665);
nand U27129 (N_27129,N_23623,N_20989);
xor U27130 (N_27130,N_20739,N_21033);
nand U27131 (N_27131,N_22465,N_23607);
or U27132 (N_27132,N_22218,N_24132);
or U27133 (N_27133,N_23639,N_20887);
nor U27134 (N_27134,N_24433,N_23895);
nor U27135 (N_27135,N_23325,N_20806);
nand U27136 (N_27136,N_24627,N_24864);
and U27137 (N_27137,N_21150,N_23727);
nand U27138 (N_27138,N_21723,N_23021);
xnor U27139 (N_27139,N_22123,N_20814);
or U27140 (N_27140,N_24950,N_24397);
xnor U27141 (N_27141,N_21194,N_24360);
xor U27142 (N_27142,N_22345,N_20810);
xor U27143 (N_27143,N_24021,N_20541);
xnor U27144 (N_27144,N_24964,N_23151);
xor U27145 (N_27145,N_21376,N_22712);
and U27146 (N_27146,N_21749,N_23620);
nor U27147 (N_27147,N_24046,N_24532);
nor U27148 (N_27148,N_22778,N_20216);
nand U27149 (N_27149,N_21599,N_20385);
and U27150 (N_27150,N_21384,N_24771);
xor U27151 (N_27151,N_23715,N_20438);
nor U27152 (N_27152,N_23176,N_20794);
nand U27153 (N_27153,N_20056,N_20525);
nor U27154 (N_27154,N_24518,N_23328);
and U27155 (N_27155,N_20747,N_24374);
nor U27156 (N_27156,N_23049,N_21691);
nand U27157 (N_27157,N_23635,N_22184);
nor U27158 (N_27158,N_24928,N_23024);
xor U27159 (N_27159,N_21319,N_24677);
and U27160 (N_27160,N_23649,N_23300);
and U27161 (N_27161,N_21969,N_23120);
nor U27162 (N_27162,N_21402,N_20161);
xnor U27163 (N_27163,N_24248,N_23905);
nor U27164 (N_27164,N_21038,N_22927);
and U27165 (N_27165,N_21247,N_23242);
or U27166 (N_27166,N_23893,N_20163);
and U27167 (N_27167,N_22267,N_23506);
and U27168 (N_27168,N_23834,N_22883);
nand U27169 (N_27169,N_23959,N_21292);
and U27170 (N_27170,N_21890,N_24321);
nand U27171 (N_27171,N_23064,N_22376);
nor U27172 (N_27172,N_21215,N_24685);
and U27173 (N_27173,N_20727,N_20082);
or U27174 (N_27174,N_24644,N_20027);
or U27175 (N_27175,N_23484,N_24196);
nor U27176 (N_27176,N_24230,N_24947);
xor U27177 (N_27177,N_21186,N_20837);
and U27178 (N_27178,N_20992,N_24165);
and U27179 (N_27179,N_22172,N_21528);
nor U27180 (N_27180,N_20844,N_24415);
nand U27181 (N_27181,N_23089,N_21300);
and U27182 (N_27182,N_23873,N_22623);
or U27183 (N_27183,N_23263,N_20341);
or U27184 (N_27184,N_24051,N_23358);
nor U27185 (N_27185,N_20754,N_20857);
nand U27186 (N_27186,N_22393,N_20441);
xnor U27187 (N_27187,N_21379,N_21016);
and U27188 (N_27188,N_24847,N_22142);
or U27189 (N_27189,N_22884,N_23213);
or U27190 (N_27190,N_23665,N_23627);
or U27191 (N_27191,N_23324,N_22328);
xor U27192 (N_27192,N_20699,N_20261);
nor U27193 (N_27193,N_23218,N_24580);
and U27194 (N_27194,N_20684,N_23856);
nand U27195 (N_27195,N_21526,N_20128);
nand U27196 (N_27196,N_24913,N_24748);
or U27197 (N_27197,N_20125,N_22288);
nand U27198 (N_27198,N_23920,N_20840);
nand U27199 (N_27199,N_21563,N_23671);
nor U27200 (N_27200,N_24687,N_23896);
nand U27201 (N_27201,N_20482,N_24586);
nand U27202 (N_27202,N_22772,N_23108);
xnor U27203 (N_27203,N_21740,N_22083);
nor U27204 (N_27204,N_24563,N_20759);
or U27205 (N_27205,N_23289,N_20504);
nand U27206 (N_27206,N_23211,N_23683);
nand U27207 (N_27207,N_24537,N_20384);
nand U27208 (N_27208,N_21613,N_24481);
or U27209 (N_27209,N_22191,N_24082);
and U27210 (N_27210,N_24031,N_22925);
and U27211 (N_27211,N_22885,N_20151);
nor U27212 (N_27212,N_23235,N_22912);
nand U27213 (N_27213,N_20966,N_22248);
nor U27214 (N_27214,N_24275,N_24049);
nand U27215 (N_27215,N_21216,N_21099);
and U27216 (N_27216,N_23497,N_23390);
xor U27217 (N_27217,N_20417,N_22346);
nor U27218 (N_27218,N_22604,N_20257);
or U27219 (N_27219,N_23619,N_20841);
xnor U27220 (N_27220,N_24446,N_24436);
nor U27221 (N_27221,N_20474,N_23257);
nand U27222 (N_27222,N_24130,N_23429);
nor U27223 (N_27223,N_24431,N_20451);
nand U27224 (N_27224,N_23091,N_24159);
nor U27225 (N_27225,N_21101,N_21505);
nand U27226 (N_27226,N_20908,N_20335);
or U27227 (N_27227,N_20394,N_24593);
nand U27228 (N_27228,N_23384,N_21598);
or U27229 (N_27229,N_23003,N_20313);
or U27230 (N_27230,N_21111,N_21530);
or U27231 (N_27231,N_21301,N_23851);
or U27232 (N_27232,N_21311,N_23709);
or U27233 (N_27233,N_20218,N_23385);
or U27234 (N_27234,N_20454,N_21794);
and U27235 (N_27235,N_21036,N_21076);
nand U27236 (N_27236,N_23136,N_23233);
nand U27237 (N_27237,N_24746,N_21228);
and U27238 (N_27238,N_22902,N_24459);
nor U27239 (N_27239,N_23313,N_20036);
nor U27240 (N_27240,N_23718,N_20233);
nand U27241 (N_27241,N_20929,N_20119);
or U27242 (N_27242,N_20018,N_22091);
xnor U27243 (N_27243,N_23304,N_24053);
and U27244 (N_27244,N_24968,N_23335);
nor U27245 (N_27245,N_24232,N_23740);
nor U27246 (N_27246,N_22620,N_22168);
nand U27247 (N_27247,N_20248,N_20144);
or U27248 (N_27248,N_20368,N_22700);
or U27249 (N_27249,N_22508,N_24121);
xnor U27250 (N_27250,N_23391,N_20995);
or U27251 (N_27251,N_24200,N_22073);
and U27252 (N_27252,N_22419,N_24353);
xnor U27253 (N_27253,N_23283,N_24363);
or U27254 (N_27254,N_22178,N_20280);
nand U27255 (N_27255,N_21933,N_20198);
xnor U27256 (N_27256,N_21079,N_23179);
or U27257 (N_27257,N_22588,N_21868);
nand U27258 (N_27258,N_20758,N_20122);
and U27259 (N_27259,N_20663,N_20129);
or U27260 (N_27260,N_20987,N_24851);
or U27261 (N_27261,N_20608,N_23137);
nand U27262 (N_27262,N_22821,N_24624);
or U27263 (N_27263,N_23031,N_23785);
nor U27264 (N_27264,N_24975,N_22160);
nand U27265 (N_27265,N_20576,N_21718);
or U27266 (N_27266,N_20492,N_21826);
xor U27267 (N_27267,N_23197,N_24209);
xor U27268 (N_27268,N_23204,N_24285);
or U27269 (N_27269,N_21798,N_23624);
xnor U27270 (N_27270,N_20288,N_21661);
xor U27271 (N_27271,N_23106,N_21109);
or U27272 (N_27272,N_24129,N_24234);
and U27273 (N_27273,N_23997,N_23835);
nand U27274 (N_27274,N_24306,N_22519);
or U27275 (N_27275,N_20776,N_23295);
nand U27276 (N_27276,N_20785,N_22293);
nand U27277 (N_27277,N_21805,N_24517);
xnor U27278 (N_27278,N_22724,N_21352);
xor U27279 (N_27279,N_20897,N_22967);
xor U27280 (N_27280,N_24222,N_20519);
xor U27281 (N_27281,N_21866,N_22764);
nand U27282 (N_27282,N_24277,N_24478);
nor U27283 (N_27283,N_21658,N_24328);
and U27284 (N_27284,N_21484,N_20191);
nor U27285 (N_27285,N_22325,N_22285);
xnor U27286 (N_27286,N_24707,N_24617);
and U27287 (N_27287,N_22844,N_22084);
nor U27288 (N_27288,N_24186,N_23053);
or U27289 (N_27289,N_23717,N_23430);
xor U27290 (N_27290,N_24506,N_24287);
nor U27291 (N_27291,N_24372,N_24043);
nor U27292 (N_27292,N_21191,N_21602);
xnor U27293 (N_27293,N_20907,N_20304);
and U27294 (N_27294,N_23332,N_21197);
nand U27295 (N_27295,N_20731,N_22822);
and U27296 (N_27296,N_24495,N_24961);
xor U27297 (N_27297,N_23622,N_22736);
or U27298 (N_27298,N_21495,N_24124);
or U27299 (N_27299,N_23163,N_24962);
nand U27300 (N_27300,N_20479,N_24791);
nor U27301 (N_27301,N_24294,N_20743);
xor U27302 (N_27302,N_21753,N_21249);
xnor U27303 (N_27303,N_24692,N_21341);
or U27304 (N_27304,N_20230,N_21474);
nand U27305 (N_27305,N_22032,N_21527);
nand U27306 (N_27306,N_23011,N_23578);
and U27307 (N_27307,N_24943,N_22072);
nor U27308 (N_27308,N_21542,N_24145);
xor U27309 (N_27309,N_20572,N_22804);
nand U27310 (N_27310,N_22127,N_22313);
nand U27311 (N_27311,N_23806,N_23210);
nor U27312 (N_27312,N_21556,N_22683);
nand U27313 (N_27313,N_24356,N_24590);
or U27314 (N_27314,N_22253,N_22636);
or U27315 (N_27315,N_24701,N_23746);
xnor U27316 (N_27316,N_20090,N_24304);
xor U27317 (N_27317,N_22614,N_22752);
or U27318 (N_27318,N_24561,N_23792);
and U27319 (N_27319,N_20954,N_23055);
or U27320 (N_27320,N_21136,N_24104);
or U27321 (N_27321,N_20465,N_23694);
nor U27322 (N_27322,N_21752,N_24102);
xor U27323 (N_27323,N_21198,N_24047);
or U27324 (N_27324,N_23278,N_24183);
and U27325 (N_27325,N_24106,N_24054);
nand U27326 (N_27326,N_24665,N_22124);
nand U27327 (N_27327,N_21715,N_21858);
or U27328 (N_27328,N_22389,N_22101);
nand U27329 (N_27329,N_24564,N_21721);
nand U27330 (N_27330,N_22480,N_21605);
nand U27331 (N_27331,N_20745,N_24239);
or U27332 (N_27332,N_22468,N_20127);
and U27333 (N_27333,N_22672,N_20084);
or U27334 (N_27334,N_21622,N_21624);
nor U27335 (N_27335,N_23371,N_21711);
xnor U27336 (N_27336,N_21163,N_24315);
or U27337 (N_27337,N_20498,N_23327);
xnor U27338 (N_27338,N_22318,N_21212);
and U27339 (N_27339,N_23028,N_21972);
nor U27340 (N_27340,N_22064,N_23005);
nand U27341 (N_27341,N_22626,N_24309);
nand U27342 (N_27342,N_22718,N_21681);
or U27343 (N_27343,N_24088,N_24882);
nor U27344 (N_27344,N_20753,N_22036);
nor U27345 (N_27345,N_20976,N_23265);
and U27346 (N_27346,N_22717,N_23234);
and U27347 (N_27347,N_23261,N_24119);
xnor U27348 (N_27348,N_23008,N_22391);
nand U27349 (N_27349,N_21639,N_24666);
nor U27350 (N_27350,N_24418,N_21433);
nor U27351 (N_27351,N_24352,N_20177);
or U27352 (N_27352,N_21488,N_24705);
nor U27353 (N_27353,N_23245,N_23651);
or U27354 (N_27354,N_20254,N_21340);
xor U27355 (N_27355,N_23334,N_21705);
xor U27356 (N_27356,N_20694,N_24158);
nand U27357 (N_27357,N_20164,N_24163);
and U27358 (N_27358,N_21358,N_20358);
and U27359 (N_27359,N_24388,N_20623);
and U27360 (N_27360,N_23695,N_20890);
and U27361 (N_27361,N_24340,N_23109);
or U27362 (N_27362,N_21664,N_22407);
xnor U27363 (N_27363,N_22913,N_24584);
or U27364 (N_27364,N_20582,N_22241);
or U27365 (N_27365,N_24022,N_20967);
xnor U27366 (N_27366,N_22373,N_20928);
and U27367 (N_27367,N_20421,N_23198);
nand U27368 (N_27368,N_20393,N_20320);
nand U27369 (N_27369,N_21097,N_20508);
and U27370 (N_27370,N_22476,N_21156);
xor U27371 (N_27371,N_22921,N_22726);
xnor U27372 (N_27372,N_23930,N_23521);
nand U27373 (N_27373,N_24926,N_24331);
nand U27374 (N_27374,N_22240,N_21656);
nand U27375 (N_27375,N_20314,N_23496);
nor U27376 (N_27376,N_22713,N_21829);
and U27377 (N_27377,N_22159,N_24020);
nor U27378 (N_27378,N_21541,N_23465);
nor U27379 (N_27379,N_20419,N_22075);
xnor U27380 (N_27380,N_20689,N_23522);
and U27381 (N_27381,N_23981,N_23672);
nor U27382 (N_27382,N_21881,N_23247);
and U27383 (N_27383,N_24151,N_22749);
xor U27384 (N_27384,N_20591,N_24547);
xnor U27385 (N_27385,N_23882,N_23122);
xnor U27386 (N_27386,N_22629,N_21130);
nor U27387 (N_27387,N_21847,N_23763);
and U27388 (N_27388,N_22795,N_23939);
nand U27389 (N_27389,N_23754,N_23252);
nand U27390 (N_27390,N_20300,N_20865);
nand U27391 (N_27391,N_21153,N_20172);
nand U27392 (N_27392,N_24056,N_23581);
nand U27393 (N_27393,N_20329,N_24533);
and U27394 (N_27394,N_21786,N_20229);
xor U27395 (N_27395,N_21270,N_23074);
and U27396 (N_27396,N_20452,N_22222);
or U27397 (N_27397,N_22936,N_24999);
nand U27398 (N_27398,N_22600,N_23829);
xor U27399 (N_27399,N_23155,N_20244);
nand U27400 (N_27400,N_24779,N_20821);
nor U27401 (N_27401,N_24274,N_21050);
and U27402 (N_27402,N_23424,N_23381);
xnor U27403 (N_27403,N_21221,N_20548);
or U27404 (N_27404,N_20165,N_24822);
xor U27405 (N_27405,N_24404,N_23352);
xnor U27406 (N_27406,N_20428,N_24219);
xor U27407 (N_27407,N_23367,N_20472);
and U27408 (N_27408,N_22706,N_20905);
xnor U27409 (N_27409,N_24193,N_20968);
or U27410 (N_27410,N_22355,N_21189);
xnor U27411 (N_27411,N_24180,N_24447);
nor U27412 (N_27412,N_21445,N_24310);
nand U27413 (N_27413,N_23152,N_21511);
nand U27414 (N_27414,N_21298,N_23965);
xnor U27415 (N_27415,N_22018,N_23891);
nor U27416 (N_27416,N_20293,N_23276);
xnor U27417 (N_27417,N_20886,N_20379);
nor U27418 (N_27418,N_21367,N_22306);
or U27419 (N_27419,N_22557,N_24057);
or U27420 (N_27420,N_22398,N_22610);
and U27421 (N_27421,N_24920,N_20279);
or U27422 (N_27422,N_21266,N_24992);
nor U27423 (N_27423,N_23461,N_21327);
nor U27424 (N_27424,N_23209,N_22314);
and U27425 (N_27425,N_22026,N_20240);
nand U27426 (N_27426,N_22977,N_23062);
and U27427 (N_27427,N_23780,N_23410);
nand U27428 (N_27428,N_24068,N_24646);
nor U27429 (N_27429,N_20635,N_22404);
nor U27430 (N_27430,N_21693,N_24904);
nor U27431 (N_27431,N_20878,N_24392);
nor U27432 (N_27432,N_22767,N_23175);
nand U27433 (N_27433,N_22635,N_22513);
xnor U27434 (N_27434,N_23057,N_23083);
nand U27435 (N_27435,N_20168,N_21918);
nand U27436 (N_27436,N_24886,N_22372);
nor U27437 (N_27437,N_23254,N_21329);
or U27438 (N_27438,N_20345,N_21733);
or U27439 (N_27439,N_24194,N_20448);
xor U27440 (N_27440,N_21648,N_20516);
and U27441 (N_27441,N_22052,N_22182);
and U27442 (N_27442,N_22851,N_23046);
xor U27443 (N_27443,N_20911,N_21687);
nand U27444 (N_27444,N_23071,N_21901);
nand U27445 (N_27445,N_22771,N_24977);
and U27446 (N_27446,N_20809,N_22062);
xnor U27447 (N_27447,N_21473,N_21841);
nand U27448 (N_27448,N_20848,N_23764);
nor U27449 (N_27449,N_20147,N_22816);
xor U27450 (N_27450,N_20536,N_21534);
xnor U27451 (N_27451,N_21925,N_24569);
nor U27452 (N_27452,N_24351,N_22998);
and U27453 (N_27453,N_23308,N_22596);
and U27454 (N_27454,N_20324,N_23095);
xor U27455 (N_27455,N_24485,N_23529);
and U27456 (N_27456,N_21220,N_24394);
or U27457 (N_27457,N_22353,N_23241);
or U27458 (N_27458,N_24760,N_20267);
nand U27459 (N_27459,N_22674,N_23345);
xor U27460 (N_27460,N_21423,N_22381);
and U27461 (N_27461,N_23407,N_23171);
nor U27462 (N_27462,N_20599,N_22585);
nand U27463 (N_27463,N_21770,N_23508);
nand U27464 (N_27464,N_21907,N_22666);
and U27465 (N_27465,N_20016,N_20940);
or U27466 (N_27466,N_22455,N_21105);
xnor U27467 (N_27467,N_20607,N_24221);
or U27468 (N_27468,N_21388,N_21362);
or U27469 (N_27469,N_24628,N_20030);
nand U27470 (N_27470,N_20132,N_23632);
nand U27471 (N_27471,N_20833,N_20407);
and U27472 (N_27472,N_24838,N_22097);
nor U27473 (N_27473,N_22941,N_20864);
nor U27474 (N_27474,N_20639,N_22466);
and U27475 (N_27475,N_20813,N_20249);
nand U27476 (N_27476,N_23376,N_22048);
and U27477 (N_27477,N_24693,N_21468);
or U27478 (N_27478,N_20564,N_24115);
or U27479 (N_27479,N_23372,N_24673);
nand U27480 (N_27480,N_24504,N_21974);
or U27481 (N_27481,N_22424,N_22213);
nor U27482 (N_27482,N_21284,N_21616);
xor U27483 (N_27483,N_21129,N_24175);
nor U27484 (N_27484,N_23688,N_23509);
xor U27485 (N_27485,N_22125,N_24625);
or U27486 (N_27486,N_23680,N_20723);
nor U27487 (N_27487,N_21072,N_24050);
nor U27488 (N_27488,N_22208,N_21287);
or U27489 (N_27489,N_20893,N_21929);
or U27490 (N_27490,N_22928,N_20962);
or U27491 (N_27491,N_21070,N_23431);
nor U27492 (N_27492,N_24405,N_22958);
xor U27493 (N_27493,N_21593,N_21985);
xor U27494 (N_27494,N_21811,N_23900);
and U27495 (N_27495,N_24583,N_23394);
or U27496 (N_27496,N_22806,N_21905);
and U27497 (N_27497,N_24251,N_21307);
or U27498 (N_27498,N_24572,N_24259);
or U27499 (N_27499,N_22974,N_22942);
nor U27500 (N_27500,N_23095,N_22623);
nor U27501 (N_27501,N_20600,N_20815);
xor U27502 (N_27502,N_21264,N_21546);
nand U27503 (N_27503,N_22088,N_21005);
xnor U27504 (N_27504,N_23314,N_20913);
xor U27505 (N_27505,N_22411,N_23035);
or U27506 (N_27506,N_21816,N_20627);
nor U27507 (N_27507,N_20913,N_22563);
xnor U27508 (N_27508,N_22485,N_22187);
xnor U27509 (N_27509,N_23785,N_24767);
nand U27510 (N_27510,N_22027,N_21004);
nor U27511 (N_27511,N_22201,N_20187);
xor U27512 (N_27512,N_24497,N_21807);
nor U27513 (N_27513,N_21440,N_24717);
nand U27514 (N_27514,N_22516,N_24014);
xnor U27515 (N_27515,N_24632,N_21835);
xnor U27516 (N_27516,N_20616,N_24350);
nand U27517 (N_27517,N_22723,N_22052);
nor U27518 (N_27518,N_20705,N_23670);
and U27519 (N_27519,N_23548,N_24763);
xnor U27520 (N_27520,N_22697,N_24249);
and U27521 (N_27521,N_22379,N_22490);
nor U27522 (N_27522,N_20256,N_23450);
nor U27523 (N_27523,N_24706,N_20499);
xor U27524 (N_27524,N_20814,N_20906);
or U27525 (N_27525,N_20652,N_22038);
nand U27526 (N_27526,N_20994,N_20602);
and U27527 (N_27527,N_24436,N_24435);
and U27528 (N_27528,N_21100,N_22470);
or U27529 (N_27529,N_24281,N_22558);
or U27530 (N_27530,N_23943,N_21621);
nand U27531 (N_27531,N_20697,N_23278);
or U27532 (N_27532,N_23667,N_22733);
xor U27533 (N_27533,N_21168,N_24617);
or U27534 (N_27534,N_20563,N_21709);
nor U27535 (N_27535,N_22401,N_22971);
or U27536 (N_27536,N_20312,N_24394);
nand U27537 (N_27537,N_23871,N_22386);
or U27538 (N_27538,N_24943,N_22144);
xnor U27539 (N_27539,N_20602,N_20273);
nand U27540 (N_27540,N_22790,N_22906);
and U27541 (N_27541,N_22938,N_22198);
xor U27542 (N_27542,N_21087,N_21462);
and U27543 (N_27543,N_22451,N_24572);
nand U27544 (N_27544,N_21119,N_22559);
xor U27545 (N_27545,N_23669,N_20160);
xnor U27546 (N_27546,N_21007,N_20540);
nor U27547 (N_27547,N_22859,N_20655);
nor U27548 (N_27548,N_20760,N_21088);
or U27549 (N_27549,N_21223,N_23629);
xnor U27550 (N_27550,N_22013,N_21573);
nand U27551 (N_27551,N_23404,N_23239);
xnor U27552 (N_27552,N_23696,N_24066);
xor U27553 (N_27553,N_21045,N_23087);
nor U27554 (N_27554,N_22346,N_23376);
or U27555 (N_27555,N_21046,N_21770);
and U27556 (N_27556,N_24417,N_23038);
or U27557 (N_27557,N_22206,N_20765);
and U27558 (N_27558,N_22313,N_24156);
and U27559 (N_27559,N_24997,N_20957);
xnor U27560 (N_27560,N_21987,N_21711);
and U27561 (N_27561,N_21389,N_21773);
nor U27562 (N_27562,N_23429,N_22995);
and U27563 (N_27563,N_21070,N_23258);
nor U27564 (N_27564,N_20721,N_20551);
or U27565 (N_27565,N_23578,N_24277);
nor U27566 (N_27566,N_24239,N_23362);
xor U27567 (N_27567,N_22116,N_21165);
and U27568 (N_27568,N_23367,N_20827);
or U27569 (N_27569,N_20382,N_24954);
and U27570 (N_27570,N_24811,N_23550);
nand U27571 (N_27571,N_24850,N_23385);
nor U27572 (N_27572,N_23596,N_23196);
nor U27573 (N_27573,N_23533,N_24020);
nand U27574 (N_27574,N_21222,N_24898);
nand U27575 (N_27575,N_23244,N_20172);
nor U27576 (N_27576,N_23235,N_24716);
or U27577 (N_27577,N_24683,N_20288);
nor U27578 (N_27578,N_24657,N_24034);
or U27579 (N_27579,N_23192,N_21110);
or U27580 (N_27580,N_20428,N_23512);
nand U27581 (N_27581,N_20246,N_23288);
xor U27582 (N_27582,N_22565,N_22090);
nand U27583 (N_27583,N_21802,N_20610);
or U27584 (N_27584,N_24173,N_24766);
xnor U27585 (N_27585,N_21912,N_22077);
or U27586 (N_27586,N_24060,N_22626);
nand U27587 (N_27587,N_21211,N_21124);
nand U27588 (N_27588,N_23547,N_20527);
nor U27589 (N_27589,N_22841,N_22665);
or U27590 (N_27590,N_24297,N_23014);
xnor U27591 (N_27591,N_20637,N_23730);
nor U27592 (N_27592,N_20322,N_22856);
nand U27593 (N_27593,N_21705,N_21092);
or U27594 (N_27594,N_23808,N_21311);
nand U27595 (N_27595,N_24819,N_22058);
nor U27596 (N_27596,N_23721,N_21475);
xnor U27597 (N_27597,N_20055,N_21395);
or U27598 (N_27598,N_22983,N_20597);
and U27599 (N_27599,N_21253,N_21630);
and U27600 (N_27600,N_21396,N_20465);
xor U27601 (N_27601,N_24786,N_20467);
xor U27602 (N_27602,N_23126,N_23693);
nand U27603 (N_27603,N_23838,N_21661);
and U27604 (N_27604,N_21981,N_23651);
or U27605 (N_27605,N_21770,N_21505);
or U27606 (N_27606,N_22281,N_22895);
or U27607 (N_27607,N_21330,N_21043);
nor U27608 (N_27608,N_22310,N_23133);
nand U27609 (N_27609,N_22223,N_24739);
nor U27610 (N_27610,N_20988,N_21935);
nand U27611 (N_27611,N_20444,N_21377);
nor U27612 (N_27612,N_21317,N_20822);
or U27613 (N_27613,N_20795,N_22440);
xnor U27614 (N_27614,N_24318,N_22090);
or U27615 (N_27615,N_23824,N_23368);
and U27616 (N_27616,N_23714,N_22048);
nand U27617 (N_27617,N_23752,N_20233);
and U27618 (N_27618,N_20309,N_21434);
or U27619 (N_27619,N_21058,N_20166);
or U27620 (N_27620,N_24707,N_21836);
nor U27621 (N_27621,N_24313,N_21636);
xnor U27622 (N_27622,N_21783,N_24723);
xnor U27623 (N_27623,N_23308,N_24815);
xnor U27624 (N_27624,N_23847,N_20128);
or U27625 (N_27625,N_24939,N_22519);
and U27626 (N_27626,N_21408,N_20315);
or U27627 (N_27627,N_21635,N_24341);
nand U27628 (N_27628,N_20758,N_24301);
and U27629 (N_27629,N_21807,N_22925);
nor U27630 (N_27630,N_23338,N_24640);
and U27631 (N_27631,N_23286,N_21878);
xnor U27632 (N_27632,N_22934,N_22881);
xnor U27633 (N_27633,N_21837,N_20697);
and U27634 (N_27634,N_22688,N_22524);
nand U27635 (N_27635,N_22228,N_23307);
nand U27636 (N_27636,N_23003,N_20561);
xnor U27637 (N_27637,N_20754,N_23954);
nand U27638 (N_27638,N_22824,N_20271);
or U27639 (N_27639,N_22994,N_24217);
or U27640 (N_27640,N_20324,N_21032);
xor U27641 (N_27641,N_24828,N_20222);
xor U27642 (N_27642,N_21428,N_22422);
nand U27643 (N_27643,N_23286,N_20544);
or U27644 (N_27644,N_20800,N_24900);
nor U27645 (N_27645,N_21063,N_21335);
xor U27646 (N_27646,N_23007,N_22262);
or U27647 (N_27647,N_22599,N_23954);
or U27648 (N_27648,N_24241,N_22661);
nand U27649 (N_27649,N_24929,N_23645);
nand U27650 (N_27650,N_21946,N_24958);
nand U27651 (N_27651,N_24518,N_23942);
and U27652 (N_27652,N_21140,N_24336);
or U27653 (N_27653,N_21895,N_23625);
nor U27654 (N_27654,N_21039,N_20414);
and U27655 (N_27655,N_20188,N_24771);
nor U27656 (N_27656,N_21235,N_21233);
nand U27657 (N_27657,N_21487,N_22377);
xnor U27658 (N_27658,N_23100,N_23414);
nor U27659 (N_27659,N_23366,N_24449);
xor U27660 (N_27660,N_20067,N_22634);
xnor U27661 (N_27661,N_23190,N_22204);
nor U27662 (N_27662,N_21551,N_23163);
and U27663 (N_27663,N_23034,N_24473);
and U27664 (N_27664,N_21340,N_22354);
nand U27665 (N_27665,N_23622,N_24323);
nor U27666 (N_27666,N_21888,N_23510);
or U27667 (N_27667,N_20346,N_22261);
nor U27668 (N_27668,N_23340,N_23116);
nand U27669 (N_27669,N_22068,N_21421);
nor U27670 (N_27670,N_23455,N_20151);
nand U27671 (N_27671,N_20739,N_21698);
and U27672 (N_27672,N_21230,N_24906);
nor U27673 (N_27673,N_22841,N_24877);
xnor U27674 (N_27674,N_23183,N_23795);
and U27675 (N_27675,N_21050,N_23398);
nand U27676 (N_27676,N_21101,N_23780);
xor U27677 (N_27677,N_22596,N_20301);
nand U27678 (N_27678,N_20428,N_20124);
and U27679 (N_27679,N_21177,N_22333);
nand U27680 (N_27680,N_24041,N_22377);
xor U27681 (N_27681,N_24791,N_21722);
nor U27682 (N_27682,N_22922,N_21065);
nor U27683 (N_27683,N_23461,N_20209);
and U27684 (N_27684,N_23285,N_23849);
and U27685 (N_27685,N_22887,N_20202);
nand U27686 (N_27686,N_20457,N_23858);
or U27687 (N_27687,N_22476,N_21414);
and U27688 (N_27688,N_21306,N_22674);
nor U27689 (N_27689,N_21398,N_20102);
nor U27690 (N_27690,N_22581,N_24377);
and U27691 (N_27691,N_23097,N_22677);
xor U27692 (N_27692,N_22226,N_22919);
or U27693 (N_27693,N_24440,N_24651);
nand U27694 (N_27694,N_23561,N_23210);
and U27695 (N_27695,N_22756,N_20050);
and U27696 (N_27696,N_21681,N_23523);
xnor U27697 (N_27697,N_23957,N_20434);
xnor U27698 (N_27698,N_23061,N_22793);
nor U27699 (N_27699,N_23126,N_21725);
or U27700 (N_27700,N_20796,N_21674);
nand U27701 (N_27701,N_24981,N_20387);
nor U27702 (N_27702,N_21069,N_22543);
and U27703 (N_27703,N_22456,N_20361);
nand U27704 (N_27704,N_21540,N_23317);
xor U27705 (N_27705,N_23350,N_21375);
and U27706 (N_27706,N_23736,N_21407);
and U27707 (N_27707,N_23776,N_22499);
nand U27708 (N_27708,N_23325,N_23034);
nand U27709 (N_27709,N_23425,N_21912);
or U27710 (N_27710,N_21652,N_23801);
and U27711 (N_27711,N_21912,N_24507);
nand U27712 (N_27712,N_22952,N_24380);
xnor U27713 (N_27713,N_20885,N_21274);
nor U27714 (N_27714,N_20202,N_22625);
and U27715 (N_27715,N_21988,N_21648);
xnor U27716 (N_27716,N_20715,N_20169);
or U27717 (N_27717,N_24713,N_21750);
nor U27718 (N_27718,N_22168,N_23547);
and U27719 (N_27719,N_22545,N_24959);
or U27720 (N_27720,N_24684,N_20664);
nor U27721 (N_27721,N_23045,N_22596);
or U27722 (N_27722,N_21571,N_22066);
or U27723 (N_27723,N_21932,N_22863);
xnor U27724 (N_27724,N_21601,N_22494);
xnor U27725 (N_27725,N_24749,N_23893);
xor U27726 (N_27726,N_20259,N_24641);
and U27727 (N_27727,N_24262,N_21236);
nor U27728 (N_27728,N_24946,N_24757);
nand U27729 (N_27729,N_22874,N_21381);
xor U27730 (N_27730,N_23746,N_24743);
nand U27731 (N_27731,N_21998,N_22940);
nand U27732 (N_27732,N_22560,N_22043);
nand U27733 (N_27733,N_23196,N_22124);
and U27734 (N_27734,N_21262,N_22207);
xor U27735 (N_27735,N_23182,N_23481);
or U27736 (N_27736,N_20450,N_21157);
or U27737 (N_27737,N_23565,N_21227);
nor U27738 (N_27738,N_20408,N_21478);
and U27739 (N_27739,N_24760,N_21869);
and U27740 (N_27740,N_24489,N_24911);
xor U27741 (N_27741,N_20921,N_23508);
or U27742 (N_27742,N_23718,N_24722);
xor U27743 (N_27743,N_22114,N_21397);
nor U27744 (N_27744,N_21880,N_24724);
and U27745 (N_27745,N_24067,N_22031);
nor U27746 (N_27746,N_23447,N_23819);
nand U27747 (N_27747,N_22342,N_23997);
nor U27748 (N_27748,N_20744,N_24202);
xnor U27749 (N_27749,N_22474,N_21034);
xor U27750 (N_27750,N_22347,N_22722);
or U27751 (N_27751,N_21375,N_23949);
nand U27752 (N_27752,N_20402,N_22057);
nand U27753 (N_27753,N_21689,N_24332);
nor U27754 (N_27754,N_20513,N_24906);
nor U27755 (N_27755,N_21965,N_22715);
nor U27756 (N_27756,N_21086,N_20932);
or U27757 (N_27757,N_23432,N_21859);
nor U27758 (N_27758,N_21976,N_20586);
and U27759 (N_27759,N_20479,N_22343);
xnor U27760 (N_27760,N_24342,N_20547);
and U27761 (N_27761,N_21113,N_20947);
nor U27762 (N_27762,N_21490,N_20886);
and U27763 (N_27763,N_21589,N_22224);
or U27764 (N_27764,N_23005,N_22845);
nor U27765 (N_27765,N_21238,N_24234);
or U27766 (N_27766,N_21638,N_23599);
or U27767 (N_27767,N_22855,N_21227);
nor U27768 (N_27768,N_21989,N_24195);
nand U27769 (N_27769,N_23285,N_20793);
nor U27770 (N_27770,N_21501,N_24513);
or U27771 (N_27771,N_21783,N_21734);
nand U27772 (N_27772,N_22982,N_24182);
and U27773 (N_27773,N_24692,N_20842);
nor U27774 (N_27774,N_24998,N_23220);
xor U27775 (N_27775,N_20310,N_21305);
or U27776 (N_27776,N_20962,N_24226);
and U27777 (N_27777,N_24623,N_24778);
nor U27778 (N_27778,N_24904,N_21733);
and U27779 (N_27779,N_22321,N_21562);
or U27780 (N_27780,N_22783,N_21929);
nand U27781 (N_27781,N_22735,N_24627);
xor U27782 (N_27782,N_22465,N_22998);
nor U27783 (N_27783,N_20016,N_23514);
nor U27784 (N_27784,N_21074,N_22134);
and U27785 (N_27785,N_22447,N_21677);
or U27786 (N_27786,N_22198,N_22565);
and U27787 (N_27787,N_24715,N_23637);
or U27788 (N_27788,N_24835,N_23398);
and U27789 (N_27789,N_24395,N_21411);
nor U27790 (N_27790,N_23115,N_20135);
and U27791 (N_27791,N_20749,N_22120);
or U27792 (N_27792,N_20008,N_22513);
nor U27793 (N_27793,N_23840,N_20486);
nand U27794 (N_27794,N_21481,N_22667);
or U27795 (N_27795,N_21374,N_24480);
and U27796 (N_27796,N_23006,N_23276);
and U27797 (N_27797,N_21142,N_21482);
xor U27798 (N_27798,N_22284,N_20973);
and U27799 (N_27799,N_21207,N_20900);
nor U27800 (N_27800,N_22539,N_24236);
or U27801 (N_27801,N_21465,N_23400);
or U27802 (N_27802,N_24996,N_22867);
and U27803 (N_27803,N_24708,N_22671);
nor U27804 (N_27804,N_23282,N_23640);
and U27805 (N_27805,N_22511,N_20662);
nand U27806 (N_27806,N_21853,N_21521);
nand U27807 (N_27807,N_20068,N_22916);
or U27808 (N_27808,N_21867,N_21918);
nor U27809 (N_27809,N_24706,N_23017);
and U27810 (N_27810,N_22162,N_20350);
and U27811 (N_27811,N_23056,N_24789);
and U27812 (N_27812,N_21482,N_23257);
nand U27813 (N_27813,N_21081,N_22008);
and U27814 (N_27814,N_23241,N_24326);
xnor U27815 (N_27815,N_24027,N_20874);
and U27816 (N_27816,N_23003,N_21849);
and U27817 (N_27817,N_20135,N_24311);
nor U27818 (N_27818,N_21097,N_24066);
or U27819 (N_27819,N_23017,N_22256);
or U27820 (N_27820,N_20560,N_24660);
or U27821 (N_27821,N_20286,N_20692);
xnor U27822 (N_27822,N_20938,N_22632);
xnor U27823 (N_27823,N_23897,N_22544);
or U27824 (N_27824,N_24925,N_24598);
nand U27825 (N_27825,N_21441,N_23452);
nor U27826 (N_27826,N_20614,N_21829);
and U27827 (N_27827,N_24273,N_24068);
or U27828 (N_27828,N_24238,N_24012);
nand U27829 (N_27829,N_21010,N_22432);
nand U27830 (N_27830,N_24213,N_22964);
and U27831 (N_27831,N_21894,N_21305);
xnor U27832 (N_27832,N_21838,N_24727);
or U27833 (N_27833,N_20160,N_21866);
nand U27834 (N_27834,N_21613,N_24315);
xnor U27835 (N_27835,N_20891,N_21952);
nand U27836 (N_27836,N_20246,N_23445);
xnor U27837 (N_27837,N_20817,N_20548);
nand U27838 (N_27838,N_22334,N_20498);
xor U27839 (N_27839,N_22336,N_21791);
or U27840 (N_27840,N_21601,N_22060);
xor U27841 (N_27841,N_23851,N_22698);
or U27842 (N_27842,N_24927,N_23637);
nand U27843 (N_27843,N_23116,N_21109);
nor U27844 (N_27844,N_22831,N_23329);
xor U27845 (N_27845,N_21366,N_21739);
or U27846 (N_27846,N_23775,N_21170);
and U27847 (N_27847,N_22734,N_24377);
xor U27848 (N_27848,N_21945,N_24474);
nand U27849 (N_27849,N_24889,N_21245);
xor U27850 (N_27850,N_23440,N_22220);
xnor U27851 (N_27851,N_24222,N_20825);
and U27852 (N_27852,N_24166,N_20180);
nand U27853 (N_27853,N_23258,N_22886);
or U27854 (N_27854,N_24480,N_24886);
and U27855 (N_27855,N_22508,N_20726);
xnor U27856 (N_27856,N_21604,N_24978);
nor U27857 (N_27857,N_20330,N_23465);
nor U27858 (N_27858,N_23292,N_22649);
xnor U27859 (N_27859,N_21390,N_20896);
and U27860 (N_27860,N_20824,N_20745);
nand U27861 (N_27861,N_22496,N_22179);
xor U27862 (N_27862,N_20229,N_23025);
nor U27863 (N_27863,N_22713,N_20396);
or U27864 (N_27864,N_21877,N_20719);
nand U27865 (N_27865,N_21905,N_21197);
nor U27866 (N_27866,N_22751,N_23840);
nand U27867 (N_27867,N_22497,N_22784);
or U27868 (N_27868,N_22876,N_23322);
nor U27869 (N_27869,N_23445,N_20346);
xnor U27870 (N_27870,N_20144,N_20138);
xnor U27871 (N_27871,N_23035,N_23010);
xor U27872 (N_27872,N_24573,N_20510);
nand U27873 (N_27873,N_21780,N_22891);
xor U27874 (N_27874,N_22053,N_24387);
and U27875 (N_27875,N_22231,N_22503);
and U27876 (N_27876,N_24680,N_22737);
nand U27877 (N_27877,N_24419,N_24694);
nand U27878 (N_27878,N_20050,N_22839);
nor U27879 (N_27879,N_22700,N_24947);
nand U27880 (N_27880,N_24754,N_21797);
or U27881 (N_27881,N_21903,N_23756);
xor U27882 (N_27882,N_23984,N_22752);
or U27883 (N_27883,N_24242,N_24280);
nor U27884 (N_27884,N_23845,N_23157);
xnor U27885 (N_27885,N_20057,N_24920);
and U27886 (N_27886,N_20011,N_21179);
or U27887 (N_27887,N_23096,N_21208);
and U27888 (N_27888,N_22507,N_23393);
or U27889 (N_27889,N_23192,N_23275);
xor U27890 (N_27890,N_21471,N_21681);
and U27891 (N_27891,N_24081,N_23563);
or U27892 (N_27892,N_21506,N_22994);
nand U27893 (N_27893,N_20736,N_20517);
or U27894 (N_27894,N_24410,N_20956);
and U27895 (N_27895,N_23644,N_24541);
nand U27896 (N_27896,N_21904,N_21549);
nand U27897 (N_27897,N_21468,N_24908);
nand U27898 (N_27898,N_24711,N_20874);
xnor U27899 (N_27899,N_21421,N_20036);
nand U27900 (N_27900,N_23730,N_21709);
or U27901 (N_27901,N_24077,N_21204);
nor U27902 (N_27902,N_24057,N_23746);
nor U27903 (N_27903,N_20821,N_22363);
nand U27904 (N_27904,N_23009,N_24142);
and U27905 (N_27905,N_23776,N_20045);
xnor U27906 (N_27906,N_24602,N_23624);
or U27907 (N_27907,N_20393,N_21014);
and U27908 (N_27908,N_22146,N_23782);
and U27909 (N_27909,N_21312,N_22584);
or U27910 (N_27910,N_20388,N_23220);
and U27911 (N_27911,N_20065,N_24786);
nor U27912 (N_27912,N_22061,N_24041);
and U27913 (N_27913,N_20248,N_21843);
nor U27914 (N_27914,N_23695,N_22973);
nand U27915 (N_27915,N_22873,N_24037);
xor U27916 (N_27916,N_23835,N_20031);
or U27917 (N_27917,N_20695,N_20304);
and U27918 (N_27918,N_24448,N_23655);
nor U27919 (N_27919,N_20158,N_24211);
nand U27920 (N_27920,N_23368,N_21477);
or U27921 (N_27921,N_20238,N_23437);
nor U27922 (N_27922,N_20922,N_20756);
nand U27923 (N_27923,N_24291,N_24837);
or U27924 (N_27924,N_22754,N_21942);
nor U27925 (N_27925,N_22731,N_24694);
nor U27926 (N_27926,N_21240,N_24749);
or U27927 (N_27927,N_20802,N_22930);
or U27928 (N_27928,N_24102,N_23220);
nor U27929 (N_27929,N_24881,N_24386);
nand U27930 (N_27930,N_22362,N_24583);
xor U27931 (N_27931,N_22419,N_24751);
nand U27932 (N_27932,N_20750,N_21892);
nor U27933 (N_27933,N_22726,N_23233);
or U27934 (N_27934,N_22352,N_21033);
xor U27935 (N_27935,N_23929,N_22498);
and U27936 (N_27936,N_21616,N_20213);
nand U27937 (N_27937,N_20558,N_21848);
xnor U27938 (N_27938,N_21857,N_24162);
or U27939 (N_27939,N_21941,N_20663);
xnor U27940 (N_27940,N_24081,N_20598);
and U27941 (N_27941,N_20021,N_24037);
nor U27942 (N_27942,N_23398,N_20760);
and U27943 (N_27943,N_23543,N_24957);
nand U27944 (N_27944,N_21224,N_21872);
and U27945 (N_27945,N_23181,N_24040);
or U27946 (N_27946,N_24893,N_24484);
and U27947 (N_27947,N_21506,N_23835);
nor U27948 (N_27948,N_23491,N_21616);
or U27949 (N_27949,N_21462,N_23832);
and U27950 (N_27950,N_22143,N_23816);
nor U27951 (N_27951,N_20197,N_23540);
nor U27952 (N_27952,N_21867,N_21007);
and U27953 (N_27953,N_20789,N_23210);
or U27954 (N_27954,N_20421,N_24277);
nand U27955 (N_27955,N_24991,N_20949);
xor U27956 (N_27956,N_23820,N_22742);
nand U27957 (N_27957,N_24442,N_23374);
nor U27958 (N_27958,N_22116,N_22439);
or U27959 (N_27959,N_20869,N_22789);
xnor U27960 (N_27960,N_22213,N_20762);
nand U27961 (N_27961,N_21661,N_21159);
nand U27962 (N_27962,N_23053,N_23189);
nor U27963 (N_27963,N_22363,N_20259);
or U27964 (N_27964,N_24137,N_20348);
nor U27965 (N_27965,N_22220,N_20247);
nand U27966 (N_27966,N_23381,N_24701);
or U27967 (N_27967,N_24929,N_24774);
and U27968 (N_27968,N_24650,N_24460);
or U27969 (N_27969,N_23094,N_23447);
or U27970 (N_27970,N_22598,N_22231);
or U27971 (N_27971,N_23973,N_24660);
or U27972 (N_27972,N_23912,N_23676);
nand U27973 (N_27973,N_24633,N_21644);
nand U27974 (N_27974,N_20244,N_23817);
and U27975 (N_27975,N_24659,N_22237);
nand U27976 (N_27976,N_23191,N_21719);
nor U27977 (N_27977,N_23870,N_24000);
xnor U27978 (N_27978,N_24017,N_21677);
nand U27979 (N_27979,N_20695,N_22871);
nand U27980 (N_27980,N_20618,N_23708);
xnor U27981 (N_27981,N_21575,N_24133);
nor U27982 (N_27982,N_20742,N_23754);
xor U27983 (N_27983,N_21808,N_21970);
nor U27984 (N_27984,N_23504,N_23997);
nand U27985 (N_27985,N_21791,N_23293);
xor U27986 (N_27986,N_21736,N_23140);
xnor U27987 (N_27987,N_21793,N_21142);
nand U27988 (N_27988,N_22958,N_22760);
xor U27989 (N_27989,N_20403,N_22659);
xor U27990 (N_27990,N_23173,N_24753);
nor U27991 (N_27991,N_23366,N_23418);
nand U27992 (N_27992,N_22495,N_23871);
xor U27993 (N_27993,N_23815,N_23622);
or U27994 (N_27994,N_24743,N_23908);
or U27995 (N_27995,N_21483,N_24165);
xor U27996 (N_27996,N_22082,N_24783);
nor U27997 (N_27997,N_24517,N_20020);
and U27998 (N_27998,N_20797,N_22406);
nor U27999 (N_27999,N_20682,N_20811);
xnor U28000 (N_28000,N_21984,N_24678);
nor U28001 (N_28001,N_21610,N_20971);
nand U28002 (N_28002,N_22358,N_21870);
and U28003 (N_28003,N_22189,N_21794);
xnor U28004 (N_28004,N_24779,N_23225);
xnor U28005 (N_28005,N_24233,N_22862);
nand U28006 (N_28006,N_22629,N_21002);
or U28007 (N_28007,N_22670,N_22409);
nand U28008 (N_28008,N_21363,N_20263);
or U28009 (N_28009,N_20014,N_23152);
nand U28010 (N_28010,N_23940,N_23056);
or U28011 (N_28011,N_23945,N_21380);
and U28012 (N_28012,N_20379,N_23966);
nor U28013 (N_28013,N_22731,N_22150);
nand U28014 (N_28014,N_23363,N_21644);
nand U28015 (N_28015,N_23919,N_23471);
xnor U28016 (N_28016,N_20235,N_20715);
nor U28017 (N_28017,N_21153,N_20153);
and U28018 (N_28018,N_23539,N_23215);
xor U28019 (N_28019,N_20722,N_23897);
nor U28020 (N_28020,N_24822,N_24622);
nand U28021 (N_28021,N_22549,N_20801);
and U28022 (N_28022,N_20609,N_20668);
or U28023 (N_28023,N_23727,N_21294);
and U28024 (N_28024,N_23909,N_20081);
or U28025 (N_28025,N_20387,N_21841);
nand U28026 (N_28026,N_22368,N_21635);
and U28027 (N_28027,N_22434,N_23832);
or U28028 (N_28028,N_21453,N_21903);
nor U28029 (N_28029,N_20853,N_23316);
or U28030 (N_28030,N_21285,N_24588);
xor U28031 (N_28031,N_20151,N_21760);
nand U28032 (N_28032,N_21556,N_20808);
xor U28033 (N_28033,N_24436,N_23058);
nor U28034 (N_28034,N_21207,N_24715);
and U28035 (N_28035,N_20566,N_24832);
nand U28036 (N_28036,N_22532,N_20660);
and U28037 (N_28037,N_20438,N_24255);
nor U28038 (N_28038,N_20501,N_20204);
xnor U28039 (N_28039,N_21309,N_21351);
xor U28040 (N_28040,N_22268,N_24650);
xor U28041 (N_28041,N_23149,N_21672);
or U28042 (N_28042,N_23219,N_23145);
and U28043 (N_28043,N_24605,N_24042);
and U28044 (N_28044,N_22871,N_21268);
or U28045 (N_28045,N_22175,N_22711);
or U28046 (N_28046,N_21501,N_21332);
xnor U28047 (N_28047,N_23815,N_20093);
or U28048 (N_28048,N_23022,N_21614);
or U28049 (N_28049,N_20368,N_21468);
and U28050 (N_28050,N_23420,N_22008);
and U28051 (N_28051,N_22337,N_22225);
xor U28052 (N_28052,N_23591,N_22567);
and U28053 (N_28053,N_22830,N_20563);
nand U28054 (N_28054,N_24751,N_22258);
nand U28055 (N_28055,N_20309,N_24323);
or U28056 (N_28056,N_24435,N_22677);
and U28057 (N_28057,N_21333,N_24006);
nor U28058 (N_28058,N_21697,N_20606);
and U28059 (N_28059,N_20184,N_22495);
and U28060 (N_28060,N_24008,N_22089);
or U28061 (N_28061,N_20672,N_20789);
nor U28062 (N_28062,N_23354,N_23819);
xnor U28063 (N_28063,N_22492,N_22583);
or U28064 (N_28064,N_24842,N_22160);
xor U28065 (N_28065,N_20604,N_20333);
nand U28066 (N_28066,N_22839,N_20764);
nor U28067 (N_28067,N_22048,N_23491);
xnor U28068 (N_28068,N_21548,N_24097);
nand U28069 (N_28069,N_21486,N_21983);
and U28070 (N_28070,N_22705,N_24321);
xnor U28071 (N_28071,N_22558,N_21674);
and U28072 (N_28072,N_24016,N_21774);
or U28073 (N_28073,N_21237,N_24157);
and U28074 (N_28074,N_23990,N_20501);
nor U28075 (N_28075,N_22819,N_20510);
and U28076 (N_28076,N_21564,N_22594);
and U28077 (N_28077,N_22085,N_24840);
nand U28078 (N_28078,N_22305,N_22461);
nor U28079 (N_28079,N_21899,N_24030);
or U28080 (N_28080,N_22914,N_20891);
xnor U28081 (N_28081,N_21650,N_24625);
and U28082 (N_28082,N_24876,N_24019);
nand U28083 (N_28083,N_23819,N_21742);
nor U28084 (N_28084,N_24347,N_23159);
nor U28085 (N_28085,N_22032,N_24573);
nand U28086 (N_28086,N_22603,N_24279);
xor U28087 (N_28087,N_20937,N_24276);
xor U28088 (N_28088,N_23577,N_24225);
or U28089 (N_28089,N_22674,N_22183);
and U28090 (N_28090,N_23074,N_23586);
xor U28091 (N_28091,N_20597,N_22098);
nor U28092 (N_28092,N_20126,N_22761);
nand U28093 (N_28093,N_24644,N_21214);
nor U28094 (N_28094,N_20839,N_23504);
nand U28095 (N_28095,N_20689,N_24416);
or U28096 (N_28096,N_23218,N_22674);
and U28097 (N_28097,N_23958,N_20537);
nor U28098 (N_28098,N_20007,N_20462);
or U28099 (N_28099,N_22879,N_23140);
and U28100 (N_28100,N_22742,N_24549);
xnor U28101 (N_28101,N_24296,N_21233);
or U28102 (N_28102,N_24359,N_23758);
or U28103 (N_28103,N_22132,N_24431);
nand U28104 (N_28104,N_21325,N_23915);
nor U28105 (N_28105,N_23618,N_22143);
nor U28106 (N_28106,N_24665,N_21078);
xnor U28107 (N_28107,N_20988,N_22292);
nand U28108 (N_28108,N_24060,N_22479);
xnor U28109 (N_28109,N_20265,N_23841);
or U28110 (N_28110,N_24231,N_21102);
nand U28111 (N_28111,N_22981,N_21778);
nor U28112 (N_28112,N_24965,N_22720);
nand U28113 (N_28113,N_23210,N_21668);
xnor U28114 (N_28114,N_20210,N_22021);
or U28115 (N_28115,N_20584,N_22799);
and U28116 (N_28116,N_20710,N_20038);
xor U28117 (N_28117,N_24737,N_20658);
and U28118 (N_28118,N_23011,N_24042);
nor U28119 (N_28119,N_21550,N_20732);
or U28120 (N_28120,N_23068,N_24719);
or U28121 (N_28121,N_21676,N_21332);
nand U28122 (N_28122,N_24583,N_24142);
nor U28123 (N_28123,N_21349,N_23044);
xor U28124 (N_28124,N_23156,N_23773);
xnor U28125 (N_28125,N_21735,N_24837);
or U28126 (N_28126,N_21929,N_21941);
xnor U28127 (N_28127,N_21096,N_23329);
xor U28128 (N_28128,N_23342,N_22955);
xnor U28129 (N_28129,N_20174,N_22113);
nor U28130 (N_28130,N_21537,N_24566);
nand U28131 (N_28131,N_24104,N_23810);
xor U28132 (N_28132,N_22443,N_23300);
xor U28133 (N_28133,N_23743,N_22766);
nor U28134 (N_28134,N_20035,N_21403);
and U28135 (N_28135,N_20368,N_20247);
and U28136 (N_28136,N_20246,N_24272);
and U28137 (N_28137,N_24222,N_21943);
xor U28138 (N_28138,N_24119,N_21952);
xor U28139 (N_28139,N_24263,N_24048);
xnor U28140 (N_28140,N_20743,N_21634);
and U28141 (N_28141,N_22632,N_21623);
and U28142 (N_28142,N_21846,N_21521);
or U28143 (N_28143,N_23234,N_20637);
nor U28144 (N_28144,N_24330,N_20157);
and U28145 (N_28145,N_23411,N_24601);
nand U28146 (N_28146,N_22408,N_21849);
nor U28147 (N_28147,N_22719,N_24943);
and U28148 (N_28148,N_23634,N_22124);
nor U28149 (N_28149,N_22481,N_23524);
xnor U28150 (N_28150,N_22115,N_20673);
xor U28151 (N_28151,N_23921,N_24903);
and U28152 (N_28152,N_22619,N_23576);
and U28153 (N_28153,N_20749,N_22056);
nor U28154 (N_28154,N_23122,N_23355);
and U28155 (N_28155,N_20519,N_21871);
or U28156 (N_28156,N_23766,N_24988);
nand U28157 (N_28157,N_20720,N_23557);
or U28158 (N_28158,N_21811,N_23876);
nor U28159 (N_28159,N_22083,N_24700);
nand U28160 (N_28160,N_24955,N_23380);
nand U28161 (N_28161,N_22996,N_23572);
nor U28162 (N_28162,N_24355,N_24771);
nand U28163 (N_28163,N_21952,N_23953);
nand U28164 (N_28164,N_20861,N_21035);
and U28165 (N_28165,N_22204,N_23923);
or U28166 (N_28166,N_21828,N_20168);
xor U28167 (N_28167,N_21344,N_22095);
nand U28168 (N_28168,N_22318,N_22216);
or U28169 (N_28169,N_22233,N_24082);
xor U28170 (N_28170,N_24695,N_22714);
and U28171 (N_28171,N_23320,N_23578);
xor U28172 (N_28172,N_24800,N_22114);
xnor U28173 (N_28173,N_23794,N_22744);
and U28174 (N_28174,N_20937,N_20516);
xnor U28175 (N_28175,N_24134,N_24550);
xor U28176 (N_28176,N_20194,N_20184);
nand U28177 (N_28177,N_20609,N_23630);
nor U28178 (N_28178,N_20192,N_22950);
nand U28179 (N_28179,N_21089,N_20728);
and U28180 (N_28180,N_22089,N_20291);
nor U28181 (N_28181,N_22954,N_20143);
nand U28182 (N_28182,N_22377,N_22992);
xor U28183 (N_28183,N_20743,N_21151);
and U28184 (N_28184,N_21993,N_20621);
nor U28185 (N_28185,N_24651,N_23225);
nand U28186 (N_28186,N_21231,N_22863);
nand U28187 (N_28187,N_22981,N_24347);
nand U28188 (N_28188,N_21081,N_20168);
and U28189 (N_28189,N_24060,N_24665);
xnor U28190 (N_28190,N_22243,N_21915);
and U28191 (N_28191,N_20644,N_24186);
nand U28192 (N_28192,N_22382,N_20993);
nor U28193 (N_28193,N_22205,N_24041);
and U28194 (N_28194,N_21687,N_23703);
xnor U28195 (N_28195,N_20757,N_24244);
nand U28196 (N_28196,N_23119,N_22325);
nor U28197 (N_28197,N_23740,N_20076);
xnor U28198 (N_28198,N_20645,N_22606);
nand U28199 (N_28199,N_23329,N_22536);
or U28200 (N_28200,N_21905,N_23854);
xor U28201 (N_28201,N_21753,N_23468);
xor U28202 (N_28202,N_22152,N_23219);
and U28203 (N_28203,N_21200,N_22095);
xnor U28204 (N_28204,N_20060,N_20507);
or U28205 (N_28205,N_20543,N_20415);
or U28206 (N_28206,N_24699,N_21655);
and U28207 (N_28207,N_23633,N_21513);
and U28208 (N_28208,N_20172,N_24119);
and U28209 (N_28209,N_22042,N_22397);
nand U28210 (N_28210,N_21800,N_21708);
and U28211 (N_28211,N_21349,N_23423);
and U28212 (N_28212,N_21814,N_24078);
or U28213 (N_28213,N_23708,N_24060);
and U28214 (N_28214,N_24223,N_21409);
and U28215 (N_28215,N_21270,N_24114);
nand U28216 (N_28216,N_21141,N_24800);
xnor U28217 (N_28217,N_21617,N_23516);
xor U28218 (N_28218,N_22548,N_20980);
nor U28219 (N_28219,N_22472,N_23348);
nor U28220 (N_28220,N_24731,N_24605);
nor U28221 (N_28221,N_23472,N_23791);
xor U28222 (N_28222,N_20528,N_21240);
and U28223 (N_28223,N_21645,N_24716);
and U28224 (N_28224,N_24807,N_24858);
nand U28225 (N_28225,N_20635,N_20712);
nand U28226 (N_28226,N_23748,N_22935);
xor U28227 (N_28227,N_23656,N_20336);
nand U28228 (N_28228,N_24286,N_21432);
nand U28229 (N_28229,N_23717,N_20818);
and U28230 (N_28230,N_24328,N_24249);
or U28231 (N_28231,N_24510,N_22645);
nand U28232 (N_28232,N_22467,N_23128);
or U28233 (N_28233,N_22013,N_20988);
xor U28234 (N_28234,N_24454,N_20360);
nor U28235 (N_28235,N_23567,N_21577);
nor U28236 (N_28236,N_23055,N_21371);
nand U28237 (N_28237,N_20857,N_22368);
nand U28238 (N_28238,N_21528,N_21514);
nor U28239 (N_28239,N_23870,N_24617);
xnor U28240 (N_28240,N_20056,N_21380);
nand U28241 (N_28241,N_24957,N_20247);
and U28242 (N_28242,N_21454,N_20986);
nor U28243 (N_28243,N_21073,N_21635);
or U28244 (N_28244,N_24669,N_20272);
nor U28245 (N_28245,N_23658,N_24338);
xor U28246 (N_28246,N_21383,N_20290);
and U28247 (N_28247,N_21970,N_24486);
or U28248 (N_28248,N_22331,N_22495);
nand U28249 (N_28249,N_21411,N_23090);
nand U28250 (N_28250,N_23957,N_21345);
or U28251 (N_28251,N_24715,N_24790);
nand U28252 (N_28252,N_23583,N_21839);
xnor U28253 (N_28253,N_24646,N_23459);
nand U28254 (N_28254,N_22348,N_20827);
nand U28255 (N_28255,N_22684,N_21927);
nand U28256 (N_28256,N_23924,N_23304);
or U28257 (N_28257,N_20168,N_22046);
nor U28258 (N_28258,N_22864,N_21474);
or U28259 (N_28259,N_20480,N_21047);
and U28260 (N_28260,N_20618,N_24922);
and U28261 (N_28261,N_20779,N_20040);
nor U28262 (N_28262,N_22897,N_20669);
nor U28263 (N_28263,N_21173,N_20404);
or U28264 (N_28264,N_22199,N_24134);
nor U28265 (N_28265,N_24167,N_22681);
xnor U28266 (N_28266,N_24807,N_23458);
and U28267 (N_28267,N_20017,N_24176);
xnor U28268 (N_28268,N_21035,N_20931);
nor U28269 (N_28269,N_24325,N_23932);
or U28270 (N_28270,N_21461,N_23311);
or U28271 (N_28271,N_24087,N_21960);
xnor U28272 (N_28272,N_24618,N_24541);
or U28273 (N_28273,N_23497,N_20049);
nand U28274 (N_28274,N_22194,N_21269);
nor U28275 (N_28275,N_23720,N_21591);
or U28276 (N_28276,N_23872,N_23981);
and U28277 (N_28277,N_22092,N_21990);
and U28278 (N_28278,N_24360,N_20727);
and U28279 (N_28279,N_20703,N_22698);
xnor U28280 (N_28280,N_24354,N_23039);
nor U28281 (N_28281,N_22447,N_22161);
and U28282 (N_28282,N_22395,N_23633);
and U28283 (N_28283,N_23879,N_20759);
xnor U28284 (N_28284,N_21765,N_20645);
nand U28285 (N_28285,N_21879,N_23654);
nand U28286 (N_28286,N_24345,N_20157);
nor U28287 (N_28287,N_22411,N_24572);
xnor U28288 (N_28288,N_20275,N_21831);
xnor U28289 (N_28289,N_20293,N_22418);
or U28290 (N_28290,N_24049,N_23889);
xnor U28291 (N_28291,N_22619,N_21043);
or U28292 (N_28292,N_22334,N_22770);
nor U28293 (N_28293,N_24702,N_22166);
nand U28294 (N_28294,N_20367,N_23226);
and U28295 (N_28295,N_21023,N_20448);
and U28296 (N_28296,N_20054,N_21183);
or U28297 (N_28297,N_21556,N_21851);
and U28298 (N_28298,N_24457,N_20045);
xor U28299 (N_28299,N_20159,N_21789);
nor U28300 (N_28300,N_21965,N_24978);
nand U28301 (N_28301,N_23924,N_20051);
xnor U28302 (N_28302,N_24691,N_22733);
nand U28303 (N_28303,N_22032,N_24168);
xnor U28304 (N_28304,N_20500,N_21954);
or U28305 (N_28305,N_20594,N_22360);
xnor U28306 (N_28306,N_21206,N_22143);
nand U28307 (N_28307,N_24004,N_20136);
or U28308 (N_28308,N_24961,N_21780);
nand U28309 (N_28309,N_22829,N_21280);
nand U28310 (N_28310,N_20926,N_23560);
and U28311 (N_28311,N_22676,N_23249);
nand U28312 (N_28312,N_24538,N_20568);
nand U28313 (N_28313,N_21645,N_22723);
nand U28314 (N_28314,N_24241,N_20909);
nor U28315 (N_28315,N_23706,N_23366);
or U28316 (N_28316,N_23902,N_24327);
nor U28317 (N_28317,N_20520,N_23790);
nand U28318 (N_28318,N_24225,N_21624);
or U28319 (N_28319,N_22267,N_21351);
or U28320 (N_28320,N_21905,N_20629);
or U28321 (N_28321,N_20606,N_21223);
xor U28322 (N_28322,N_24514,N_23326);
and U28323 (N_28323,N_24582,N_24657);
or U28324 (N_28324,N_22540,N_23255);
xnor U28325 (N_28325,N_23472,N_20034);
nor U28326 (N_28326,N_22831,N_22286);
and U28327 (N_28327,N_21489,N_20070);
nor U28328 (N_28328,N_20177,N_20869);
or U28329 (N_28329,N_22447,N_21195);
nand U28330 (N_28330,N_23623,N_23990);
nand U28331 (N_28331,N_23300,N_21995);
xnor U28332 (N_28332,N_22898,N_21014);
and U28333 (N_28333,N_24142,N_24851);
and U28334 (N_28334,N_21617,N_20489);
nor U28335 (N_28335,N_24856,N_22555);
nand U28336 (N_28336,N_23124,N_21251);
and U28337 (N_28337,N_23404,N_24890);
nor U28338 (N_28338,N_20784,N_23532);
or U28339 (N_28339,N_20159,N_23207);
and U28340 (N_28340,N_20321,N_20673);
or U28341 (N_28341,N_21981,N_20996);
xor U28342 (N_28342,N_23554,N_24809);
nor U28343 (N_28343,N_20345,N_22305);
and U28344 (N_28344,N_23856,N_22140);
nor U28345 (N_28345,N_23168,N_20817);
xor U28346 (N_28346,N_21917,N_20295);
or U28347 (N_28347,N_21232,N_23171);
nand U28348 (N_28348,N_21735,N_20248);
xor U28349 (N_28349,N_20769,N_21535);
nand U28350 (N_28350,N_21029,N_20978);
nand U28351 (N_28351,N_23714,N_20902);
xor U28352 (N_28352,N_22599,N_22749);
xor U28353 (N_28353,N_21653,N_21198);
nand U28354 (N_28354,N_21235,N_24994);
xor U28355 (N_28355,N_20110,N_24636);
and U28356 (N_28356,N_20647,N_21076);
nand U28357 (N_28357,N_22249,N_22859);
nor U28358 (N_28358,N_21432,N_20454);
nand U28359 (N_28359,N_23992,N_23478);
nand U28360 (N_28360,N_20471,N_22372);
nor U28361 (N_28361,N_20308,N_22977);
xor U28362 (N_28362,N_20609,N_21053);
and U28363 (N_28363,N_23465,N_20002);
or U28364 (N_28364,N_21712,N_20118);
and U28365 (N_28365,N_24529,N_22753);
xor U28366 (N_28366,N_21450,N_23441);
nor U28367 (N_28367,N_20604,N_23453);
nand U28368 (N_28368,N_24432,N_24608);
xnor U28369 (N_28369,N_20994,N_22991);
and U28370 (N_28370,N_21604,N_20335);
xnor U28371 (N_28371,N_20172,N_24773);
nor U28372 (N_28372,N_21938,N_22037);
or U28373 (N_28373,N_24452,N_20026);
xnor U28374 (N_28374,N_24699,N_21071);
nor U28375 (N_28375,N_22793,N_23358);
xor U28376 (N_28376,N_20181,N_23021);
or U28377 (N_28377,N_21563,N_21212);
xor U28378 (N_28378,N_20963,N_23572);
or U28379 (N_28379,N_24726,N_24949);
xor U28380 (N_28380,N_23442,N_22453);
or U28381 (N_28381,N_24702,N_22523);
nor U28382 (N_28382,N_24142,N_21478);
and U28383 (N_28383,N_24305,N_22677);
xor U28384 (N_28384,N_20665,N_21891);
xor U28385 (N_28385,N_22183,N_24385);
xnor U28386 (N_28386,N_22343,N_20417);
and U28387 (N_28387,N_23510,N_23340);
nand U28388 (N_28388,N_21655,N_20569);
nand U28389 (N_28389,N_23820,N_23931);
xnor U28390 (N_28390,N_22609,N_23801);
nand U28391 (N_28391,N_24829,N_24838);
xor U28392 (N_28392,N_21541,N_22804);
nor U28393 (N_28393,N_24388,N_20287);
and U28394 (N_28394,N_22498,N_24900);
nand U28395 (N_28395,N_23921,N_21106);
nand U28396 (N_28396,N_21260,N_24613);
nand U28397 (N_28397,N_24831,N_24691);
and U28398 (N_28398,N_20370,N_21902);
or U28399 (N_28399,N_24475,N_20675);
or U28400 (N_28400,N_24639,N_20573);
xor U28401 (N_28401,N_21040,N_22079);
xnor U28402 (N_28402,N_21014,N_24836);
xnor U28403 (N_28403,N_21486,N_22957);
and U28404 (N_28404,N_23847,N_20676);
or U28405 (N_28405,N_24295,N_23291);
nand U28406 (N_28406,N_23659,N_24469);
xnor U28407 (N_28407,N_21473,N_23309);
and U28408 (N_28408,N_21687,N_22234);
nor U28409 (N_28409,N_23935,N_24461);
and U28410 (N_28410,N_21119,N_21691);
or U28411 (N_28411,N_22590,N_21014);
nor U28412 (N_28412,N_23247,N_24006);
and U28413 (N_28413,N_20785,N_21722);
xor U28414 (N_28414,N_22783,N_21578);
xnor U28415 (N_28415,N_21927,N_22081);
and U28416 (N_28416,N_23754,N_21858);
or U28417 (N_28417,N_22587,N_23928);
nor U28418 (N_28418,N_23967,N_21698);
and U28419 (N_28419,N_21701,N_22848);
xnor U28420 (N_28420,N_23599,N_24166);
nand U28421 (N_28421,N_21451,N_23773);
xor U28422 (N_28422,N_24987,N_22068);
nand U28423 (N_28423,N_21971,N_23654);
xnor U28424 (N_28424,N_23767,N_24032);
xnor U28425 (N_28425,N_21685,N_23875);
nand U28426 (N_28426,N_22291,N_22710);
xnor U28427 (N_28427,N_22810,N_23343);
nor U28428 (N_28428,N_20197,N_24150);
xnor U28429 (N_28429,N_20880,N_24682);
or U28430 (N_28430,N_23525,N_20319);
nor U28431 (N_28431,N_21989,N_20056);
xnor U28432 (N_28432,N_20665,N_24393);
and U28433 (N_28433,N_23363,N_22811);
xor U28434 (N_28434,N_21506,N_23907);
xnor U28435 (N_28435,N_23887,N_22506);
nor U28436 (N_28436,N_21021,N_24391);
xor U28437 (N_28437,N_21539,N_22987);
nand U28438 (N_28438,N_20438,N_21516);
or U28439 (N_28439,N_20331,N_20790);
nand U28440 (N_28440,N_24573,N_23918);
nand U28441 (N_28441,N_22247,N_24269);
and U28442 (N_28442,N_21338,N_21635);
or U28443 (N_28443,N_20491,N_24371);
or U28444 (N_28444,N_24372,N_21906);
nand U28445 (N_28445,N_21277,N_23104);
and U28446 (N_28446,N_23434,N_24211);
nor U28447 (N_28447,N_22134,N_20853);
and U28448 (N_28448,N_20392,N_24260);
and U28449 (N_28449,N_23997,N_21442);
nand U28450 (N_28450,N_23307,N_23629);
nor U28451 (N_28451,N_21533,N_24577);
nand U28452 (N_28452,N_22786,N_24233);
nor U28453 (N_28453,N_22419,N_24919);
xnor U28454 (N_28454,N_24320,N_21736);
or U28455 (N_28455,N_22257,N_24146);
nor U28456 (N_28456,N_21966,N_21270);
nand U28457 (N_28457,N_20489,N_24094);
nor U28458 (N_28458,N_21304,N_24503);
xnor U28459 (N_28459,N_24649,N_22821);
nor U28460 (N_28460,N_24179,N_21868);
xnor U28461 (N_28461,N_22429,N_23827);
nor U28462 (N_28462,N_22924,N_24067);
nand U28463 (N_28463,N_23021,N_20699);
xor U28464 (N_28464,N_21597,N_21961);
nor U28465 (N_28465,N_20496,N_24815);
nor U28466 (N_28466,N_24666,N_20002);
xnor U28467 (N_28467,N_20735,N_21099);
nor U28468 (N_28468,N_21991,N_20739);
and U28469 (N_28469,N_21485,N_20507);
nor U28470 (N_28470,N_22610,N_22403);
nor U28471 (N_28471,N_24890,N_23428);
or U28472 (N_28472,N_23581,N_24959);
nand U28473 (N_28473,N_22432,N_21945);
xor U28474 (N_28474,N_20448,N_20452);
xnor U28475 (N_28475,N_23933,N_23721);
xor U28476 (N_28476,N_20983,N_23877);
nor U28477 (N_28477,N_23158,N_20892);
or U28478 (N_28478,N_21003,N_24785);
and U28479 (N_28479,N_23261,N_24551);
and U28480 (N_28480,N_21568,N_20741);
or U28481 (N_28481,N_22869,N_24974);
or U28482 (N_28482,N_21895,N_22934);
nor U28483 (N_28483,N_24657,N_20794);
and U28484 (N_28484,N_23141,N_22864);
or U28485 (N_28485,N_20644,N_21230);
or U28486 (N_28486,N_23761,N_21625);
or U28487 (N_28487,N_24019,N_20871);
nand U28488 (N_28488,N_21329,N_20978);
or U28489 (N_28489,N_22653,N_24137);
nand U28490 (N_28490,N_23821,N_20400);
or U28491 (N_28491,N_23277,N_22966);
nand U28492 (N_28492,N_20058,N_24364);
nor U28493 (N_28493,N_20147,N_23860);
or U28494 (N_28494,N_23304,N_21114);
or U28495 (N_28495,N_24140,N_22062);
xnor U28496 (N_28496,N_20517,N_24787);
or U28497 (N_28497,N_21330,N_20856);
nor U28498 (N_28498,N_24538,N_21786);
and U28499 (N_28499,N_23007,N_23398);
nor U28500 (N_28500,N_20271,N_21999);
and U28501 (N_28501,N_23974,N_20832);
nor U28502 (N_28502,N_22690,N_20249);
nor U28503 (N_28503,N_23381,N_20214);
xor U28504 (N_28504,N_23593,N_22410);
and U28505 (N_28505,N_24108,N_20227);
nor U28506 (N_28506,N_22493,N_22585);
nor U28507 (N_28507,N_20054,N_24863);
nor U28508 (N_28508,N_20158,N_24424);
xnor U28509 (N_28509,N_20643,N_22563);
xor U28510 (N_28510,N_22315,N_21232);
nor U28511 (N_28511,N_23148,N_20411);
xor U28512 (N_28512,N_23648,N_24819);
nor U28513 (N_28513,N_24832,N_20223);
and U28514 (N_28514,N_20953,N_22826);
nand U28515 (N_28515,N_21029,N_23812);
nand U28516 (N_28516,N_22368,N_20780);
xor U28517 (N_28517,N_22913,N_24096);
and U28518 (N_28518,N_22606,N_21990);
nor U28519 (N_28519,N_24755,N_21153);
or U28520 (N_28520,N_24803,N_23133);
or U28521 (N_28521,N_20222,N_23358);
nor U28522 (N_28522,N_21077,N_21478);
or U28523 (N_28523,N_24924,N_23286);
nand U28524 (N_28524,N_22514,N_20476);
nor U28525 (N_28525,N_21337,N_21766);
and U28526 (N_28526,N_24647,N_24527);
or U28527 (N_28527,N_22474,N_20602);
or U28528 (N_28528,N_23653,N_21932);
xnor U28529 (N_28529,N_21806,N_22932);
or U28530 (N_28530,N_20592,N_22757);
nor U28531 (N_28531,N_20460,N_21919);
xor U28532 (N_28532,N_23210,N_24754);
nor U28533 (N_28533,N_23869,N_22680);
xnor U28534 (N_28534,N_22295,N_23306);
or U28535 (N_28535,N_21294,N_22373);
nor U28536 (N_28536,N_22854,N_22065);
nand U28537 (N_28537,N_21793,N_21203);
xor U28538 (N_28538,N_21396,N_23765);
nor U28539 (N_28539,N_22353,N_23369);
or U28540 (N_28540,N_20731,N_23909);
nor U28541 (N_28541,N_21605,N_20225);
and U28542 (N_28542,N_24154,N_22318);
nor U28543 (N_28543,N_21599,N_22921);
nand U28544 (N_28544,N_23288,N_23808);
xnor U28545 (N_28545,N_24224,N_20802);
nand U28546 (N_28546,N_21083,N_24849);
and U28547 (N_28547,N_22468,N_22233);
nand U28548 (N_28548,N_20271,N_20748);
or U28549 (N_28549,N_21813,N_24369);
or U28550 (N_28550,N_20830,N_21563);
or U28551 (N_28551,N_22146,N_22024);
and U28552 (N_28552,N_23488,N_20545);
xnor U28553 (N_28553,N_24704,N_21458);
or U28554 (N_28554,N_20964,N_20657);
xor U28555 (N_28555,N_20088,N_22151);
or U28556 (N_28556,N_21513,N_21731);
and U28557 (N_28557,N_21614,N_21703);
or U28558 (N_28558,N_22976,N_24388);
nand U28559 (N_28559,N_23175,N_22117);
or U28560 (N_28560,N_20952,N_23481);
xor U28561 (N_28561,N_20737,N_24457);
and U28562 (N_28562,N_21172,N_20605);
nand U28563 (N_28563,N_22237,N_20480);
xnor U28564 (N_28564,N_23486,N_22839);
and U28565 (N_28565,N_20028,N_23930);
nor U28566 (N_28566,N_23346,N_22488);
or U28567 (N_28567,N_20444,N_24196);
nand U28568 (N_28568,N_21825,N_24791);
and U28569 (N_28569,N_21370,N_23913);
xor U28570 (N_28570,N_24431,N_21581);
xnor U28571 (N_28571,N_23653,N_22162);
nor U28572 (N_28572,N_23828,N_22732);
and U28573 (N_28573,N_23691,N_24908);
and U28574 (N_28574,N_24794,N_21352);
xnor U28575 (N_28575,N_24009,N_21113);
xnor U28576 (N_28576,N_21922,N_20695);
nor U28577 (N_28577,N_24260,N_24902);
xnor U28578 (N_28578,N_20820,N_24782);
or U28579 (N_28579,N_20758,N_24588);
nor U28580 (N_28580,N_24863,N_22764);
nand U28581 (N_28581,N_21054,N_21991);
nor U28582 (N_28582,N_21225,N_21743);
nand U28583 (N_28583,N_21076,N_23569);
nand U28584 (N_28584,N_21543,N_22827);
or U28585 (N_28585,N_23018,N_23213);
xor U28586 (N_28586,N_21925,N_23013);
and U28587 (N_28587,N_21539,N_23989);
or U28588 (N_28588,N_20413,N_21346);
nand U28589 (N_28589,N_23641,N_21686);
and U28590 (N_28590,N_23495,N_22353);
nor U28591 (N_28591,N_21967,N_20163);
or U28592 (N_28592,N_20253,N_23373);
nand U28593 (N_28593,N_20843,N_20409);
and U28594 (N_28594,N_23925,N_20904);
and U28595 (N_28595,N_21283,N_22393);
nand U28596 (N_28596,N_20880,N_22146);
xnor U28597 (N_28597,N_24463,N_21278);
and U28598 (N_28598,N_20572,N_22203);
or U28599 (N_28599,N_24809,N_22843);
nand U28600 (N_28600,N_22882,N_24985);
or U28601 (N_28601,N_24051,N_21008);
or U28602 (N_28602,N_22488,N_20171);
nand U28603 (N_28603,N_20892,N_22245);
xnor U28604 (N_28604,N_21316,N_23228);
xor U28605 (N_28605,N_24229,N_24242);
nand U28606 (N_28606,N_21790,N_23856);
or U28607 (N_28607,N_22293,N_23432);
or U28608 (N_28608,N_23351,N_23040);
and U28609 (N_28609,N_20342,N_23990);
and U28610 (N_28610,N_22916,N_20345);
or U28611 (N_28611,N_22510,N_22014);
or U28612 (N_28612,N_20567,N_20885);
xor U28613 (N_28613,N_24045,N_24738);
and U28614 (N_28614,N_24932,N_20375);
xor U28615 (N_28615,N_23687,N_21263);
and U28616 (N_28616,N_24318,N_23151);
and U28617 (N_28617,N_22919,N_22779);
or U28618 (N_28618,N_22012,N_21915);
nor U28619 (N_28619,N_21116,N_20182);
xnor U28620 (N_28620,N_24435,N_24151);
nand U28621 (N_28621,N_22603,N_24870);
nor U28622 (N_28622,N_22375,N_22269);
nand U28623 (N_28623,N_21542,N_20116);
nand U28624 (N_28624,N_20267,N_23563);
xnor U28625 (N_28625,N_23405,N_24497);
xor U28626 (N_28626,N_22151,N_20939);
and U28627 (N_28627,N_20306,N_21436);
and U28628 (N_28628,N_23771,N_24582);
xnor U28629 (N_28629,N_20012,N_24627);
and U28630 (N_28630,N_21371,N_24002);
nand U28631 (N_28631,N_23214,N_20138);
and U28632 (N_28632,N_21560,N_22134);
xor U28633 (N_28633,N_20309,N_21449);
xnor U28634 (N_28634,N_21427,N_23622);
xnor U28635 (N_28635,N_21133,N_22762);
or U28636 (N_28636,N_23577,N_24097);
or U28637 (N_28637,N_24643,N_23924);
or U28638 (N_28638,N_24759,N_22996);
nand U28639 (N_28639,N_24029,N_21971);
or U28640 (N_28640,N_21101,N_24751);
nand U28641 (N_28641,N_21583,N_24661);
nor U28642 (N_28642,N_21189,N_23977);
nor U28643 (N_28643,N_20892,N_21114);
and U28644 (N_28644,N_20606,N_22340);
or U28645 (N_28645,N_24941,N_22150);
and U28646 (N_28646,N_23198,N_23995);
nor U28647 (N_28647,N_20656,N_21333);
nor U28648 (N_28648,N_21530,N_23318);
nor U28649 (N_28649,N_24124,N_22817);
nor U28650 (N_28650,N_21276,N_23989);
and U28651 (N_28651,N_24581,N_23553);
nor U28652 (N_28652,N_20305,N_24316);
nand U28653 (N_28653,N_20922,N_20284);
xor U28654 (N_28654,N_23653,N_20298);
nor U28655 (N_28655,N_20443,N_23307);
and U28656 (N_28656,N_20686,N_20682);
nand U28657 (N_28657,N_22592,N_21211);
or U28658 (N_28658,N_20623,N_23654);
xor U28659 (N_28659,N_23955,N_21052);
nor U28660 (N_28660,N_24069,N_24400);
nand U28661 (N_28661,N_21666,N_22728);
and U28662 (N_28662,N_22180,N_24653);
or U28663 (N_28663,N_24386,N_21093);
or U28664 (N_28664,N_20620,N_22198);
or U28665 (N_28665,N_24856,N_21072);
nor U28666 (N_28666,N_23965,N_22342);
and U28667 (N_28667,N_21747,N_24130);
nand U28668 (N_28668,N_22110,N_21654);
xor U28669 (N_28669,N_21179,N_20654);
and U28670 (N_28670,N_24474,N_20841);
xor U28671 (N_28671,N_21590,N_21816);
xnor U28672 (N_28672,N_24889,N_21111);
nand U28673 (N_28673,N_21152,N_21331);
or U28674 (N_28674,N_22937,N_22370);
and U28675 (N_28675,N_24217,N_21131);
and U28676 (N_28676,N_20405,N_22379);
and U28677 (N_28677,N_23163,N_24458);
nor U28678 (N_28678,N_23716,N_22066);
or U28679 (N_28679,N_20817,N_21855);
and U28680 (N_28680,N_24787,N_24549);
nand U28681 (N_28681,N_23820,N_22115);
nand U28682 (N_28682,N_22662,N_24904);
nand U28683 (N_28683,N_21368,N_20840);
nor U28684 (N_28684,N_20063,N_24542);
or U28685 (N_28685,N_20962,N_20587);
nand U28686 (N_28686,N_22012,N_24270);
nor U28687 (N_28687,N_24278,N_23897);
and U28688 (N_28688,N_21193,N_21032);
nor U28689 (N_28689,N_21344,N_23674);
or U28690 (N_28690,N_22496,N_21009);
xnor U28691 (N_28691,N_23167,N_24482);
nand U28692 (N_28692,N_24495,N_24320);
nor U28693 (N_28693,N_20240,N_23444);
xnor U28694 (N_28694,N_23567,N_24644);
or U28695 (N_28695,N_20474,N_20042);
or U28696 (N_28696,N_20356,N_21665);
xor U28697 (N_28697,N_24674,N_24104);
nand U28698 (N_28698,N_21614,N_21874);
nand U28699 (N_28699,N_23413,N_23747);
nor U28700 (N_28700,N_21297,N_24755);
nor U28701 (N_28701,N_21901,N_24180);
xnor U28702 (N_28702,N_20285,N_24079);
nor U28703 (N_28703,N_24761,N_21775);
nand U28704 (N_28704,N_24000,N_22584);
nand U28705 (N_28705,N_24212,N_22715);
xnor U28706 (N_28706,N_21632,N_22125);
nand U28707 (N_28707,N_23312,N_24645);
or U28708 (N_28708,N_23527,N_21282);
or U28709 (N_28709,N_21634,N_23311);
and U28710 (N_28710,N_21294,N_23015);
xor U28711 (N_28711,N_20635,N_20564);
nor U28712 (N_28712,N_22618,N_24304);
and U28713 (N_28713,N_23312,N_21900);
or U28714 (N_28714,N_20511,N_20170);
or U28715 (N_28715,N_23768,N_20310);
nor U28716 (N_28716,N_22482,N_23914);
nand U28717 (N_28717,N_20329,N_22346);
xor U28718 (N_28718,N_21291,N_23367);
nand U28719 (N_28719,N_22796,N_23248);
nor U28720 (N_28720,N_22402,N_20868);
and U28721 (N_28721,N_20176,N_24267);
or U28722 (N_28722,N_20951,N_24134);
and U28723 (N_28723,N_23795,N_24613);
xnor U28724 (N_28724,N_22245,N_23841);
nor U28725 (N_28725,N_20158,N_21971);
xor U28726 (N_28726,N_23385,N_22714);
nand U28727 (N_28727,N_23008,N_24172);
xor U28728 (N_28728,N_20192,N_20584);
or U28729 (N_28729,N_22450,N_20131);
nor U28730 (N_28730,N_21357,N_23747);
xor U28731 (N_28731,N_21559,N_21719);
and U28732 (N_28732,N_23997,N_21123);
nand U28733 (N_28733,N_21867,N_20228);
xnor U28734 (N_28734,N_22488,N_21985);
xor U28735 (N_28735,N_21665,N_21235);
nor U28736 (N_28736,N_24905,N_20097);
and U28737 (N_28737,N_23599,N_20741);
and U28738 (N_28738,N_24069,N_21137);
and U28739 (N_28739,N_21172,N_22415);
nor U28740 (N_28740,N_21618,N_21525);
or U28741 (N_28741,N_23899,N_24636);
and U28742 (N_28742,N_23733,N_23003);
nor U28743 (N_28743,N_22940,N_21048);
or U28744 (N_28744,N_21403,N_23237);
nor U28745 (N_28745,N_21817,N_23982);
or U28746 (N_28746,N_22868,N_21672);
or U28747 (N_28747,N_21766,N_24285);
and U28748 (N_28748,N_24270,N_21103);
or U28749 (N_28749,N_24886,N_20972);
and U28750 (N_28750,N_23087,N_22187);
xnor U28751 (N_28751,N_22426,N_21705);
nor U28752 (N_28752,N_23852,N_23682);
nand U28753 (N_28753,N_21504,N_24813);
or U28754 (N_28754,N_21237,N_22616);
or U28755 (N_28755,N_22545,N_21993);
xor U28756 (N_28756,N_22278,N_24101);
nand U28757 (N_28757,N_21064,N_22541);
xor U28758 (N_28758,N_23278,N_20477);
nand U28759 (N_28759,N_23446,N_22859);
and U28760 (N_28760,N_23031,N_23456);
nor U28761 (N_28761,N_20191,N_22640);
nor U28762 (N_28762,N_23836,N_22200);
nor U28763 (N_28763,N_24308,N_22888);
or U28764 (N_28764,N_20828,N_24479);
and U28765 (N_28765,N_22912,N_23153);
nand U28766 (N_28766,N_22326,N_21717);
nand U28767 (N_28767,N_21589,N_21474);
or U28768 (N_28768,N_23615,N_20472);
nor U28769 (N_28769,N_23988,N_22467);
xor U28770 (N_28770,N_21786,N_21679);
and U28771 (N_28771,N_22614,N_21727);
xor U28772 (N_28772,N_23969,N_23988);
nor U28773 (N_28773,N_20197,N_20533);
and U28774 (N_28774,N_24705,N_23258);
and U28775 (N_28775,N_20709,N_23773);
nor U28776 (N_28776,N_22999,N_24731);
and U28777 (N_28777,N_23557,N_22503);
or U28778 (N_28778,N_24592,N_20915);
nor U28779 (N_28779,N_20011,N_21773);
xor U28780 (N_28780,N_21664,N_22634);
nand U28781 (N_28781,N_23896,N_20215);
and U28782 (N_28782,N_20587,N_22220);
or U28783 (N_28783,N_21834,N_21562);
nand U28784 (N_28784,N_22039,N_20564);
nor U28785 (N_28785,N_21457,N_21074);
and U28786 (N_28786,N_24846,N_22882);
nand U28787 (N_28787,N_20610,N_23423);
nor U28788 (N_28788,N_23303,N_22665);
and U28789 (N_28789,N_23513,N_21449);
and U28790 (N_28790,N_21809,N_20218);
nor U28791 (N_28791,N_21445,N_21152);
nand U28792 (N_28792,N_20790,N_21855);
or U28793 (N_28793,N_23489,N_21584);
and U28794 (N_28794,N_23320,N_24947);
and U28795 (N_28795,N_22183,N_23157);
xor U28796 (N_28796,N_24577,N_21275);
xor U28797 (N_28797,N_24178,N_22193);
or U28798 (N_28798,N_23912,N_22212);
nand U28799 (N_28799,N_23016,N_20388);
or U28800 (N_28800,N_23233,N_22764);
and U28801 (N_28801,N_23622,N_23349);
nor U28802 (N_28802,N_21019,N_22802);
nor U28803 (N_28803,N_21380,N_22675);
or U28804 (N_28804,N_24330,N_24908);
and U28805 (N_28805,N_21842,N_21782);
and U28806 (N_28806,N_24668,N_23005);
or U28807 (N_28807,N_22479,N_20790);
and U28808 (N_28808,N_21612,N_24258);
nand U28809 (N_28809,N_21813,N_23679);
xor U28810 (N_28810,N_20695,N_22767);
or U28811 (N_28811,N_24503,N_21324);
nor U28812 (N_28812,N_22326,N_23655);
nor U28813 (N_28813,N_23288,N_21216);
or U28814 (N_28814,N_22540,N_22809);
nand U28815 (N_28815,N_20531,N_23200);
and U28816 (N_28816,N_24362,N_24807);
and U28817 (N_28817,N_21177,N_22056);
and U28818 (N_28818,N_20370,N_21105);
nand U28819 (N_28819,N_23642,N_22260);
xor U28820 (N_28820,N_20203,N_24863);
or U28821 (N_28821,N_22502,N_22322);
xor U28822 (N_28822,N_23192,N_20216);
and U28823 (N_28823,N_21346,N_23139);
nand U28824 (N_28824,N_20551,N_24101);
xnor U28825 (N_28825,N_22741,N_20005);
or U28826 (N_28826,N_24477,N_23280);
nand U28827 (N_28827,N_21950,N_24602);
and U28828 (N_28828,N_22993,N_24660);
nand U28829 (N_28829,N_23175,N_21728);
or U28830 (N_28830,N_21017,N_24074);
nand U28831 (N_28831,N_22322,N_24230);
nand U28832 (N_28832,N_24099,N_23389);
and U28833 (N_28833,N_23332,N_23585);
and U28834 (N_28834,N_23525,N_21749);
and U28835 (N_28835,N_24928,N_20620);
or U28836 (N_28836,N_24109,N_20025);
or U28837 (N_28837,N_21492,N_22049);
and U28838 (N_28838,N_22922,N_23370);
nor U28839 (N_28839,N_22098,N_21000);
and U28840 (N_28840,N_20893,N_21274);
xor U28841 (N_28841,N_20231,N_22381);
or U28842 (N_28842,N_24846,N_21712);
nand U28843 (N_28843,N_23691,N_22717);
nand U28844 (N_28844,N_21895,N_23454);
or U28845 (N_28845,N_23736,N_24116);
nand U28846 (N_28846,N_23513,N_20967);
nor U28847 (N_28847,N_22308,N_21719);
or U28848 (N_28848,N_22953,N_21420);
and U28849 (N_28849,N_23145,N_24420);
xor U28850 (N_28850,N_23292,N_22880);
xnor U28851 (N_28851,N_24809,N_22689);
nand U28852 (N_28852,N_20349,N_24708);
and U28853 (N_28853,N_22460,N_20574);
nand U28854 (N_28854,N_22387,N_21994);
nand U28855 (N_28855,N_23506,N_20345);
and U28856 (N_28856,N_21071,N_23008);
nor U28857 (N_28857,N_20367,N_22656);
nand U28858 (N_28858,N_24275,N_24205);
or U28859 (N_28859,N_24632,N_20549);
nor U28860 (N_28860,N_22907,N_20691);
nand U28861 (N_28861,N_22491,N_24242);
nor U28862 (N_28862,N_22097,N_21104);
or U28863 (N_28863,N_20540,N_23273);
and U28864 (N_28864,N_22964,N_20128);
and U28865 (N_28865,N_23841,N_22854);
nor U28866 (N_28866,N_22101,N_21491);
or U28867 (N_28867,N_21612,N_24851);
nand U28868 (N_28868,N_22798,N_20605);
xnor U28869 (N_28869,N_20717,N_23021);
and U28870 (N_28870,N_23046,N_22126);
nor U28871 (N_28871,N_22870,N_20783);
nor U28872 (N_28872,N_24625,N_24545);
or U28873 (N_28873,N_21450,N_22929);
and U28874 (N_28874,N_21972,N_20589);
nor U28875 (N_28875,N_22682,N_24878);
and U28876 (N_28876,N_23290,N_24790);
xor U28877 (N_28877,N_22242,N_23305);
nand U28878 (N_28878,N_21139,N_23611);
nand U28879 (N_28879,N_24798,N_20927);
nor U28880 (N_28880,N_21810,N_23867);
and U28881 (N_28881,N_24140,N_21722);
nand U28882 (N_28882,N_21478,N_21836);
nand U28883 (N_28883,N_21318,N_20345);
xnor U28884 (N_28884,N_23557,N_20423);
or U28885 (N_28885,N_22455,N_22368);
and U28886 (N_28886,N_23980,N_21246);
or U28887 (N_28887,N_23405,N_21598);
and U28888 (N_28888,N_24579,N_21266);
nand U28889 (N_28889,N_23897,N_24978);
nand U28890 (N_28890,N_24458,N_21099);
nand U28891 (N_28891,N_20667,N_20940);
and U28892 (N_28892,N_22288,N_23567);
nor U28893 (N_28893,N_23880,N_24749);
and U28894 (N_28894,N_21805,N_23659);
nand U28895 (N_28895,N_22859,N_22491);
nand U28896 (N_28896,N_20669,N_23620);
or U28897 (N_28897,N_21026,N_21860);
nor U28898 (N_28898,N_23028,N_23048);
nor U28899 (N_28899,N_22145,N_24280);
and U28900 (N_28900,N_23167,N_22164);
nor U28901 (N_28901,N_21901,N_20637);
xor U28902 (N_28902,N_21916,N_23982);
nor U28903 (N_28903,N_23172,N_20714);
xor U28904 (N_28904,N_20695,N_20113);
nand U28905 (N_28905,N_24826,N_24206);
xnor U28906 (N_28906,N_24524,N_20347);
and U28907 (N_28907,N_24903,N_22586);
or U28908 (N_28908,N_22260,N_20943);
or U28909 (N_28909,N_22072,N_20102);
or U28910 (N_28910,N_23310,N_22950);
or U28911 (N_28911,N_24793,N_24422);
nor U28912 (N_28912,N_22691,N_20209);
xnor U28913 (N_28913,N_23389,N_23709);
nor U28914 (N_28914,N_24566,N_21458);
xnor U28915 (N_28915,N_22346,N_20806);
and U28916 (N_28916,N_21819,N_21952);
and U28917 (N_28917,N_22842,N_23055);
and U28918 (N_28918,N_24389,N_21120);
nand U28919 (N_28919,N_22455,N_23988);
nand U28920 (N_28920,N_23965,N_23581);
xnor U28921 (N_28921,N_20512,N_20202);
nand U28922 (N_28922,N_22016,N_23764);
nand U28923 (N_28923,N_21376,N_20439);
or U28924 (N_28924,N_23392,N_24678);
nand U28925 (N_28925,N_24073,N_20614);
or U28926 (N_28926,N_21226,N_22344);
xnor U28927 (N_28927,N_23199,N_23830);
or U28928 (N_28928,N_22104,N_21296);
nor U28929 (N_28929,N_24348,N_21229);
or U28930 (N_28930,N_24026,N_22883);
nand U28931 (N_28931,N_20720,N_21486);
nand U28932 (N_28932,N_23337,N_22923);
nor U28933 (N_28933,N_23552,N_23582);
and U28934 (N_28934,N_20212,N_24829);
and U28935 (N_28935,N_24207,N_23947);
and U28936 (N_28936,N_24615,N_21736);
xor U28937 (N_28937,N_20515,N_20316);
nand U28938 (N_28938,N_20989,N_20847);
nor U28939 (N_28939,N_20075,N_23775);
xnor U28940 (N_28940,N_20142,N_22503);
nor U28941 (N_28941,N_20361,N_21708);
xnor U28942 (N_28942,N_22662,N_24771);
xnor U28943 (N_28943,N_22844,N_22456);
nor U28944 (N_28944,N_23282,N_22965);
and U28945 (N_28945,N_23218,N_21672);
nand U28946 (N_28946,N_23732,N_22805);
nand U28947 (N_28947,N_24806,N_20036);
nand U28948 (N_28948,N_20356,N_20235);
or U28949 (N_28949,N_21628,N_22720);
and U28950 (N_28950,N_20250,N_24233);
and U28951 (N_28951,N_22851,N_20840);
xor U28952 (N_28952,N_21587,N_20572);
xor U28953 (N_28953,N_23843,N_22016);
or U28954 (N_28954,N_22602,N_24843);
xnor U28955 (N_28955,N_20272,N_22441);
nand U28956 (N_28956,N_24270,N_24535);
nor U28957 (N_28957,N_20003,N_22083);
and U28958 (N_28958,N_23939,N_21381);
or U28959 (N_28959,N_22229,N_24999);
xor U28960 (N_28960,N_23890,N_23277);
nor U28961 (N_28961,N_23569,N_21071);
xnor U28962 (N_28962,N_22484,N_23332);
nand U28963 (N_28963,N_24286,N_23193);
nand U28964 (N_28964,N_20655,N_22313);
and U28965 (N_28965,N_21961,N_23931);
or U28966 (N_28966,N_24740,N_20198);
nand U28967 (N_28967,N_21193,N_23397);
nor U28968 (N_28968,N_22395,N_20277);
and U28969 (N_28969,N_21283,N_20261);
xnor U28970 (N_28970,N_22032,N_22951);
xnor U28971 (N_28971,N_24220,N_23298);
or U28972 (N_28972,N_23170,N_24316);
xnor U28973 (N_28973,N_20692,N_22660);
xnor U28974 (N_28974,N_22548,N_24477);
and U28975 (N_28975,N_20734,N_20763);
nor U28976 (N_28976,N_22802,N_20566);
and U28977 (N_28977,N_20812,N_22497);
and U28978 (N_28978,N_22600,N_23839);
xor U28979 (N_28979,N_22277,N_23745);
or U28980 (N_28980,N_24908,N_23699);
xnor U28981 (N_28981,N_23756,N_20936);
xor U28982 (N_28982,N_21270,N_20617);
nor U28983 (N_28983,N_21892,N_22471);
nor U28984 (N_28984,N_23363,N_22825);
and U28985 (N_28985,N_20829,N_21145);
and U28986 (N_28986,N_21347,N_24626);
and U28987 (N_28987,N_20127,N_23883);
nand U28988 (N_28988,N_23752,N_23694);
or U28989 (N_28989,N_20587,N_24117);
xor U28990 (N_28990,N_21076,N_22519);
xor U28991 (N_28991,N_20654,N_22076);
and U28992 (N_28992,N_23693,N_23934);
or U28993 (N_28993,N_22608,N_22559);
or U28994 (N_28994,N_24309,N_24708);
nand U28995 (N_28995,N_24203,N_24293);
or U28996 (N_28996,N_24485,N_21400);
xor U28997 (N_28997,N_20352,N_22860);
and U28998 (N_28998,N_20908,N_24991);
and U28999 (N_28999,N_22580,N_20847);
and U29000 (N_29000,N_23735,N_21852);
nor U29001 (N_29001,N_22822,N_23568);
or U29002 (N_29002,N_20350,N_21978);
xnor U29003 (N_29003,N_23988,N_21691);
nor U29004 (N_29004,N_20317,N_20329);
or U29005 (N_29005,N_24678,N_21123);
nand U29006 (N_29006,N_22466,N_23067);
and U29007 (N_29007,N_23656,N_24658);
nand U29008 (N_29008,N_24024,N_21499);
nand U29009 (N_29009,N_24008,N_21491);
or U29010 (N_29010,N_22131,N_23244);
or U29011 (N_29011,N_24026,N_24806);
nor U29012 (N_29012,N_21698,N_21861);
or U29013 (N_29013,N_24343,N_22025);
nand U29014 (N_29014,N_23351,N_22503);
and U29015 (N_29015,N_21771,N_22773);
nand U29016 (N_29016,N_23788,N_24451);
nand U29017 (N_29017,N_20569,N_22776);
nand U29018 (N_29018,N_22269,N_20211);
nand U29019 (N_29019,N_21908,N_21211);
and U29020 (N_29020,N_24633,N_24296);
nand U29021 (N_29021,N_21436,N_24019);
and U29022 (N_29022,N_21604,N_24425);
xnor U29023 (N_29023,N_22357,N_22805);
or U29024 (N_29024,N_23926,N_20780);
and U29025 (N_29025,N_24976,N_21487);
and U29026 (N_29026,N_22469,N_24206);
xnor U29027 (N_29027,N_21566,N_23752);
xor U29028 (N_29028,N_22257,N_20720);
and U29029 (N_29029,N_22896,N_23201);
nand U29030 (N_29030,N_20895,N_22303);
xor U29031 (N_29031,N_20234,N_23635);
nor U29032 (N_29032,N_21885,N_24095);
xnor U29033 (N_29033,N_24190,N_22695);
nand U29034 (N_29034,N_21874,N_21983);
and U29035 (N_29035,N_23490,N_20364);
or U29036 (N_29036,N_24315,N_20157);
nor U29037 (N_29037,N_24619,N_23702);
nor U29038 (N_29038,N_24962,N_22092);
xor U29039 (N_29039,N_20666,N_23684);
or U29040 (N_29040,N_23138,N_21173);
nor U29041 (N_29041,N_24001,N_23217);
and U29042 (N_29042,N_22311,N_20278);
and U29043 (N_29043,N_20754,N_23006);
xnor U29044 (N_29044,N_24801,N_21130);
or U29045 (N_29045,N_24773,N_20262);
nand U29046 (N_29046,N_20370,N_22649);
and U29047 (N_29047,N_21982,N_20095);
nand U29048 (N_29048,N_23317,N_20045);
nand U29049 (N_29049,N_20843,N_24922);
and U29050 (N_29050,N_21176,N_21507);
xor U29051 (N_29051,N_22414,N_23295);
and U29052 (N_29052,N_20121,N_23889);
xor U29053 (N_29053,N_22564,N_20303);
and U29054 (N_29054,N_23806,N_23858);
nand U29055 (N_29055,N_21510,N_23173);
or U29056 (N_29056,N_21405,N_24793);
nor U29057 (N_29057,N_22691,N_23217);
and U29058 (N_29058,N_23317,N_24441);
nand U29059 (N_29059,N_20794,N_22593);
nand U29060 (N_29060,N_22871,N_22142);
nand U29061 (N_29061,N_21887,N_21021);
nand U29062 (N_29062,N_22895,N_21195);
or U29063 (N_29063,N_23101,N_22620);
nor U29064 (N_29064,N_22657,N_20104);
nand U29065 (N_29065,N_20533,N_23486);
and U29066 (N_29066,N_23308,N_24179);
xnor U29067 (N_29067,N_23974,N_20127);
nor U29068 (N_29068,N_23536,N_20310);
nand U29069 (N_29069,N_23559,N_24325);
or U29070 (N_29070,N_22726,N_22177);
nor U29071 (N_29071,N_22599,N_20849);
and U29072 (N_29072,N_23364,N_22497);
and U29073 (N_29073,N_23048,N_24127);
nand U29074 (N_29074,N_20540,N_24120);
nor U29075 (N_29075,N_20237,N_22638);
nand U29076 (N_29076,N_20054,N_24908);
nand U29077 (N_29077,N_24586,N_24144);
nand U29078 (N_29078,N_22388,N_21260);
nand U29079 (N_29079,N_24893,N_22637);
nand U29080 (N_29080,N_23246,N_21720);
or U29081 (N_29081,N_21130,N_20901);
or U29082 (N_29082,N_21113,N_23834);
and U29083 (N_29083,N_23711,N_24417);
nand U29084 (N_29084,N_21713,N_21867);
and U29085 (N_29085,N_23844,N_20888);
or U29086 (N_29086,N_22961,N_20764);
xnor U29087 (N_29087,N_23707,N_24518);
nor U29088 (N_29088,N_21278,N_23959);
nor U29089 (N_29089,N_20020,N_24927);
or U29090 (N_29090,N_21574,N_20900);
or U29091 (N_29091,N_21750,N_22278);
nor U29092 (N_29092,N_24808,N_23976);
and U29093 (N_29093,N_21470,N_24914);
or U29094 (N_29094,N_24349,N_21661);
nand U29095 (N_29095,N_23790,N_21701);
xor U29096 (N_29096,N_21914,N_24492);
or U29097 (N_29097,N_24308,N_21751);
and U29098 (N_29098,N_24538,N_20640);
nand U29099 (N_29099,N_20792,N_21389);
xnor U29100 (N_29100,N_22730,N_22399);
xor U29101 (N_29101,N_24877,N_24925);
nor U29102 (N_29102,N_23444,N_23792);
xnor U29103 (N_29103,N_21422,N_21065);
nor U29104 (N_29104,N_20408,N_24767);
nand U29105 (N_29105,N_24736,N_22678);
or U29106 (N_29106,N_20904,N_21962);
nand U29107 (N_29107,N_23296,N_21599);
and U29108 (N_29108,N_21426,N_20988);
nor U29109 (N_29109,N_23617,N_22187);
or U29110 (N_29110,N_22889,N_20383);
xor U29111 (N_29111,N_20544,N_23758);
nand U29112 (N_29112,N_20100,N_21628);
xnor U29113 (N_29113,N_23223,N_22265);
nand U29114 (N_29114,N_22382,N_21411);
xnor U29115 (N_29115,N_24474,N_24514);
or U29116 (N_29116,N_23166,N_21540);
xor U29117 (N_29117,N_21482,N_24015);
and U29118 (N_29118,N_22497,N_23956);
and U29119 (N_29119,N_20507,N_20266);
or U29120 (N_29120,N_20981,N_21783);
xor U29121 (N_29121,N_22410,N_22672);
nor U29122 (N_29122,N_20535,N_24406);
or U29123 (N_29123,N_21345,N_22414);
nor U29124 (N_29124,N_23834,N_22330);
xnor U29125 (N_29125,N_22765,N_20095);
xor U29126 (N_29126,N_23996,N_24282);
and U29127 (N_29127,N_21262,N_21303);
xnor U29128 (N_29128,N_22025,N_24358);
and U29129 (N_29129,N_24035,N_22892);
nor U29130 (N_29130,N_23766,N_24317);
xnor U29131 (N_29131,N_23248,N_21288);
or U29132 (N_29132,N_22160,N_20055);
and U29133 (N_29133,N_22620,N_22424);
nor U29134 (N_29134,N_22765,N_22885);
nand U29135 (N_29135,N_20007,N_20720);
nand U29136 (N_29136,N_20942,N_24727);
nand U29137 (N_29137,N_20264,N_22962);
nor U29138 (N_29138,N_24761,N_22274);
xor U29139 (N_29139,N_20703,N_24057);
and U29140 (N_29140,N_22753,N_24284);
and U29141 (N_29141,N_23310,N_21875);
xor U29142 (N_29142,N_21118,N_20838);
nor U29143 (N_29143,N_24864,N_21105);
or U29144 (N_29144,N_23105,N_23937);
xnor U29145 (N_29145,N_22297,N_20503);
nand U29146 (N_29146,N_23380,N_21218);
and U29147 (N_29147,N_22101,N_20032);
xor U29148 (N_29148,N_21195,N_24072);
or U29149 (N_29149,N_23837,N_23632);
or U29150 (N_29150,N_24411,N_20776);
nor U29151 (N_29151,N_24238,N_23260);
xor U29152 (N_29152,N_24326,N_23339);
nor U29153 (N_29153,N_22777,N_21613);
nand U29154 (N_29154,N_22121,N_23235);
nor U29155 (N_29155,N_22798,N_22752);
nor U29156 (N_29156,N_22062,N_23501);
xor U29157 (N_29157,N_21317,N_22736);
or U29158 (N_29158,N_22071,N_23340);
xnor U29159 (N_29159,N_22316,N_22211);
nand U29160 (N_29160,N_23324,N_22697);
and U29161 (N_29161,N_23397,N_20135);
or U29162 (N_29162,N_20131,N_23364);
nand U29163 (N_29163,N_21666,N_20463);
xor U29164 (N_29164,N_21011,N_21523);
nand U29165 (N_29165,N_23218,N_20167);
xor U29166 (N_29166,N_20930,N_21504);
and U29167 (N_29167,N_21921,N_22245);
nor U29168 (N_29168,N_24421,N_20389);
xnor U29169 (N_29169,N_21434,N_24292);
xnor U29170 (N_29170,N_24293,N_21045);
xor U29171 (N_29171,N_20054,N_21592);
xnor U29172 (N_29172,N_22289,N_20574);
nor U29173 (N_29173,N_24272,N_21521);
and U29174 (N_29174,N_23783,N_22342);
nand U29175 (N_29175,N_21378,N_21328);
or U29176 (N_29176,N_21235,N_20211);
nand U29177 (N_29177,N_23665,N_22394);
xor U29178 (N_29178,N_23448,N_23056);
nand U29179 (N_29179,N_21231,N_21405);
xnor U29180 (N_29180,N_23110,N_23055);
nand U29181 (N_29181,N_24342,N_20982);
nand U29182 (N_29182,N_21898,N_23179);
nor U29183 (N_29183,N_21351,N_20690);
nor U29184 (N_29184,N_21870,N_22204);
or U29185 (N_29185,N_21006,N_24212);
nand U29186 (N_29186,N_21787,N_23036);
xnor U29187 (N_29187,N_21628,N_24118);
or U29188 (N_29188,N_22006,N_23385);
xor U29189 (N_29189,N_21235,N_21696);
or U29190 (N_29190,N_22344,N_22411);
nor U29191 (N_29191,N_21464,N_22309);
or U29192 (N_29192,N_21862,N_24501);
or U29193 (N_29193,N_22341,N_21074);
or U29194 (N_29194,N_21095,N_23871);
nand U29195 (N_29195,N_21199,N_23131);
nand U29196 (N_29196,N_22879,N_21694);
xnor U29197 (N_29197,N_21223,N_24370);
or U29198 (N_29198,N_20672,N_24390);
nand U29199 (N_29199,N_24667,N_23857);
or U29200 (N_29200,N_20856,N_22327);
or U29201 (N_29201,N_23424,N_23902);
xor U29202 (N_29202,N_22901,N_22050);
nand U29203 (N_29203,N_21769,N_22920);
or U29204 (N_29204,N_24913,N_22673);
nor U29205 (N_29205,N_23103,N_23398);
and U29206 (N_29206,N_22000,N_21357);
nor U29207 (N_29207,N_22990,N_22723);
xor U29208 (N_29208,N_22675,N_21881);
and U29209 (N_29209,N_24816,N_20179);
and U29210 (N_29210,N_24871,N_23795);
nor U29211 (N_29211,N_22049,N_23493);
or U29212 (N_29212,N_22473,N_22021);
nor U29213 (N_29213,N_24356,N_22952);
or U29214 (N_29214,N_23303,N_22319);
nor U29215 (N_29215,N_24008,N_21823);
nor U29216 (N_29216,N_20235,N_21320);
xor U29217 (N_29217,N_20873,N_23362);
nor U29218 (N_29218,N_20079,N_23203);
nor U29219 (N_29219,N_21560,N_23527);
or U29220 (N_29220,N_23759,N_22649);
nor U29221 (N_29221,N_20039,N_24424);
xor U29222 (N_29222,N_20794,N_24705);
nor U29223 (N_29223,N_23957,N_20296);
xnor U29224 (N_29224,N_21956,N_23180);
nand U29225 (N_29225,N_23897,N_24309);
and U29226 (N_29226,N_23683,N_22498);
or U29227 (N_29227,N_23691,N_21963);
and U29228 (N_29228,N_22779,N_24821);
or U29229 (N_29229,N_22716,N_22290);
or U29230 (N_29230,N_23035,N_23877);
or U29231 (N_29231,N_22972,N_24391);
and U29232 (N_29232,N_21131,N_20931);
or U29233 (N_29233,N_24014,N_23543);
xnor U29234 (N_29234,N_24230,N_21838);
and U29235 (N_29235,N_20605,N_23360);
or U29236 (N_29236,N_23234,N_23590);
xor U29237 (N_29237,N_21129,N_20716);
nand U29238 (N_29238,N_21740,N_24253);
or U29239 (N_29239,N_23660,N_24831);
nor U29240 (N_29240,N_23623,N_21948);
nand U29241 (N_29241,N_21945,N_22638);
or U29242 (N_29242,N_21976,N_23316);
nor U29243 (N_29243,N_22323,N_24505);
and U29244 (N_29244,N_24338,N_20581);
xor U29245 (N_29245,N_21907,N_24406);
xnor U29246 (N_29246,N_24485,N_21222);
and U29247 (N_29247,N_23364,N_23618);
or U29248 (N_29248,N_24455,N_24493);
or U29249 (N_29249,N_23024,N_20772);
and U29250 (N_29250,N_20739,N_23946);
and U29251 (N_29251,N_20866,N_22922);
and U29252 (N_29252,N_24591,N_21801);
and U29253 (N_29253,N_24242,N_20853);
nor U29254 (N_29254,N_21103,N_21512);
or U29255 (N_29255,N_24218,N_22833);
and U29256 (N_29256,N_23468,N_20679);
and U29257 (N_29257,N_23337,N_23348);
or U29258 (N_29258,N_24712,N_23381);
xor U29259 (N_29259,N_22796,N_22898);
and U29260 (N_29260,N_20087,N_23707);
xor U29261 (N_29261,N_22593,N_23142);
nand U29262 (N_29262,N_21290,N_23273);
and U29263 (N_29263,N_21925,N_22112);
nor U29264 (N_29264,N_21830,N_21314);
xor U29265 (N_29265,N_23733,N_23832);
or U29266 (N_29266,N_24221,N_20777);
xnor U29267 (N_29267,N_21276,N_23744);
nand U29268 (N_29268,N_23857,N_20501);
and U29269 (N_29269,N_23743,N_22738);
nor U29270 (N_29270,N_20432,N_20352);
nand U29271 (N_29271,N_20291,N_23615);
nand U29272 (N_29272,N_23152,N_20170);
or U29273 (N_29273,N_23504,N_21281);
or U29274 (N_29274,N_20453,N_21515);
xnor U29275 (N_29275,N_20007,N_23233);
nor U29276 (N_29276,N_22796,N_22290);
or U29277 (N_29277,N_22716,N_20077);
xnor U29278 (N_29278,N_20809,N_22464);
xor U29279 (N_29279,N_24494,N_20585);
nand U29280 (N_29280,N_23286,N_23442);
xnor U29281 (N_29281,N_20589,N_21983);
and U29282 (N_29282,N_21680,N_24066);
xor U29283 (N_29283,N_21646,N_20244);
nor U29284 (N_29284,N_24419,N_21453);
nand U29285 (N_29285,N_23720,N_21396);
nand U29286 (N_29286,N_24100,N_22858);
nor U29287 (N_29287,N_20912,N_21681);
and U29288 (N_29288,N_23124,N_21488);
and U29289 (N_29289,N_23238,N_21976);
nand U29290 (N_29290,N_21751,N_23136);
xor U29291 (N_29291,N_24642,N_20374);
nor U29292 (N_29292,N_23261,N_21297);
and U29293 (N_29293,N_23474,N_22297);
nor U29294 (N_29294,N_24802,N_20126);
nand U29295 (N_29295,N_23402,N_21901);
or U29296 (N_29296,N_20268,N_23058);
nand U29297 (N_29297,N_22212,N_21522);
nor U29298 (N_29298,N_21653,N_21643);
nor U29299 (N_29299,N_24736,N_22120);
and U29300 (N_29300,N_24866,N_22556);
xor U29301 (N_29301,N_20324,N_22393);
or U29302 (N_29302,N_20327,N_24258);
nor U29303 (N_29303,N_20479,N_20844);
and U29304 (N_29304,N_20568,N_22103);
nor U29305 (N_29305,N_24379,N_22251);
nand U29306 (N_29306,N_23014,N_23043);
and U29307 (N_29307,N_22171,N_22461);
nand U29308 (N_29308,N_20867,N_22228);
xor U29309 (N_29309,N_22594,N_21074);
nor U29310 (N_29310,N_22092,N_23790);
and U29311 (N_29311,N_24119,N_20817);
nor U29312 (N_29312,N_22219,N_23746);
or U29313 (N_29313,N_24769,N_21733);
nor U29314 (N_29314,N_23381,N_20157);
nand U29315 (N_29315,N_21152,N_24847);
nor U29316 (N_29316,N_22325,N_20948);
and U29317 (N_29317,N_23728,N_22248);
or U29318 (N_29318,N_24865,N_23022);
nor U29319 (N_29319,N_23902,N_21113);
nor U29320 (N_29320,N_24425,N_23584);
and U29321 (N_29321,N_23013,N_20659);
nand U29322 (N_29322,N_23850,N_24118);
or U29323 (N_29323,N_24242,N_22500);
nand U29324 (N_29324,N_21113,N_24261);
nand U29325 (N_29325,N_24732,N_20504);
xnor U29326 (N_29326,N_22572,N_22206);
nand U29327 (N_29327,N_24402,N_20346);
nor U29328 (N_29328,N_24160,N_22218);
nor U29329 (N_29329,N_22253,N_24270);
and U29330 (N_29330,N_21167,N_21440);
nor U29331 (N_29331,N_23375,N_24033);
nor U29332 (N_29332,N_20635,N_22119);
or U29333 (N_29333,N_23311,N_24202);
nor U29334 (N_29334,N_22737,N_23076);
nor U29335 (N_29335,N_23018,N_23684);
nor U29336 (N_29336,N_21294,N_22268);
nand U29337 (N_29337,N_22427,N_21667);
nand U29338 (N_29338,N_20581,N_23004);
nor U29339 (N_29339,N_24900,N_21467);
or U29340 (N_29340,N_20102,N_21825);
and U29341 (N_29341,N_22916,N_20664);
nor U29342 (N_29342,N_21867,N_22760);
nor U29343 (N_29343,N_23175,N_23484);
nor U29344 (N_29344,N_22849,N_23235);
nor U29345 (N_29345,N_22182,N_22540);
or U29346 (N_29346,N_23687,N_22029);
or U29347 (N_29347,N_24999,N_23014);
xor U29348 (N_29348,N_23756,N_24403);
and U29349 (N_29349,N_22091,N_20489);
and U29350 (N_29350,N_22082,N_23778);
xnor U29351 (N_29351,N_21081,N_21624);
nor U29352 (N_29352,N_20745,N_23027);
nand U29353 (N_29353,N_23645,N_22138);
or U29354 (N_29354,N_21641,N_23191);
xnor U29355 (N_29355,N_24912,N_23812);
nor U29356 (N_29356,N_22941,N_22711);
nand U29357 (N_29357,N_24962,N_20846);
and U29358 (N_29358,N_22415,N_23728);
or U29359 (N_29359,N_20986,N_23332);
nor U29360 (N_29360,N_21023,N_23741);
nor U29361 (N_29361,N_22214,N_24400);
and U29362 (N_29362,N_21104,N_23389);
or U29363 (N_29363,N_23303,N_21048);
nand U29364 (N_29364,N_24826,N_22910);
nor U29365 (N_29365,N_23334,N_21587);
nor U29366 (N_29366,N_23371,N_23993);
and U29367 (N_29367,N_24116,N_23847);
xor U29368 (N_29368,N_23141,N_22518);
xor U29369 (N_29369,N_23982,N_24908);
and U29370 (N_29370,N_20194,N_24883);
or U29371 (N_29371,N_22575,N_20917);
and U29372 (N_29372,N_22109,N_23258);
and U29373 (N_29373,N_24760,N_22612);
xor U29374 (N_29374,N_22806,N_21308);
or U29375 (N_29375,N_21496,N_22459);
nand U29376 (N_29376,N_24612,N_22834);
xnor U29377 (N_29377,N_20866,N_22298);
xnor U29378 (N_29378,N_20128,N_24676);
nand U29379 (N_29379,N_21981,N_23927);
or U29380 (N_29380,N_24237,N_21079);
xor U29381 (N_29381,N_21265,N_24313);
and U29382 (N_29382,N_24087,N_20870);
xnor U29383 (N_29383,N_20530,N_21238);
and U29384 (N_29384,N_20414,N_21916);
xnor U29385 (N_29385,N_22547,N_24250);
or U29386 (N_29386,N_23951,N_23059);
nor U29387 (N_29387,N_22143,N_23109);
or U29388 (N_29388,N_20451,N_24585);
nor U29389 (N_29389,N_20748,N_23270);
nor U29390 (N_29390,N_24870,N_23814);
xnor U29391 (N_29391,N_23320,N_23334);
and U29392 (N_29392,N_22201,N_24685);
nand U29393 (N_29393,N_20259,N_22341);
and U29394 (N_29394,N_20478,N_21197);
xnor U29395 (N_29395,N_22029,N_20774);
nor U29396 (N_29396,N_22351,N_20039);
nor U29397 (N_29397,N_21479,N_20317);
or U29398 (N_29398,N_24445,N_23299);
nand U29399 (N_29399,N_22995,N_21709);
nor U29400 (N_29400,N_23018,N_23563);
or U29401 (N_29401,N_22982,N_24504);
and U29402 (N_29402,N_24595,N_21214);
nor U29403 (N_29403,N_22950,N_22499);
or U29404 (N_29404,N_22749,N_21201);
xor U29405 (N_29405,N_24246,N_24666);
nor U29406 (N_29406,N_23282,N_23868);
or U29407 (N_29407,N_24529,N_21517);
and U29408 (N_29408,N_21379,N_22484);
nor U29409 (N_29409,N_24415,N_24756);
and U29410 (N_29410,N_24103,N_24236);
and U29411 (N_29411,N_21841,N_24487);
nand U29412 (N_29412,N_21817,N_21465);
and U29413 (N_29413,N_23517,N_20614);
nand U29414 (N_29414,N_21410,N_24583);
xor U29415 (N_29415,N_21459,N_24027);
nand U29416 (N_29416,N_21968,N_24542);
nand U29417 (N_29417,N_20802,N_23586);
nor U29418 (N_29418,N_20185,N_22014);
or U29419 (N_29419,N_22704,N_23026);
and U29420 (N_29420,N_24653,N_21451);
nand U29421 (N_29421,N_23826,N_24430);
nor U29422 (N_29422,N_20793,N_24021);
and U29423 (N_29423,N_24519,N_21499);
nor U29424 (N_29424,N_21167,N_21556);
and U29425 (N_29425,N_23620,N_23227);
and U29426 (N_29426,N_20893,N_23102);
nand U29427 (N_29427,N_20156,N_22130);
nand U29428 (N_29428,N_21573,N_21232);
and U29429 (N_29429,N_24079,N_23580);
or U29430 (N_29430,N_20045,N_20916);
nand U29431 (N_29431,N_20524,N_21491);
nor U29432 (N_29432,N_20952,N_21251);
and U29433 (N_29433,N_24418,N_23249);
nand U29434 (N_29434,N_23008,N_21871);
nand U29435 (N_29435,N_20674,N_23342);
nand U29436 (N_29436,N_20144,N_22219);
xor U29437 (N_29437,N_23967,N_24934);
nand U29438 (N_29438,N_23239,N_24591);
nor U29439 (N_29439,N_21835,N_20287);
or U29440 (N_29440,N_21373,N_22725);
xnor U29441 (N_29441,N_24120,N_20360);
or U29442 (N_29442,N_24386,N_22640);
xor U29443 (N_29443,N_23524,N_22704);
nor U29444 (N_29444,N_21928,N_24337);
xor U29445 (N_29445,N_23808,N_20575);
nand U29446 (N_29446,N_23454,N_23325);
and U29447 (N_29447,N_20680,N_24908);
xnor U29448 (N_29448,N_21709,N_21038);
nor U29449 (N_29449,N_21211,N_21119);
and U29450 (N_29450,N_23694,N_20959);
and U29451 (N_29451,N_22518,N_20382);
xor U29452 (N_29452,N_23681,N_22954);
nand U29453 (N_29453,N_21766,N_21556);
nand U29454 (N_29454,N_20555,N_20735);
xor U29455 (N_29455,N_21487,N_24070);
or U29456 (N_29456,N_21653,N_22312);
or U29457 (N_29457,N_21294,N_23345);
and U29458 (N_29458,N_20429,N_22701);
nor U29459 (N_29459,N_24534,N_21960);
and U29460 (N_29460,N_23754,N_20856);
or U29461 (N_29461,N_21157,N_21286);
nand U29462 (N_29462,N_22067,N_21935);
nand U29463 (N_29463,N_22457,N_21359);
xor U29464 (N_29464,N_20638,N_21078);
and U29465 (N_29465,N_23630,N_20065);
and U29466 (N_29466,N_22500,N_22405);
nand U29467 (N_29467,N_22295,N_21770);
nand U29468 (N_29468,N_23685,N_23321);
or U29469 (N_29469,N_23371,N_22344);
and U29470 (N_29470,N_23898,N_24927);
or U29471 (N_29471,N_23800,N_20299);
or U29472 (N_29472,N_23977,N_23991);
nand U29473 (N_29473,N_20016,N_22513);
xor U29474 (N_29474,N_24280,N_22396);
nor U29475 (N_29475,N_21544,N_22673);
and U29476 (N_29476,N_21256,N_23731);
xnor U29477 (N_29477,N_20234,N_22487);
nor U29478 (N_29478,N_22426,N_23326);
or U29479 (N_29479,N_22008,N_22388);
or U29480 (N_29480,N_20945,N_21865);
nand U29481 (N_29481,N_23788,N_20604);
nand U29482 (N_29482,N_24161,N_24691);
or U29483 (N_29483,N_20400,N_20391);
or U29484 (N_29484,N_24056,N_23688);
nand U29485 (N_29485,N_20435,N_21880);
nand U29486 (N_29486,N_23039,N_21080);
nor U29487 (N_29487,N_23728,N_21946);
and U29488 (N_29488,N_22157,N_24721);
or U29489 (N_29489,N_22935,N_23220);
and U29490 (N_29490,N_24990,N_23281);
or U29491 (N_29491,N_24447,N_23015);
xor U29492 (N_29492,N_20809,N_23701);
nor U29493 (N_29493,N_23099,N_23561);
xor U29494 (N_29494,N_22008,N_24443);
and U29495 (N_29495,N_21878,N_22076);
nor U29496 (N_29496,N_24449,N_20396);
nand U29497 (N_29497,N_21794,N_24132);
xnor U29498 (N_29498,N_23086,N_22118);
or U29499 (N_29499,N_21847,N_20675);
or U29500 (N_29500,N_20581,N_20630);
nand U29501 (N_29501,N_24454,N_21419);
xor U29502 (N_29502,N_22935,N_21006);
or U29503 (N_29503,N_20929,N_22484);
nand U29504 (N_29504,N_24273,N_21262);
or U29505 (N_29505,N_20666,N_20423);
nor U29506 (N_29506,N_20428,N_22519);
nor U29507 (N_29507,N_20508,N_20665);
xnor U29508 (N_29508,N_22684,N_22564);
nor U29509 (N_29509,N_22840,N_21016);
xor U29510 (N_29510,N_20727,N_20622);
and U29511 (N_29511,N_21556,N_21715);
or U29512 (N_29512,N_24323,N_21746);
nor U29513 (N_29513,N_21336,N_21354);
xor U29514 (N_29514,N_22404,N_21606);
and U29515 (N_29515,N_23602,N_24837);
xnor U29516 (N_29516,N_21523,N_20775);
xnor U29517 (N_29517,N_21051,N_21217);
xnor U29518 (N_29518,N_20775,N_20448);
nand U29519 (N_29519,N_23425,N_20158);
xor U29520 (N_29520,N_23446,N_20871);
and U29521 (N_29521,N_20861,N_22710);
nor U29522 (N_29522,N_21689,N_24126);
nor U29523 (N_29523,N_21245,N_23904);
and U29524 (N_29524,N_20088,N_24651);
nor U29525 (N_29525,N_24700,N_20744);
nand U29526 (N_29526,N_24752,N_22161);
xnor U29527 (N_29527,N_22709,N_20926);
xor U29528 (N_29528,N_20225,N_22698);
or U29529 (N_29529,N_24696,N_20206);
and U29530 (N_29530,N_20255,N_22428);
xor U29531 (N_29531,N_20417,N_22638);
nor U29532 (N_29532,N_21368,N_23392);
xor U29533 (N_29533,N_21290,N_20873);
xor U29534 (N_29534,N_22294,N_23334);
nor U29535 (N_29535,N_24860,N_21357);
or U29536 (N_29536,N_21855,N_20307);
or U29537 (N_29537,N_23766,N_20703);
nor U29538 (N_29538,N_20580,N_22212);
nor U29539 (N_29539,N_20323,N_24362);
nand U29540 (N_29540,N_21143,N_22226);
nor U29541 (N_29541,N_22599,N_24739);
and U29542 (N_29542,N_23222,N_24607);
or U29543 (N_29543,N_20982,N_23105);
and U29544 (N_29544,N_21510,N_24035);
xnor U29545 (N_29545,N_22083,N_20938);
and U29546 (N_29546,N_22356,N_21635);
xnor U29547 (N_29547,N_20366,N_23135);
or U29548 (N_29548,N_22496,N_24363);
nor U29549 (N_29549,N_22468,N_22937);
xor U29550 (N_29550,N_21437,N_20793);
or U29551 (N_29551,N_24743,N_24719);
and U29552 (N_29552,N_23657,N_20431);
nand U29553 (N_29553,N_22307,N_21834);
nor U29554 (N_29554,N_24985,N_20398);
or U29555 (N_29555,N_22813,N_21610);
xor U29556 (N_29556,N_21378,N_23755);
xnor U29557 (N_29557,N_21718,N_21702);
xor U29558 (N_29558,N_24969,N_21224);
or U29559 (N_29559,N_24585,N_22094);
xnor U29560 (N_29560,N_20557,N_23453);
nor U29561 (N_29561,N_23787,N_22810);
xnor U29562 (N_29562,N_23688,N_23279);
nor U29563 (N_29563,N_22080,N_21107);
xor U29564 (N_29564,N_21515,N_22924);
nor U29565 (N_29565,N_20359,N_24639);
nand U29566 (N_29566,N_24475,N_23956);
and U29567 (N_29567,N_22651,N_23328);
or U29568 (N_29568,N_24396,N_22556);
nand U29569 (N_29569,N_21443,N_22579);
nor U29570 (N_29570,N_20516,N_22457);
or U29571 (N_29571,N_23054,N_20572);
xor U29572 (N_29572,N_21248,N_24218);
nor U29573 (N_29573,N_22020,N_20568);
nand U29574 (N_29574,N_22934,N_23208);
xor U29575 (N_29575,N_23353,N_21904);
nand U29576 (N_29576,N_21719,N_23200);
and U29577 (N_29577,N_22626,N_24238);
and U29578 (N_29578,N_20751,N_23986);
nor U29579 (N_29579,N_23586,N_24056);
nor U29580 (N_29580,N_22102,N_23139);
nor U29581 (N_29581,N_22318,N_23554);
xnor U29582 (N_29582,N_24309,N_24282);
nand U29583 (N_29583,N_22421,N_20869);
nor U29584 (N_29584,N_24908,N_23154);
nor U29585 (N_29585,N_24362,N_24837);
xnor U29586 (N_29586,N_20066,N_20985);
nand U29587 (N_29587,N_23161,N_21066);
or U29588 (N_29588,N_20153,N_21582);
nor U29589 (N_29589,N_22501,N_24311);
xnor U29590 (N_29590,N_22478,N_21985);
and U29591 (N_29591,N_21892,N_24080);
nand U29592 (N_29592,N_24122,N_23423);
and U29593 (N_29593,N_20543,N_23361);
or U29594 (N_29594,N_24007,N_23918);
nand U29595 (N_29595,N_20753,N_20166);
or U29596 (N_29596,N_20697,N_20100);
and U29597 (N_29597,N_22510,N_20245);
nor U29598 (N_29598,N_20588,N_22311);
nor U29599 (N_29599,N_23597,N_21671);
or U29600 (N_29600,N_23190,N_22082);
nand U29601 (N_29601,N_23096,N_21316);
xor U29602 (N_29602,N_20102,N_21613);
nand U29603 (N_29603,N_24714,N_20776);
nand U29604 (N_29604,N_24797,N_22982);
nor U29605 (N_29605,N_22364,N_24919);
or U29606 (N_29606,N_24513,N_24431);
and U29607 (N_29607,N_20398,N_22191);
nand U29608 (N_29608,N_22256,N_21673);
and U29609 (N_29609,N_20642,N_21086);
nor U29610 (N_29610,N_21592,N_24557);
or U29611 (N_29611,N_22603,N_23787);
and U29612 (N_29612,N_21367,N_21621);
and U29613 (N_29613,N_22612,N_20253);
nor U29614 (N_29614,N_22347,N_24971);
xor U29615 (N_29615,N_21303,N_22945);
or U29616 (N_29616,N_23699,N_24425);
nor U29617 (N_29617,N_21688,N_22035);
nor U29618 (N_29618,N_24224,N_20070);
xnor U29619 (N_29619,N_22340,N_24914);
nand U29620 (N_29620,N_20254,N_23473);
or U29621 (N_29621,N_20587,N_21002);
nor U29622 (N_29622,N_22686,N_24596);
nand U29623 (N_29623,N_20463,N_24561);
nor U29624 (N_29624,N_24542,N_24130);
xnor U29625 (N_29625,N_22944,N_20953);
or U29626 (N_29626,N_22104,N_20274);
and U29627 (N_29627,N_20587,N_20553);
nor U29628 (N_29628,N_20104,N_23938);
nand U29629 (N_29629,N_20230,N_24242);
and U29630 (N_29630,N_21821,N_24074);
and U29631 (N_29631,N_23847,N_24792);
and U29632 (N_29632,N_23872,N_23212);
nor U29633 (N_29633,N_23790,N_23886);
xnor U29634 (N_29634,N_22730,N_24512);
or U29635 (N_29635,N_21999,N_24105);
nor U29636 (N_29636,N_22101,N_22670);
xor U29637 (N_29637,N_21806,N_23194);
or U29638 (N_29638,N_20262,N_23561);
xnor U29639 (N_29639,N_22552,N_21306);
and U29640 (N_29640,N_21498,N_21829);
xnor U29641 (N_29641,N_23562,N_21564);
or U29642 (N_29642,N_22439,N_20163);
nand U29643 (N_29643,N_21519,N_23187);
xor U29644 (N_29644,N_22213,N_21499);
or U29645 (N_29645,N_24643,N_24519);
nand U29646 (N_29646,N_23154,N_20692);
nor U29647 (N_29647,N_21458,N_21395);
and U29648 (N_29648,N_20806,N_23476);
and U29649 (N_29649,N_20445,N_23612);
nor U29650 (N_29650,N_21725,N_23459);
nor U29651 (N_29651,N_20252,N_23496);
nor U29652 (N_29652,N_23978,N_21944);
or U29653 (N_29653,N_23219,N_23367);
nor U29654 (N_29654,N_23096,N_23598);
xnor U29655 (N_29655,N_22807,N_23366);
nor U29656 (N_29656,N_20817,N_21347);
nand U29657 (N_29657,N_20785,N_24157);
nor U29658 (N_29658,N_24988,N_21088);
nand U29659 (N_29659,N_22467,N_22706);
nand U29660 (N_29660,N_23107,N_21329);
nor U29661 (N_29661,N_22079,N_20255);
nor U29662 (N_29662,N_22816,N_24417);
and U29663 (N_29663,N_23717,N_20775);
and U29664 (N_29664,N_24336,N_23151);
or U29665 (N_29665,N_21271,N_22429);
nand U29666 (N_29666,N_22927,N_20859);
and U29667 (N_29667,N_21917,N_21101);
nor U29668 (N_29668,N_23036,N_24309);
nor U29669 (N_29669,N_20996,N_24623);
or U29670 (N_29670,N_24566,N_24938);
nor U29671 (N_29671,N_20433,N_21604);
and U29672 (N_29672,N_24791,N_21594);
nand U29673 (N_29673,N_24164,N_22451);
nand U29674 (N_29674,N_24610,N_24371);
nand U29675 (N_29675,N_24272,N_22013);
or U29676 (N_29676,N_22399,N_21924);
and U29677 (N_29677,N_22121,N_20276);
nand U29678 (N_29678,N_24918,N_24201);
nand U29679 (N_29679,N_24135,N_23052);
nor U29680 (N_29680,N_21569,N_24265);
nand U29681 (N_29681,N_24194,N_23277);
and U29682 (N_29682,N_22147,N_24890);
or U29683 (N_29683,N_23843,N_21328);
or U29684 (N_29684,N_24190,N_20776);
xor U29685 (N_29685,N_21211,N_22022);
nor U29686 (N_29686,N_24868,N_20820);
xor U29687 (N_29687,N_21930,N_22733);
or U29688 (N_29688,N_24879,N_20320);
or U29689 (N_29689,N_22530,N_21993);
nor U29690 (N_29690,N_20762,N_21523);
nand U29691 (N_29691,N_24758,N_21859);
xnor U29692 (N_29692,N_21629,N_23216);
xor U29693 (N_29693,N_24487,N_20949);
and U29694 (N_29694,N_24311,N_20203);
xor U29695 (N_29695,N_24138,N_24931);
nor U29696 (N_29696,N_23413,N_20294);
and U29697 (N_29697,N_23307,N_23430);
nand U29698 (N_29698,N_22985,N_23280);
nand U29699 (N_29699,N_21913,N_23729);
or U29700 (N_29700,N_22052,N_23782);
or U29701 (N_29701,N_24182,N_20671);
and U29702 (N_29702,N_20885,N_21439);
nor U29703 (N_29703,N_21754,N_22074);
nor U29704 (N_29704,N_22951,N_24661);
nor U29705 (N_29705,N_24392,N_23039);
nand U29706 (N_29706,N_24012,N_20019);
nand U29707 (N_29707,N_22531,N_24104);
nand U29708 (N_29708,N_23807,N_23655);
nor U29709 (N_29709,N_24656,N_20960);
xor U29710 (N_29710,N_24992,N_22054);
nand U29711 (N_29711,N_24280,N_23949);
nor U29712 (N_29712,N_24257,N_21119);
nand U29713 (N_29713,N_23067,N_24168);
nand U29714 (N_29714,N_24280,N_20484);
or U29715 (N_29715,N_20079,N_22128);
xor U29716 (N_29716,N_24033,N_24402);
and U29717 (N_29717,N_24245,N_24913);
nor U29718 (N_29718,N_21830,N_23984);
nand U29719 (N_29719,N_22045,N_22819);
nand U29720 (N_29720,N_22828,N_21772);
and U29721 (N_29721,N_24822,N_20366);
nand U29722 (N_29722,N_22508,N_24419);
nor U29723 (N_29723,N_24488,N_21871);
nand U29724 (N_29724,N_21240,N_23292);
nand U29725 (N_29725,N_24337,N_22524);
nor U29726 (N_29726,N_20185,N_23450);
xor U29727 (N_29727,N_24556,N_22850);
nor U29728 (N_29728,N_20987,N_24439);
nor U29729 (N_29729,N_22056,N_24838);
or U29730 (N_29730,N_21573,N_21248);
nor U29731 (N_29731,N_24530,N_20667);
or U29732 (N_29732,N_23482,N_22622);
nor U29733 (N_29733,N_21325,N_20047);
nand U29734 (N_29734,N_20731,N_24033);
nand U29735 (N_29735,N_22524,N_24455);
xor U29736 (N_29736,N_23617,N_21496);
nand U29737 (N_29737,N_24251,N_20886);
nand U29738 (N_29738,N_21645,N_22796);
and U29739 (N_29739,N_24543,N_23382);
or U29740 (N_29740,N_21737,N_23186);
or U29741 (N_29741,N_20004,N_23568);
and U29742 (N_29742,N_22082,N_24798);
nor U29743 (N_29743,N_24071,N_22717);
or U29744 (N_29744,N_20232,N_23176);
nand U29745 (N_29745,N_21218,N_24387);
xnor U29746 (N_29746,N_24461,N_23238);
and U29747 (N_29747,N_23769,N_22761);
and U29748 (N_29748,N_20926,N_23793);
and U29749 (N_29749,N_23265,N_21136);
nor U29750 (N_29750,N_24265,N_20585);
nand U29751 (N_29751,N_21343,N_21587);
nand U29752 (N_29752,N_24314,N_20774);
xnor U29753 (N_29753,N_22263,N_22232);
or U29754 (N_29754,N_22643,N_20572);
and U29755 (N_29755,N_23589,N_21442);
nand U29756 (N_29756,N_24972,N_24924);
and U29757 (N_29757,N_24001,N_20996);
xnor U29758 (N_29758,N_20309,N_21387);
and U29759 (N_29759,N_23316,N_22522);
or U29760 (N_29760,N_21329,N_24175);
xnor U29761 (N_29761,N_20984,N_24085);
and U29762 (N_29762,N_23948,N_21981);
nand U29763 (N_29763,N_21430,N_21491);
and U29764 (N_29764,N_23939,N_21644);
and U29765 (N_29765,N_24446,N_21185);
or U29766 (N_29766,N_21688,N_23054);
nor U29767 (N_29767,N_24546,N_24804);
or U29768 (N_29768,N_23905,N_24096);
or U29769 (N_29769,N_21733,N_20899);
and U29770 (N_29770,N_24981,N_22889);
nor U29771 (N_29771,N_20897,N_23286);
xor U29772 (N_29772,N_24872,N_24346);
and U29773 (N_29773,N_21315,N_22373);
and U29774 (N_29774,N_22957,N_20220);
nand U29775 (N_29775,N_20753,N_24929);
and U29776 (N_29776,N_22671,N_23851);
xnor U29777 (N_29777,N_24656,N_22038);
or U29778 (N_29778,N_21432,N_22445);
and U29779 (N_29779,N_23005,N_23873);
and U29780 (N_29780,N_24586,N_22161);
xnor U29781 (N_29781,N_21958,N_23164);
nor U29782 (N_29782,N_23976,N_20936);
nor U29783 (N_29783,N_21830,N_22211);
nor U29784 (N_29784,N_22629,N_24400);
and U29785 (N_29785,N_21604,N_24356);
nor U29786 (N_29786,N_21652,N_23461);
xor U29787 (N_29787,N_20697,N_24872);
or U29788 (N_29788,N_20844,N_22278);
xnor U29789 (N_29789,N_23254,N_20395);
nor U29790 (N_29790,N_21386,N_21039);
xnor U29791 (N_29791,N_21866,N_23610);
xor U29792 (N_29792,N_20854,N_20990);
and U29793 (N_29793,N_21126,N_24059);
xor U29794 (N_29794,N_23532,N_23795);
xnor U29795 (N_29795,N_24356,N_24523);
and U29796 (N_29796,N_23789,N_22768);
and U29797 (N_29797,N_20344,N_24234);
or U29798 (N_29798,N_23488,N_24827);
and U29799 (N_29799,N_20381,N_22332);
nand U29800 (N_29800,N_22419,N_21726);
nand U29801 (N_29801,N_21329,N_22493);
or U29802 (N_29802,N_20201,N_24885);
nand U29803 (N_29803,N_23778,N_22265);
nand U29804 (N_29804,N_23604,N_21454);
nor U29805 (N_29805,N_20055,N_20573);
nor U29806 (N_29806,N_22404,N_21091);
or U29807 (N_29807,N_23831,N_24435);
or U29808 (N_29808,N_22615,N_20725);
and U29809 (N_29809,N_20279,N_20396);
xnor U29810 (N_29810,N_23594,N_20351);
or U29811 (N_29811,N_24092,N_23737);
or U29812 (N_29812,N_23373,N_22748);
nand U29813 (N_29813,N_20467,N_21537);
nand U29814 (N_29814,N_23650,N_23834);
or U29815 (N_29815,N_22110,N_23019);
and U29816 (N_29816,N_24119,N_24192);
nor U29817 (N_29817,N_20047,N_23387);
nand U29818 (N_29818,N_24406,N_20051);
nand U29819 (N_29819,N_21058,N_23230);
xor U29820 (N_29820,N_22299,N_22353);
nand U29821 (N_29821,N_22139,N_20137);
or U29822 (N_29822,N_21349,N_20138);
or U29823 (N_29823,N_22665,N_23577);
and U29824 (N_29824,N_21641,N_24198);
nand U29825 (N_29825,N_20602,N_22923);
or U29826 (N_29826,N_23151,N_21560);
or U29827 (N_29827,N_21891,N_23502);
or U29828 (N_29828,N_23615,N_21091);
xnor U29829 (N_29829,N_21218,N_24388);
and U29830 (N_29830,N_23891,N_24485);
nor U29831 (N_29831,N_21181,N_20045);
xor U29832 (N_29832,N_22524,N_22439);
xnor U29833 (N_29833,N_22305,N_20133);
nand U29834 (N_29834,N_22205,N_22055);
nand U29835 (N_29835,N_23100,N_21472);
and U29836 (N_29836,N_24951,N_23605);
xnor U29837 (N_29837,N_24134,N_23798);
xor U29838 (N_29838,N_21002,N_20819);
or U29839 (N_29839,N_22440,N_22557);
or U29840 (N_29840,N_22467,N_21384);
and U29841 (N_29841,N_20535,N_23097);
xor U29842 (N_29842,N_22370,N_22196);
and U29843 (N_29843,N_21871,N_23612);
and U29844 (N_29844,N_20080,N_20142);
nor U29845 (N_29845,N_23942,N_22483);
or U29846 (N_29846,N_20088,N_22146);
and U29847 (N_29847,N_24458,N_21652);
nand U29848 (N_29848,N_22658,N_22044);
nor U29849 (N_29849,N_23861,N_22017);
and U29850 (N_29850,N_21644,N_20827);
nor U29851 (N_29851,N_23874,N_21195);
or U29852 (N_29852,N_22069,N_23939);
nor U29853 (N_29853,N_21496,N_21153);
or U29854 (N_29854,N_20094,N_22746);
xnor U29855 (N_29855,N_23582,N_23419);
and U29856 (N_29856,N_20736,N_20891);
nor U29857 (N_29857,N_24868,N_24269);
nor U29858 (N_29858,N_20824,N_22144);
nand U29859 (N_29859,N_22490,N_21975);
and U29860 (N_29860,N_23536,N_22612);
and U29861 (N_29861,N_24946,N_22498);
nor U29862 (N_29862,N_23629,N_21633);
nand U29863 (N_29863,N_23795,N_24891);
xor U29864 (N_29864,N_24848,N_21576);
and U29865 (N_29865,N_20338,N_20209);
nor U29866 (N_29866,N_20517,N_22801);
nor U29867 (N_29867,N_21945,N_23868);
xor U29868 (N_29868,N_23764,N_21895);
nand U29869 (N_29869,N_22497,N_24491);
or U29870 (N_29870,N_20126,N_23082);
nor U29871 (N_29871,N_22203,N_22010);
or U29872 (N_29872,N_24011,N_24326);
xor U29873 (N_29873,N_20209,N_22422);
or U29874 (N_29874,N_21111,N_22265);
or U29875 (N_29875,N_22444,N_21748);
nand U29876 (N_29876,N_20151,N_22911);
nand U29877 (N_29877,N_23300,N_24016);
or U29878 (N_29878,N_22689,N_22939);
and U29879 (N_29879,N_21625,N_24499);
or U29880 (N_29880,N_24798,N_21204);
nor U29881 (N_29881,N_23435,N_20739);
nor U29882 (N_29882,N_24819,N_23517);
and U29883 (N_29883,N_24325,N_20962);
or U29884 (N_29884,N_22111,N_24520);
nand U29885 (N_29885,N_23721,N_21646);
nand U29886 (N_29886,N_20059,N_20160);
xnor U29887 (N_29887,N_20826,N_20231);
or U29888 (N_29888,N_21035,N_22819);
or U29889 (N_29889,N_24500,N_22187);
or U29890 (N_29890,N_22262,N_22035);
nand U29891 (N_29891,N_21940,N_20155);
nor U29892 (N_29892,N_24455,N_20926);
and U29893 (N_29893,N_24005,N_20589);
nor U29894 (N_29894,N_23084,N_21622);
and U29895 (N_29895,N_21812,N_22289);
and U29896 (N_29896,N_22976,N_22841);
xnor U29897 (N_29897,N_22007,N_24262);
or U29898 (N_29898,N_22792,N_23134);
xor U29899 (N_29899,N_21617,N_20014);
nor U29900 (N_29900,N_21290,N_21804);
nand U29901 (N_29901,N_22835,N_22135);
nand U29902 (N_29902,N_22761,N_21332);
or U29903 (N_29903,N_21615,N_24792);
or U29904 (N_29904,N_23714,N_21621);
xor U29905 (N_29905,N_20473,N_22815);
nor U29906 (N_29906,N_20806,N_23802);
nand U29907 (N_29907,N_21599,N_22806);
xor U29908 (N_29908,N_24046,N_21804);
nor U29909 (N_29909,N_22514,N_20383);
or U29910 (N_29910,N_24806,N_21260);
nor U29911 (N_29911,N_22628,N_23455);
nor U29912 (N_29912,N_24678,N_20924);
xnor U29913 (N_29913,N_24746,N_23455);
nor U29914 (N_29914,N_22468,N_21437);
xnor U29915 (N_29915,N_20472,N_22917);
xnor U29916 (N_29916,N_20630,N_20714);
nor U29917 (N_29917,N_20880,N_21176);
or U29918 (N_29918,N_22319,N_24966);
or U29919 (N_29919,N_21743,N_21493);
or U29920 (N_29920,N_22036,N_22392);
nand U29921 (N_29921,N_23836,N_21228);
nor U29922 (N_29922,N_24563,N_23381);
or U29923 (N_29923,N_21701,N_23660);
xor U29924 (N_29924,N_22624,N_23022);
and U29925 (N_29925,N_22423,N_23730);
or U29926 (N_29926,N_24324,N_21375);
nor U29927 (N_29927,N_22545,N_24968);
nand U29928 (N_29928,N_20839,N_22977);
xnor U29929 (N_29929,N_24668,N_20957);
nand U29930 (N_29930,N_22152,N_21591);
nand U29931 (N_29931,N_20681,N_21624);
nand U29932 (N_29932,N_21629,N_23903);
and U29933 (N_29933,N_21337,N_24727);
or U29934 (N_29934,N_24589,N_23413);
nor U29935 (N_29935,N_22872,N_23730);
nand U29936 (N_29936,N_24119,N_21817);
or U29937 (N_29937,N_24571,N_23580);
or U29938 (N_29938,N_21620,N_21084);
nand U29939 (N_29939,N_20973,N_24601);
nor U29940 (N_29940,N_20535,N_24428);
or U29941 (N_29941,N_22557,N_22050);
nand U29942 (N_29942,N_23695,N_24236);
or U29943 (N_29943,N_20105,N_23741);
or U29944 (N_29944,N_20072,N_22871);
or U29945 (N_29945,N_20978,N_23009);
nor U29946 (N_29946,N_20367,N_24996);
nor U29947 (N_29947,N_22833,N_24162);
nor U29948 (N_29948,N_22059,N_23230);
or U29949 (N_29949,N_23941,N_22060);
or U29950 (N_29950,N_22102,N_23398);
or U29951 (N_29951,N_20230,N_21074);
or U29952 (N_29952,N_22190,N_24916);
and U29953 (N_29953,N_24454,N_23866);
nand U29954 (N_29954,N_21340,N_20367);
nand U29955 (N_29955,N_23371,N_20708);
or U29956 (N_29956,N_21940,N_21147);
xnor U29957 (N_29957,N_23790,N_21096);
or U29958 (N_29958,N_23375,N_23964);
nand U29959 (N_29959,N_20965,N_24418);
nor U29960 (N_29960,N_24484,N_22065);
or U29961 (N_29961,N_24898,N_21724);
or U29962 (N_29962,N_22906,N_20869);
and U29963 (N_29963,N_22751,N_22180);
and U29964 (N_29964,N_23055,N_24059);
and U29965 (N_29965,N_24934,N_22809);
nor U29966 (N_29966,N_20741,N_23067);
xor U29967 (N_29967,N_24274,N_20452);
or U29968 (N_29968,N_24592,N_23260);
nor U29969 (N_29969,N_24528,N_21137);
nand U29970 (N_29970,N_20294,N_22091);
or U29971 (N_29971,N_22527,N_21730);
or U29972 (N_29972,N_23268,N_22482);
nand U29973 (N_29973,N_21944,N_21675);
nor U29974 (N_29974,N_20652,N_20779);
or U29975 (N_29975,N_24712,N_22818);
or U29976 (N_29976,N_20037,N_20755);
and U29977 (N_29977,N_22090,N_24211);
and U29978 (N_29978,N_22815,N_20893);
or U29979 (N_29979,N_23266,N_24657);
or U29980 (N_29980,N_21097,N_23462);
and U29981 (N_29981,N_21350,N_22093);
or U29982 (N_29982,N_23696,N_24271);
xor U29983 (N_29983,N_20486,N_21249);
xor U29984 (N_29984,N_23813,N_23944);
nand U29985 (N_29985,N_23106,N_22007);
xor U29986 (N_29986,N_22891,N_22775);
xor U29987 (N_29987,N_20287,N_22975);
nor U29988 (N_29988,N_20037,N_20605);
nor U29989 (N_29989,N_24674,N_23236);
xor U29990 (N_29990,N_20427,N_22452);
nor U29991 (N_29991,N_22051,N_23519);
or U29992 (N_29992,N_21115,N_22562);
and U29993 (N_29993,N_24663,N_22014);
or U29994 (N_29994,N_24262,N_22044);
and U29995 (N_29995,N_24998,N_20464);
nand U29996 (N_29996,N_21999,N_24885);
or U29997 (N_29997,N_20290,N_20160);
or U29998 (N_29998,N_21623,N_21217);
xnor U29999 (N_29999,N_24687,N_24791);
or U30000 (N_30000,N_26286,N_29916);
and U30001 (N_30001,N_26554,N_25863);
and U30002 (N_30002,N_27816,N_26068);
nand U30003 (N_30003,N_26866,N_25575);
xor U30004 (N_30004,N_29126,N_25809);
and U30005 (N_30005,N_25642,N_26531);
nand U30006 (N_30006,N_29704,N_29194);
and U30007 (N_30007,N_25308,N_26894);
nor U30008 (N_30008,N_25462,N_27895);
nor U30009 (N_30009,N_26895,N_29355);
and U30010 (N_30010,N_28385,N_27728);
xor U30011 (N_30011,N_29939,N_29018);
nor U30012 (N_30012,N_26253,N_28278);
or U30013 (N_30013,N_28657,N_26745);
nor U30014 (N_30014,N_26376,N_27509);
and U30015 (N_30015,N_26901,N_26267);
nor U30016 (N_30016,N_25457,N_27575);
nor U30017 (N_30017,N_26299,N_25606);
nand U30018 (N_30018,N_27944,N_29236);
or U30019 (N_30019,N_25071,N_26400);
or U30020 (N_30020,N_29424,N_25368);
or U30021 (N_30021,N_27857,N_25986);
nand U30022 (N_30022,N_26443,N_26606);
and U30023 (N_30023,N_28665,N_27440);
nor U30024 (N_30024,N_27809,N_25278);
nor U30025 (N_30025,N_27841,N_28750);
or U30026 (N_30026,N_26645,N_25820);
nand U30027 (N_30027,N_29652,N_25310);
and U30028 (N_30028,N_26278,N_27349);
nand U30029 (N_30029,N_26808,N_28238);
nor U30030 (N_30030,N_28712,N_29395);
nand U30031 (N_30031,N_28601,N_27780);
nor U30032 (N_30032,N_27913,N_29245);
or U30033 (N_30033,N_27386,N_27388);
nor U30034 (N_30034,N_29712,N_25243);
xnor U30035 (N_30035,N_25586,N_27149);
nor U30036 (N_30036,N_28367,N_25136);
or U30037 (N_30037,N_25211,N_27287);
nor U30038 (N_30038,N_27639,N_26572);
or U30039 (N_30039,N_26625,N_28841);
xnor U30040 (N_30040,N_25132,N_27945);
and U30041 (N_30041,N_29799,N_28247);
nor U30042 (N_30042,N_28793,N_29407);
xor U30043 (N_30043,N_28880,N_29670);
nor U30044 (N_30044,N_28637,N_29388);
nor U30045 (N_30045,N_29452,N_27993);
nand U30046 (N_30046,N_29467,N_25500);
and U30047 (N_30047,N_26817,N_26450);
or U30048 (N_30048,N_29621,N_27422);
or U30049 (N_30049,N_28873,N_28212);
nand U30050 (N_30050,N_29515,N_28130);
nor U30051 (N_30051,N_25572,N_29443);
xnor U30052 (N_30052,N_27500,N_29171);
nor U30053 (N_30053,N_25679,N_26371);
nand U30054 (N_30054,N_29199,N_26779);
and U30055 (N_30055,N_27581,N_25355);
xor U30056 (N_30056,N_25821,N_27492);
or U30057 (N_30057,N_29461,N_27960);
xor U30058 (N_30058,N_26004,N_25294);
nand U30059 (N_30059,N_29569,N_28127);
and U30060 (N_30060,N_26141,N_25527);
nor U30061 (N_30061,N_25413,N_25522);
or U30062 (N_30062,N_26571,N_28609);
nor U30063 (N_30063,N_25142,N_28610);
nor U30064 (N_30064,N_29910,N_29160);
and U30065 (N_30065,N_29383,N_29660);
nand U30066 (N_30066,N_29787,N_28423);
or U30067 (N_30067,N_25823,N_28962);
xor U30068 (N_30068,N_25026,N_28320);
xnor U30069 (N_30069,N_27455,N_29694);
or U30070 (N_30070,N_28046,N_29516);
or U30071 (N_30071,N_29863,N_25836);
xor U30072 (N_30072,N_25540,N_28583);
and U30073 (N_30073,N_28080,N_26188);
nand U30074 (N_30074,N_26784,N_27361);
nor U30075 (N_30075,N_28525,N_26463);
or U30076 (N_30076,N_29542,N_27112);
nand U30077 (N_30077,N_28124,N_28202);
nand U30078 (N_30078,N_27057,N_27401);
nor U30079 (N_30079,N_26219,N_29172);
xnor U30080 (N_30080,N_27878,N_29336);
xor U30081 (N_30081,N_28459,N_27070);
nand U30082 (N_30082,N_27048,N_28613);
nor U30083 (N_30083,N_26142,N_25541);
nor U30084 (N_30084,N_27000,N_27820);
or U30085 (N_30085,N_26934,N_29492);
or U30086 (N_30086,N_26962,N_29153);
nand U30087 (N_30087,N_28984,N_28058);
xor U30088 (N_30088,N_28940,N_26398);
or U30089 (N_30089,N_28932,N_28431);
xnor U30090 (N_30090,N_29350,N_27027);
xor U30091 (N_30091,N_25009,N_29124);
and U30092 (N_30092,N_25359,N_26546);
and U30093 (N_30093,N_26911,N_26041);
nand U30094 (N_30094,N_25099,N_26378);
xor U30095 (N_30095,N_25502,N_28888);
xnor U30096 (N_30096,N_26172,N_28980);
xnor U30097 (N_30097,N_27962,N_29938);
nand U30098 (N_30098,N_29000,N_26467);
and U30099 (N_30099,N_28799,N_29005);
nand U30100 (N_30100,N_25912,N_25323);
nand U30101 (N_30101,N_25934,N_28507);
nor U30102 (N_30102,N_29330,N_25810);
nand U30103 (N_30103,N_26447,N_26790);
and U30104 (N_30104,N_25017,N_28322);
nor U30105 (N_30105,N_28344,N_26920);
and U30106 (N_30106,N_29796,N_29511);
xnor U30107 (N_30107,N_28981,N_25474);
or U30108 (N_30108,N_26643,N_28312);
nor U30109 (N_30109,N_29357,N_29514);
or U30110 (N_30110,N_29664,N_25037);
nor U30111 (N_30111,N_29014,N_27197);
xnor U30112 (N_30112,N_26140,N_29300);
nor U30113 (N_30113,N_27733,N_25720);
xor U30114 (N_30114,N_26291,N_29249);
nor U30115 (N_30115,N_28305,N_26823);
or U30116 (N_30116,N_27556,N_26013);
nor U30117 (N_30117,N_25415,N_25241);
nor U30118 (N_30118,N_25232,N_29051);
nand U30119 (N_30119,N_27647,N_27050);
nand U30120 (N_30120,N_29317,N_27496);
or U30121 (N_30121,N_25531,N_28267);
nor U30122 (N_30122,N_27548,N_25234);
or U30123 (N_30123,N_28397,N_29689);
or U30124 (N_30124,N_25941,N_25712);
nor U30125 (N_30125,N_29354,N_29417);
nand U30126 (N_30126,N_25125,N_29952);
xnor U30127 (N_30127,N_26787,N_28713);
xnor U30128 (N_30128,N_28653,N_28786);
or U30129 (N_30129,N_26707,N_25746);
or U30130 (N_30130,N_25162,N_27054);
nor U30131 (N_30131,N_25429,N_29861);
and U30132 (N_30132,N_26063,N_25370);
and U30133 (N_30133,N_29656,N_28812);
and U30134 (N_30134,N_25425,N_28033);
xnor U30135 (N_30135,N_29472,N_26154);
xnor U30136 (N_30136,N_28438,N_28389);
xnor U30137 (N_30137,N_26012,N_27844);
xnor U30138 (N_30138,N_29296,N_27209);
or U30139 (N_30139,N_29699,N_27906);
xor U30140 (N_30140,N_28952,N_25560);
xor U30141 (N_30141,N_26101,N_29303);
nand U30142 (N_30142,N_25604,N_27465);
or U30143 (N_30143,N_26608,N_27371);
xor U30144 (N_30144,N_25752,N_29364);
or U30145 (N_30145,N_26337,N_26747);
and U30146 (N_30146,N_25690,N_25840);
nand U30147 (N_30147,N_25350,N_28970);
or U30148 (N_30148,N_29585,N_28417);
and U30149 (N_30149,N_26048,N_25143);
nand U30150 (N_30150,N_25641,N_29009);
and U30151 (N_30151,N_28086,N_27606);
or U30152 (N_30152,N_27546,N_27310);
nand U30153 (N_30153,N_27311,N_25906);
and U30154 (N_30154,N_27708,N_26650);
or U30155 (N_30155,N_28023,N_25126);
xnor U30156 (N_30156,N_26201,N_26964);
xor U30157 (N_30157,N_26959,N_26290);
and U30158 (N_30158,N_28376,N_26046);
nand U30159 (N_30159,N_26610,N_28430);
or U30160 (N_30160,N_29304,N_28769);
or U30161 (N_30161,N_25302,N_28135);
nor U30162 (N_30162,N_26277,N_29725);
nand U30163 (N_30163,N_29456,N_29220);
nand U30164 (N_30164,N_26739,N_29015);
xnor U30165 (N_30165,N_25061,N_29095);
nand U30166 (N_30166,N_26247,N_29162);
xnor U30167 (N_30167,N_25373,N_28805);
nand U30168 (N_30168,N_26327,N_26311);
or U30169 (N_30169,N_27420,N_25051);
and U30170 (N_30170,N_29958,N_28266);
nor U30171 (N_30171,N_26859,N_28233);
xnor U30172 (N_30172,N_28097,N_26899);
nor U30173 (N_30173,N_27023,N_27397);
nand U30174 (N_30174,N_26539,N_28439);
and U30175 (N_30175,N_29818,N_25782);
and U30176 (N_30176,N_25842,N_29113);
and U30177 (N_30177,N_25191,N_29648);
or U30178 (N_30178,N_28626,N_29468);
and U30179 (N_30179,N_26027,N_28783);
or U30180 (N_30180,N_26213,N_28722);
nor U30181 (N_30181,N_25552,N_26434);
or U30182 (N_30182,N_29310,N_29106);
nand U30183 (N_30183,N_26854,N_26344);
nor U30184 (N_30184,N_27037,N_26953);
nand U30185 (N_30185,N_26474,N_28522);
nand U30186 (N_30186,N_28508,N_25683);
and U30187 (N_30187,N_28040,N_25616);
or U30188 (N_30188,N_25284,N_28270);
and U30189 (N_30189,N_26726,N_26574);
xor U30190 (N_30190,N_25307,N_28067);
and U30191 (N_30191,N_27785,N_29842);
nand U30192 (N_30192,N_29596,N_28916);
xor U30193 (N_30193,N_27744,N_28304);
and U30194 (N_30194,N_28502,N_26150);
or U30195 (N_30195,N_25776,N_28147);
and U30196 (N_30196,N_27421,N_29845);
nand U30197 (N_30197,N_27199,N_25729);
or U30198 (N_30198,N_27924,N_28704);
nand U30199 (N_30199,N_27796,N_28093);
nand U30200 (N_30200,N_25834,N_26364);
or U30201 (N_30201,N_25334,N_25257);
nand U30202 (N_30202,N_27097,N_27398);
nor U30203 (N_30203,N_26016,N_29993);
nand U30204 (N_30204,N_29804,N_26518);
and U30205 (N_30205,N_26521,N_28628);
and U30206 (N_30206,N_25212,N_27846);
and U30207 (N_30207,N_27467,N_27890);
or U30208 (N_30208,N_28745,N_28616);
or U30209 (N_30209,N_27712,N_26026);
and U30210 (N_30210,N_26465,N_25240);
or U30211 (N_30211,N_29021,N_29161);
xor U30212 (N_30212,N_25837,N_25794);
nand U30213 (N_30213,N_29368,N_26613);
or U30214 (N_30214,N_27497,N_28677);
nor U30215 (N_30215,N_26452,N_26743);
nor U30216 (N_30216,N_26662,N_26082);
nand U30217 (N_30217,N_29375,N_25832);
nand U30218 (N_30218,N_27760,N_27264);
nand U30219 (N_30219,N_27534,N_25301);
nor U30220 (N_30220,N_26544,N_29742);
or U30221 (N_30221,N_26744,N_27474);
or U30222 (N_30222,N_27995,N_27787);
nor U30223 (N_30223,N_25317,N_28638);
xor U30224 (N_30224,N_27304,N_29159);
xnor U30225 (N_30225,N_25236,N_26054);
nand U30226 (N_30226,N_25981,N_28811);
nand U30227 (N_30227,N_25290,N_27735);
xor U30228 (N_30228,N_27550,N_29555);
nor U30229 (N_30229,N_25808,N_26918);
and U30230 (N_30230,N_26017,N_26120);
and U30231 (N_30231,N_27437,N_29687);
nand U30232 (N_30232,N_25033,N_29566);
nor U30233 (N_30233,N_28243,N_26462);
xnor U30234 (N_30234,N_26672,N_27459);
nor U30235 (N_30235,N_26352,N_27130);
xor U30236 (N_30236,N_26634,N_25313);
or U30237 (N_30237,N_25392,N_28864);
and U30238 (N_30238,N_28333,N_27797);
nand U30239 (N_30239,N_27162,N_29672);
nor U30240 (N_30240,N_28772,N_27638);
nor U30241 (N_30241,N_26635,N_25733);
or U30242 (N_30242,N_26604,N_27210);
or U30243 (N_30243,N_29572,N_29372);
nand U30244 (N_30244,N_25872,N_28785);
nor U30245 (N_30245,N_29911,N_28910);
xor U30246 (N_30246,N_28106,N_27717);
or U30247 (N_30247,N_27636,N_26783);
and U30248 (N_30248,N_27980,N_29004);
and U30249 (N_30249,N_27768,N_27279);
and U30250 (N_30250,N_26514,N_27525);
nand U30251 (N_30251,N_28540,N_26942);
and U30252 (N_30252,N_29949,N_29554);
nor U30253 (N_30253,N_26761,N_27183);
and U30254 (N_30254,N_26674,N_25396);
and U30255 (N_30255,N_29411,N_28061);
xnor U30256 (N_30256,N_27964,N_25882);
xnor U30257 (N_30257,N_27681,N_29077);
nor U30258 (N_30258,N_29537,N_26758);
nor U30259 (N_30259,N_28001,N_29274);
xnor U30260 (N_30260,N_28699,N_29844);
nand U30261 (N_30261,N_29504,N_29586);
nor U30262 (N_30262,N_28440,N_25996);
nand U30263 (N_30263,N_26878,N_29001);
nor U30264 (N_30264,N_28530,N_27602);
xnor U30265 (N_30265,N_26086,N_28487);
nor U30266 (N_30266,N_27439,N_29565);
nand U30267 (N_30267,N_26475,N_28101);
xor U30268 (N_30268,N_26035,N_26076);
or U30269 (N_30269,N_28565,N_28907);
nand U30270 (N_30270,N_27894,N_28707);
nand U30271 (N_30271,N_29995,N_27207);
xnor U30272 (N_30272,N_29540,N_27561);
and U30273 (N_30273,N_28598,N_29260);
and U30274 (N_30274,N_25957,N_28314);
or U30275 (N_30275,N_26717,N_25884);
nor U30276 (N_30276,N_29921,N_27021);
nand U30277 (N_30277,N_28108,N_25685);
and U30278 (N_30278,N_26487,N_29616);
nand U30279 (N_30279,N_29392,N_26751);
nand U30280 (N_30280,N_25760,N_27375);
xor U30281 (N_30281,N_27700,N_27128);
xor U30282 (N_30282,N_27483,N_28371);
or U30283 (N_30283,N_25770,N_25183);
or U30284 (N_30284,N_28009,N_29603);
nand U30285 (N_30285,N_28072,N_28643);
and U30286 (N_30286,N_25804,N_28291);
nor U30287 (N_30287,N_25473,N_28770);
nand U30288 (N_30288,N_27516,N_29746);
or U30289 (N_30289,N_25175,N_28410);
nand U30290 (N_30290,N_25452,N_26910);
xnor U30291 (N_30291,N_27551,N_26641);
nor U30292 (N_30292,N_25377,N_29299);
nor U30293 (N_30293,N_25592,N_29717);
xor U30294 (N_30294,N_26621,N_26782);
and U30295 (N_30295,N_27940,N_27389);
nor U30296 (N_30296,N_26484,N_25015);
and U30297 (N_30297,N_29080,N_26904);
nand U30298 (N_30298,N_28412,N_26670);
or U30299 (N_30299,N_27030,N_26191);
and U30300 (N_30300,N_26537,N_28154);
xor U30301 (N_30301,N_29577,N_26297);
or U30302 (N_30302,N_25815,N_26906);
or U30303 (N_30303,N_27547,N_27903);
nand U30304 (N_30304,N_28350,N_29747);
or U30305 (N_30305,N_26470,N_25653);
or U30306 (N_30306,N_29319,N_28373);
xnor U30307 (N_30307,N_25978,N_29063);
and U30308 (N_30308,N_25795,N_25580);
and U30309 (N_30309,N_27661,N_28162);
or U30310 (N_30310,N_29881,N_29235);
and U30311 (N_30311,N_25476,N_25072);
nor U30312 (N_30312,N_25847,N_25495);
nand U30313 (N_30313,N_28338,N_26214);
and U30314 (N_30314,N_28639,N_27189);
and U30315 (N_30315,N_28470,N_26809);
or U30316 (N_30316,N_27416,N_25948);
or U30317 (N_30317,N_26373,N_25657);
and U30318 (N_30318,N_28809,N_27049);
nor U30319 (N_30319,N_29255,N_27196);
or U30320 (N_30320,N_28355,N_27658);
nand U30321 (N_30321,N_29494,N_29186);
xnor U30322 (N_30322,N_25329,N_29700);
nor U30323 (N_30323,N_29943,N_29091);
and U30324 (N_30324,N_27594,N_29849);
and U30325 (N_30325,N_25264,N_26951);
nand U30326 (N_30326,N_28946,N_28190);
xor U30327 (N_30327,N_25702,N_26689);
xor U30328 (N_30328,N_27979,N_27665);
xnor U30329 (N_30329,N_26679,N_27019);
nor U30330 (N_30330,N_29047,N_25496);
nor U30331 (N_30331,N_26656,N_28457);
or U30332 (N_30332,N_28273,N_25715);
nor U30333 (N_30333,N_28422,N_29244);
nor U30334 (N_30334,N_26128,N_25738);
or U30335 (N_30335,N_28330,N_25238);
or U30336 (N_30336,N_27089,N_29036);
or U30337 (N_30337,N_26198,N_28425);
nand U30338 (N_30338,N_26081,N_27634);
and U30339 (N_30339,N_25116,N_29207);
nor U30340 (N_30340,N_26697,N_25983);
and U30341 (N_30341,N_27641,N_25154);
xor U30342 (N_30342,N_28436,N_27449);
xor U30343 (N_30343,N_26456,N_26137);
xnor U30344 (N_30344,N_26304,N_28052);
or U30345 (N_30345,N_28949,N_26535);
xor U30346 (N_30346,N_27732,N_26764);
and U30347 (N_30347,N_28803,N_28670);
nor U30348 (N_30348,N_29795,N_25638);
nand U30349 (N_30349,N_25724,N_25521);
or U30350 (N_30350,N_25732,N_25726);
nor U30351 (N_30351,N_28697,N_28201);
and U30352 (N_30352,N_29730,N_28794);
nor U30353 (N_30353,N_29120,N_29705);
nor U30354 (N_30354,N_27839,N_29608);
or U30355 (N_30355,N_28361,N_27985);
xnor U30356 (N_30356,N_27410,N_29810);
or U30357 (N_30357,N_27445,N_29779);
and U30358 (N_30358,N_28095,N_28323);
xnor U30359 (N_30359,N_29924,N_26788);
nor U30360 (N_30360,N_29164,N_25841);
and U30361 (N_30361,N_28790,N_27374);
or U30362 (N_30362,N_25216,N_26956);
xor U30363 (N_30363,N_27499,N_27519);
xor U30364 (N_30364,N_27303,N_27758);
or U30365 (N_30365,N_27669,N_28928);
xnor U30366 (N_30366,N_26636,N_26098);
nand U30367 (N_30367,N_28945,N_28240);
nor U30368 (N_30368,N_28335,N_26412);
or U30369 (N_30369,N_29283,N_27400);
nor U30370 (N_30370,N_27317,N_27265);
xor U30371 (N_30371,N_29366,N_28078);
or U30372 (N_30372,N_26181,N_27243);
or U30373 (N_30373,N_28363,N_26178);
nor U30374 (N_30374,N_26317,N_26777);
or U30375 (N_30375,N_26960,N_27013);
or U30376 (N_30376,N_25750,N_26970);
nand U30377 (N_30377,N_28332,N_27329);
xnor U30378 (N_30378,N_25293,N_29729);
nand U30379 (N_30379,N_27380,N_27868);
or U30380 (N_30380,N_25202,N_26361);
nor U30381 (N_30381,N_26440,N_28586);
nand U30382 (N_30382,N_25169,N_25239);
nand U30383 (N_30383,N_27932,N_28982);
nor U30384 (N_30384,N_25588,N_25997);
xor U30385 (N_30385,N_29848,N_29931);
nand U30386 (N_30386,N_28571,N_27542);
or U30387 (N_30387,N_26569,N_28137);
nor U30388 (N_30388,N_27975,N_29815);
and U30389 (N_30389,N_28223,N_29377);
nor U30390 (N_30390,N_29913,N_25148);
xor U30391 (N_30391,N_26603,N_29308);
xor U30392 (N_30392,N_26728,N_29528);
xnor U30393 (N_30393,N_26167,N_28319);
nor U30394 (N_30394,N_27336,N_26731);
or U30395 (N_30395,N_26583,N_28953);
or U30396 (N_30396,N_28475,N_29751);
nand U30397 (N_30397,N_25073,N_29797);
or U30398 (N_30398,N_25484,N_29216);
or U30399 (N_30399,N_29465,N_26925);
or U30400 (N_30400,N_26966,N_29398);
xnor U30401 (N_30401,N_28587,N_27452);
xnor U30402 (N_30402,N_29509,N_27295);
nor U30403 (N_30403,N_27362,N_28694);
nor U30404 (N_30404,N_25043,N_26413);
xnor U30405 (N_30405,N_28105,N_29885);
xnor U30406 (N_30406,N_29755,N_26426);
and U30407 (N_30407,N_28123,N_27505);
nand U30408 (N_30408,N_28004,N_26691);
nor U30409 (N_30409,N_28661,N_26981);
nor U30410 (N_30410,N_25545,N_26202);
or U30411 (N_30411,N_25023,N_29192);
nor U30412 (N_30412,N_28405,N_25371);
xnor U30413 (N_30413,N_28235,N_28007);
xor U30414 (N_30414,N_26365,N_27280);
and U30415 (N_30415,N_27201,N_25263);
xnor U30416 (N_30416,N_26459,N_29728);
or U30417 (N_30417,N_28964,N_27862);
xnor U30418 (N_30418,N_28452,N_29264);
xnor U30419 (N_30419,N_29482,N_29583);
nor U30420 (N_30420,N_29788,N_29447);
xnor U30421 (N_30421,N_28229,N_27079);
nand U30422 (N_30422,N_26008,N_25999);
or U30423 (N_30423,N_29320,N_28280);
nand U30424 (N_30424,N_28069,N_29778);
nor U30425 (N_30425,N_27907,N_26179);
or U30426 (N_30426,N_27494,N_29935);
nand U30427 (N_30427,N_27897,N_26489);
nand U30428 (N_30428,N_27348,N_25698);
nor U30429 (N_30429,N_27729,N_26534);
nand U30430 (N_30430,N_25910,N_28163);
and U30431 (N_30431,N_27076,N_28044);
and U30432 (N_30432,N_29534,N_26381);
nand U30433 (N_30433,N_28680,N_28943);
nand U30434 (N_30434,N_29790,N_26271);
and U30435 (N_30435,N_26543,N_26194);
or U30436 (N_30436,N_27224,N_25439);
xor U30437 (N_30437,N_26284,N_27052);
nor U30438 (N_30438,N_26388,N_27424);
nor U30439 (N_30439,N_28682,N_26169);
nand U30440 (N_30440,N_28060,N_28726);
and U30441 (N_30441,N_29217,N_25774);
nor U30442 (N_30442,N_29064,N_29551);
nor U30443 (N_30443,N_27704,N_29582);
and U30444 (N_30444,N_29553,N_27671);
nor U30445 (N_30445,N_25155,N_29466);
nor U30446 (N_30446,N_29741,N_28399);
xnor U30447 (N_30447,N_26767,N_28537);
and U30448 (N_30448,N_27538,N_29977);
nor U30449 (N_30449,N_28924,N_25489);
nand U30450 (N_30450,N_29812,N_28559);
xor U30451 (N_30451,N_28370,N_25442);
nor U30452 (N_30452,N_27709,N_29762);
or U30453 (N_30453,N_25137,N_28492);
nor U30454 (N_30454,N_29181,N_28277);
nand U30455 (N_30455,N_27042,N_25319);
nand U30456 (N_30456,N_25800,N_27369);
xor U30457 (N_30457,N_29400,N_25059);
nand U30458 (N_30458,N_27378,N_26362);
xor U30459 (N_30459,N_27316,N_25469);
and U30460 (N_30460,N_28780,N_28250);
nor U30461 (N_30461,N_28819,N_25945);
nor U30462 (N_30462,N_26858,N_28658);
nor U30463 (N_30463,N_28538,N_26733);
nand U30464 (N_30464,N_26312,N_28855);
nor U30465 (N_30465,N_28892,N_25708);
nand U30466 (N_30466,N_25594,N_25922);
xnor U30467 (N_30467,N_28224,N_27242);
and U30468 (N_30468,N_28447,N_27627);
nor U30469 (N_30469,N_28210,N_27033);
and U30470 (N_30470,N_26346,N_26917);
nand U30471 (N_30471,N_25088,N_27554);
xor U30472 (N_30472,N_27678,N_28729);
and U30473 (N_30473,N_27481,N_27012);
nor U30474 (N_30474,N_26748,N_28757);
xor U30475 (N_30475,N_28527,N_26308);
and U30476 (N_30476,N_29108,N_26668);
nor U30477 (N_30477,N_28420,N_26841);
xor U30478 (N_30478,N_27833,N_26108);
and U30479 (N_30479,N_27240,N_29232);
and U30480 (N_30480,N_29381,N_28258);
xor U30481 (N_30481,N_27355,N_29195);
nor U30482 (N_30482,N_26228,N_25816);
and U30483 (N_30483,N_25485,N_27664);
nor U30484 (N_30484,N_25060,N_29662);
or U30485 (N_30485,N_28092,N_26494);
nand U30486 (N_30486,N_29546,N_26123);
nand U30487 (N_30487,N_29632,N_28797);
or U30488 (N_30488,N_26153,N_28546);
nor U30489 (N_30489,N_28554,N_25851);
nand U30490 (N_30490,N_27078,N_27902);
xor U30491 (N_30491,N_25303,N_26216);
and U30492 (N_30492,N_25607,N_28303);
or U30493 (N_30493,N_28979,N_28611);
nand U30494 (N_30494,N_26044,N_26722);
or U30495 (N_30495,N_28282,N_28364);
nor U30496 (N_30496,N_28696,N_29635);
xor U30497 (N_30497,N_26309,N_26824);
xnor U30498 (N_30498,N_25354,N_25460);
xnor U30499 (N_30499,N_25564,N_27165);
and U30500 (N_30500,N_25864,N_29624);
nor U30501 (N_30501,N_26057,N_27859);
nor U30502 (N_30502,N_25237,N_26673);
xor U30503 (N_30503,N_26495,N_26792);
and U30504 (N_30504,N_26741,N_28861);
and U30505 (N_30505,N_28890,N_26713);
nor U30506 (N_30506,N_29805,N_26061);
or U30507 (N_30507,N_26993,N_29558);
xor U30508 (N_30508,N_25523,N_28967);
xor U30509 (N_30509,N_26240,N_26667);
or U30510 (N_30510,N_28723,N_25718);
or U30511 (N_30511,N_25001,N_25477);
xnor U30512 (N_30512,N_26457,N_26159);
nand U30513 (N_30513,N_26814,N_29607);
nand U30514 (N_30514,N_28302,N_26454);
nand U30515 (N_30515,N_26302,N_28996);
or U30516 (N_30516,N_27107,N_25189);
and U30517 (N_30517,N_28264,N_25411);
or U30518 (N_30518,N_27693,N_25897);
or U30519 (N_30519,N_26112,N_25372);
and U30520 (N_30520,N_28489,N_25601);
xor U30521 (N_30521,N_25493,N_28839);
nor U30522 (N_30522,N_28030,N_28602);
or U30523 (N_30523,N_28384,N_29180);
xnor U30524 (N_30524,N_28776,N_27766);
xor U30525 (N_30525,N_25393,N_29972);
nor U30526 (N_30526,N_29745,N_28169);
and U30527 (N_30527,N_28121,N_28215);
and U30528 (N_30528,N_27954,N_29107);
nand U30529 (N_30529,N_26839,N_27281);
or U30530 (N_30530,N_27482,N_26551);
xnor U30531 (N_30531,N_27167,N_28594);
and U30532 (N_30532,N_26220,N_25406);
nor U30533 (N_30533,N_28019,N_26998);
xnor U30534 (N_30534,N_29275,N_28039);
xnor U30535 (N_30535,N_29619,N_27751);
or U30536 (N_30536,N_28835,N_25672);
or U30537 (N_30537,N_26190,N_27640);
and U30538 (N_30538,N_29785,N_27943);
xor U30539 (N_30539,N_25204,N_25384);
nor U30540 (N_30540,N_28189,N_27094);
nand U30541 (N_30541,N_27777,N_25867);
xor U30542 (N_30542,N_26813,N_29587);
and U30543 (N_30543,N_26533,N_27599);
xnor U30544 (N_30544,N_28418,N_26106);
or U30545 (N_30545,N_26131,N_29448);
or U30546 (N_30546,N_27829,N_27628);
and U30547 (N_30547,N_27314,N_29010);
and U30548 (N_30548,N_25987,N_25727);
nor U30549 (N_30549,N_28500,N_28881);
nand U30550 (N_30550,N_28013,N_27702);
nor U30551 (N_30551,N_26876,N_29899);
nand U30552 (N_30552,N_26146,N_26006);
xor U30553 (N_30553,N_27179,N_28824);
and U30554 (N_30554,N_27046,N_26916);
and U30555 (N_30555,N_29523,N_26760);
xnor U30556 (N_30556,N_29423,N_25200);
and U30557 (N_30557,N_26197,N_28008);
and U30558 (N_30558,N_26113,N_25246);
and U30559 (N_30559,N_28719,N_26562);
nand U30560 (N_30560,N_25146,N_25669);
xor U30561 (N_30561,N_26114,N_29824);
or U30562 (N_30562,N_28591,N_25120);
nand U30563 (N_30563,N_27423,N_26132);
nor U30564 (N_30564,N_27866,N_26620);
xnor U30565 (N_30565,N_27477,N_28736);
nor U30566 (N_30566,N_26002,N_29433);
nand U30567 (N_30567,N_26303,N_28836);
and U30568 (N_30568,N_29322,N_26607);
nor U30569 (N_30569,N_25269,N_28299);
or U30570 (N_30570,N_25258,N_26774);
xor U30571 (N_30571,N_29478,N_29127);
nor U30572 (N_30572,N_28756,N_27438);
nand U30573 (N_30573,N_26585,N_29271);
nand U30574 (N_30574,N_25084,N_27790);
and U30575 (N_30575,N_28274,N_28568);
xnor U30576 (N_30576,N_25519,N_25348);
nand U30577 (N_30577,N_27589,N_26385);
xnor U30578 (N_30578,N_26025,N_27428);
and U30579 (N_30579,N_26504,N_27436);
nor U30580 (N_30580,N_29968,N_27419);
or U30581 (N_30581,N_26601,N_29333);
or U30582 (N_30582,N_25045,N_26433);
or U30583 (N_30583,N_28331,N_28950);
xor U30584 (N_30584,N_25844,N_28467);
nor U30585 (N_30585,N_29370,N_28755);
nor U30586 (N_30586,N_27727,N_27684);
xnor U30587 (N_30587,N_28377,N_26992);
nor U30588 (N_30588,N_26595,N_25207);
xor U30589 (N_30589,N_28795,N_27101);
nor U30590 (N_30590,N_29771,N_29581);
nand U30591 (N_30591,N_29757,N_28068);
or U30592 (N_30592,N_28931,N_29871);
and U30593 (N_30593,N_27691,N_29518);
and U30594 (N_30594,N_25118,N_25065);
nand U30595 (N_30595,N_26754,N_25353);
nand U30596 (N_30596,N_29535,N_29786);
or U30597 (N_30597,N_26182,N_25160);
or U30598 (N_30598,N_26896,N_26584);
nand U30599 (N_30599,N_27532,N_26955);
xor U30600 (N_30600,N_27241,N_28778);
and U30601 (N_30601,N_29281,N_29976);
or U30602 (N_30602,N_26037,N_28186);
nand U30603 (N_30603,N_25547,N_27901);
or U30604 (N_30604,N_25375,N_27450);
nor U30605 (N_30605,N_26567,N_26078);
xor U30606 (N_30606,N_25217,N_28133);
and U30607 (N_30607,N_29859,N_25608);
xor U30608 (N_30608,N_29289,N_27715);
nor U30609 (N_30609,N_25673,N_27978);
or U30610 (N_30610,N_27882,N_27723);
or U30611 (N_30611,N_27138,N_28652);
xor U30612 (N_30612,N_25193,N_29096);
nor U30613 (N_30613,N_25721,N_28182);
xnor U30614 (N_30614,N_28029,N_27479);
xnor U30615 (N_30615,N_27114,N_29083);
nor U30616 (N_30616,N_25528,N_28830);
nand U30617 (N_30617,N_25706,N_28968);
xnor U30618 (N_30618,N_29816,N_27004);
or U30619 (N_30619,N_29453,N_28110);
or U30620 (N_30620,N_29168,N_28585);
nor U30621 (N_30621,N_26517,N_25011);
nor U30622 (N_30622,N_29069,N_25042);
or U30623 (N_30623,N_29408,N_29793);
xor U30624 (N_30624,N_26614,N_26939);
nor U30625 (N_30625,N_29698,N_28545);
or U30626 (N_30626,N_29888,N_29144);
and U30627 (N_30627,N_25984,N_26499);
xnor U30628 (N_30628,N_29832,N_26407);
xnor U30629 (N_30629,N_28262,N_28372);
or U30630 (N_30630,N_27706,N_28209);
nand U30631 (N_30631,N_29072,N_27738);
or U30632 (N_30632,N_25870,N_27236);
nand U30633 (N_30633,N_25916,N_29519);
nor U30634 (N_30634,N_29946,N_28343);
nand U30635 (N_30635,N_28972,N_28326);
and U30636 (N_30636,N_27929,N_27812);
and U30637 (N_30637,N_29291,N_29838);
or U30638 (N_30638,N_27889,N_29893);
xnor U30639 (N_30639,N_25111,N_25838);
and U30640 (N_30640,N_29915,N_25487);
nor U30641 (N_30641,N_27966,N_25376);
xnor U30642 (N_30642,N_29716,N_25762);
or U30643 (N_30643,N_29645,N_27576);
and U30644 (N_30644,N_27177,N_25789);
and U30645 (N_30645,N_27016,N_26196);
and U30646 (N_30646,N_28779,N_29020);
xnor U30647 (N_30647,N_27540,N_27904);
nor U30648 (N_30648,N_28166,N_28094);
and U30649 (N_30649,N_28187,N_29313);
nor U30650 (N_30650,N_27813,N_29343);
nor U30651 (N_30651,N_27867,N_28152);
nor U30652 (N_30652,N_27623,N_28381);
or U30653 (N_30653,N_26599,N_25190);
nor U30654 (N_30654,N_27838,N_29369);
and U30655 (N_30655,N_27896,N_29834);
xnor U30656 (N_30656,N_28768,N_25002);
nor U30657 (N_30657,N_25298,N_28845);
nor U30658 (N_30658,N_25499,N_25389);
nor U30659 (N_30659,N_26207,N_28177);
nand U30660 (N_30660,N_28742,N_26596);
and U30661 (N_30661,N_26021,N_29013);
or U30662 (N_30662,N_29432,N_26357);
nor U30663 (N_30663,N_27257,N_29287);
or U30664 (N_30664,N_27769,N_25184);
and U30665 (N_30665,N_27582,N_28485);
and U30666 (N_30666,N_28112,N_27515);
nand U30667 (N_30667,N_25188,N_29580);
and U30668 (N_30668,N_27997,N_27806);
xor U30669 (N_30669,N_25709,N_29722);
nand U30670 (N_30670,N_29394,N_26262);
or U30671 (N_30671,N_25509,N_29763);
xor U30672 (N_30672,N_29631,N_28838);
and U30673 (N_30673,N_27132,N_29695);
or U30674 (N_30674,N_29415,N_25149);
nand U30675 (N_30675,N_25972,N_28672);
and U30676 (N_30676,N_26785,N_25448);
nand U30677 (N_30677,N_29965,N_28128);
and U30678 (N_30678,N_25314,N_25617);
nand U30679 (N_30679,N_26898,N_25322);
or U30680 (N_30680,N_27874,N_28462);
nor U30681 (N_30681,N_25032,N_25028);
nand U30682 (N_30682,N_25883,N_27802);
xor U30683 (N_30683,N_25643,N_26420);
or U30684 (N_30684,N_29640,N_26305);
nor U30685 (N_30685,N_25173,N_25859);
and U30686 (N_30686,N_25968,N_28226);
nand U30687 (N_30687,N_29265,N_29484);
and U30688 (N_30688,N_27963,N_29820);
xor U30689 (N_30689,N_25426,N_25573);
and U30690 (N_30690,N_29601,N_27612);
nand U30691 (N_30691,N_26822,N_26289);
and U30692 (N_30692,N_25078,N_25518);
nor U30693 (N_30693,N_26941,N_28192);
and U30694 (N_30694,N_25080,N_28577);
xnor U30695 (N_30695,N_27195,N_28035);
nor U30696 (N_30696,N_25455,N_26232);
nor U30697 (N_30697,N_27292,N_26501);
or U30698 (N_30698,N_28925,N_25854);
or U30699 (N_30699,N_26694,N_29724);
or U30700 (N_30700,N_25058,N_25913);
or U30701 (N_30701,N_27286,N_28196);
nand U30702 (N_30702,N_27725,N_29944);
nand U30703 (N_30703,N_25262,N_25513);
xor U30704 (N_30704,N_25279,N_26710);
nand U30705 (N_30705,N_29464,N_25796);
and U30706 (N_30706,N_25013,N_29520);
nor U30707 (N_30707,N_29496,N_27990);
and U30708 (N_30708,N_29869,N_29637);
nor U30709 (N_30709,N_29152,N_25849);
xnor U30710 (N_30710,N_29883,N_28296);
or U30711 (N_30711,N_25765,N_28818);
xnor U30712 (N_30712,N_29145,N_26630);
and U30713 (N_30713,N_27677,N_27382);
nor U30714 (N_30714,N_27463,N_26756);
xor U30715 (N_30715,N_28476,N_25339);
nor U30716 (N_30716,N_25097,N_29851);
and U30717 (N_30717,N_26453,N_28241);
xor U30718 (N_30718,N_28334,N_27776);
xnor U30719 (N_30719,N_25105,N_28869);
and U30720 (N_30720,N_29007,N_28056);
nand U30721 (N_30721,N_25611,N_27625);
or U30722 (N_30722,N_25719,N_28674);
or U30723 (N_30723,N_27151,N_27524);
nand U30724 (N_30724,N_25276,N_26211);
nand U30725 (N_30725,N_26102,N_25128);
or U30726 (N_30726,N_27476,N_27160);
or U30727 (N_30727,N_25918,N_26780);
nand U30728 (N_30728,N_29775,N_29226);
xnor U30729 (N_30729,N_28091,N_27617);
or U30730 (N_30730,N_26836,N_25548);
and U30731 (N_30731,N_25558,N_29657);
or U30732 (N_30732,N_28342,N_26200);
xor U30733 (N_30733,N_26410,N_25492);
nor U30734 (N_30734,N_25963,N_29327);
nand U30735 (N_30735,N_28821,N_26295);
and U30736 (N_30736,N_28689,N_25511);
nor U30737 (N_30737,N_29463,N_29389);
nor U30738 (N_30738,N_27487,N_26056);
or U30739 (N_30739,N_26359,N_26244);
or U30740 (N_30740,N_25312,N_26272);
nor U30741 (N_30741,N_29098,N_29685);
nand U30742 (N_30742,N_26696,N_27544);
nor U30743 (N_30743,N_29428,N_28870);
or U30744 (N_30744,N_28715,N_27536);
or U30745 (N_30745,N_25902,N_25428);
xnor U30746 (N_30746,N_29748,N_29634);
nor U30747 (N_30747,N_25292,N_27066);
nor U30748 (N_30748,N_28927,N_27003);
or U30749 (N_30749,N_29073,N_29500);
xor U30750 (N_30750,N_29030,N_27583);
and U30751 (N_30751,N_29223,N_28254);
nand U30752 (N_30752,N_25759,N_27667);
nand U30753 (N_30753,N_28074,N_26540);
and U30754 (N_30754,N_25555,N_29446);
or U30755 (N_30755,N_28404,N_25430);
nor U30756 (N_30756,N_26575,N_25123);
and U30757 (N_30757,N_27731,N_26819);
and U30758 (N_30758,N_25739,N_28180);
nand U30759 (N_30759,N_25704,N_25114);
nor U30760 (N_30760,N_29710,N_26711);
xnor U30761 (N_30761,N_26394,N_26294);
nand U30762 (N_30762,N_28896,N_26622);
nor U30763 (N_30763,N_26655,N_26511);
xnor U30764 (N_30764,N_29868,N_27754);
nand U30765 (N_30765,N_26322,N_29920);
nand U30766 (N_30766,N_26699,N_25054);
and U30767 (N_30767,N_25093,N_28073);
nand U30768 (N_30768,N_25827,N_27850);
and U30769 (N_30769,N_28022,N_28903);
nor U30770 (N_30770,N_26425,N_29891);
nand U30771 (N_30771,N_28876,N_28107);
or U30772 (N_30772,N_27180,N_26929);
or U30773 (N_30773,N_29046,N_29019);
nor U30774 (N_30774,N_26652,N_27937);
and U30775 (N_30775,N_25075,N_26935);
or U30776 (N_30776,N_27322,N_27950);
xor U30777 (N_30777,N_25367,N_26639);
nor U30778 (N_30778,N_29808,N_25289);
or U30779 (N_30779,N_27136,N_26045);
nor U30780 (N_30780,N_28804,N_25129);
or U30781 (N_30781,N_26979,N_27067);
and U30782 (N_30782,N_26781,N_25134);
and U30783 (N_30783,N_29578,N_29092);
nor U30784 (N_30784,N_25950,N_25424);
or U30785 (N_30785,N_25605,N_26512);
xor U30786 (N_30786,N_29268,N_25004);
and U30787 (N_30787,N_29835,N_25196);
or U30788 (N_30788,N_29817,N_25713);
nand U30789 (N_30789,N_29156,N_25621);
xor U30790 (N_30790,N_26503,N_28564);
xor U30791 (N_30791,N_27852,N_25352);
and U30792 (N_30792,N_27126,N_29777);
nand U30793 (N_30793,N_27883,N_25494);
nor U30794 (N_30794,N_29688,N_28663);
nor U30795 (N_30795,N_28310,N_29174);
and U30796 (N_30796,N_29807,N_28308);
or U30797 (N_30797,N_27767,N_28259);
or U30798 (N_30798,N_29344,N_26427);
xnor U30799 (N_30799,N_25773,N_27456);
nor U30800 (N_30800,N_26349,N_25803);
or U30801 (N_30801,N_27170,N_29385);
nor U30802 (N_30802,N_26264,N_25378);
nor U30803 (N_30803,N_25098,N_26251);
xor U30804 (N_30804,N_27872,N_27148);
and U30805 (N_30805,N_26903,N_28145);
and U30806 (N_30806,N_25335,N_29609);
nor U30807 (N_30807,N_26328,N_27772);
nor U30808 (N_30808,N_27285,N_28624);
nand U30809 (N_30809,N_28194,N_27453);
nand U30810 (N_30810,N_27968,N_28050);
nand U30811 (N_30811,N_25788,N_27668);
and U30812 (N_30812,N_27560,N_28205);
xor U30813 (N_30813,N_28641,N_27173);
or U30814 (N_30814,N_25671,N_28047);
nand U30815 (N_30815,N_25390,N_28286);
xnor U30816 (N_30816,N_27092,N_28390);
xor U30817 (N_30817,N_25208,N_29349);
nor U30818 (N_30818,N_27597,N_28884);
nand U30819 (N_30819,N_27102,N_28175);
nor U30820 (N_30820,N_25094,N_25403);
nor U30821 (N_30821,N_26341,N_26406);
and U30822 (N_30822,N_27338,N_29919);
nand U30823 (N_30823,N_27294,N_25824);
nand U30824 (N_30824,N_26804,N_28214);
or U30825 (N_30825,N_27284,N_28386);
nor U30826 (N_30826,N_25338,N_29948);
and U30827 (N_30827,N_26830,N_26266);
xnor U30828 (N_30828,N_28679,N_26033);
xor U30829 (N_30829,N_26187,N_28807);
xnor U30830 (N_30830,N_26753,N_27247);
xor U30831 (N_30831,N_26666,N_26446);
or U30832 (N_30832,N_26891,N_29951);
xnor U30833 (N_30833,N_26403,N_27328);
nand U30834 (N_30834,N_25636,N_27091);
nor U30835 (N_30835,N_26241,N_29139);
xor U30836 (N_30836,N_29099,N_26015);
or U30837 (N_30837,N_28894,N_29963);
xnor U30838 (N_30838,N_28754,N_29384);
and U30839 (N_30839,N_29614,N_28176);
or U30840 (N_30840,N_29629,N_26342);
nor U30841 (N_30841,N_25412,N_27942);
and U30842 (N_30842,N_25695,N_26769);
nor U30843 (N_30843,N_27134,N_28236);
or U30844 (N_30844,N_29479,N_29830);
and U30845 (N_30845,N_29622,N_27824);
or U30846 (N_30846,N_29675,N_28010);
or U30847 (N_30847,N_25900,N_26924);
xor U30848 (N_30848,N_25614,N_29679);
nor U30849 (N_30849,N_28151,N_28710);
and U30850 (N_30850,N_26144,N_26215);
and U30851 (N_30851,N_26909,N_27185);
or U30852 (N_30852,N_28695,N_28178);
nor U30853 (N_30853,N_26409,N_25923);
or U30854 (N_30854,N_29595,N_27131);
or U30855 (N_30855,N_27899,N_29006);
nand U30856 (N_30856,N_27200,N_27031);
nand U30857 (N_30857,N_25052,N_27523);
nand U30858 (N_30858,N_29297,N_28607);
or U30859 (N_30859,N_27637,N_26867);
nand U30860 (N_30860,N_28801,N_25907);
nor U30861 (N_30861,N_26556,N_29016);
nor U30862 (N_30862,N_28576,N_27543);
nand U30863 (N_30863,N_29208,N_26589);
and U30864 (N_30864,N_26541,N_25470);
nand U30865 (N_30865,N_25975,N_25660);
nor U30866 (N_30866,N_28368,N_25791);
nor U30867 (N_30867,N_29034,N_26887);
xor U30868 (N_30868,N_28579,N_28963);
nor U30869 (N_30869,N_26773,N_27085);
nand U30870 (N_30870,N_28498,N_25340);
nor U30871 (N_30871,N_25909,N_28668);
nand U30872 (N_30872,N_27584,N_29800);
nand U30873 (N_30873,N_29731,N_25506);
and U30874 (N_30874,N_29766,N_27334);
xnor U30875 (N_30875,N_26180,N_28142);
nand U30876 (N_30876,N_25772,N_26292);
xor U30877 (N_30877,N_26332,N_27988);
nand U30878 (N_30878,N_28791,N_27512);
xor U30879 (N_30879,N_25675,N_28461);
nand U30880 (N_30880,N_28796,N_29571);
nand U30881 (N_30881,N_25230,N_28248);
nor U30882 (N_30882,N_26893,N_29678);
nor U30883 (N_30883,N_25697,N_28325);
and U30884 (N_30884,N_27941,N_27662);
nand U30885 (N_30885,N_27144,N_28463);
or U30886 (N_30886,N_28437,N_28798);
and U30887 (N_30887,N_29132,N_25482);
nand U30888 (N_30888,N_25351,N_25938);
nor U30889 (N_30889,N_28636,N_29163);
and U30890 (N_30890,N_26837,N_25942);
and U30891 (N_30891,N_28041,N_28617);
nand U30892 (N_30892,N_26509,N_26671);
xnor U30893 (N_30893,N_29332,N_26372);
nand U30894 (N_30894,N_28349,N_26174);
or U30895 (N_30895,N_27522,N_25273);
nand U30896 (N_30896,N_28427,N_28253);
nor U30897 (N_30897,N_29512,N_27799);
xor U30898 (N_30898,N_26031,N_28588);
nor U30899 (N_30899,N_28913,N_29658);
and U30900 (N_30900,N_29732,N_25976);
xnor U30901 (N_30901,N_26351,N_27996);
nand U30902 (N_30902,N_25964,N_27504);
or U30903 (N_30903,N_29773,N_29964);
nor U30904 (N_30904,N_28165,N_25753);
and U30905 (N_30905,N_27624,N_29454);
nand U30906 (N_30906,N_26800,N_27485);
nor U30907 (N_30907,N_28134,N_27153);
nor U30908 (N_30908,N_29860,N_29474);
xor U30909 (N_30909,N_29959,N_27804);
nor U30910 (N_30910,N_29937,N_29123);
xnor U30911 (N_30911,N_25268,N_27002);
nand U30912 (N_30912,N_28398,N_27272);
or U30913 (N_30913,N_26138,N_25680);
nand U30914 (N_30914,N_25543,N_29112);
nor U30915 (N_30915,N_29416,N_29241);
and U30916 (N_30916,N_29175,N_25530);
nor U30917 (N_30917,N_28647,N_25958);
nand U30918 (N_30918,N_26273,N_28081);
nor U30919 (N_30919,N_26160,N_29352);
or U30920 (N_30920,N_27959,N_29238);
and U30921 (N_30921,N_25932,N_26912);
xnor U30922 (N_30922,N_29991,N_28895);
or U30923 (N_30923,N_25661,N_28111);
xnor U30924 (N_30924,N_29142,N_27557);
and U30925 (N_30925,N_29821,N_29197);
and U30926 (N_30926,N_29875,N_28702);
and U30927 (N_30927,N_26384,N_26254);
and U30928 (N_30928,N_25525,N_26762);
or U30929 (N_30929,N_26038,N_29783);
xnor U30930 (N_30930,N_28929,N_27620);
or U30931 (N_30931,N_26805,N_29600);
nor U30932 (N_30932,N_25024,N_25542);
and U30933 (N_30933,N_26612,N_26177);
or U30934 (N_30934,N_25326,N_25281);
xor U30935 (N_30935,N_27480,N_25503);
xnor U30936 (N_30936,N_25801,N_29012);
and U30937 (N_30937,N_27433,N_27958);
xnor U30938 (N_30938,N_28168,N_27300);
nor U30939 (N_30939,N_27568,N_29059);
and U30940 (N_30940,N_29772,N_29683);
or U30941 (N_30941,N_25887,N_25461);
xor U30942 (N_30942,N_28558,N_28179);
or U30943 (N_30943,N_27644,N_25878);
nand U30944 (N_30944,N_28909,N_26498);
or U30945 (N_30945,N_25091,N_28645);
or U30946 (N_30946,N_29980,N_27853);
or U30947 (N_30947,N_25895,N_26840);
xnor U30948 (N_30948,N_26158,N_26864);
nand U30949 (N_30949,N_26121,N_29840);
and U30950 (N_30950,N_25647,N_26334);
nor U30951 (N_30951,N_26598,N_25057);
and U30952 (N_30952,N_27204,N_27849);
xnor U30953 (N_30953,N_26036,N_28941);
and U30954 (N_30954,N_26869,N_27720);
xnor U30955 (N_30955,N_27006,N_26049);
nand U30956 (N_30956,N_26246,N_26083);
nor U30957 (N_30957,N_27673,N_28408);
and U30958 (N_30958,N_27381,N_25596);
or U30959 (N_30959,N_29305,N_26847);
xnor U30960 (N_30960,N_29999,N_27961);
nand U30961 (N_30961,N_29211,N_29508);
nand U30962 (N_30962,N_28450,N_26863);
nand U30963 (N_30963,N_26724,N_26664);
or U30964 (N_30964,N_27282,N_27154);
xor U30965 (N_30965,N_28784,N_29781);
or U30966 (N_30966,N_29024,N_29727);
nand U30967 (N_30967,N_29550,N_26772);
xor U30968 (N_30968,N_27426,N_25242);
xnor U30969 (N_30969,N_27887,N_28922);
nor U30970 (N_30970,N_27028,N_27460);
xnor U30971 (N_30971,N_25185,N_27044);
nand U30972 (N_30972,N_25745,N_25949);
nor U30973 (N_30973,N_29050,N_29338);
or U30974 (N_30974,N_28771,N_27685);
xor U30975 (N_30975,N_28850,N_29536);
or U30976 (N_30976,N_29703,N_29653);
nand U30977 (N_30977,N_29989,N_26091);
xor U30978 (N_30978,N_28415,N_26852);
or U30979 (N_30979,N_27350,N_29872);
nand U30980 (N_30980,N_28442,N_27619);
xnor U30981 (N_30981,N_26192,N_25819);
nand U30982 (N_30982,N_28403,N_29351);
and U30983 (N_30983,N_26600,N_29008);
or U30984 (N_30984,N_26257,N_27161);
nand U30985 (N_30985,N_25865,N_28990);
or U30986 (N_30986,N_26646,N_25036);
nor U30987 (N_30987,N_26520,N_29676);
or U30988 (N_30988,N_27069,N_28283);
nor U30989 (N_30989,N_28849,N_27041);
and U30990 (N_30990,N_29182,N_25571);
and U30991 (N_30991,N_29539,N_29301);
xnor U30992 (N_30992,N_29337,N_29251);
and U30993 (N_30993,N_26530,N_27251);
or U30994 (N_30994,N_27155,N_25920);
and U30995 (N_30995,N_28173,N_25570);
xor U30996 (N_30996,N_25297,N_28064);
or U30997 (N_30997,N_26161,N_28222);
or U30998 (N_30998,N_28294,N_27110);
xnor U30999 (N_30999,N_26005,N_28954);
nand U31000 (N_31000,N_26382,N_29237);
or U31001 (N_31001,N_28488,N_29191);
nand U31002 (N_31002,N_27805,N_28444);
nand U31003 (N_31003,N_26709,N_25046);
or U31004 (N_31004,N_28474,N_26285);
xor U31005 (N_31005,N_26519,N_25341);
xnor U31006 (N_31006,N_27268,N_26926);
nand U31007 (N_31007,N_27585,N_29003);
or U31008 (N_31008,N_25436,N_27698);
or U31009 (N_31009,N_27193,N_29298);
nand U31010 (N_31010,N_26527,N_28012);
nand U31011 (N_31011,N_26555,N_29420);
xor U31012 (N_31012,N_27090,N_28230);
nand U31013 (N_31013,N_26070,N_26092);
nor U31014 (N_31014,N_28451,N_25176);
nor U31015 (N_31015,N_29597,N_27129);
nor U31016 (N_31016,N_25618,N_29538);
nand U31017 (N_31017,N_28837,N_27342);
xor U31018 (N_31018,N_27590,N_26757);
nand U31019 (N_31019,N_25535,N_25087);
or U31020 (N_31020,N_28119,N_26226);
nor U31021 (N_31021,N_27526,N_29611);
nand U31022 (N_31022,N_25214,N_29032);
or U31023 (N_31023,N_27934,N_28787);
xnor U31024 (N_31024,N_28195,N_27234);
and U31025 (N_31025,N_27119,N_26552);
and U31026 (N_31026,N_27133,N_28816);
nand U31027 (N_31027,N_26715,N_29713);
or U31028 (N_31028,N_29789,N_27253);
nand U31029 (N_31029,N_28552,N_26810);
nand U31030 (N_31030,N_28172,N_29318);
or U31031 (N_31031,N_27250,N_26249);
nand U31032 (N_31032,N_26961,N_25288);
nand U31033 (N_31033,N_29234,N_29334);
nand U31034 (N_31034,N_26714,N_28197);
nor U31035 (N_31035,N_26441,N_27588);
nor U31036 (N_31036,N_27675,N_26631);
or U31037 (N_31037,N_29760,N_28813);
or U31038 (N_31038,N_27366,N_25320);
or U31039 (N_31039,N_29708,N_25904);
nor U31040 (N_31040,N_29434,N_28279);
nor U31041 (N_31041,N_29561,N_27081);
xnor U31042 (N_31042,N_29341,N_25741);
xnor U31043 (N_31043,N_28345,N_25174);
nand U31044 (N_31044,N_29973,N_25512);
xor U31045 (N_31045,N_27104,N_26445);
and U31046 (N_31046,N_26806,N_27212);
nand U31047 (N_31047,N_25347,N_28879);
nand U31048 (N_31048,N_28146,N_25437);
nor U31049 (N_31049,N_27198,N_28365);
nand U31050 (N_31050,N_27596,N_28011);
nand U31051 (N_31051,N_29887,N_26437);
nand U31052 (N_31052,N_27466,N_27578);
or U31053 (N_31053,N_25282,N_28520);
xor U31054 (N_31054,N_28635,N_25182);
or U31055 (N_31055,N_27045,N_25402);
and U31056 (N_31056,N_28116,N_27856);
nand U31057 (N_31057,N_25928,N_25082);
and U31058 (N_31058,N_26050,N_26293);
nor U31059 (N_31059,N_25684,N_25096);
nand U31060 (N_31060,N_28318,N_29498);
and U31061 (N_31061,N_25843,N_29936);
xnor U31062 (N_31062,N_26497,N_27666);
or U31063 (N_31063,N_28139,N_25113);
xnor U31064 (N_31064,N_25599,N_28631);
nor U31065 (N_31065,N_27111,N_27221);
nand U31066 (N_31066,N_28848,N_27580);
xnor U31067 (N_31067,N_27490,N_25852);
xor U31068 (N_31068,N_27024,N_27176);
and U31069 (N_31069,N_28618,N_28882);
and U31070 (N_31070,N_25454,N_29023);
nor U31071 (N_31071,N_28782,N_25551);
and U31072 (N_31072,N_25549,N_26391);
nand U31073 (N_31073,N_27194,N_25985);
nor U31074 (N_31074,N_28481,N_28792);
xor U31075 (N_31075,N_25769,N_27290);
and U31076 (N_31076,N_28829,N_28084);
nor U31077 (N_31077,N_26084,N_25956);
nor U31078 (N_31078,N_27773,N_27337);
nand U31079 (N_31079,N_28265,N_26282);
nor U31080 (N_31080,N_25049,N_28622);
nand U31081 (N_31081,N_29691,N_29642);
and U31082 (N_31082,N_28446,N_29043);
or U31083 (N_31083,N_29259,N_27029);
nor U31084 (N_31084,N_29819,N_28534);
and U31085 (N_31085,N_26268,N_26834);
xnor U31086 (N_31086,N_26884,N_26095);
or U31087 (N_31087,N_25034,N_25775);
nand U31088 (N_31088,N_28207,N_25730);
or U31089 (N_31089,N_29459,N_29425);
nor U31090 (N_31090,N_28307,N_26611);
and U31091 (N_31091,N_29686,N_27593);
nor U31092 (N_31092,N_29470,N_26369);
or U31093 (N_31093,N_28902,N_25283);
and U31094 (N_31094,N_27214,N_29079);
or U31095 (N_31095,N_26701,N_29978);
or U31096 (N_31096,N_26375,N_26438);
xnor U31097 (N_31097,N_28746,N_25977);
nor U31098 (N_31098,N_28573,N_28375);
nand U31099 (N_31099,N_27233,N_29462);
xor U31100 (N_31100,N_25793,N_26139);
xnor U31101 (N_31101,N_26580,N_26963);
nor U31102 (N_31102,N_26173,N_29987);
xnor U31103 (N_31103,N_29770,N_25806);
and U31104 (N_31104,N_28521,N_27699);
and U31105 (N_31105,N_29233,N_27071);
nand U31106 (N_31106,N_25271,N_28859);
xnor U31107 (N_31107,N_29552,N_25799);
nor U31108 (N_31108,N_25180,N_25885);
xor U31109 (N_31109,N_25625,N_27365);
nand U31110 (N_31110,N_28826,N_25076);
and U31111 (N_31111,N_25797,N_27252);
or U31112 (N_31112,N_27977,N_25085);
nor U31113 (N_31113,N_28872,N_25056);
nor U31114 (N_31114,N_26913,N_29853);
nor U31115 (N_31115,N_26493,N_25891);
xnor U31116 (N_31116,N_28592,N_29179);
or U31117 (N_31117,N_26548,N_26042);
and U31118 (N_31118,N_26592,N_25166);
and U31119 (N_31119,N_27225,N_26997);
or U31120 (N_31120,N_25705,N_29451);
or U31121 (N_31121,N_28862,N_25717);
xnor U31122 (N_31122,N_25546,N_28353);
and U31123 (N_31123,N_26073,N_25361);
nand U31124 (N_31124,N_28912,N_28031);
or U31125 (N_31125,N_27762,N_26651);
nand U31126 (N_31126,N_28024,N_25860);
nand U31127 (N_31127,N_25561,N_29711);
and U31128 (N_31128,N_26148,N_25771);
or U31129 (N_31129,N_25645,N_28999);
and U31130 (N_31130,N_26421,N_25893);
nand U31131 (N_31131,N_28292,N_27795);
nor U31132 (N_31132,N_27586,N_26164);
and U31133 (N_31133,N_29460,N_26340);
nand U31134 (N_31134,N_28802,N_26632);
nand U31135 (N_31135,N_28063,N_27622);
xor U31136 (N_31136,N_29898,N_28524);
nor U31137 (N_31137,N_27475,N_28042);
or U31138 (N_31138,N_29435,N_29413);
or U31139 (N_31139,N_27786,N_26729);
nor U31140 (N_31140,N_26218,N_25171);
or U31141 (N_31141,N_27905,N_26976);
xnor U31142 (N_31142,N_28810,N_25205);
or U31143 (N_31143,N_28599,N_29100);
nor U31144 (N_31144,N_27384,N_27925);
or U31145 (N_31145,N_26461,N_28295);
and U31146 (N_31146,N_29476,N_26321);
nor U31147 (N_31147,N_28883,N_25168);
xnor U31148 (N_31148,N_27642,N_27145);
xor U31149 (N_31149,N_27724,N_25853);
nand U31150 (N_31150,N_25229,N_27084);
and U31151 (N_31151,N_25491,N_29961);
nand U31152 (N_31152,N_26816,N_26107);
nand U31153 (N_31153,N_27232,N_25600);
nand U31154 (N_31154,N_27900,N_25995);
xor U31155 (N_31155,N_28070,N_27123);
nand U31156 (N_31156,N_29709,N_27357);
and U31157 (N_31157,N_25266,N_29403);
and U31158 (N_31158,N_28079,N_27313);
nor U31159 (N_31159,N_28132,N_29579);
nor U31160 (N_31160,N_28566,N_27682);
or U31161 (N_31161,N_26473,N_29348);
and U31162 (N_31162,N_27356,N_29870);
and U31163 (N_31163,N_25533,N_29405);
and U31164 (N_31164,N_28160,N_25880);
xor U31165 (N_31165,N_26105,N_29440);
and U31166 (N_31166,N_26802,N_25270);
or U31167 (N_31167,N_28654,N_26127);
nor U31168 (N_31168,N_25901,N_27748);
or U31169 (N_31169,N_27826,N_27158);
or U31170 (N_31170,N_25090,N_27230);
nand U31171 (N_31171,N_28298,N_25311);
nand U31172 (N_31172,N_28563,N_26414);
xor U31173 (N_31173,N_28218,N_26706);
nand U31174 (N_31174,N_25007,N_25016);
nand U31175 (N_31175,N_25164,N_25598);
or U31176 (N_31176,N_29576,N_29984);
nand U31177 (N_31177,N_26857,N_28866);
nor U31178 (N_31178,N_29353,N_25676);
nand U31179 (N_31179,N_26115,N_25408);
or U31180 (N_31180,N_27001,N_25998);
xnor U31181 (N_31181,N_28394,N_26209);
or U31182 (N_31182,N_27345,N_26478);
nor U31183 (N_31183,N_25663,N_27759);
nand U31184 (N_31184,N_27863,N_26402);
xnor U31185 (N_31185,N_27755,N_28028);
nor U31186 (N_31186,N_28170,N_28471);
or U31187 (N_31187,N_25404,N_25488);
and U31188 (N_31188,N_28865,N_27370);
xnor U31189 (N_31189,N_28083,N_26492);
xor U31190 (N_31190,N_25532,N_28919);
and U31191 (N_31191,N_28506,N_28868);
or U31192 (N_31192,N_27855,N_28843);
and U31193 (N_31193,N_25931,N_29025);
xor U31194 (N_31194,N_26659,N_27510);
or U31195 (N_31195,N_27643,N_28455);
xnor U31196 (N_31196,N_29567,N_29049);
or U31197 (N_31197,N_27068,N_25107);
or U31198 (N_31198,N_27927,N_27387);
or U31199 (N_31199,N_26675,N_25346);
nor U31200 (N_31200,N_26977,N_28698);
or U31201 (N_31201,N_27689,N_29626);
nand U31202 (N_31202,N_29419,N_27520);
or U31203 (N_31203,N_25163,N_29279);
and U31204 (N_31204,N_29894,N_27840);
or U31205 (N_31205,N_26829,N_25325);
xnor U31206 (N_31206,N_28490,N_26801);
xnor U31207 (N_31207,N_27245,N_25812);
or U31208 (N_31208,N_29272,N_25508);
or U31209 (N_31209,N_25659,N_28542);
nand U31210 (N_31210,N_29681,N_25410);
or U31211 (N_31211,N_29480,N_27660);
or U31212 (N_31212,N_27150,N_28985);
nor U31213 (N_31213,N_26296,N_25559);
nor U31214 (N_31214,N_25754,N_26602);
xor U31215 (N_31215,N_29102,N_28414);
xor U31216 (N_31216,N_28705,N_29306);
nand U31217 (N_31217,N_29128,N_25763);
and U31218 (N_31218,N_29602,N_28686);
nand U31219 (N_31219,N_27274,N_25894);
xor U31220 (N_31220,N_26367,N_27368);
or U31221 (N_31221,N_28992,N_26795);
or U31222 (N_31222,N_28076,N_27649);
nor U31223 (N_31223,N_28728,N_29125);
xor U31224 (N_31224,N_28526,N_28486);
xor U31225 (N_31225,N_25466,N_26320);
and U31226 (N_31226,N_28988,N_29202);
xnor U31227 (N_31227,N_25479,N_26444);
and U31228 (N_31228,N_25554,N_27539);
nor U31229 (N_31229,N_29022,N_29137);
or U31230 (N_31230,N_28117,N_29165);
nor U31231 (N_31231,N_27711,N_25419);
and U31232 (N_31232,N_25414,N_29225);
nand U31233 (N_31233,N_25131,N_29292);
xor U31234 (N_31234,N_26301,N_27565);
and U31235 (N_31235,N_27405,N_27854);
xnor U31236 (N_31236,N_29230,N_28468);
nand U31237 (N_31237,N_28102,N_28905);
or U31238 (N_31238,N_29078,N_25197);
nand U31239 (N_31239,N_25265,N_26597);
or U31240 (N_31240,N_29721,N_28923);
xnor U31241 (N_31241,N_28814,N_27060);
nor U31242 (N_31242,N_27938,N_29205);
and U31243 (N_31243,N_28660,N_29282);
nand U31244 (N_31244,N_26937,N_28969);
nand U31245 (N_31245,N_25846,N_25515);
nand U31246 (N_31246,N_26205,N_28561);
or U31247 (N_31247,N_29543,N_26550);
and U31248 (N_31248,N_26439,N_28454);
and U31249 (N_31249,N_29839,N_27992);
nor U31250 (N_31250,N_26151,N_25936);
nor U31251 (N_31251,N_29527,N_27870);
nand U31252 (N_31252,N_27503,N_27710);
or U31253 (N_31253,N_28673,N_27679);
xor U31254 (N_31254,N_25104,N_29386);
or U31255 (N_31255,N_26170,N_27174);
nor U31256 (N_31256,N_27235,N_28138);
xor U31257 (N_31257,N_26256,N_28556);
or U31258 (N_31258,N_29115,N_27047);
nor U31259 (N_31259,N_26695,N_26570);
nand U31260 (N_31260,N_26325,N_26307);
or U31261 (N_31261,N_28396,N_27987);
or U31262 (N_31262,N_27478,N_28519);
xor U31263 (N_31263,N_26647,N_26356);
nand U31264 (N_31264,N_28560,N_28466);
nor U31265 (N_31265,N_28360,N_25688);
nand U31266 (N_31266,N_26060,N_26133);
or U31267 (N_31267,N_29792,N_29488);
nand U31268 (N_31268,N_26360,N_25914);
or U31269 (N_31269,N_25839,N_25139);
or U31270 (N_31270,N_28926,N_25119);
xnor U31271 (N_31271,N_25652,N_27886);
or U31272 (N_31272,N_28272,N_27358);
nand U31273 (N_31273,N_26199,N_29039);
and U31274 (N_31274,N_28400,N_26059);
nor U31275 (N_31275,N_25451,N_28025);
xnor U31276 (N_31276,N_26243,N_25961);
and U31277 (N_31277,N_25627,N_27270);
xor U31278 (N_31278,N_26746,N_26513);
or U31279 (N_31279,N_26411,N_28469);
nor U31280 (N_31280,N_29715,N_26163);
or U31281 (N_31281,N_25584,N_27648);
xnor U31282 (N_31282,N_25286,N_27753);
nand U31283 (N_31283,N_29599,N_25664);
or U31284 (N_31284,N_29950,N_25386);
nand U31285 (N_31285,N_28853,N_27931);
nor U31286 (N_31286,N_28021,N_27026);
nor U31287 (N_31287,N_25526,N_26018);
or U31288 (N_31288,N_28109,N_29146);
nor U31289 (N_31289,N_29864,N_25693);
xnor U31290 (N_31290,N_27451,N_27077);
xnor U31291 (N_31291,N_29339,N_25363);
xor U31292 (N_31292,N_28149,N_28339);
nor U31293 (N_31293,N_25395,N_26919);
nor U31294 (N_31294,N_27553,N_26609);
nand U31295 (N_31295,N_29421,N_29618);
nand U31296 (N_31296,N_25889,N_28574);
or U31297 (N_31297,N_28478,N_25194);
nand U31298 (N_31298,N_25192,N_27734);
nor U31299 (N_31299,N_25632,N_25658);
nand U31300 (N_31300,N_28297,N_29720);
and U31301 (N_31301,N_27312,N_25332);
nand U31302 (N_31302,N_29677,N_28539);
nor U31303 (N_31303,N_25813,N_26217);
nand U31304 (N_31304,N_29203,N_28681);
nand U31305 (N_31305,N_26110,N_27783);
nor U31306 (N_31306,N_28832,N_26330);
nor U31307 (N_31307,N_25337,N_29390);
xnor U31308 (N_31308,N_25399,N_25591);
xnor U31309 (N_31309,N_29074,N_28834);
or U31310 (N_31310,N_29105,N_27278);
nor U31311 (N_31311,N_25349,N_26306);
or U31312 (N_31312,N_29206,N_26386);
nand U31313 (N_31313,N_27953,N_26827);
or U31314 (N_31314,N_26523,N_28441);
xor U31315 (N_31315,N_28015,N_25609);
and U31316 (N_31316,N_26122,N_27442);
or U31317 (N_31317,N_27994,N_29794);
nor U31318 (N_31318,N_25694,N_28453);
nor U31319 (N_31319,N_29185,N_29969);
or U31320 (N_31320,N_29638,N_27383);
or U31321 (N_31321,N_25538,N_26424);
or U31322 (N_31322,N_29904,N_27914);
nand U31323 (N_31323,N_26529,N_26040);
xnor U31324 (N_31324,N_26594,N_26775);
and U31325 (N_31325,N_26740,N_27053);
nand U31326 (N_31326,N_27629,N_27810);
nor U31327 (N_31327,N_25734,N_27043);
nor U31328 (N_31328,N_27025,N_29430);
or U31329 (N_31329,N_27818,N_28690);
and U31330 (N_31330,N_27752,N_28581);
nor U31331 (N_31331,N_27875,N_26923);
or U31332 (N_31332,N_29324,N_27823);
nand U31333 (N_31333,N_27486,N_25100);
nor U31334 (N_31334,N_25012,N_29122);
nor U31335 (N_31335,N_28336,N_25662);
or U31336 (N_31336,N_29630,N_26028);
nor U31337 (N_31337,N_26558,N_28143);
xor U31338 (N_31338,N_29053,N_29347);
and U31339 (N_31339,N_28017,N_26995);
xnor U31340 (N_31340,N_29734,N_29329);
nand U31341 (N_31341,N_29469,N_27791);
or U31342 (N_31342,N_25965,N_28337);
xnor U31343 (N_31343,N_28324,N_28732);
xnor U31344 (N_31344,N_29735,N_25550);
and U31345 (N_31345,N_28604,N_29896);
and U31346 (N_31346,N_28944,N_27191);
nor U31347 (N_31347,N_25227,N_29776);
and U31348 (N_31348,N_27794,N_29391);
xnor U31349 (N_31349,N_27821,N_29402);
and U31350 (N_31350,N_28721,N_25478);
nand U31351 (N_31351,N_26855,N_26980);
nand U31352 (N_31352,N_28606,N_29659);
and U31353 (N_31353,N_28252,N_26507);
nand U31354 (N_31354,N_26496,N_28393);
nor U31355 (N_31355,N_26897,N_25925);
nor U31356 (N_31356,N_27828,N_27530);
nor U31357 (N_31357,N_27869,N_26516);
xnor U31358 (N_31358,N_27498,N_28605);
xor U31359 (N_31359,N_28842,N_29490);
or U31360 (N_31360,N_27848,N_28181);
and U31361 (N_31361,N_28002,N_29038);
nor U31362 (N_31362,N_28103,N_27211);
and U31363 (N_31363,N_27701,N_28650);
or U31364 (N_31364,N_27489,N_27425);
nor U31365 (N_31365,N_27696,N_28036);
nand U31366 (N_31366,N_25362,N_25514);
nor U31367 (N_31367,N_26835,N_28634);
nand U31368 (N_31368,N_27099,N_25150);
xor U31369 (N_31369,N_29342,N_26931);
or U31370 (N_31370,N_26401,N_28148);
nor U31371 (N_31371,N_26538,N_26458);
nand U31372 (N_31372,N_25858,N_27694);
xnor U31373 (N_31373,N_26838,N_25215);
nor U31374 (N_31374,N_25201,N_25602);
or U31375 (N_31375,N_29723,N_28947);
xnor U31376 (N_31376,N_26957,N_29071);
or U31377 (N_31377,N_28374,N_26011);
xnor U31378 (N_31378,N_27566,N_27618);
xnor U31379 (N_31379,N_28366,N_29491);
nand U31380 (N_31380,N_28327,N_29639);
or U31381 (N_31381,N_25210,N_28667);
nor U31382 (N_31382,N_25391,N_27740);
nor U31383 (N_31383,N_26432,N_29895);
nand U31384 (N_31384,N_27893,N_25345);
and U31385 (N_31385,N_27858,N_25644);
xnor U31386 (N_31386,N_26665,N_25318);
xnor U31387 (N_31387,N_27320,N_28034);
nor U31388 (N_31388,N_28448,N_26564);
nor U31389 (N_31389,N_26255,N_29647);
nor U31390 (N_31390,N_29136,N_29166);
or U31391 (N_31391,N_25879,N_29992);
and U31392 (N_31392,N_26237,N_29151);
or U31393 (N_31393,N_27142,N_28957);
nand U31394 (N_31394,N_28288,N_27392);
and U31395 (N_31395,N_27972,N_25590);
nand U31396 (N_31396,N_29200,N_25666);
nand U31397 (N_31397,N_25030,N_25562);
or U31398 (N_31398,N_26982,N_27892);
or U31399 (N_31399,N_27491,N_25955);
nand U31400 (N_31400,N_26700,N_27471);
nand U31401 (N_31401,N_29791,N_28516);
nand U31402 (N_31402,N_29769,N_26654);
nand U31403 (N_31403,N_25678,N_28948);
nor U31404 (N_31404,N_25649,N_27122);
and U31405 (N_31405,N_29229,N_29588);
xor U31406 (N_31406,N_27663,N_25199);
or U31407 (N_31407,N_25156,N_26627);
xor U31408 (N_31408,N_29231,N_26698);
and U31409 (N_31409,N_26938,N_28773);
nand U31410 (N_31410,N_29933,N_29438);
and U31411 (N_31411,N_28760,N_28978);
nand U31412 (N_31412,N_29487,N_25101);
xnor U31413 (N_31413,N_28484,N_27088);
nand U31414 (N_31414,N_26971,N_28185);
xnor U31415 (N_31415,N_28066,N_29221);
xor U31416 (N_31416,N_26526,N_25583);
and U31417 (N_31417,N_28051,N_26193);
and U31418 (N_31418,N_28548,N_29764);
nor U31419 (N_31419,N_29087,N_27984);
xor U31420 (N_31420,N_27800,N_29442);
xor U31421 (N_31421,N_28043,N_27326);
nor U31422 (N_31422,N_26972,N_28649);
nand U31423 (N_31423,N_26766,N_25802);
and U31424 (N_31424,N_25416,N_27074);
xnor U31425 (N_31425,N_28823,N_25711);
xnor U31426 (N_31426,N_28666,N_28171);
nand U31427 (N_31427,N_27059,N_28567);
nand U31428 (N_31428,N_25665,N_25291);
xor U31429 (N_31429,N_29590,N_27062);
xnor U31430 (N_31430,N_29667,N_26944);
or U31431 (N_31431,N_29284,N_29323);
nor U31432 (N_31432,N_25761,N_27372);
nand U31433 (N_31433,N_28648,N_27157);
or U31434 (N_31434,N_28827,N_27163);
or U31435 (N_31435,N_27344,N_29457);
and U31436 (N_31436,N_29399,N_28535);
nor U31437 (N_31437,N_29070,N_28293);
and U31438 (N_31438,N_27141,N_29598);
and U31439 (N_31439,N_26648,N_29831);
or U31440 (N_31440,N_27093,N_26074);
nor U31441 (N_31441,N_25568,N_29365);
nor U31442 (N_31442,N_26615,N_25151);
or U31443 (N_31443,N_28460,N_28833);
xnor U31444 (N_31444,N_29513,N_26616);
nor U31445 (N_31445,N_27315,N_25714);
nor U31446 (N_31446,N_29620,N_25053);
nand U31447 (N_31447,N_26629,N_29380);
or U31448 (N_31448,N_27918,N_28159);
and U31449 (N_31449,N_26077,N_28014);
and U31450 (N_31450,N_28261,N_26383);
nand U31451 (N_31451,N_29923,N_28510);
and U31452 (N_31452,N_25031,N_27178);
xnor U31453 (N_31453,N_29669,N_27714);
nand U31454 (N_31454,N_26591,N_26536);
nor U31455 (N_31455,N_25041,N_28993);
and U31456 (N_31456,N_25141,N_25835);
xnor U31457 (N_31457,N_29222,N_29002);
nor U31458 (N_31458,N_28974,N_29167);
or U31459 (N_31459,N_29836,N_28627);
nand U31460 (N_31460,N_27537,N_26853);
nor U31461 (N_31461,N_27393,N_25619);
or U31462 (N_31462,N_25875,N_25177);
and U31463 (N_31463,N_25465,N_28246);
xnor U31464 (N_31464,N_25102,N_26062);
or U31465 (N_31465,N_27434,N_26259);
xnor U31466 (N_31466,N_28268,N_25556);
xor U31467 (N_31467,N_25475,N_28998);
nand U31468 (N_31468,N_28456,N_28659);
xnor U31469 (N_31469,N_28406,N_29359);
xnor U31470 (N_31470,N_29356,N_26843);
and U31471 (N_31471,N_27659,N_26390);
nor U31472 (N_31472,N_26617,N_25768);
nor U31473 (N_31473,N_25954,N_27507);
or U31474 (N_31474,N_25044,N_27493);
or U31475 (N_31475,N_29605,N_29592);
nor U31476 (N_31476,N_28886,N_27014);
nor U31477 (N_31477,N_26099,N_27655);
nand U31478 (N_31478,N_25035,N_29690);
and U31479 (N_31479,N_28897,N_25962);
or U31480 (N_31480,N_27427,N_27670);
or U31481 (N_31481,N_28505,N_25777);
nand U31482 (N_31482,N_25947,N_26849);
nor U31483 (N_31483,N_27763,N_27171);
or U31484 (N_31484,N_25579,N_29560);
xor U31485 (N_31485,N_25066,N_28482);
or U31486 (N_31486,N_27227,N_25203);
or U31487 (N_31487,N_29604,N_28994);
nor U31488 (N_31488,N_26799,N_26803);
xnor U31489 (N_31489,N_25445,N_29066);
nor U31490 (N_31490,N_25387,N_29613);
xnor U31491 (N_31491,N_29086,N_26486);
nand U31492 (N_31492,N_25857,N_26428);
or U31493 (N_31493,N_29651,N_26354);
nand U31494 (N_31494,N_29646,N_27654);
and U31495 (N_31495,N_26771,N_29262);
nor U31496 (N_31496,N_26208,N_26134);
and U31497 (N_31497,N_25825,N_25927);
and U31498 (N_31498,N_28198,N_29215);
xnor U31499 (N_31499,N_28640,N_26234);
nand U31500 (N_31500,N_26129,N_26003);
xnor U31501 (N_31501,N_27514,N_29097);
nand U31502 (N_31502,N_26649,N_26983);
or U31503 (N_31503,N_26883,N_28906);
xor U31504 (N_31504,N_29953,N_26793);
nand U31505 (N_31505,N_26103,N_28740);
and U31506 (N_31506,N_29549,N_29767);
nand U31507 (N_31507,N_29176,N_26549);
and U31508 (N_31508,N_25868,N_26418);
nand U31509 (N_31509,N_28038,N_29906);
or U31510 (N_31510,N_27346,N_29183);
or U31511 (N_31511,N_26231,N_27650);
xor U31512 (N_31512,N_29131,N_29362);
or U31513 (N_31513,N_29905,N_27928);
xnor U31514 (N_31514,N_26408,N_27275);
or U31515 (N_31515,N_27103,N_26377);
and U31516 (N_31516,N_28570,N_29917);
xor U31517 (N_31517,N_27409,N_29661);
nand U31518 (N_31518,N_28416,N_27435);
or U31519 (N_31519,N_26940,N_27873);
nor U31520 (N_31520,N_28642,N_28199);
nand U31521 (N_31521,N_26999,N_29878);
nand U31522 (N_31522,N_27333,N_27871);
and U31523 (N_31523,N_26206,N_27324);
nand U31524 (N_31524,N_29267,N_28515);
and U31525 (N_31525,N_25070,N_28260);
xnor U31526 (N_31526,N_29547,N_27965);
nand U31527 (N_31527,N_26547,N_28781);
xnor U31528 (N_31528,N_25138,N_29882);
and U31529 (N_31529,N_28503,N_28491);
or U31530 (N_31530,N_25450,N_26736);
and U31531 (N_31531,N_27601,N_25122);
nand U31532 (N_31532,N_28806,N_27626);
xor U31533 (N_31533,N_29307,N_26605);
and U31534 (N_31534,N_27827,N_29155);
nor U31535 (N_31535,N_26318,N_29856);
or U31536 (N_31536,N_25400,N_26735);
nor U31537 (N_31537,N_26593,N_26677);
xor U31538 (N_31538,N_28517,N_28237);
nor U31539 (N_31539,N_26366,N_28664);
or U31540 (N_31540,N_29506,N_28874);
nand U31541 (N_31541,N_25628,N_28582);
nor U31542 (N_31542,N_29455,N_26776);
or U31543 (N_31543,N_27613,N_27402);
nor U31544 (N_31544,N_27926,N_26882);
nand U31545 (N_31545,N_26832,N_26111);
and U31546 (N_31546,N_26657,N_27674);
or U31547 (N_31547,N_25577,N_27860);
nor U31548 (N_31548,N_25595,N_25458);
or U31549 (N_31549,N_27321,N_26628);
nand U31550 (N_31550,N_28930,N_26752);
nand U31551 (N_31551,N_28309,N_26483);
nand U31552 (N_31552,N_29363,N_26708);
nand U31553 (N_31553,N_29148,N_28191);
xnor U31554 (N_31554,N_28817,N_29493);
and U31555 (N_31555,N_26147,N_28157);
nand U31556 (N_31556,N_28889,N_26828);
nor U31557 (N_31557,N_28762,N_25152);
and U31558 (N_31558,N_29945,N_26058);
or U31559 (N_31559,N_26245,N_26637);
xnor U31560 (N_31560,N_26946,N_27577);
or U31561 (N_31561,N_29422,N_25943);
nor U31562 (N_31562,N_28921,N_27169);
and U31563 (N_31563,N_29031,N_25766);
nand U31564 (N_31564,N_28615,N_26577);
nor U31565 (N_31565,N_26431,N_25108);
xnor U31566 (N_31566,N_28914,N_26900);
or U31567 (N_31567,N_27215,N_26860);
nor U31568 (N_31568,N_27446,N_27096);
nand U31569 (N_31569,N_26069,N_26488);
xor U31570 (N_31570,N_26684,N_28765);
and U31571 (N_31571,N_29374,N_28433);
nand U31572 (N_31572,N_29044,N_29696);
nor U31573 (N_31573,N_25187,N_29886);
nor U31574 (N_31574,N_28977,N_28840);
xnor U31575 (N_31575,N_28662,N_27807);
nor U31576 (N_31576,N_29316,N_27182);
and U31577 (N_31577,N_28211,N_27687);
and U31578 (N_31578,N_28716,N_25767);
or U31579 (N_31579,N_28878,N_26914);
xnor U31580 (N_31580,N_25077,N_25274);
xor U31581 (N_31581,N_29035,N_25063);
nor U31582 (N_31582,N_29219,N_27414);
nor U31583 (N_31583,N_27363,N_29502);
xnor U31584 (N_31584,N_26094,N_29955);
xor U31585 (N_31585,N_26269,N_27746);
nor U31586 (N_31586,N_26921,N_29784);
nor U31587 (N_31587,N_29692,N_25358);
xor U31588 (N_31588,N_27947,N_25464);
xor U31589 (N_31589,N_25449,N_26166);
nor U31590 (N_31590,N_28090,N_27880);
xnor U31591 (N_31591,N_26954,N_27595);
nor U31592 (N_31592,N_27429,N_27415);
or U31593 (N_31593,N_26449,N_27444);
xnor U31594 (N_31594,N_26553,N_26379);
or U31595 (N_31595,N_27635,N_28382);
nor U31596 (N_31596,N_25380,N_25256);
or U31597 (N_31597,N_27690,N_27244);
and U31598 (N_31598,N_25498,N_27367);
and U31599 (N_31599,N_25939,N_26343);
nor U31600 (N_31600,N_26430,N_29346);
nor U31601 (N_31601,N_29445,N_29149);
and U31602 (N_31602,N_25327,N_28717);
and U31603 (N_31603,N_29737,N_26089);
nor U31604 (N_31604,N_26319,N_25251);
nand U31605 (N_31605,N_25620,N_25127);
xnor U31606 (N_31606,N_26314,N_28518);
or U31607 (N_31607,N_25441,N_26258);
xnor U31608 (N_31608,N_27653,N_27837);
and U31609 (N_31609,N_29198,N_27065);
xnor U31610 (N_31610,N_29068,N_29743);
or U31611 (N_31611,N_29559,N_28358);
or U31612 (N_31612,N_28987,N_28701);
nor U31613 (N_31613,N_27335,N_29623);
and U31614 (N_31614,N_29429,N_26633);
xnor U31615 (N_31615,N_28543,N_29045);
nand U31616 (N_31616,N_29981,N_27957);
and U31617 (N_31617,N_25018,N_29266);
and U31618 (N_31618,N_27527,N_27231);
or U31619 (N_31619,N_29532,N_28937);
or U31620 (N_31620,N_25423,N_26506);
xor U31621 (N_31621,N_25112,N_29909);
nand U31622 (N_31622,N_28115,N_28020);
nand U31623 (N_31623,N_26323,N_27686);
and U31624 (N_31624,N_28596,N_26355);
xnor U31625 (N_31625,N_29701,N_25681);
or U31626 (N_31626,N_25140,N_29627);
nand U31627 (N_31627,N_25117,N_25544);
nor U31628 (N_31628,N_28753,N_29088);
xor U31629 (N_31629,N_29170,N_25899);
nand U31630 (N_31630,N_25674,N_28059);
nor U31631 (N_31631,N_28735,N_25022);
xnor U31632 (N_31632,N_29253,N_25006);
nand U31633 (N_31633,N_28419,N_27447);
nor U31634 (N_31634,N_27359,N_26195);
xor U31635 (N_31635,N_29873,N_25817);
and U31636 (N_31636,N_27501,N_25991);
xor U31637 (N_31637,N_26203,N_29042);
and U31638 (N_31638,N_26491,N_27579);
nand U31639 (N_31639,N_29497,N_27535);
nor U31640 (N_31640,N_25381,N_29636);
nand U31641 (N_31641,N_26124,N_26568);
xnor U31642 (N_31642,N_27249,N_28395);
nand U31643 (N_31643,N_28464,N_27216);
xnor U31644 (N_31644,N_29507,N_28276);
nand U31645 (N_31645,N_27587,N_26014);
and U31646 (N_31646,N_25764,N_29048);
nor U31647 (N_31647,N_27203,N_27418);
and U31648 (N_31648,N_28316,N_29903);
xnor U31649 (N_31649,N_27879,N_27506);
or U31650 (N_31650,N_25397,N_25435);
nor U31651 (N_31651,N_25687,N_26393);
or U31652 (N_31652,N_29277,N_25779);
and U31653 (N_31653,N_25418,N_29473);
nor U31654 (N_31654,N_28269,N_29649);
or U31655 (N_31655,N_28435,N_26143);
xor U31656 (N_31656,N_26902,N_26233);
or U31657 (N_31657,N_27139,N_29239);
and U31658 (N_31658,N_25328,N_25124);
or U31659 (N_31659,N_25463,N_26324);
and U31660 (N_31660,N_29054,N_28608);
and U31661 (N_31661,N_27952,N_25737);
xor U31662 (N_31662,N_28409,N_28630);
or U31663 (N_31663,N_28445,N_27458);
nand U31664 (N_31664,N_25749,N_29089);
or U31665 (N_31665,N_25453,N_29843);
nor U31666 (N_31666,N_25287,N_26778);
nor U31667 (N_31667,N_29475,N_29084);
nand U31668 (N_31668,N_29204,N_28875);
xnor U31669 (N_31669,N_26879,N_28989);
and U31670 (N_31670,N_25567,N_25224);
and U31671 (N_31671,N_29037,N_25471);
xor U31672 (N_31672,N_27558,N_28737);
and U31673 (N_31673,N_28725,N_27408);
or U31674 (N_31674,N_25635,N_28341);
xor U31675 (N_31675,N_28217,N_25634);
nor U31676 (N_31676,N_29907,N_25062);
nand U31677 (N_31677,N_27339,N_27226);
xnor U31678 (N_31678,N_29918,N_26720);
nor U31679 (N_31679,N_25728,N_28651);
xor U31680 (N_31680,N_28144,N_26236);
nand U31681 (N_31681,N_28477,N_26175);
and U31682 (N_31682,N_25845,N_28100);
xor U31683 (N_31683,N_27256,N_27127);
xor U31684 (N_31684,N_25055,N_27105);
or U31685 (N_31685,N_28529,N_25873);
nor U31686 (N_31686,N_28597,N_27528);
and U31687 (N_31687,N_29650,N_26624);
and U31688 (N_31688,N_28788,N_29340);
nor U31689 (N_31689,N_26565,N_28465);
and U31690 (N_31690,N_26130,N_25157);
nand U31691 (N_31691,N_29256,N_25929);
xor U31692 (N_31692,N_26136,N_25989);
and U31693 (N_31693,N_29485,N_28458);
nor U31694 (N_31694,N_25869,N_28509);
or U31695 (N_31695,N_25218,N_29129);
nor U31696 (N_31696,N_26363,N_26097);
xor U31697 (N_31697,N_26067,N_28228);
and U31698 (N_31698,N_27721,N_28158);
or U31699 (N_31699,N_27351,N_26395);
xor U31700 (N_31700,N_27319,N_29278);
and U31701 (N_31701,N_29736,N_26230);
or U31702 (N_31702,N_25534,N_27877);
nor U31703 (N_31703,N_27771,N_26716);
or U31704 (N_31704,N_29261,N_27770);
and U31705 (N_31705,N_27443,N_27152);
or U31706 (N_31706,N_29057,N_27018);
or U31707 (N_31707,N_29501,N_27412);
nor U31708 (N_31708,N_28239,N_27325);
or U31709 (N_31709,N_27100,N_29837);
or U31710 (N_31710,N_26149,N_29822);
and U31711 (N_31711,N_26587,N_25170);
or U31712 (N_31712,N_27555,N_26238);
xnor U31713 (N_31713,N_25145,N_27956);
xnor U31714 (N_31714,N_27377,N_26283);
or U31715 (N_31715,N_26022,N_28893);
nor U31716 (N_31716,N_29589,N_27217);
nand U31717 (N_31717,N_26024,N_27288);
nor U31718 (N_31718,N_26479,N_25743);
nand U31719 (N_31719,N_25008,N_26669);
xnor U31720 (N_31720,N_27238,N_27991);
and U31721 (N_31721,N_28752,N_26476);
nor U31722 (N_31722,N_29302,N_26930);
or U31723 (N_31723,N_25228,N_28340);
nand U31724 (N_31724,N_29154,N_26986);
nor U31725 (N_31725,N_25382,N_28449);
or U31726 (N_31726,N_25497,N_27269);
nand U31727 (N_31727,N_27884,N_29184);
and U31728 (N_31728,N_26235,N_27082);
nand U31729 (N_31729,N_25433,N_26846);
and U31730 (N_31730,N_27834,N_27469);
and U31731 (N_31731,N_27168,N_29908);
and U31732 (N_31732,N_26023,N_28939);
nor U31733 (N_31733,N_29458,N_25871);
or U31734 (N_31734,N_25110,N_25585);
and U31735 (N_31735,N_29971,N_27808);
xnor U31736 (N_31736,N_28311,N_27289);
nor U31737 (N_31737,N_26985,N_27747);
or U31738 (N_31738,N_25158,N_29315);
or U31739 (N_31739,N_29410,N_28578);
xnor U31740 (N_31740,N_26618,N_25081);
and U31741 (N_31741,N_28497,N_26000);
or U31742 (N_31742,N_28687,N_25784);
nand U31743 (N_31743,N_25905,N_28917);
xor U31744 (N_31744,N_28098,N_28871);
xor U31745 (N_31745,N_26890,N_28544);
nor U31746 (N_31746,N_29061,N_29956);
xor U31747 (N_31747,N_26973,N_27989);
nor U31748 (N_31748,N_27390,N_26798);
nor U31749 (N_31749,N_26508,N_26313);
or U31750 (N_31750,N_29926,N_25915);
and U31751 (N_31751,N_27517,N_29524);
or U31752 (N_31752,N_26370,N_27106);
or U31753 (N_31753,N_26945,N_28306);
nor U31754 (N_31754,N_28216,N_25014);
or U31755 (N_31755,N_27332,N_26034);
nand U31756 (N_31756,N_26532,N_27632);
nand U31757 (N_31757,N_27955,N_25581);
nand U31758 (N_31758,N_27598,N_25569);
xnor U31759 (N_31759,N_26252,N_28472);
nand U31760 (N_31760,N_27705,N_26119);
nand U31761 (N_31761,N_25195,N_25862);
and U31762 (N_31762,N_25700,N_29665);
and U31763 (N_31763,N_26020,N_25483);
nand U31764 (N_31764,N_28287,N_29827);
xnor U31765 (N_31765,N_26464,N_25751);
xor U31766 (N_31766,N_27011,N_25255);
nor U31767 (N_31767,N_29246,N_28764);
or U31768 (N_31768,N_28691,N_25780);
xnor U31769 (N_31769,N_29393,N_25407);
and U31770 (N_31770,N_29927,N_26749);
and U31771 (N_31771,N_29643,N_27273);
and U31772 (N_31772,N_27352,N_28054);
or U31773 (N_31773,N_25086,N_25064);
or U31774 (N_31774,N_27888,N_28961);
and U31775 (N_31775,N_25039,N_26156);
nor U31776 (N_31776,N_26090,N_28120);
and U31777 (N_31777,N_29814,N_27246);
and U31778 (N_31778,N_27464,N_29985);
nand U31779 (N_31779,N_28620,N_26051);
xor U31780 (N_31780,N_25946,N_25219);
and U31781 (N_31781,N_26315,N_26087);
nor U31782 (N_31782,N_29111,N_27939);
nand U31783 (N_31783,N_27297,N_27020);
nor U31784 (N_31784,N_26644,N_28348);
or U31785 (N_31785,N_25172,N_26316);
xor U31786 (N_31786,N_29285,N_27591);
and U31787 (N_31787,N_26417,N_28671);
xor U31788 (N_31788,N_27202,N_26480);
and U31789 (N_31789,N_27098,N_25517);
or U31790 (N_31790,N_26873,N_29803);
nor U31791 (N_31791,N_28995,N_25486);
xor U31792 (N_31792,N_25856,N_27909);
nand U31793 (N_31793,N_26104,N_26165);
nand U31794 (N_31794,N_26734,N_27219);
and U31795 (N_31795,N_27039,N_27117);
nand U31796 (N_31796,N_27756,N_27801);
nand U31797 (N_31797,N_28317,N_26135);
or U31798 (N_31798,N_26704,N_29177);
and U31799 (N_31799,N_25133,N_29573);
or U31800 (N_31800,N_28580,N_29193);
nand U31801 (N_31801,N_26466,N_28800);
nor U31802 (N_31802,N_28575,N_26270);
and U31803 (N_31803,N_25029,N_29811);
or U31804 (N_31804,N_28495,N_29584);
nand U31805 (N_31805,N_28053,N_27086);
nor U31806 (N_31806,N_27571,N_29387);
nand U31807 (N_31807,N_29666,N_27657);
nand U31808 (N_31808,N_27842,N_26658);
nor U31809 (N_31809,N_29998,N_25855);
or U31810 (N_31810,N_28656,N_28986);
nor U31811 (N_31811,N_27614,N_27917);
or U31812 (N_31812,N_25401,N_26933);
nand U31813 (N_31813,N_27529,N_28595);
xnor U31814 (N_31814,N_28378,N_29158);
or U31815 (N_31815,N_25047,N_27986);
or U31816 (N_31816,N_25383,N_26789);
nor U31817 (N_31817,N_29544,N_26221);
or U31818 (N_31818,N_28289,N_28733);
nor U31819 (N_31819,N_26712,N_28867);
nand U31820 (N_31820,N_28744,N_25667);
and U31821 (N_31821,N_28555,N_25092);
or U31822 (N_31822,N_27343,N_25725);
xor U31823 (N_31823,N_27159,N_29865);
nor U31824 (N_31824,N_25631,N_27680);
and U31825 (N_31825,N_27364,N_28533);
and U31826 (N_31826,N_28572,N_26047);
or U31827 (N_31827,N_26275,N_25792);
nor U31828 (N_31828,N_28300,N_29744);
or U31829 (N_31829,N_26721,N_25296);
nand U31830 (N_31830,N_29986,N_25364);
nand U31831 (N_31831,N_28898,N_29201);
nand U31832 (N_31832,N_25505,N_28075);
xnor U31833 (N_31833,N_29979,N_27765);
xor U31834 (N_31834,N_25756,N_29228);
nor U31835 (N_31835,N_27970,N_25300);
nor U31836 (N_31836,N_29780,N_27683);
and U31837 (N_31837,N_26528,N_27822);
xnor U31838 (N_31838,N_28612,N_26472);
nor U31839 (N_31839,N_27034,N_26419);
nor U31840 (N_31840,N_29813,N_29190);
or U31841 (N_31841,N_27058,N_28027);
and U31842 (N_31842,N_26280,N_27737);
nand U31843 (N_31843,N_26126,N_26738);
or U31844 (N_31844,N_25828,N_28828);
nor U31845 (N_31845,N_28854,N_29311);
nor U31846 (N_31846,N_28104,N_26389);
xnor U31847 (N_31847,N_25755,N_25438);
xnor U31848 (N_31848,N_29093,N_25186);
nand U31849 (N_31849,N_28045,N_25083);
xnor U31850 (N_31850,N_29862,N_25892);
xnor U31851 (N_31851,N_27610,N_25626);
xor U31852 (N_31852,N_28938,N_25612);
and U31853 (N_31853,N_29752,N_28328);
and U31854 (N_31854,N_29437,N_29471);
and U31855 (N_31855,N_28789,N_28711);
nand U31856 (N_31856,N_28851,N_25459);
or U31857 (N_31857,N_27298,N_25421);
and U31858 (N_31858,N_25888,N_25648);
xnor U31859 (N_31859,N_27213,N_27920);
and U31860 (N_31860,N_28523,N_26007);
or U31861 (N_31861,N_26422,N_25692);
xnor U31862 (N_31862,N_25536,N_27008);
or U31863 (N_31863,N_28724,N_26796);
xnor U31864 (N_31864,N_26093,N_26742);
or U31865 (N_31865,N_25930,N_27080);
or U31866 (N_31866,N_27951,N_29426);
xnor U31867 (N_31867,N_28718,N_26223);
or U31868 (N_31868,N_29702,N_26224);
nand U31869 (N_31869,N_29495,N_27891);
xnor U31870 (N_31870,N_26515,N_27600);
nor U31871 (N_31871,N_27574,N_27248);
nor U31872 (N_31872,N_25356,N_29081);
xor U31873 (N_31873,N_27793,N_26276);
nand U31874 (N_31874,N_28623,N_25342);
or U31875 (N_31875,N_29286,N_28632);
or U31876 (N_31876,N_29877,N_28899);
or U31877 (N_31877,N_25079,N_25510);
xor U31878 (N_31878,N_27407,N_28584);
xor U31879 (N_31879,N_29749,N_28933);
nand U31880 (N_31880,N_29930,N_26435);
nand U31881 (N_31881,N_25398,N_25587);
or U31882 (N_31882,N_28747,N_29331);
nor U31883 (N_31883,N_28512,N_29902);
nand U31884 (N_31884,N_29564,N_27592);
and U31885 (N_31885,N_26500,N_27819);
xnor U31886 (N_31886,N_26477,N_26682);
or U31887 (N_31887,N_27607,N_28734);
and U31888 (N_31888,N_25144,N_29802);
and U31889 (N_31889,N_27306,N_26392);
xor U31890 (N_31890,N_26281,N_27745);
and U31891 (N_31891,N_29412,N_26831);
nor U31892 (N_31892,N_28118,N_25309);
and U31893 (N_31893,N_27260,N_28763);
nor U31894 (N_31894,N_27441,N_26811);
and U31895 (N_31895,N_29133,N_26871);
nor U31896 (N_31896,N_29116,N_25003);
xor U31897 (N_31897,N_28016,N_25722);
xnor U31898 (N_31898,N_25306,N_29914);
xor U31899 (N_31899,N_25365,N_26310);
and U31900 (N_31900,N_28863,N_29188);
nor U31901 (N_31901,N_26725,N_29706);
nor U31902 (N_31902,N_29925,N_26229);
nor U31903 (N_31903,N_27742,N_29449);
xnor U31904 (N_31904,N_28256,N_26183);
and U31905 (N_31905,N_27688,N_29673);
or U31906 (N_31906,N_26967,N_29510);
xnor U31907 (N_31907,N_25235,N_26640);
and U31908 (N_31908,N_29436,N_29655);
nand U31909 (N_31909,N_29884,N_29570);
and U31910 (N_31910,N_25830,N_29118);
xnor U31911 (N_31911,N_28831,N_27229);
or U31912 (N_31912,N_28407,N_26663);
or U31913 (N_31913,N_26586,N_27726);
xnor U31914 (N_31914,N_26922,N_29257);
or U31915 (N_31915,N_25622,N_28026);
or U31916 (N_31916,N_26326,N_26100);
xor U31917 (N_31917,N_25405,N_29563);
nand U31918 (N_31918,N_26212,N_26227);
nand U31919 (N_31919,N_28877,N_28329);
nand U31920 (N_31920,N_29361,N_25748);
xor U31921 (N_31921,N_26681,N_27396);
and U31922 (N_31922,N_26088,N_25434);
and U31923 (N_31923,N_28313,N_29947);
and U31924 (N_31924,N_25980,N_27299);
nand U31925 (N_31925,N_28532,N_28706);
xor U31926 (N_31926,N_27399,N_27255);
nand U31927 (N_31927,N_28071,N_25736);
nor U31928 (N_31928,N_26833,N_29990);
or U31929 (N_31929,N_25206,N_27220);
nand U31930 (N_31930,N_27533,N_26250);
or U31931 (N_31931,N_25966,N_26989);
xnor U31932 (N_31932,N_26485,N_28380);
nand U31933 (N_31933,N_27373,N_27208);
or U31934 (N_31934,N_25333,N_29382);
and U31935 (N_31935,N_26661,N_29309);
nor U31936 (N_31936,N_27946,N_27969);
xor U31937 (N_31937,N_25280,N_28633);
xor U31938 (N_31938,N_29997,N_25898);
xnor U31939 (N_31939,N_25747,N_29065);
xnor U31940 (N_31940,N_25940,N_29058);
or U31941 (N_31941,N_26189,N_29852);
nand U31942 (N_31942,N_26705,N_25069);
nor U31943 (N_31943,N_27064,N_28275);
nand U31944 (N_31944,N_26502,N_26947);
or U31945 (N_31945,N_25701,N_26396);
nor U31946 (N_31946,N_28401,N_27461);
nand U31947 (N_31947,N_28685,N_28183);
nand U31948 (N_31948,N_26686,N_27277);
nand U31949 (N_31949,N_25603,N_27266);
or U31950 (N_31950,N_27413,N_25874);
nand U31951 (N_31951,N_26055,N_28669);
and U31952 (N_31952,N_25633,N_29975);
nand U31953 (N_31953,N_25811,N_26072);
nor U31954 (N_31954,N_26885,N_25369);
nand U31955 (N_31955,N_25798,N_26579);
or U31956 (N_31956,N_25357,N_29529);
or U31957 (N_31957,N_29373,N_28614);
xnor U31958 (N_31958,N_25781,N_26274);
and U31959 (N_31959,N_29850,N_27331);
nor U31960 (N_31960,N_26936,N_29912);
or U31961 (N_31961,N_25089,N_29693);
nor U31962 (N_31962,N_25025,N_25833);
nor U31963 (N_31963,N_26204,N_26590);
or U31964 (N_31964,N_28129,N_29210);
nor U31965 (N_31965,N_26768,N_27761);
or U31966 (N_31966,N_26043,N_27190);
or U31967 (N_31967,N_29052,N_29828);
xnor U31968 (N_31968,N_27187,N_26797);
and U31969 (N_31969,N_28619,N_26387);
nand U31970 (N_31970,N_28494,N_27798);
or U31971 (N_31971,N_28048,N_29240);
xnor U31972 (N_31972,N_27116,N_29942);
or U31973 (N_31973,N_28846,N_25005);
or U31974 (N_31974,N_25213,N_25953);
and U31975 (N_31975,N_27508,N_27676);
xnor U31976 (N_31976,N_29857,N_27774);
nor U31977 (N_31977,N_26566,N_26265);
xnor U31978 (N_31978,N_27376,N_27567);
or U31979 (N_31979,N_25490,N_27933);
and U31980 (N_31980,N_29187,N_27228);
nor U31981 (N_31981,N_29121,N_29147);
nor U31982 (N_31982,N_27120,N_29866);
or U31983 (N_31983,N_26436,N_25691);
and U31984 (N_31984,N_29371,N_28751);
and U31985 (N_31985,N_25221,N_29625);
nor U31986 (N_31986,N_27815,N_27341);
and U31987 (N_31987,N_29801,N_29101);
nor U31988 (N_31988,N_28774,N_29556);
nor U31989 (N_31989,N_29258,N_25988);
nor U31990 (N_31990,N_25967,N_28141);
nor U31991 (N_31991,N_28775,N_25637);
or U31992 (N_31992,N_27572,N_26222);
and U31993 (N_31993,N_28720,N_25336);
nor U31994 (N_31994,N_27005,N_25443);
xor U31995 (N_31995,N_27811,N_27307);
or U31996 (N_31996,N_25249,N_26505);
xnor U31997 (N_31997,N_27616,N_28684);
nand U31998 (N_31998,N_28688,N_29196);
nand U31999 (N_31999,N_25501,N_25814);
nor U32000 (N_32000,N_28167,N_27007);
nand U32001 (N_32001,N_26877,N_28321);
nor U32002 (N_32002,N_25593,N_28646);
and U32003 (N_32003,N_26907,N_29270);
or U32004 (N_32004,N_29548,N_27999);
or U32005 (N_32005,N_29970,N_27223);
or U32006 (N_32006,N_27347,N_25480);
nor U32007 (N_32007,N_26949,N_28531);
or U32008 (N_32008,N_27395,N_25529);
nand U32009 (N_32009,N_27146,N_28479);
and U32010 (N_32010,N_27184,N_28708);
and U32011 (N_32011,N_25385,N_29739);
and U32012 (N_32012,N_29892,N_27573);
and U32013 (N_32013,N_28551,N_29017);
and U32014 (N_32014,N_26176,N_29606);
nand U32015 (N_32015,N_25153,N_29358);
xor U32016 (N_32016,N_29750,N_27125);
or U32017 (N_32017,N_28315,N_26807);
nand U32018 (N_32018,N_29243,N_26066);
and U32019 (N_32019,N_25109,N_25253);
nor U32020 (N_32020,N_25639,N_28193);
nand U32021 (N_32021,N_28759,N_27784);
nor U32022 (N_32022,N_28965,N_29809);
or U32023 (N_32023,N_28346,N_27218);
nor U32024 (N_32024,N_25881,N_27707);
nor U32025 (N_32025,N_28920,N_26162);
nor U32026 (N_32026,N_25038,N_29085);
xor U32027 (N_32027,N_29269,N_28136);
and U32028 (N_32028,N_25000,N_26676);
and U32029 (N_32029,N_27656,N_26850);
xnor U32030 (N_32030,N_26875,N_25589);
nor U32031 (N_32031,N_28037,N_28767);
nor U32032 (N_32032,N_28126,N_26118);
xnor U32033 (N_32033,N_25121,N_25516);
or U32034 (N_32034,N_28727,N_29525);
nor U32035 (N_32035,N_26872,N_25507);
nand U32036 (N_32036,N_26791,N_28501);
nor U32037 (N_32037,N_25563,N_29982);
nor U32038 (N_32038,N_26952,N_29444);
or U32039 (N_32039,N_26542,N_25447);
and U32040 (N_32040,N_27454,N_28852);
or U32041 (N_32041,N_26727,N_29040);
or U32042 (N_32042,N_28369,N_28847);
xnor U32043 (N_32043,N_29119,N_29404);
nor U32044 (N_32044,N_27559,N_29738);
or U32045 (N_32045,N_29273,N_27549);
and U32046 (N_32046,N_29954,N_25316);
nor U32047 (N_32047,N_29489,N_25818);
xnor U32048 (N_32048,N_26693,N_27186);
xor U32049 (N_32049,N_25244,N_26723);
nand U32050 (N_32050,N_26889,N_28625);
nand U32051 (N_32051,N_28428,N_25731);
or U32052 (N_32052,N_27124,N_25161);
or U32053 (N_32053,N_25723,N_28983);
nand U32054 (N_32054,N_29594,N_27404);
xor U32055 (N_32055,N_29929,N_28860);
or U32056 (N_32056,N_28766,N_26415);
xnor U32057 (N_32057,N_25504,N_26071);
or U32058 (N_32058,N_25650,N_26009);
and U32059 (N_32059,N_26576,N_28131);
xor U32060 (N_32060,N_29033,N_27910);
nand U32061 (N_32061,N_29409,N_29753);
and U32062 (N_32062,N_28200,N_29522);
xor U32063 (N_32063,N_28749,N_27293);
or U32064 (N_32064,N_29214,N_27615);
xor U32065 (N_32065,N_27083,N_28204);
and U32066 (N_32066,N_27118,N_25344);
and U32067 (N_32067,N_25233,N_27502);
or U32068 (N_32068,N_28231,N_26703);
and U32069 (N_32069,N_27009,N_27403);
xnor U32070 (N_32070,N_25223,N_29876);
and U32071 (N_32071,N_26347,N_27851);
xor U32072 (N_32072,N_26397,N_26794);
or U32073 (N_32073,N_27832,N_29401);
xor U32074 (N_32074,N_26848,N_28392);
and U32075 (N_32075,N_26030,N_27609);
nand U32076 (N_32076,N_29076,N_27604);
nand U32077 (N_32077,N_29104,N_25304);
and U32078 (N_32078,N_26335,N_29759);
nor U32079 (N_32079,N_27912,N_29889);
xor U32080 (N_32080,N_28220,N_27495);
nor U32081 (N_32081,N_27263,N_26116);
and U32082 (N_32082,N_29114,N_28156);
xnor U32083 (N_32083,N_25074,N_27353);
nand U32084 (N_32084,N_27121,N_28603);
or U32085 (N_32085,N_28099,N_27462);
nor U32086 (N_32086,N_25343,N_25285);
xnor U32087 (N_32087,N_28113,N_27175);
xor U32088 (N_32088,N_25165,N_26248);
nand U32089 (N_32089,N_29774,N_29067);
or U32090 (N_32090,N_25209,N_29901);
or U32091 (N_32091,N_27825,N_28891);
and U32092 (N_32092,N_25040,N_29847);
nor U32093 (N_32093,N_28018,N_28206);
nand U32094 (N_32094,N_29140,N_29248);
or U32095 (N_32095,N_28242,N_25646);
and U32096 (N_32096,N_25974,N_25917);
nor U32097 (N_32097,N_26125,N_28971);
or U32098 (N_32098,N_29612,N_27140);
and U32099 (N_32099,N_25446,N_29477);
nor U32100 (N_32100,N_29684,N_29932);
or U32101 (N_32101,N_25252,N_26880);
and U32102 (N_32102,N_27695,N_28547);
nand U32103 (N_32103,N_27716,N_25689);
xor U32104 (N_32104,N_27239,N_26638);
nor U32105 (N_32105,N_29173,N_27448);
or U32106 (N_32106,N_27743,N_27922);
xor U32107 (N_32107,N_27713,N_27051);
nor U32108 (N_32108,N_26287,N_25926);
or U32109 (N_32109,N_27861,N_27739);
or U32110 (N_32110,N_28255,N_26619);
xnor U32111 (N_32111,N_26405,N_27038);
nor U32112 (N_32112,N_27327,N_25805);
nand U32113 (N_32113,N_28188,N_28402);
nand U32114 (N_32114,N_27472,N_27431);
and U32115 (N_32115,N_29940,N_25472);
nand U32116 (N_32116,N_29028,N_29376);
xnor U32117 (N_32117,N_25710,N_29545);
nor U32118 (N_32118,N_27876,N_26263);
xnor U32119 (N_32119,N_29295,N_27360);
or U32120 (N_32120,N_25682,N_26145);
nand U32121 (N_32121,N_27976,N_27531);
nor U32122 (N_32122,N_28956,N_29396);
and U32123 (N_32123,N_29541,N_25807);
nand U32124 (N_32124,N_25565,N_29218);
and U32125 (N_32125,N_28991,N_28942);
nand U32126 (N_32126,N_29293,N_25432);
or U32127 (N_32127,N_25826,N_25640);
and U32128 (N_32128,N_26019,N_28935);
nor U32129 (N_32129,N_25267,N_29082);
and U32130 (N_32130,N_28424,N_26416);
or U32131 (N_32131,N_27473,N_25566);
nor U32132 (N_32132,N_26168,N_25758);
or U32133 (N_32133,N_27258,N_26581);
or U32134 (N_32134,N_27967,N_26152);
xnor U32135 (N_32135,N_29697,N_28085);
nor U32136 (N_32136,N_29733,N_28421);
and U32137 (N_32137,N_29213,N_26927);
nor U32138 (N_32138,N_25067,N_26460);
xor U32139 (N_32139,N_25557,N_25877);
nor U32140 (N_32140,N_29224,N_26481);
and U32141 (N_32141,N_27672,N_29758);
xor U32142 (N_32142,N_27845,N_28815);
nor U32143 (N_32143,N_27718,N_27983);
nand U32144 (N_32144,N_26825,N_27552);
or U32145 (N_32145,N_25757,N_26336);
nor U32146 (N_32146,N_26560,N_27323);
xor U32147 (N_32147,N_28541,N_28049);
nand U32148 (N_32148,N_26812,N_28125);
xor U32149 (N_32149,N_25115,N_26687);
nand U32150 (N_32150,N_27521,N_25440);
xnor U32151 (N_32151,N_26374,N_25951);
nand U32152 (N_32152,N_28301,N_28114);
xor U32153 (N_32153,N_27541,N_25651);
or U32154 (N_32154,N_27930,N_26932);
nor U32155 (N_32155,N_26861,N_28227);
xnor U32156 (N_32156,N_29825,N_25275);
nand U32157 (N_32157,N_27206,N_29575);
xor U32158 (N_32158,N_27722,N_27847);
nor U32159 (N_32159,N_27072,N_28391);
nor U32160 (N_32160,N_29846,N_27843);
nor U32161 (N_32161,N_26080,N_28676);
nand U32162 (N_32162,N_29874,N_26851);
and U32163 (N_32163,N_26561,N_28411);
or U32164 (N_32164,N_29110,N_25027);
and U32165 (N_32165,N_26821,N_26052);
or U32166 (N_32166,N_29439,N_27782);
xnor U32167 (N_32167,N_28359,N_28232);
xor U32168 (N_32168,N_29499,N_26818);
and U32169 (N_32169,N_28208,N_29157);
and U32170 (N_32170,N_26888,N_28161);
nand U32171 (N_32171,N_26010,N_29526);
nand U32172 (N_32172,N_28955,N_28709);
nor U32173 (N_32173,N_26786,N_29928);
nand U32174 (N_32174,N_27075,N_25742);
nand U32175 (N_32175,N_27222,N_27147);
nand U32176 (N_32176,N_25520,N_29517);
and U32177 (N_32177,N_25226,N_29591);
xnor U32178 (N_32178,N_29617,N_28219);
nand U32179 (N_32179,N_27330,N_29867);
or U32180 (N_32180,N_29922,N_27830);
nand U32181 (N_32181,N_29768,N_27645);
or U32182 (N_32182,N_26870,N_26353);
nor U32183 (N_32183,N_26642,N_28959);
and U32184 (N_32184,N_28973,N_26856);
and U32185 (N_32185,N_27916,N_28904);
nand U32186 (N_32186,N_28150,N_28493);
nand U32187 (N_32187,N_25578,N_25539);
nand U32188 (N_32188,N_25822,N_27703);
and U32189 (N_32189,N_28155,N_28975);
and U32190 (N_32190,N_25994,N_28249);
or U32191 (N_32191,N_25324,N_27056);
nand U32192 (N_32192,N_29974,N_29209);
nand U32193 (N_32193,N_29707,N_28743);
xor U32194 (N_32194,N_29117,N_27411);
nor U32195 (N_32195,N_25394,N_26185);
and U32196 (N_32196,N_27788,N_29628);
nand U32197 (N_32197,N_25924,N_29481);
or U32198 (N_32198,N_25247,N_28887);
xnor U32199 (N_32199,N_27936,N_29325);
or U32200 (N_32200,N_26965,N_25010);
nand U32201 (N_32201,N_25656,N_26001);
nor U32202 (N_32202,N_28082,N_27262);
and U32203 (N_32203,N_29531,N_27652);
nor U32204 (N_32204,N_25850,N_29254);
nand U32205 (N_32205,N_26820,N_25886);
xor U32206 (N_32206,N_29134,N_25696);
or U32207 (N_32207,N_28285,N_26683);
or U32208 (N_32208,N_28822,N_25716);
and U32209 (N_32209,N_25785,N_26186);
or U32210 (N_32210,N_26842,N_25876);
xor U32211 (N_32211,N_27484,N_29060);
or U32212 (N_32212,N_25050,N_27470);
xor U32213 (N_32213,N_28164,N_27137);
and U32214 (N_32214,N_29227,N_26685);
xnor U32215 (N_32215,N_27741,N_25919);
and U32216 (N_32216,N_29505,N_27156);
nor U32217 (N_32217,N_26260,N_25374);
xor U32218 (N_32218,N_26770,N_26991);
nor U32219 (N_32219,N_28621,N_27135);
nand U32220 (N_32220,N_28087,N_25615);
nand U32221 (N_32221,N_29568,N_26950);
or U32222 (N_32222,N_26988,N_29855);
and U32223 (N_32223,N_26039,N_26623);
nor U32224 (N_32224,N_27254,N_26065);
xnor U32225 (N_32225,N_26588,N_25272);
nand U32226 (N_32226,N_26892,N_29833);
xnor U32227 (N_32227,N_25231,N_28244);
xnor U32228 (N_32228,N_28483,N_25933);
and U32229 (N_32229,N_27885,N_27417);
xor U32230 (N_32230,N_29143,N_26755);
nand U32231 (N_32231,N_28549,N_27835);
or U32232 (N_32232,N_25935,N_27750);
nor U32233 (N_32233,N_26737,N_25744);
nor U32234 (N_32234,N_28383,N_28005);
and U32235 (N_32235,N_26064,N_26210);
or U32236 (N_32236,N_25979,N_25982);
xor U32237 (N_32237,N_28777,N_28908);
and U32238 (N_32238,N_27563,N_27457);
nand U32239 (N_32239,N_29826,N_26678);
and U32240 (N_32240,N_28589,N_25686);
nand U32241 (N_32241,N_27919,N_28590);
nor U32242 (N_32242,N_26578,N_29130);
nor U32243 (N_32243,N_26075,N_29450);
xor U32244 (N_32244,N_29854,N_27764);
nand U32245 (N_32245,N_27789,N_29075);
nor U32246 (N_32246,N_28077,N_26399);
or U32247 (N_32247,N_29314,N_27259);
or U32248 (N_32248,N_29680,N_29029);
xor U32249 (N_32249,N_29056,N_28434);
nand U32250 (N_32250,N_27570,N_28976);
nor U32251 (N_32251,N_28550,N_28379);
nand U32252 (N_32252,N_27291,N_26482);
and U32253 (N_32253,N_28089,N_28918);
or U32254 (N_32254,N_28213,N_25147);
nor U32255 (N_32255,N_27309,N_29806);
nand U32256 (N_32256,N_27831,N_25890);
nand U32257 (N_32257,N_29503,N_27205);
nand U32258 (N_32258,N_29782,N_29719);
and U32259 (N_32259,N_25315,N_28528);
and U32260 (N_32260,N_26881,N_25707);
nand U32261 (N_32261,N_26117,N_29212);
nand U32262 (N_32262,N_29754,N_28693);
or U32263 (N_32263,N_28140,N_28496);
nand U32264 (N_32264,N_28499,N_29367);
nor U32265 (N_32265,N_28088,N_29321);
or U32266 (N_32266,N_26688,N_27792);
nor U32267 (N_32267,N_27109,N_29335);
nor U32268 (N_32268,N_26732,N_28739);
nand U32269 (N_32269,N_28432,N_29294);
xor U32270 (N_32270,N_27379,N_27261);
and U32271 (N_32271,N_28245,N_26471);
or U32272 (N_32272,N_27055,N_25831);
nor U32273 (N_32273,N_26948,N_27468);
xnor U32274 (N_32274,N_26928,N_29486);
nor U32275 (N_32275,N_25740,N_26905);
and U32276 (N_32276,N_28958,N_26974);
nor U32277 (N_32277,N_28825,N_29610);
xor U32278 (N_32278,N_27308,N_29841);
or U32279 (N_32279,N_25481,N_28857);
nor U32280 (N_32280,N_25911,N_27164);
nor U32281 (N_32281,N_26339,N_29765);
and U32282 (N_32282,N_26996,N_26975);
or U32283 (N_32283,N_29090,N_27982);
or U32284 (N_32284,N_25248,N_28678);
or U32285 (N_32285,N_28655,N_25220);
or U32286 (N_32286,N_25467,N_27115);
xnor U32287 (N_32287,N_27015,N_26908);
nor U32288 (N_32288,N_25417,N_27633);
or U32289 (N_32289,N_28504,N_26380);
or U32290 (N_32290,N_29718,N_27998);
or U32291 (N_32291,N_27340,N_27908);
or U32292 (N_32292,N_29026,N_28856);
nor U32293 (N_32293,N_25971,N_29027);
and U32294 (N_32294,N_25305,N_27391);
nor U32295 (N_32295,N_25159,N_28357);
nor U32296 (N_32296,N_26333,N_27948);
and U32297 (N_32297,N_28443,N_29562);
nor U32298 (N_32298,N_26338,N_28032);
and U32299 (N_32299,N_27301,N_29714);
xor U32300 (N_32300,N_29055,N_25179);
and U32301 (N_32301,N_27181,N_25330);
xor U32302 (N_32302,N_29934,N_26171);
and U32303 (N_32303,N_29103,N_27511);
nor U32304 (N_32304,N_29247,N_26763);
or U32305 (N_32305,N_28284,N_29062);
nor U32306 (N_32306,N_25260,N_26573);
and U32307 (N_32307,N_27488,N_26451);
and U32308 (N_32308,N_25908,N_25582);
nor U32309 (N_32309,N_29141,N_28761);
nor U32310 (N_32310,N_29996,N_29312);
xnor U32311 (N_32311,N_25261,N_29967);
and U32312 (N_32312,N_26225,N_26969);
or U32313 (N_32313,N_25623,N_26085);
nor U32314 (N_32314,N_29674,N_27608);
nor U32315 (N_32315,N_27923,N_27935);
xnor U32316 (N_32316,N_26844,N_27817);
nor U32317 (N_32317,N_27692,N_27814);
xnor U32318 (N_32318,N_28703,N_28356);
and U32319 (N_32319,N_27108,N_26692);
xnor U32320 (N_32320,N_28290,N_27562);
xnor U32321 (N_32321,N_28271,N_29879);
and U32322 (N_32322,N_27981,N_29397);
xor U32323 (N_32323,N_25019,N_27063);
or U32324 (N_32324,N_26155,N_28426);
or U32325 (N_32325,N_29966,N_28569);
xnor U32326 (N_32326,N_29530,N_28644);
xor U32327 (N_32327,N_27113,N_26702);
nand U32328 (N_32328,N_28513,N_26442);
and U32329 (N_32329,N_25896,N_25735);
xor U32330 (N_32330,N_29829,N_25130);
nor U32331 (N_32331,N_28714,N_26331);
nand U32332 (N_32332,N_29858,N_26109);
or U32333 (N_32333,N_29941,N_28997);
and U32334 (N_32334,N_26990,N_27305);
and U32335 (N_32335,N_26968,N_25366);
xnor U32336 (N_32336,N_27385,N_26522);
nand U32337 (N_32337,N_29726,N_27697);
nor U32338 (N_32338,N_26298,N_25921);
nand U32339 (N_32339,N_26730,N_27032);
or U32340 (N_32340,N_25944,N_27881);
xnor U32341 (N_32341,N_29574,N_27749);
xnor U32342 (N_32342,N_27188,N_25624);
nand U32343 (N_32343,N_26865,N_28221);
and U32344 (N_32344,N_27394,N_27836);
or U32345 (N_32345,N_27779,N_26029);
and U32346 (N_32346,N_26468,N_26448);
nor U32347 (N_32347,N_26559,N_27803);
nand U32348 (N_32348,N_29169,N_25295);
nand U32349 (N_32349,N_27569,N_25973);
nand U32350 (N_32350,N_25331,N_25468);
nand U32351 (N_32351,N_25379,N_28257);
xor U32352 (N_32352,N_26765,N_27318);
nand U32353 (N_32353,N_25537,N_29250);
or U32354 (N_32354,N_25654,N_27898);
xnor U32355 (N_32355,N_27719,N_28966);
or U32356 (N_32356,N_29138,N_27603);
nand U32357 (N_32357,N_26653,N_29644);
nand U32358 (N_32358,N_25574,N_26239);
and U32359 (N_32359,N_25668,N_27974);
or U32360 (N_32360,N_25277,N_28885);
xnor U32361 (N_32361,N_28808,N_26660);
nand U32362 (N_32362,N_29431,N_29682);
nand U32363 (N_32363,N_29406,N_25952);
and U32364 (N_32364,N_25048,N_25553);
nand U32365 (N_32365,N_26348,N_28562);
and U32366 (N_32366,N_26524,N_25778);
nor U32367 (N_32367,N_25786,N_29483);
nand U32368 (N_32368,N_26987,N_29427);
and U32369 (N_32369,N_27017,N_26242);
and U32370 (N_32370,N_25135,N_27296);
and U32371 (N_32371,N_26874,N_25250);
xnor U32372 (N_32372,N_29593,N_28844);
nor U32373 (N_32373,N_29290,N_25630);
nand U32374 (N_32374,N_28153,N_27172);
nor U32375 (N_32375,N_26429,N_28758);
nand U32376 (N_32376,N_28184,N_28055);
and U32377 (N_32377,N_26300,N_28514);
or U32378 (N_32378,N_25866,N_29740);
nand U32379 (N_32379,N_27545,N_29663);
or U32380 (N_32380,N_27865,N_28683);
or U32381 (N_32381,N_25992,N_25597);
xor U32382 (N_32382,N_29276,N_26958);
or U32383 (N_32383,N_28960,N_26680);
or U32384 (N_32384,N_28352,N_28096);
xnor U32385 (N_32385,N_25103,N_27035);
nor U32386 (N_32386,N_28936,N_26490);
nor U32387 (N_32387,N_29189,N_27430);
and U32388 (N_32388,N_26404,N_29521);
or U32389 (N_32389,N_29345,N_26329);
nor U32390 (N_32390,N_27036,N_25937);
nand U32391 (N_32391,N_28675,N_25970);
xnor U32392 (N_32392,N_25299,N_26563);
xor U32393 (N_32393,N_28234,N_27781);
nor U32394 (N_32394,N_28901,N_28203);
nor U32395 (N_32395,N_28692,N_25198);
and U32396 (N_32396,N_27631,N_27513);
nor U32397 (N_32397,N_25095,N_29798);
and U32398 (N_32398,N_29379,N_27192);
or U32399 (N_32399,N_29041,N_29326);
nand U32400 (N_32400,N_29897,N_27736);
or U32401 (N_32401,N_27864,N_27757);
nand U32402 (N_32402,N_27432,N_28934);
nor U32403 (N_32403,N_26510,N_28741);
xnor U32404 (N_32404,N_28281,N_28900);
xnor U32405 (N_32405,N_28057,N_27276);
and U32406 (N_32406,N_26994,N_28065);
nand U32407 (N_32407,N_25360,N_27166);
nand U32408 (N_32408,N_25699,N_28387);
or U32409 (N_32409,N_25783,N_29328);
nor U32410 (N_32410,N_27061,N_25861);
xor U32411 (N_32411,N_26719,N_25787);
or U32412 (N_32412,N_27518,N_29823);
nand U32413 (N_32413,N_25409,N_25613);
xnor U32414 (N_32414,N_25677,N_25629);
or U32415 (N_32415,N_27915,N_25790);
nand U32416 (N_32416,N_26184,N_25960);
nor U32417 (N_32417,N_25068,N_26358);
and U32418 (N_32418,N_29418,N_26690);
xnor U32419 (N_32419,N_28122,N_29263);
xor U32420 (N_32420,N_28003,N_25427);
nand U32421 (N_32421,N_28006,N_29900);
nor U32422 (N_32422,N_28473,N_29633);
or U32423 (N_32423,N_28413,N_29880);
nor U32424 (N_32424,N_29668,N_28362);
nor U32425 (N_32425,N_29280,N_28251);
nor U32426 (N_32426,N_27143,N_26545);
xor U32427 (N_32427,N_29671,N_26288);
or U32428 (N_32428,N_28263,N_26423);
or U32429 (N_32429,N_29983,N_28553);
or U32430 (N_32430,N_25222,N_27605);
nand U32431 (N_32431,N_25167,N_25456);
nor U32432 (N_32432,N_29761,N_29109);
or U32433 (N_32433,N_26350,N_25388);
and U32434 (N_32434,N_28748,N_27730);
or U32435 (N_32435,N_25422,N_29178);
nor U32436 (N_32436,N_25259,N_26261);
xnor U32437 (N_32437,N_25225,N_27911);
nand U32438 (N_32438,N_28429,N_26868);
or U32439 (N_32439,N_28730,N_27949);
nor U32440 (N_32440,N_27775,N_25670);
or U32441 (N_32441,N_29378,N_27087);
and U32442 (N_32442,N_25655,N_28731);
nor U32443 (N_32443,N_28629,N_26984);
nor U32444 (N_32444,N_28511,N_28820);
nor U32445 (N_32445,N_29988,N_27621);
nor U32446 (N_32446,N_26368,N_29242);
nand U32447 (N_32447,N_26915,N_26886);
and U32448 (N_32448,N_29135,N_29441);
and U32449 (N_32449,N_29360,N_28593);
and U32450 (N_32450,N_25321,N_27271);
nor U32451 (N_32451,N_29615,N_29654);
or U32452 (N_32452,N_26815,N_25610);
nand U32453 (N_32453,N_26557,N_26750);
and U32454 (N_32454,N_28062,N_27564);
nand U32455 (N_32455,N_27267,N_28225);
and U32456 (N_32456,N_29011,N_26626);
or U32457 (N_32457,N_26525,N_29756);
and U32458 (N_32458,N_25020,N_29094);
xor U32459 (N_32459,N_27283,N_29960);
and U32460 (N_32460,N_28351,N_26053);
or U32461 (N_32461,N_28480,N_29288);
nor U32462 (N_32462,N_28738,N_27022);
xor U32463 (N_32463,N_29533,N_27040);
or U32464 (N_32464,N_27237,N_28915);
nor U32465 (N_32465,N_29957,N_29890);
xnor U32466 (N_32466,N_25990,N_25829);
and U32467 (N_32467,N_25181,N_27354);
xor U32468 (N_32468,N_27073,N_27973);
nor U32469 (N_32469,N_28557,N_26279);
xnor U32470 (N_32470,N_26862,N_28174);
and U32471 (N_32471,N_27651,N_26943);
nor U32472 (N_32472,N_27095,N_26157);
xnor U32473 (N_32473,N_27921,N_29962);
and U32474 (N_32474,N_26826,N_25254);
or U32475 (N_32475,N_29252,N_29641);
nand U32476 (N_32476,N_26582,N_26469);
and U32477 (N_32477,N_28951,N_25848);
and U32478 (N_32478,N_27646,N_25969);
or U32479 (N_32479,N_25993,N_27611);
and U32480 (N_32480,N_26079,N_25106);
or U32481 (N_32481,N_26845,N_25703);
xnor U32482 (N_32482,N_28600,N_28536);
nor U32483 (N_32483,N_26032,N_25903);
nor U32484 (N_32484,N_27971,N_28354);
nor U32485 (N_32485,N_26345,N_26096);
or U32486 (N_32486,N_29150,N_26759);
or U32487 (N_32487,N_25178,N_25245);
nor U32488 (N_32488,N_26978,N_29414);
xnor U32489 (N_32489,N_27302,N_29557);
xor U32490 (N_32490,N_28347,N_26718);
nor U32491 (N_32491,N_27778,N_25021);
nand U32492 (N_32492,N_27630,N_28858);
xor U32493 (N_32493,N_25431,N_29994);
xnor U32494 (N_32494,N_28700,N_28000);
and U32495 (N_32495,N_25524,N_25576);
nor U32496 (N_32496,N_27010,N_25420);
or U32497 (N_32497,N_27406,N_28388);
and U32498 (N_32498,N_28911,N_26455);
nor U32499 (N_32499,N_25959,N_25444);
and U32500 (N_32500,N_29004,N_27810);
and U32501 (N_32501,N_29907,N_25401);
or U32502 (N_32502,N_26714,N_26893);
nor U32503 (N_32503,N_27205,N_29054);
or U32504 (N_32504,N_27724,N_29656);
xnor U32505 (N_32505,N_27293,N_29751);
xnor U32506 (N_32506,N_28927,N_27173);
and U32507 (N_32507,N_28306,N_28127);
nand U32508 (N_32508,N_27912,N_26000);
nand U32509 (N_32509,N_28273,N_27719);
and U32510 (N_32510,N_29703,N_29430);
nor U32511 (N_32511,N_26778,N_26611);
and U32512 (N_32512,N_29782,N_26254);
xor U32513 (N_32513,N_29634,N_28189);
nor U32514 (N_32514,N_29916,N_29773);
or U32515 (N_32515,N_26527,N_26779);
xor U32516 (N_32516,N_28995,N_28160);
nor U32517 (N_32517,N_29093,N_28183);
xnor U32518 (N_32518,N_27690,N_29655);
xor U32519 (N_32519,N_28140,N_29839);
xnor U32520 (N_32520,N_28037,N_29820);
nand U32521 (N_32521,N_27995,N_27563);
and U32522 (N_32522,N_27154,N_25925);
nor U32523 (N_32523,N_27036,N_28011);
nand U32524 (N_32524,N_27733,N_27929);
nand U32525 (N_32525,N_25706,N_25311);
nor U32526 (N_32526,N_27858,N_25994);
nor U32527 (N_32527,N_27640,N_29254);
or U32528 (N_32528,N_26145,N_27368);
or U32529 (N_32529,N_29153,N_26744);
nand U32530 (N_32530,N_28812,N_28357);
xnor U32531 (N_32531,N_27645,N_28265);
nand U32532 (N_32532,N_28523,N_28051);
xor U32533 (N_32533,N_28428,N_25346);
and U32534 (N_32534,N_26870,N_29849);
nor U32535 (N_32535,N_25926,N_27049);
and U32536 (N_32536,N_25110,N_28658);
or U32537 (N_32537,N_27353,N_26166);
xor U32538 (N_32538,N_29893,N_29124);
xnor U32539 (N_32539,N_25023,N_27853);
xor U32540 (N_32540,N_26453,N_26503);
or U32541 (N_32541,N_29032,N_26075);
nand U32542 (N_32542,N_25113,N_27839);
nor U32543 (N_32543,N_26884,N_27439);
xor U32544 (N_32544,N_28686,N_29321);
xnor U32545 (N_32545,N_29961,N_26790);
xor U32546 (N_32546,N_25142,N_25758);
nor U32547 (N_32547,N_28576,N_28783);
and U32548 (N_32548,N_26757,N_29729);
nand U32549 (N_32549,N_25548,N_25421);
xnor U32550 (N_32550,N_27848,N_29410);
nand U32551 (N_32551,N_28240,N_25288);
and U32552 (N_32552,N_26427,N_28263);
or U32553 (N_32553,N_29313,N_26404);
nand U32554 (N_32554,N_28423,N_27433);
and U32555 (N_32555,N_29691,N_26927);
or U32556 (N_32556,N_25476,N_29782);
and U32557 (N_32557,N_26866,N_28118);
nor U32558 (N_32558,N_28483,N_28953);
and U32559 (N_32559,N_29678,N_27514);
or U32560 (N_32560,N_28374,N_26003);
xnor U32561 (N_32561,N_27849,N_25762);
and U32562 (N_32562,N_27879,N_29037);
or U32563 (N_32563,N_27342,N_28526);
nand U32564 (N_32564,N_28470,N_29265);
or U32565 (N_32565,N_25407,N_26887);
xnor U32566 (N_32566,N_28094,N_26910);
xnor U32567 (N_32567,N_27791,N_25011);
xor U32568 (N_32568,N_27931,N_27631);
nand U32569 (N_32569,N_26747,N_27325);
nor U32570 (N_32570,N_25951,N_26902);
and U32571 (N_32571,N_28611,N_26747);
nand U32572 (N_32572,N_26355,N_25862);
nand U32573 (N_32573,N_29255,N_25335);
or U32574 (N_32574,N_25821,N_29533);
nor U32575 (N_32575,N_25305,N_28073);
and U32576 (N_32576,N_28073,N_29703);
or U32577 (N_32577,N_27765,N_25083);
xor U32578 (N_32578,N_27147,N_25233);
and U32579 (N_32579,N_28024,N_29009);
and U32580 (N_32580,N_29906,N_27307);
nand U32581 (N_32581,N_26417,N_29523);
nand U32582 (N_32582,N_28589,N_29337);
or U32583 (N_32583,N_27918,N_29270);
or U32584 (N_32584,N_25040,N_28991);
nand U32585 (N_32585,N_25781,N_29688);
and U32586 (N_32586,N_25210,N_26475);
nor U32587 (N_32587,N_25841,N_26506);
nand U32588 (N_32588,N_25985,N_28606);
nand U32589 (N_32589,N_28317,N_27986);
or U32590 (N_32590,N_28677,N_27733);
or U32591 (N_32591,N_25432,N_27324);
nand U32592 (N_32592,N_29244,N_28152);
nor U32593 (N_32593,N_28304,N_25018);
nand U32594 (N_32594,N_29975,N_28347);
xor U32595 (N_32595,N_29326,N_28415);
xor U32596 (N_32596,N_25714,N_29543);
nor U32597 (N_32597,N_29796,N_27119);
and U32598 (N_32598,N_27966,N_27972);
or U32599 (N_32599,N_28509,N_28972);
nor U32600 (N_32600,N_25529,N_29754);
or U32601 (N_32601,N_28130,N_27786);
and U32602 (N_32602,N_27312,N_28650);
xor U32603 (N_32603,N_26224,N_27231);
or U32604 (N_32604,N_25226,N_25436);
or U32605 (N_32605,N_28399,N_26661);
nor U32606 (N_32606,N_28020,N_26748);
or U32607 (N_32607,N_29266,N_29307);
nand U32608 (N_32608,N_26456,N_29902);
or U32609 (N_32609,N_26945,N_27682);
xor U32610 (N_32610,N_29888,N_28879);
nand U32611 (N_32611,N_28700,N_25100);
and U32612 (N_32612,N_27890,N_29945);
nand U32613 (N_32613,N_25400,N_25248);
xor U32614 (N_32614,N_26249,N_26981);
or U32615 (N_32615,N_27911,N_26370);
and U32616 (N_32616,N_25168,N_26375);
and U32617 (N_32617,N_29347,N_26352);
nor U32618 (N_32618,N_25646,N_27806);
xor U32619 (N_32619,N_29341,N_29600);
xnor U32620 (N_32620,N_28460,N_27783);
nor U32621 (N_32621,N_25800,N_28307);
and U32622 (N_32622,N_29616,N_29477);
nand U32623 (N_32623,N_29014,N_26260);
xor U32624 (N_32624,N_26512,N_26016);
nand U32625 (N_32625,N_27202,N_28074);
xnor U32626 (N_32626,N_26775,N_25595);
nand U32627 (N_32627,N_25360,N_26498);
nor U32628 (N_32628,N_26185,N_25462);
nor U32629 (N_32629,N_25036,N_28714);
and U32630 (N_32630,N_29964,N_28672);
nor U32631 (N_32631,N_25629,N_27800);
nand U32632 (N_32632,N_25582,N_28071);
and U32633 (N_32633,N_29460,N_27531);
and U32634 (N_32634,N_25055,N_26852);
nand U32635 (N_32635,N_25887,N_25963);
xnor U32636 (N_32636,N_28302,N_26113);
xnor U32637 (N_32637,N_29014,N_26848);
nand U32638 (N_32638,N_27864,N_26796);
nor U32639 (N_32639,N_29120,N_25090);
and U32640 (N_32640,N_27447,N_29097);
or U32641 (N_32641,N_28366,N_29375);
and U32642 (N_32642,N_28102,N_27161);
xor U32643 (N_32643,N_26312,N_25552);
xor U32644 (N_32644,N_25519,N_28784);
or U32645 (N_32645,N_29540,N_29527);
nand U32646 (N_32646,N_25282,N_26693);
nand U32647 (N_32647,N_28348,N_27476);
or U32648 (N_32648,N_26158,N_26375);
nor U32649 (N_32649,N_28382,N_27126);
or U32650 (N_32650,N_25307,N_27153);
nand U32651 (N_32651,N_25574,N_29191);
nor U32652 (N_32652,N_25727,N_25121);
or U32653 (N_32653,N_25263,N_25106);
nand U32654 (N_32654,N_26674,N_25487);
xor U32655 (N_32655,N_25711,N_29852);
xor U32656 (N_32656,N_28096,N_28691);
nor U32657 (N_32657,N_27889,N_25553);
xor U32658 (N_32658,N_26876,N_25391);
or U32659 (N_32659,N_28293,N_28567);
and U32660 (N_32660,N_27081,N_29590);
and U32661 (N_32661,N_26838,N_29007);
xnor U32662 (N_32662,N_29307,N_25084);
nor U32663 (N_32663,N_27802,N_28648);
xnor U32664 (N_32664,N_29828,N_27984);
xnor U32665 (N_32665,N_25833,N_28393);
and U32666 (N_32666,N_25744,N_27540);
and U32667 (N_32667,N_25028,N_29882);
nor U32668 (N_32668,N_26464,N_25635);
nor U32669 (N_32669,N_29661,N_26364);
nor U32670 (N_32670,N_28859,N_26521);
xnor U32671 (N_32671,N_26407,N_27878);
nor U32672 (N_32672,N_26290,N_26838);
nor U32673 (N_32673,N_28346,N_25728);
nand U32674 (N_32674,N_29851,N_29354);
or U32675 (N_32675,N_29446,N_27664);
xor U32676 (N_32676,N_26155,N_26299);
nand U32677 (N_32677,N_29660,N_27019);
and U32678 (N_32678,N_26746,N_27321);
nand U32679 (N_32679,N_29025,N_25313);
xor U32680 (N_32680,N_29721,N_25885);
nor U32681 (N_32681,N_28803,N_28753);
or U32682 (N_32682,N_25776,N_27886);
nor U32683 (N_32683,N_29695,N_29630);
nand U32684 (N_32684,N_27871,N_25465);
nand U32685 (N_32685,N_29328,N_28484);
nor U32686 (N_32686,N_29222,N_29261);
nand U32687 (N_32687,N_27718,N_27618);
or U32688 (N_32688,N_26534,N_25209);
and U32689 (N_32689,N_29490,N_27488);
xnor U32690 (N_32690,N_29226,N_26271);
or U32691 (N_32691,N_25705,N_29481);
and U32692 (N_32692,N_28675,N_28024);
and U32693 (N_32693,N_29707,N_27557);
or U32694 (N_32694,N_29478,N_27752);
nand U32695 (N_32695,N_26534,N_29974);
or U32696 (N_32696,N_26975,N_28492);
nor U32697 (N_32697,N_25874,N_27407);
nor U32698 (N_32698,N_27373,N_26773);
nand U32699 (N_32699,N_29807,N_27847);
and U32700 (N_32700,N_27091,N_25743);
or U32701 (N_32701,N_29058,N_27691);
xor U32702 (N_32702,N_25497,N_29839);
xor U32703 (N_32703,N_28162,N_27039);
nand U32704 (N_32704,N_25177,N_29380);
nand U32705 (N_32705,N_26406,N_29929);
and U32706 (N_32706,N_29061,N_28819);
nand U32707 (N_32707,N_27712,N_29695);
xnor U32708 (N_32708,N_28358,N_27210);
or U32709 (N_32709,N_29771,N_28858);
nand U32710 (N_32710,N_25888,N_28065);
nor U32711 (N_32711,N_29082,N_28272);
nor U32712 (N_32712,N_28876,N_29372);
nor U32713 (N_32713,N_28088,N_25531);
xor U32714 (N_32714,N_25378,N_26760);
xor U32715 (N_32715,N_29198,N_29788);
nor U32716 (N_32716,N_29756,N_25132);
nand U32717 (N_32717,N_28635,N_29631);
or U32718 (N_32718,N_28536,N_29500);
or U32719 (N_32719,N_29957,N_25275);
and U32720 (N_32720,N_29004,N_26490);
xor U32721 (N_32721,N_25887,N_29474);
nand U32722 (N_32722,N_26692,N_26371);
and U32723 (N_32723,N_26069,N_28217);
nand U32724 (N_32724,N_29810,N_25965);
nor U32725 (N_32725,N_29245,N_28470);
or U32726 (N_32726,N_25232,N_28193);
xnor U32727 (N_32727,N_25221,N_28209);
and U32728 (N_32728,N_25792,N_29764);
or U32729 (N_32729,N_25184,N_26294);
nor U32730 (N_32730,N_26360,N_25395);
nor U32731 (N_32731,N_29000,N_28889);
xnor U32732 (N_32732,N_26261,N_26203);
nor U32733 (N_32733,N_27504,N_29288);
and U32734 (N_32734,N_28553,N_26996);
xor U32735 (N_32735,N_26795,N_25682);
nand U32736 (N_32736,N_27851,N_25091);
nand U32737 (N_32737,N_26784,N_28587);
nand U32738 (N_32738,N_25217,N_25360);
nor U32739 (N_32739,N_26818,N_26805);
nand U32740 (N_32740,N_27623,N_28938);
and U32741 (N_32741,N_25905,N_28884);
and U32742 (N_32742,N_25210,N_29844);
or U32743 (N_32743,N_29943,N_29215);
or U32744 (N_32744,N_25720,N_25054);
xnor U32745 (N_32745,N_28101,N_29395);
or U32746 (N_32746,N_26865,N_25922);
nor U32747 (N_32747,N_25033,N_26622);
or U32748 (N_32748,N_29376,N_28496);
or U32749 (N_32749,N_29318,N_27149);
or U32750 (N_32750,N_25456,N_28120);
or U32751 (N_32751,N_25943,N_26657);
nand U32752 (N_32752,N_26045,N_27173);
and U32753 (N_32753,N_29866,N_28411);
or U32754 (N_32754,N_25040,N_26166);
and U32755 (N_32755,N_26182,N_28479);
xnor U32756 (N_32756,N_25432,N_28875);
nand U32757 (N_32757,N_25900,N_27962);
nor U32758 (N_32758,N_26452,N_27649);
nand U32759 (N_32759,N_25172,N_29520);
xnor U32760 (N_32760,N_29090,N_29523);
and U32761 (N_32761,N_25951,N_29603);
and U32762 (N_32762,N_25177,N_26192);
nor U32763 (N_32763,N_27321,N_28893);
xor U32764 (N_32764,N_28129,N_25471);
xnor U32765 (N_32765,N_27458,N_27650);
or U32766 (N_32766,N_29785,N_27142);
nand U32767 (N_32767,N_29251,N_27747);
or U32768 (N_32768,N_27605,N_26167);
xnor U32769 (N_32769,N_26196,N_25202);
and U32770 (N_32770,N_29251,N_27000);
or U32771 (N_32771,N_27593,N_29884);
and U32772 (N_32772,N_27137,N_28970);
xor U32773 (N_32773,N_28310,N_26838);
xor U32774 (N_32774,N_28867,N_29044);
xnor U32775 (N_32775,N_27797,N_28172);
nand U32776 (N_32776,N_26166,N_28637);
xor U32777 (N_32777,N_25594,N_25271);
nor U32778 (N_32778,N_27889,N_28057);
nand U32779 (N_32779,N_26511,N_29172);
xnor U32780 (N_32780,N_25483,N_29234);
or U32781 (N_32781,N_27148,N_29866);
nand U32782 (N_32782,N_26638,N_25958);
nor U32783 (N_32783,N_29107,N_27146);
nor U32784 (N_32784,N_26276,N_27844);
nand U32785 (N_32785,N_29653,N_27846);
nor U32786 (N_32786,N_27385,N_28472);
or U32787 (N_32787,N_26419,N_26097);
nand U32788 (N_32788,N_28442,N_26273);
nor U32789 (N_32789,N_26618,N_26298);
or U32790 (N_32790,N_28987,N_25991);
or U32791 (N_32791,N_27613,N_29683);
and U32792 (N_32792,N_27578,N_25082);
nor U32793 (N_32793,N_27007,N_26973);
nor U32794 (N_32794,N_26761,N_26150);
nand U32795 (N_32795,N_28674,N_29265);
or U32796 (N_32796,N_27123,N_28152);
nor U32797 (N_32797,N_29728,N_29820);
or U32798 (N_32798,N_27666,N_29361);
or U32799 (N_32799,N_26772,N_26678);
and U32800 (N_32800,N_28667,N_29377);
xnor U32801 (N_32801,N_26420,N_26652);
xnor U32802 (N_32802,N_26018,N_28527);
nand U32803 (N_32803,N_25115,N_27782);
nand U32804 (N_32804,N_27864,N_26159);
nor U32805 (N_32805,N_25822,N_26779);
nand U32806 (N_32806,N_28267,N_28190);
and U32807 (N_32807,N_28794,N_27255);
nand U32808 (N_32808,N_26795,N_28639);
xnor U32809 (N_32809,N_26310,N_26200);
nand U32810 (N_32810,N_25104,N_28670);
nor U32811 (N_32811,N_29173,N_28864);
nor U32812 (N_32812,N_27593,N_27528);
and U32813 (N_32813,N_27437,N_29801);
nand U32814 (N_32814,N_29762,N_27505);
or U32815 (N_32815,N_25801,N_27942);
nand U32816 (N_32816,N_27486,N_27021);
nand U32817 (N_32817,N_27647,N_27677);
and U32818 (N_32818,N_26391,N_27674);
nor U32819 (N_32819,N_28027,N_27557);
or U32820 (N_32820,N_27629,N_25077);
and U32821 (N_32821,N_29040,N_27930);
nor U32822 (N_32822,N_28936,N_28777);
or U32823 (N_32823,N_29712,N_26613);
nor U32824 (N_32824,N_27183,N_28711);
nor U32825 (N_32825,N_25867,N_26895);
nand U32826 (N_32826,N_29539,N_29003);
nor U32827 (N_32827,N_29819,N_25194);
or U32828 (N_32828,N_29193,N_27340);
nor U32829 (N_32829,N_29235,N_28695);
nand U32830 (N_32830,N_29914,N_28211);
xnor U32831 (N_32831,N_26555,N_26549);
and U32832 (N_32832,N_27891,N_25680);
nand U32833 (N_32833,N_25401,N_29204);
nor U32834 (N_32834,N_25623,N_25202);
xor U32835 (N_32835,N_29769,N_27806);
nor U32836 (N_32836,N_25353,N_29300);
nand U32837 (N_32837,N_29274,N_29902);
nor U32838 (N_32838,N_28673,N_27626);
nor U32839 (N_32839,N_29430,N_27430);
and U32840 (N_32840,N_26148,N_26579);
or U32841 (N_32841,N_28453,N_28785);
or U32842 (N_32842,N_27415,N_29778);
nand U32843 (N_32843,N_27297,N_27409);
nand U32844 (N_32844,N_26961,N_27887);
or U32845 (N_32845,N_26907,N_25692);
nor U32846 (N_32846,N_26222,N_29688);
nor U32847 (N_32847,N_27774,N_25063);
nand U32848 (N_32848,N_25207,N_28963);
nor U32849 (N_32849,N_29454,N_27349);
nand U32850 (N_32850,N_27953,N_25036);
and U32851 (N_32851,N_25149,N_28888);
or U32852 (N_32852,N_29506,N_28677);
nor U32853 (N_32853,N_29003,N_28930);
xnor U32854 (N_32854,N_29764,N_28680);
nor U32855 (N_32855,N_28652,N_29382);
or U32856 (N_32856,N_25646,N_28983);
xor U32857 (N_32857,N_28456,N_26033);
nand U32858 (N_32858,N_27587,N_28440);
nand U32859 (N_32859,N_26030,N_28040);
nor U32860 (N_32860,N_29921,N_26991);
xor U32861 (N_32861,N_27183,N_26954);
nand U32862 (N_32862,N_29255,N_28037);
xor U32863 (N_32863,N_29413,N_27892);
or U32864 (N_32864,N_27952,N_25402);
and U32865 (N_32865,N_29269,N_25303);
nand U32866 (N_32866,N_26444,N_28804);
nand U32867 (N_32867,N_26237,N_25808);
xnor U32868 (N_32868,N_28735,N_25224);
nor U32869 (N_32869,N_25022,N_29626);
or U32870 (N_32870,N_25134,N_25731);
or U32871 (N_32871,N_28345,N_26689);
or U32872 (N_32872,N_28017,N_27600);
or U32873 (N_32873,N_26210,N_28020);
nand U32874 (N_32874,N_27856,N_25599);
nand U32875 (N_32875,N_26049,N_29953);
xnor U32876 (N_32876,N_25419,N_27437);
or U32877 (N_32877,N_27110,N_26644);
nor U32878 (N_32878,N_26797,N_25847);
nor U32879 (N_32879,N_26098,N_25421);
nand U32880 (N_32880,N_29198,N_26108);
or U32881 (N_32881,N_29271,N_26672);
nor U32882 (N_32882,N_29714,N_28423);
xnor U32883 (N_32883,N_28584,N_27900);
nand U32884 (N_32884,N_26961,N_29476);
or U32885 (N_32885,N_25776,N_29027);
nand U32886 (N_32886,N_25306,N_26573);
and U32887 (N_32887,N_29924,N_27008);
or U32888 (N_32888,N_25310,N_29438);
nor U32889 (N_32889,N_29145,N_25356);
nor U32890 (N_32890,N_27533,N_28465);
nor U32891 (N_32891,N_26428,N_29073);
or U32892 (N_32892,N_26633,N_29938);
or U32893 (N_32893,N_29820,N_25766);
nand U32894 (N_32894,N_27708,N_28991);
and U32895 (N_32895,N_27048,N_28083);
and U32896 (N_32896,N_27258,N_26853);
or U32897 (N_32897,N_26572,N_26457);
and U32898 (N_32898,N_27027,N_26707);
nor U32899 (N_32899,N_25732,N_25063);
and U32900 (N_32900,N_27713,N_27196);
or U32901 (N_32901,N_28914,N_25189);
nor U32902 (N_32902,N_29554,N_25525);
and U32903 (N_32903,N_27008,N_28064);
or U32904 (N_32904,N_29454,N_28851);
xor U32905 (N_32905,N_29997,N_27586);
xnor U32906 (N_32906,N_29033,N_29380);
or U32907 (N_32907,N_26217,N_27947);
nand U32908 (N_32908,N_27027,N_27312);
or U32909 (N_32909,N_27716,N_25284);
nor U32910 (N_32910,N_27401,N_28684);
or U32911 (N_32911,N_29606,N_27831);
nor U32912 (N_32912,N_25346,N_27157);
and U32913 (N_32913,N_28708,N_25208);
and U32914 (N_32914,N_29280,N_25323);
nor U32915 (N_32915,N_27477,N_28761);
nor U32916 (N_32916,N_25769,N_28751);
and U32917 (N_32917,N_27274,N_26752);
and U32918 (N_32918,N_28043,N_25260);
nor U32919 (N_32919,N_25445,N_27272);
nand U32920 (N_32920,N_28711,N_27571);
nand U32921 (N_32921,N_29522,N_28407);
and U32922 (N_32922,N_29931,N_28998);
xnor U32923 (N_32923,N_29470,N_26259);
and U32924 (N_32924,N_27774,N_27565);
nor U32925 (N_32925,N_25081,N_26153);
xor U32926 (N_32926,N_27134,N_29811);
nand U32927 (N_32927,N_27382,N_25040);
and U32928 (N_32928,N_25147,N_28713);
nand U32929 (N_32929,N_29030,N_27634);
nor U32930 (N_32930,N_28454,N_28602);
nor U32931 (N_32931,N_28801,N_25938);
xor U32932 (N_32932,N_29118,N_25975);
or U32933 (N_32933,N_28238,N_29342);
nand U32934 (N_32934,N_29867,N_25481);
or U32935 (N_32935,N_25744,N_29976);
nand U32936 (N_32936,N_28612,N_29076);
xnor U32937 (N_32937,N_26192,N_26816);
nand U32938 (N_32938,N_27246,N_28807);
xor U32939 (N_32939,N_26673,N_26602);
nand U32940 (N_32940,N_25631,N_27578);
and U32941 (N_32941,N_29933,N_25709);
or U32942 (N_32942,N_27534,N_27933);
or U32943 (N_32943,N_29095,N_28848);
nor U32944 (N_32944,N_27836,N_27401);
or U32945 (N_32945,N_25653,N_26639);
xnor U32946 (N_32946,N_25495,N_28375);
nand U32947 (N_32947,N_25321,N_25527);
and U32948 (N_32948,N_29216,N_25058);
or U32949 (N_32949,N_27652,N_27694);
and U32950 (N_32950,N_28866,N_27845);
or U32951 (N_32951,N_29588,N_25546);
nand U32952 (N_32952,N_27638,N_25579);
or U32953 (N_32953,N_25549,N_25773);
nor U32954 (N_32954,N_28338,N_26118);
nand U32955 (N_32955,N_28353,N_27438);
nor U32956 (N_32956,N_25495,N_27747);
xnor U32957 (N_32957,N_25336,N_25417);
xor U32958 (N_32958,N_28935,N_27848);
xor U32959 (N_32959,N_27182,N_28371);
and U32960 (N_32960,N_26283,N_25017);
or U32961 (N_32961,N_28206,N_27883);
nand U32962 (N_32962,N_27381,N_28199);
nand U32963 (N_32963,N_27639,N_26833);
or U32964 (N_32964,N_26933,N_28394);
nand U32965 (N_32965,N_27046,N_26907);
nor U32966 (N_32966,N_28163,N_28158);
nand U32967 (N_32967,N_27770,N_25716);
and U32968 (N_32968,N_25071,N_26432);
nand U32969 (N_32969,N_29152,N_29594);
nand U32970 (N_32970,N_28524,N_29529);
or U32971 (N_32971,N_25048,N_27341);
or U32972 (N_32972,N_28645,N_28260);
xor U32973 (N_32973,N_27803,N_26029);
nor U32974 (N_32974,N_29630,N_25129);
or U32975 (N_32975,N_28291,N_26524);
nor U32976 (N_32976,N_29884,N_26118);
nand U32977 (N_32977,N_27044,N_26480);
or U32978 (N_32978,N_26702,N_25960);
nand U32979 (N_32979,N_26125,N_29802);
nor U32980 (N_32980,N_26940,N_26390);
nor U32981 (N_32981,N_29743,N_27499);
or U32982 (N_32982,N_29949,N_28496);
nor U32983 (N_32983,N_26981,N_26191);
or U32984 (N_32984,N_27633,N_29921);
xnor U32985 (N_32985,N_25914,N_27894);
xnor U32986 (N_32986,N_27938,N_29771);
nor U32987 (N_32987,N_29973,N_28423);
or U32988 (N_32988,N_25716,N_26850);
nor U32989 (N_32989,N_29101,N_27971);
and U32990 (N_32990,N_29280,N_26502);
xor U32991 (N_32991,N_26282,N_28493);
and U32992 (N_32992,N_29504,N_29958);
xor U32993 (N_32993,N_26930,N_28573);
or U32994 (N_32994,N_26921,N_28242);
or U32995 (N_32995,N_26468,N_28140);
and U32996 (N_32996,N_26451,N_28272);
nand U32997 (N_32997,N_25531,N_29475);
nand U32998 (N_32998,N_26212,N_27598);
nor U32999 (N_32999,N_29920,N_28882);
or U33000 (N_33000,N_25186,N_28729);
and U33001 (N_33001,N_29909,N_29241);
xor U33002 (N_33002,N_25309,N_27194);
xnor U33003 (N_33003,N_29509,N_27744);
or U33004 (N_33004,N_26050,N_29174);
or U33005 (N_33005,N_28608,N_28829);
and U33006 (N_33006,N_25188,N_25704);
nor U33007 (N_33007,N_28915,N_26806);
nor U33008 (N_33008,N_26238,N_29392);
nand U33009 (N_33009,N_26185,N_27030);
or U33010 (N_33010,N_26211,N_25584);
nor U33011 (N_33011,N_28012,N_26191);
nor U33012 (N_33012,N_26734,N_28277);
and U33013 (N_33013,N_25819,N_26569);
and U33014 (N_33014,N_27613,N_27656);
nand U33015 (N_33015,N_27215,N_26267);
and U33016 (N_33016,N_28034,N_26850);
nor U33017 (N_33017,N_27425,N_29934);
and U33018 (N_33018,N_27147,N_28776);
nand U33019 (N_33019,N_26149,N_25759);
nand U33020 (N_33020,N_29013,N_25239);
nand U33021 (N_33021,N_27256,N_26014);
or U33022 (N_33022,N_25338,N_25723);
or U33023 (N_33023,N_29514,N_26961);
nor U33024 (N_33024,N_28800,N_27553);
xnor U33025 (N_33025,N_29081,N_29594);
and U33026 (N_33026,N_26618,N_29587);
and U33027 (N_33027,N_25882,N_29931);
nand U33028 (N_33028,N_27807,N_26109);
or U33029 (N_33029,N_27937,N_28832);
nand U33030 (N_33030,N_27490,N_28062);
nand U33031 (N_33031,N_28359,N_25025);
nand U33032 (N_33032,N_28406,N_25700);
nand U33033 (N_33033,N_26169,N_29684);
or U33034 (N_33034,N_25660,N_28974);
and U33035 (N_33035,N_28463,N_25255);
and U33036 (N_33036,N_29012,N_29487);
nor U33037 (N_33037,N_27744,N_25939);
nand U33038 (N_33038,N_27949,N_27690);
and U33039 (N_33039,N_29137,N_29876);
or U33040 (N_33040,N_29580,N_29941);
xor U33041 (N_33041,N_28842,N_28814);
and U33042 (N_33042,N_25836,N_27645);
xnor U33043 (N_33043,N_25333,N_26649);
nor U33044 (N_33044,N_25233,N_28970);
or U33045 (N_33045,N_26552,N_29957);
xnor U33046 (N_33046,N_25070,N_29512);
xnor U33047 (N_33047,N_25767,N_26134);
nor U33048 (N_33048,N_28831,N_26395);
nor U33049 (N_33049,N_28151,N_27023);
nand U33050 (N_33050,N_27759,N_26152);
or U33051 (N_33051,N_27786,N_28322);
or U33052 (N_33052,N_29969,N_25222);
xnor U33053 (N_33053,N_29908,N_29686);
xnor U33054 (N_33054,N_29571,N_26391);
nor U33055 (N_33055,N_29767,N_29586);
xnor U33056 (N_33056,N_28575,N_29220);
nand U33057 (N_33057,N_25540,N_29217);
nand U33058 (N_33058,N_26063,N_26136);
xnor U33059 (N_33059,N_28453,N_26699);
nand U33060 (N_33060,N_27860,N_26472);
nor U33061 (N_33061,N_28214,N_25191);
xor U33062 (N_33062,N_29111,N_27076);
nor U33063 (N_33063,N_29961,N_28557);
nor U33064 (N_33064,N_25478,N_27575);
xnor U33065 (N_33065,N_28854,N_27895);
nand U33066 (N_33066,N_25456,N_27657);
nand U33067 (N_33067,N_29208,N_25232);
or U33068 (N_33068,N_26977,N_25030);
nand U33069 (N_33069,N_27952,N_26888);
and U33070 (N_33070,N_26994,N_25075);
nand U33071 (N_33071,N_25696,N_27051);
xnor U33072 (N_33072,N_29967,N_28833);
xor U33073 (N_33073,N_25274,N_25909);
nor U33074 (N_33074,N_25140,N_27336);
nand U33075 (N_33075,N_26285,N_27350);
or U33076 (N_33076,N_29710,N_28967);
or U33077 (N_33077,N_26745,N_26096);
and U33078 (N_33078,N_28909,N_25148);
xor U33079 (N_33079,N_28921,N_28142);
and U33080 (N_33080,N_25692,N_25885);
nand U33081 (N_33081,N_29919,N_26803);
nand U33082 (N_33082,N_27601,N_27667);
or U33083 (N_33083,N_29109,N_27592);
nor U33084 (N_33084,N_28253,N_29855);
or U33085 (N_33085,N_27128,N_29725);
or U33086 (N_33086,N_28499,N_29047);
and U33087 (N_33087,N_28947,N_25807);
nand U33088 (N_33088,N_25287,N_25014);
and U33089 (N_33089,N_26476,N_26303);
or U33090 (N_33090,N_26625,N_26701);
and U33091 (N_33091,N_25654,N_28163);
xor U33092 (N_33092,N_26770,N_25827);
nor U33093 (N_33093,N_25519,N_27681);
or U33094 (N_33094,N_26572,N_26564);
or U33095 (N_33095,N_28676,N_26672);
xor U33096 (N_33096,N_26190,N_25130);
xnor U33097 (N_33097,N_29006,N_28123);
or U33098 (N_33098,N_27046,N_28089);
or U33099 (N_33099,N_26118,N_28096);
xnor U33100 (N_33100,N_28269,N_28492);
or U33101 (N_33101,N_29342,N_27214);
nand U33102 (N_33102,N_28093,N_25734);
nor U33103 (N_33103,N_26239,N_26124);
nor U33104 (N_33104,N_28699,N_25927);
nor U33105 (N_33105,N_29114,N_26955);
xnor U33106 (N_33106,N_26861,N_26343);
nor U33107 (N_33107,N_25989,N_28680);
or U33108 (N_33108,N_25554,N_25095);
or U33109 (N_33109,N_26171,N_26134);
nor U33110 (N_33110,N_26404,N_26618);
and U33111 (N_33111,N_25556,N_29255);
or U33112 (N_33112,N_27402,N_26523);
nand U33113 (N_33113,N_28052,N_28803);
nand U33114 (N_33114,N_26656,N_26605);
or U33115 (N_33115,N_28335,N_27994);
and U33116 (N_33116,N_25603,N_25380);
nor U33117 (N_33117,N_27341,N_26212);
nor U33118 (N_33118,N_27546,N_29689);
and U33119 (N_33119,N_26971,N_29560);
nor U33120 (N_33120,N_27888,N_25339);
or U33121 (N_33121,N_29983,N_26567);
nor U33122 (N_33122,N_25836,N_25592);
nor U33123 (N_33123,N_25796,N_25772);
and U33124 (N_33124,N_26936,N_28478);
nand U33125 (N_33125,N_28691,N_26453);
nand U33126 (N_33126,N_28239,N_25707);
nor U33127 (N_33127,N_25380,N_28737);
or U33128 (N_33128,N_29531,N_26983);
nand U33129 (N_33129,N_26921,N_29322);
nand U33130 (N_33130,N_27768,N_28778);
xnor U33131 (N_33131,N_25879,N_29742);
xnor U33132 (N_33132,N_26414,N_25995);
or U33133 (N_33133,N_25576,N_29478);
nand U33134 (N_33134,N_27589,N_25271);
nand U33135 (N_33135,N_26543,N_28715);
xor U33136 (N_33136,N_28132,N_28375);
and U33137 (N_33137,N_25275,N_28210);
xnor U33138 (N_33138,N_28355,N_29420);
or U33139 (N_33139,N_28035,N_25306);
xnor U33140 (N_33140,N_25266,N_28634);
nor U33141 (N_33141,N_28309,N_25973);
xnor U33142 (N_33142,N_28952,N_28370);
nor U33143 (N_33143,N_25265,N_28892);
nor U33144 (N_33144,N_25390,N_28094);
xnor U33145 (N_33145,N_29728,N_27067);
or U33146 (N_33146,N_26897,N_28435);
and U33147 (N_33147,N_27474,N_27250);
nor U33148 (N_33148,N_25015,N_29572);
and U33149 (N_33149,N_26047,N_28513);
or U33150 (N_33150,N_27049,N_25334);
nand U33151 (N_33151,N_29592,N_25013);
or U33152 (N_33152,N_26497,N_29085);
nand U33153 (N_33153,N_28961,N_29129);
nor U33154 (N_33154,N_28516,N_25391);
nand U33155 (N_33155,N_28811,N_26733);
nand U33156 (N_33156,N_29212,N_29293);
nand U33157 (N_33157,N_29915,N_26535);
nor U33158 (N_33158,N_29171,N_25019);
and U33159 (N_33159,N_28617,N_27412);
nand U33160 (N_33160,N_29275,N_27607);
and U33161 (N_33161,N_25218,N_25878);
xor U33162 (N_33162,N_25855,N_27226);
or U33163 (N_33163,N_27760,N_27319);
xnor U33164 (N_33164,N_27483,N_26347);
xnor U33165 (N_33165,N_26336,N_25956);
xnor U33166 (N_33166,N_29406,N_26655);
and U33167 (N_33167,N_29985,N_29539);
or U33168 (N_33168,N_25914,N_27985);
xor U33169 (N_33169,N_25673,N_25768);
xor U33170 (N_33170,N_26316,N_25167);
or U33171 (N_33171,N_29516,N_27046);
nor U33172 (N_33172,N_27420,N_25570);
nand U33173 (N_33173,N_27189,N_29549);
nor U33174 (N_33174,N_26795,N_28428);
nor U33175 (N_33175,N_26111,N_28296);
nand U33176 (N_33176,N_29920,N_28844);
and U33177 (N_33177,N_25282,N_25171);
xnor U33178 (N_33178,N_29492,N_25142);
or U33179 (N_33179,N_27664,N_29328);
or U33180 (N_33180,N_29730,N_28588);
nor U33181 (N_33181,N_25115,N_25124);
nand U33182 (N_33182,N_28106,N_27627);
nor U33183 (N_33183,N_26619,N_25879);
nand U33184 (N_33184,N_27386,N_25086);
and U33185 (N_33185,N_27412,N_25636);
and U33186 (N_33186,N_29454,N_27119);
or U33187 (N_33187,N_28652,N_25946);
nor U33188 (N_33188,N_26389,N_26267);
or U33189 (N_33189,N_25613,N_25798);
and U33190 (N_33190,N_26133,N_27032);
and U33191 (N_33191,N_29635,N_29305);
and U33192 (N_33192,N_28185,N_28230);
nand U33193 (N_33193,N_27620,N_26067);
and U33194 (N_33194,N_28363,N_27713);
or U33195 (N_33195,N_26029,N_26328);
and U33196 (N_33196,N_27232,N_26227);
nor U33197 (N_33197,N_27639,N_25474);
or U33198 (N_33198,N_26041,N_26998);
nor U33199 (N_33199,N_25061,N_27189);
or U33200 (N_33200,N_27405,N_27677);
nand U33201 (N_33201,N_29643,N_27893);
or U33202 (N_33202,N_26279,N_27765);
and U33203 (N_33203,N_28058,N_25453);
nand U33204 (N_33204,N_26749,N_25458);
xor U33205 (N_33205,N_27547,N_26460);
nor U33206 (N_33206,N_29329,N_25355);
nor U33207 (N_33207,N_27201,N_27848);
xnor U33208 (N_33208,N_25919,N_25774);
and U33209 (N_33209,N_27938,N_26710);
and U33210 (N_33210,N_28702,N_28090);
nand U33211 (N_33211,N_25995,N_27299);
or U33212 (N_33212,N_28634,N_28150);
nor U33213 (N_33213,N_26441,N_26431);
or U33214 (N_33214,N_25863,N_26032);
and U33215 (N_33215,N_26120,N_25201);
nor U33216 (N_33216,N_29379,N_26300);
nand U33217 (N_33217,N_25590,N_28138);
nor U33218 (N_33218,N_26698,N_25577);
nor U33219 (N_33219,N_28686,N_26509);
nand U33220 (N_33220,N_26836,N_25998);
nor U33221 (N_33221,N_28704,N_25376);
nand U33222 (N_33222,N_25721,N_28284);
nand U33223 (N_33223,N_27741,N_26904);
nor U33224 (N_33224,N_29534,N_25074);
or U33225 (N_33225,N_25752,N_25270);
or U33226 (N_33226,N_25253,N_25660);
or U33227 (N_33227,N_28192,N_28738);
xor U33228 (N_33228,N_26393,N_26801);
or U33229 (N_33229,N_29536,N_25584);
xnor U33230 (N_33230,N_25608,N_25778);
nor U33231 (N_33231,N_26349,N_29221);
nor U33232 (N_33232,N_29696,N_27819);
nor U33233 (N_33233,N_25533,N_28464);
nand U33234 (N_33234,N_27186,N_27106);
xnor U33235 (N_33235,N_29963,N_25912);
xor U33236 (N_33236,N_27393,N_27783);
nor U33237 (N_33237,N_29971,N_29892);
or U33238 (N_33238,N_25250,N_26564);
nor U33239 (N_33239,N_29179,N_26863);
nand U33240 (N_33240,N_29904,N_26654);
and U33241 (N_33241,N_25674,N_27288);
nand U33242 (N_33242,N_26562,N_26372);
or U33243 (N_33243,N_27352,N_28377);
xnor U33244 (N_33244,N_29567,N_25383);
xor U33245 (N_33245,N_29930,N_27176);
xor U33246 (N_33246,N_27560,N_28156);
xnor U33247 (N_33247,N_28653,N_28713);
or U33248 (N_33248,N_29046,N_28764);
nor U33249 (N_33249,N_28717,N_27790);
xnor U33250 (N_33250,N_26155,N_26914);
or U33251 (N_33251,N_28863,N_26276);
xnor U33252 (N_33252,N_28214,N_29049);
and U33253 (N_33253,N_29803,N_25649);
or U33254 (N_33254,N_27258,N_27597);
nor U33255 (N_33255,N_26674,N_26915);
nand U33256 (N_33256,N_27521,N_27223);
or U33257 (N_33257,N_28520,N_27480);
nand U33258 (N_33258,N_27088,N_25505);
and U33259 (N_33259,N_29746,N_25437);
nand U33260 (N_33260,N_25045,N_25536);
nor U33261 (N_33261,N_29708,N_26212);
and U33262 (N_33262,N_25917,N_28144);
or U33263 (N_33263,N_28417,N_26357);
or U33264 (N_33264,N_26809,N_25589);
or U33265 (N_33265,N_26089,N_26694);
or U33266 (N_33266,N_25534,N_25540);
xor U33267 (N_33267,N_26722,N_25045);
nor U33268 (N_33268,N_29197,N_29684);
nand U33269 (N_33269,N_25491,N_27557);
or U33270 (N_33270,N_27527,N_27432);
xor U33271 (N_33271,N_25826,N_27139);
and U33272 (N_33272,N_28417,N_25471);
and U33273 (N_33273,N_25808,N_26389);
or U33274 (N_33274,N_28549,N_25531);
or U33275 (N_33275,N_29310,N_29102);
or U33276 (N_33276,N_25537,N_26736);
or U33277 (N_33277,N_29450,N_25694);
nand U33278 (N_33278,N_26942,N_28079);
xnor U33279 (N_33279,N_26252,N_26779);
and U33280 (N_33280,N_28272,N_29974);
nor U33281 (N_33281,N_28928,N_25641);
nor U33282 (N_33282,N_26129,N_27885);
and U33283 (N_33283,N_27304,N_29731);
xnor U33284 (N_33284,N_25916,N_25301);
and U33285 (N_33285,N_27769,N_29493);
nor U33286 (N_33286,N_25462,N_27510);
xnor U33287 (N_33287,N_27559,N_26717);
and U33288 (N_33288,N_25347,N_28149);
or U33289 (N_33289,N_28054,N_25874);
nand U33290 (N_33290,N_26025,N_28202);
nor U33291 (N_33291,N_27935,N_29844);
and U33292 (N_33292,N_25550,N_26203);
or U33293 (N_33293,N_27291,N_25586);
xnor U33294 (N_33294,N_27253,N_28930);
or U33295 (N_33295,N_25155,N_25929);
xnor U33296 (N_33296,N_25903,N_27614);
or U33297 (N_33297,N_26451,N_26984);
nor U33298 (N_33298,N_29651,N_26939);
and U33299 (N_33299,N_27966,N_29096);
or U33300 (N_33300,N_28284,N_28241);
or U33301 (N_33301,N_25326,N_29797);
xor U33302 (N_33302,N_29001,N_26349);
nor U33303 (N_33303,N_28673,N_26949);
and U33304 (N_33304,N_25465,N_25893);
nor U33305 (N_33305,N_27681,N_28201);
xor U33306 (N_33306,N_29371,N_25155);
nand U33307 (N_33307,N_28315,N_25868);
nand U33308 (N_33308,N_25711,N_27281);
xnor U33309 (N_33309,N_29069,N_27031);
and U33310 (N_33310,N_25907,N_29956);
or U33311 (N_33311,N_27897,N_25127);
and U33312 (N_33312,N_27264,N_29880);
nor U33313 (N_33313,N_27809,N_27282);
nor U33314 (N_33314,N_27191,N_29934);
and U33315 (N_33315,N_27529,N_28798);
and U33316 (N_33316,N_29756,N_28987);
xnor U33317 (N_33317,N_25513,N_26058);
and U33318 (N_33318,N_26275,N_29790);
nor U33319 (N_33319,N_25953,N_29421);
and U33320 (N_33320,N_26567,N_28434);
nor U33321 (N_33321,N_28487,N_27005);
and U33322 (N_33322,N_28526,N_28348);
xnor U33323 (N_33323,N_29296,N_28218);
nand U33324 (N_33324,N_27951,N_27027);
or U33325 (N_33325,N_26760,N_26683);
nand U33326 (N_33326,N_29239,N_27606);
nand U33327 (N_33327,N_25555,N_25270);
xnor U33328 (N_33328,N_28684,N_28138);
or U33329 (N_33329,N_29496,N_26331);
nor U33330 (N_33330,N_27599,N_29310);
nor U33331 (N_33331,N_28312,N_25513);
or U33332 (N_33332,N_26388,N_27399);
nand U33333 (N_33333,N_26244,N_26106);
or U33334 (N_33334,N_28430,N_25810);
and U33335 (N_33335,N_25673,N_25345);
nand U33336 (N_33336,N_28650,N_29906);
nand U33337 (N_33337,N_27387,N_27733);
nand U33338 (N_33338,N_28453,N_25240);
and U33339 (N_33339,N_29007,N_25003);
nor U33340 (N_33340,N_27451,N_29205);
and U33341 (N_33341,N_26345,N_27799);
nor U33342 (N_33342,N_25152,N_25359);
and U33343 (N_33343,N_27151,N_29242);
or U33344 (N_33344,N_26878,N_25070);
nand U33345 (N_33345,N_26500,N_29494);
xor U33346 (N_33346,N_26090,N_26440);
nor U33347 (N_33347,N_29743,N_29512);
and U33348 (N_33348,N_29567,N_25804);
xnor U33349 (N_33349,N_25508,N_25718);
and U33350 (N_33350,N_29689,N_28251);
xor U33351 (N_33351,N_27952,N_26306);
nor U33352 (N_33352,N_28254,N_28096);
nor U33353 (N_33353,N_25082,N_28091);
nand U33354 (N_33354,N_27075,N_29217);
and U33355 (N_33355,N_28521,N_25430);
nor U33356 (N_33356,N_27966,N_25971);
and U33357 (N_33357,N_25339,N_28338);
or U33358 (N_33358,N_27146,N_26233);
and U33359 (N_33359,N_28879,N_28604);
nor U33360 (N_33360,N_25129,N_29203);
or U33361 (N_33361,N_26180,N_27680);
and U33362 (N_33362,N_29181,N_28976);
and U33363 (N_33363,N_29836,N_25545);
nand U33364 (N_33364,N_26800,N_27518);
nand U33365 (N_33365,N_29146,N_25817);
xor U33366 (N_33366,N_27898,N_27291);
nor U33367 (N_33367,N_27273,N_27260);
xor U33368 (N_33368,N_29447,N_27008);
or U33369 (N_33369,N_25107,N_25378);
nand U33370 (N_33370,N_26038,N_25446);
or U33371 (N_33371,N_29634,N_28795);
nand U33372 (N_33372,N_26265,N_27492);
and U33373 (N_33373,N_25660,N_29326);
nor U33374 (N_33374,N_25021,N_28469);
and U33375 (N_33375,N_26025,N_27635);
xor U33376 (N_33376,N_25586,N_27172);
and U33377 (N_33377,N_25402,N_25111);
xor U33378 (N_33378,N_29442,N_27243);
nor U33379 (N_33379,N_29596,N_29100);
nor U33380 (N_33380,N_29105,N_26965);
nor U33381 (N_33381,N_26705,N_26177);
or U33382 (N_33382,N_28204,N_28597);
or U33383 (N_33383,N_26796,N_27058);
and U33384 (N_33384,N_28868,N_28790);
nand U33385 (N_33385,N_28762,N_27394);
nor U33386 (N_33386,N_28856,N_29270);
nor U33387 (N_33387,N_28204,N_29783);
nor U33388 (N_33388,N_25425,N_26387);
nor U33389 (N_33389,N_29337,N_26620);
and U33390 (N_33390,N_25395,N_26018);
xor U33391 (N_33391,N_27757,N_28770);
xnor U33392 (N_33392,N_28396,N_29300);
nand U33393 (N_33393,N_28566,N_28363);
xnor U33394 (N_33394,N_29235,N_27576);
nor U33395 (N_33395,N_26337,N_28251);
or U33396 (N_33396,N_28709,N_28369);
nand U33397 (N_33397,N_29375,N_29283);
xnor U33398 (N_33398,N_25753,N_26237);
nor U33399 (N_33399,N_27749,N_26066);
xnor U33400 (N_33400,N_26224,N_25752);
nand U33401 (N_33401,N_25324,N_28114);
and U33402 (N_33402,N_28305,N_29131);
and U33403 (N_33403,N_28872,N_29233);
and U33404 (N_33404,N_26299,N_25081);
or U33405 (N_33405,N_25274,N_27334);
nor U33406 (N_33406,N_28704,N_26209);
and U33407 (N_33407,N_25618,N_26775);
and U33408 (N_33408,N_27161,N_25603);
and U33409 (N_33409,N_26112,N_29880);
nand U33410 (N_33410,N_28122,N_26399);
xor U33411 (N_33411,N_29905,N_29848);
or U33412 (N_33412,N_29730,N_29237);
xnor U33413 (N_33413,N_28483,N_28072);
and U33414 (N_33414,N_28342,N_25507);
or U33415 (N_33415,N_27719,N_29539);
nand U33416 (N_33416,N_28011,N_26636);
and U33417 (N_33417,N_26148,N_28250);
nand U33418 (N_33418,N_25430,N_28254);
xnor U33419 (N_33419,N_28216,N_28957);
nand U33420 (N_33420,N_29224,N_27052);
and U33421 (N_33421,N_25419,N_25980);
nor U33422 (N_33422,N_28581,N_28483);
xnor U33423 (N_33423,N_27840,N_26930);
xor U33424 (N_33424,N_27181,N_25662);
nor U33425 (N_33425,N_29778,N_27470);
or U33426 (N_33426,N_29112,N_28144);
and U33427 (N_33427,N_25567,N_27877);
nand U33428 (N_33428,N_27521,N_27800);
nor U33429 (N_33429,N_26065,N_25943);
nand U33430 (N_33430,N_25492,N_26309);
nand U33431 (N_33431,N_26645,N_29526);
xor U33432 (N_33432,N_29378,N_27716);
xor U33433 (N_33433,N_28734,N_27953);
xnor U33434 (N_33434,N_25627,N_29836);
nor U33435 (N_33435,N_28300,N_27636);
xnor U33436 (N_33436,N_29081,N_25889);
nand U33437 (N_33437,N_28144,N_29012);
nor U33438 (N_33438,N_27170,N_27962);
nand U33439 (N_33439,N_26814,N_29162);
nand U33440 (N_33440,N_28444,N_29722);
xnor U33441 (N_33441,N_27463,N_27974);
and U33442 (N_33442,N_29913,N_26679);
xor U33443 (N_33443,N_28802,N_28011);
or U33444 (N_33444,N_29217,N_28577);
and U33445 (N_33445,N_29535,N_28323);
nor U33446 (N_33446,N_28562,N_27179);
xnor U33447 (N_33447,N_26464,N_28799);
nand U33448 (N_33448,N_28565,N_25404);
or U33449 (N_33449,N_27391,N_25945);
nand U33450 (N_33450,N_27956,N_25486);
and U33451 (N_33451,N_26959,N_27700);
and U33452 (N_33452,N_28188,N_28217);
nand U33453 (N_33453,N_26482,N_27909);
nor U33454 (N_33454,N_25585,N_26342);
xnor U33455 (N_33455,N_29660,N_28630);
or U33456 (N_33456,N_26864,N_26453);
nand U33457 (N_33457,N_26721,N_26804);
and U33458 (N_33458,N_26059,N_29871);
xor U33459 (N_33459,N_26686,N_28743);
nand U33460 (N_33460,N_26987,N_29079);
and U33461 (N_33461,N_26182,N_26951);
and U33462 (N_33462,N_28238,N_25125);
xnor U33463 (N_33463,N_27539,N_25675);
or U33464 (N_33464,N_27884,N_28412);
and U33465 (N_33465,N_26618,N_28494);
xnor U33466 (N_33466,N_29832,N_28338);
nor U33467 (N_33467,N_26443,N_25286);
or U33468 (N_33468,N_26921,N_29668);
xor U33469 (N_33469,N_27494,N_27184);
nand U33470 (N_33470,N_29988,N_29479);
and U33471 (N_33471,N_26525,N_25139);
and U33472 (N_33472,N_27327,N_25414);
nand U33473 (N_33473,N_29857,N_27094);
and U33474 (N_33474,N_29714,N_29534);
and U33475 (N_33475,N_29397,N_28242);
and U33476 (N_33476,N_27716,N_27803);
nand U33477 (N_33477,N_28911,N_26664);
nand U33478 (N_33478,N_25656,N_27302);
xnor U33479 (N_33479,N_28246,N_27051);
and U33480 (N_33480,N_28293,N_28635);
or U33481 (N_33481,N_29252,N_27378);
and U33482 (N_33482,N_29661,N_28770);
or U33483 (N_33483,N_29422,N_26201);
and U33484 (N_33484,N_26647,N_26363);
xnor U33485 (N_33485,N_27977,N_27397);
nor U33486 (N_33486,N_25972,N_27541);
nand U33487 (N_33487,N_29633,N_25007);
nor U33488 (N_33488,N_27050,N_25126);
and U33489 (N_33489,N_29909,N_25122);
and U33490 (N_33490,N_25948,N_28862);
nor U33491 (N_33491,N_27991,N_27387);
and U33492 (N_33492,N_27863,N_26437);
and U33493 (N_33493,N_28507,N_28524);
nor U33494 (N_33494,N_29045,N_25262);
nor U33495 (N_33495,N_27695,N_27936);
nand U33496 (N_33496,N_29163,N_28689);
xor U33497 (N_33497,N_29719,N_25713);
and U33498 (N_33498,N_25582,N_29297);
or U33499 (N_33499,N_25493,N_28467);
nor U33500 (N_33500,N_28086,N_25474);
xnor U33501 (N_33501,N_27611,N_25109);
nor U33502 (N_33502,N_28730,N_27695);
nand U33503 (N_33503,N_27454,N_29138);
and U33504 (N_33504,N_25193,N_28088);
or U33505 (N_33505,N_26686,N_29842);
and U33506 (N_33506,N_29619,N_27954);
nor U33507 (N_33507,N_28285,N_27841);
or U33508 (N_33508,N_28495,N_27432);
and U33509 (N_33509,N_27277,N_25879);
or U33510 (N_33510,N_29279,N_26646);
xnor U33511 (N_33511,N_26873,N_26335);
and U33512 (N_33512,N_28290,N_28887);
nor U33513 (N_33513,N_28753,N_26750);
nor U33514 (N_33514,N_25444,N_26223);
or U33515 (N_33515,N_25263,N_27797);
nand U33516 (N_33516,N_28434,N_26951);
or U33517 (N_33517,N_25527,N_28215);
and U33518 (N_33518,N_25518,N_25206);
and U33519 (N_33519,N_29331,N_27407);
nor U33520 (N_33520,N_29381,N_25171);
nor U33521 (N_33521,N_27376,N_29813);
or U33522 (N_33522,N_27466,N_27671);
and U33523 (N_33523,N_27280,N_28838);
nand U33524 (N_33524,N_25569,N_29140);
or U33525 (N_33525,N_25492,N_27945);
xnor U33526 (N_33526,N_25643,N_26600);
or U33527 (N_33527,N_27766,N_29558);
and U33528 (N_33528,N_25992,N_29379);
and U33529 (N_33529,N_25592,N_28511);
or U33530 (N_33530,N_26738,N_28585);
xor U33531 (N_33531,N_29480,N_25845);
and U33532 (N_33532,N_26328,N_28405);
xor U33533 (N_33533,N_26242,N_29913);
xnor U33534 (N_33534,N_28746,N_28585);
xor U33535 (N_33535,N_26556,N_28981);
xnor U33536 (N_33536,N_29022,N_27935);
nor U33537 (N_33537,N_25331,N_26567);
nor U33538 (N_33538,N_26963,N_27640);
xor U33539 (N_33539,N_25446,N_27056);
and U33540 (N_33540,N_27121,N_26045);
nand U33541 (N_33541,N_27776,N_27191);
nor U33542 (N_33542,N_26399,N_29796);
or U33543 (N_33543,N_28848,N_27784);
nand U33544 (N_33544,N_25282,N_28588);
nor U33545 (N_33545,N_27624,N_28659);
nand U33546 (N_33546,N_25474,N_25327);
nor U33547 (N_33547,N_29845,N_26584);
nor U33548 (N_33548,N_25319,N_26033);
nand U33549 (N_33549,N_25219,N_25707);
and U33550 (N_33550,N_29575,N_26161);
xor U33551 (N_33551,N_27231,N_26432);
and U33552 (N_33552,N_25584,N_29623);
or U33553 (N_33553,N_26754,N_29115);
xnor U33554 (N_33554,N_27674,N_25258);
and U33555 (N_33555,N_29763,N_29950);
nor U33556 (N_33556,N_26021,N_25265);
and U33557 (N_33557,N_27310,N_29490);
nor U33558 (N_33558,N_28396,N_29600);
or U33559 (N_33559,N_27212,N_26208);
nand U33560 (N_33560,N_28518,N_29947);
or U33561 (N_33561,N_25970,N_28150);
nand U33562 (N_33562,N_29879,N_26651);
nor U33563 (N_33563,N_25078,N_29802);
nor U33564 (N_33564,N_25973,N_28023);
xnor U33565 (N_33565,N_25187,N_27120);
xor U33566 (N_33566,N_27907,N_27243);
or U33567 (N_33567,N_25932,N_28017);
nand U33568 (N_33568,N_29788,N_26251);
nand U33569 (N_33569,N_27495,N_27238);
xnor U33570 (N_33570,N_25832,N_25454);
xor U33571 (N_33571,N_25697,N_26642);
and U33572 (N_33572,N_26569,N_29008);
nor U33573 (N_33573,N_28438,N_27318);
or U33574 (N_33574,N_25074,N_25991);
or U33575 (N_33575,N_26690,N_27321);
nand U33576 (N_33576,N_29061,N_25305);
nand U33577 (N_33577,N_27214,N_27919);
nor U33578 (N_33578,N_28100,N_29345);
nor U33579 (N_33579,N_27066,N_26140);
and U33580 (N_33580,N_28523,N_28265);
nand U33581 (N_33581,N_26285,N_27568);
or U33582 (N_33582,N_27738,N_28759);
xor U33583 (N_33583,N_26174,N_27637);
nand U33584 (N_33584,N_29129,N_26652);
xnor U33585 (N_33585,N_26231,N_25526);
and U33586 (N_33586,N_26424,N_26520);
and U33587 (N_33587,N_27869,N_28819);
or U33588 (N_33588,N_26421,N_29004);
nor U33589 (N_33589,N_28006,N_28502);
nand U33590 (N_33590,N_25608,N_27363);
nor U33591 (N_33591,N_28606,N_28567);
and U33592 (N_33592,N_27232,N_29511);
and U33593 (N_33593,N_25619,N_25754);
nand U33594 (N_33594,N_25753,N_25591);
or U33595 (N_33595,N_25144,N_29441);
and U33596 (N_33596,N_25601,N_27335);
or U33597 (N_33597,N_26645,N_26007);
xor U33598 (N_33598,N_27432,N_27276);
nor U33599 (N_33599,N_29764,N_25024);
nand U33600 (N_33600,N_28552,N_28729);
xnor U33601 (N_33601,N_27341,N_26546);
nand U33602 (N_33602,N_26087,N_25766);
xnor U33603 (N_33603,N_25153,N_25347);
nand U33604 (N_33604,N_26020,N_25317);
and U33605 (N_33605,N_25337,N_26689);
or U33606 (N_33606,N_27763,N_26186);
nor U33607 (N_33607,N_28710,N_27514);
xor U33608 (N_33608,N_29647,N_25868);
nand U33609 (N_33609,N_29364,N_27437);
and U33610 (N_33610,N_27091,N_29955);
nor U33611 (N_33611,N_27751,N_29074);
or U33612 (N_33612,N_28309,N_27245);
or U33613 (N_33613,N_25406,N_28730);
or U33614 (N_33614,N_25321,N_25425);
nand U33615 (N_33615,N_27421,N_25888);
nand U33616 (N_33616,N_25313,N_26932);
and U33617 (N_33617,N_28083,N_28454);
nor U33618 (N_33618,N_25638,N_25718);
or U33619 (N_33619,N_25782,N_26781);
and U33620 (N_33620,N_26588,N_28173);
or U33621 (N_33621,N_27399,N_26585);
nor U33622 (N_33622,N_27699,N_27648);
xnor U33623 (N_33623,N_25097,N_29530);
nor U33624 (N_33624,N_28658,N_28635);
nor U33625 (N_33625,N_28444,N_25075);
nand U33626 (N_33626,N_29367,N_28314);
nand U33627 (N_33627,N_29702,N_27127);
nor U33628 (N_33628,N_25967,N_25485);
nand U33629 (N_33629,N_28320,N_25334);
nand U33630 (N_33630,N_25796,N_29052);
nor U33631 (N_33631,N_27606,N_29857);
and U33632 (N_33632,N_28362,N_28178);
nand U33633 (N_33633,N_26032,N_26042);
and U33634 (N_33634,N_25134,N_26613);
nor U33635 (N_33635,N_25758,N_28914);
and U33636 (N_33636,N_28346,N_26463);
nor U33637 (N_33637,N_29279,N_26851);
and U33638 (N_33638,N_28592,N_29131);
nor U33639 (N_33639,N_28617,N_28452);
nor U33640 (N_33640,N_28406,N_25696);
nor U33641 (N_33641,N_29826,N_27243);
nand U33642 (N_33642,N_25230,N_25140);
and U33643 (N_33643,N_28774,N_28213);
nor U33644 (N_33644,N_25921,N_28687);
or U33645 (N_33645,N_29414,N_28064);
and U33646 (N_33646,N_28823,N_26779);
xnor U33647 (N_33647,N_28232,N_26330);
or U33648 (N_33648,N_25821,N_25107);
and U33649 (N_33649,N_27933,N_25767);
xnor U33650 (N_33650,N_28222,N_26848);
nor U33651 (N_33651,N_26154,N_29023);
and U33652 (N_33652,N_29750,N_28300);
xor U33653 (N_33653,N_25321,N_28726);
nor U33654 (N_33654,N_25102,N_29187);
or U33655 (N_33655,N_25904,N_28139);
or U33656 (N_33656,N_25098,N_29652);
nand U33657 (N_33657,N_29679,N_29542);
xor U33658 (N_33658,N_27976,N_26874);
nand U33659 (N_33659,N_26129,N_27818);
nand U33660 (N_33660,N_29277,N_29111);
and U33661 (N_33661,N_26699,N_27739);
xnor U33662 (N_33662,N_25605,N_26331);
or U33663 (N_33663,N_28633,N_26019);
xnor U33664 (N_33664,N_29692,N_27307);
nand U33665 (N_33665,N_26859,N_25080);
nand U33666 (N_33666,N_26740,N_29822);
nor U33667 (N_33667,N_26923,N_25129);
nand U33668 (N_33668,N_25872,N_25614);
xor U33669 (N_33669,N_29348,N_25530);
xor U33670 (N_33670,N_26642,N_25868);
xor U33671 (N_33671,N_26405,N_29713);
or U33672 (N_33672,N_29754,N_26876);
xnor U33673 (N_33673,N_29217,N_29020);
xor U33674 (N_33674,N_29622,N_25820);
or U33675 (N_33675,N_28780,N_28786);
or U33676 (N_33676,N_28071,N_28584);
nand U33677 (N_33677,N_28686,N_25097);
nor U33678 (N_33678,N_28674,N_25345);
xnor U33679 (N_33679,N_29407,N_25343);
nor U33680 (N_33680,N_26464,N_25504);
and U33681 (N_33681,N_28405,N_26068);
or U33682 (N_33682,N_26477,N_25120);
nor U33683 (N_33683,N_26093,N_25473);
and U33684 (N_33684,N_29356,N_26856);
xor U33685 (N_33685,N_26453,N_27659);
and U33686 (N_33686,N_28753,N_27108);
nor U33687 (N_33687,N_27303,N_29372);
and U33688 (N_33688,N_27934,N_27234);
xor U33689 (N_33689,N_28778,N_28214);
xor U33690 (N_33690,N_29697,N_28073);
and U33691 (N_33691,N_26088,N_25592);
nand U33692 (N_33692,N_29604,N_28498);
nor U33693 (N_33693,N_28775,N_28640);
or U33694 (N_33694,N_26510,N_25367);
nor U33695 (N_33695,N_28884,N_29869);
nor U33696 (N_33696,N_26109,N_28585);
xnor U33697 (N_33697,N_27223,N_27353);
and U33698 (N_33698,N_28840,N_25152);
nand U33699 (N_33699,N_26507,N_29966);
and U33700 (N_33700,N_28872,N_26539);
nand U33701 (N_33701,N_25819,N_29694);
or U33702 (N_33702,N_26781,N_26724);
or U33703 (N_33703,N_29742,N_25819);
and U33704 (N_33704,N_27383,N_26495);
or U33705 (N_33705,N_28786,N_26320);
xnor U33706 (N_33706,N_25026,N_26180);
xnor U33707 (N_33707,N_29614,N_27717);
or U33708 (N_33708,N_28996,N_29878);
xnor U33709 (N_33709,N_28043,N_28780);
nor U33710 (N_33710,N_29200,N_25769);
xnor U33711 (N_33711,N_29274,N_25722);
and U33712 (N_33712,N_26096,N_28507);
and U33713 (N_33713,N_29712,N_29593);
and U33714 (N_33714,N_28863,N_25191);
and U33715 (N_33715,N_25853,N_26229);
and U33716 (N_33716,N_27905,N_25039);
xnor U33717 (N_33717,N_28298,N_26283);
nor U33718 (N_33718,N_29830,N_25042);
nor U33719 (N_33719,N_27086,N_27712);
nor U33720 (N_33720,N_29380,N_28177);
nor U33721 (N_33721,N_26337,N_25842);
or U33722 (N_33722,N_27753,N_29980);
or U33723 (N_33723,N_26329,N_26504);
or U33724 (N_33724,N_28031,N_25656);
or U33725 (N_33725,N_28108,N_25326);
or U33726 (N_33726,N_29526,N_27181);
nor U33727 (N_33727,N_26495,N_27392);
nor U33728 (N_33728,N_26992,N_28023);
or U33729 (N_33729,N_28434,N_28010);
or U33730 (N_33730,N_25681,N_27418);
xnor U33731 (N_33731,N_26884,N_29661);
and U33732 (N_33732,N_28926,N_25666);
nand U33733 (N_33733,N_29612,N_29638);
or U33734 (N_33734,N_25465,N_26809);
xor U33735 (N_33735,N_25094,N_26063);
and U33736 (N_33736,N_26840,N_25582);
nand U33737 (N_33737,N_27322,N_25601);
xnor U33738 (N_33738,N_25821,N_28914);
xnor U33739 (N_33739,N_27144,N_27479);
nand U33740 (N_33740,N_26459,N_25123);
nor U33741 (N_33741,N_26338,N_29581);
nand U33742 (N_33742,N_25337,N_25207);
or U33743 (N_33743,N_28938,N_26530);
xnor U33744 (N_33744,N_25660,N_28408);
nand U33745 (N_33745,N_25769,N_25930);
or U33746 (N_33746,N_29820,N_27269);
or U33747 (N_33747,N_25079,N_25132);
nand U33748 (N_33748,N_29529,N_29072);
xnor U33749 (N_33749,N_27715,N_28738);
nand U33750 (N_33750,N_28944,N_29967);
nand U33751 (N_33751,N_26524,N_28653);
xor U33752 (N_33752,N_27897,N_28466);
and U33753 (N_33753,N_29566,N_26397);
nand U33754 (N_33754,N_28806,N_27033);
and U33755 (N_33755,N_27438,N_29558);
and U33756 (N_33756,N_29354,N_25350);
nor U33757 (N_33757,N_26898,N_26887);
and U33758 (N_33758,N_26999,N_27016);
and U33759 (N_33759,N_25140,N_26547);
or U33760 (N_33760,N_28065,N_29978);
and U33761 (N_33761,N_29491,N_28904);
xor U33762 (N_33762,N_27161,N_27863);
xnor U33763 (N_33763,N_29047,N_29525);
and U33764 (N_33764,N_28983,N_29841);
and U33765 (N_33765,N_26732,N_25560);
nor U33766 (N_33766,N_28970,N_25182);
or U33767 (N_33767,N_26247,N_28688);
or U33768 (N_33768,N_28603,N_28499);
nand U33769 (N_33769,N_26020,N_28884);
nand U33770 (N_33770,N_26030,N_29756);
nor U33771 (N_33771,N_27736,N_29571);
and U33772 (N_33772,N_26837,N_25747);
nor U33773 (N_33773,N_25457,N_27061);
xor U33774 (N_33774,N_26463,N_25665);
nor U33775 (N_33775,N_25875,N_25225);
xor U33776 (N_33776,N_29510,N_26490);
nor U33777 (N_33777,N_26660,N_27655);
xor U33778 (N_33778,N_26123,N_26729);
nand U33779 (N_33779,N_29621,N_25591);
or U33780 (N_33780,N_26307,N_26299);
and U33781 (N_33781,N_25308,N_29836);
or U33782 (N_33782,N_27466,N_29603);
xor U33783 (N_33783,N_27538,N_28937);
xor U33784 (N_33784,N_25368,N_27339);
nand U33785 (N_33785,N_25800,N_27849);
xor U33786 (N_33786,N_25809,N_28733);
nor U33787 (N_33787,N_28050,N_28594);
nand U33788 (N_33788,N_28430,N_29465);
and U33789 (N_33789,N_29941,N_25165);
and U33790 (N_33790,N_29122,N_25844);
and U33791 (N_33791,N_29581,N_29169);
nand U33792 (N_33792,N_28363,N_27414);
or U33793 (N_33793,N_29284,N_26684);
or U33794 (N_33794,N_29368,N_25267);
xor U33795 (N_33795,N_25287,N_26719);
and U33796 (N_33796,N_27243,N_26974);
nand U33797 (N_33797,N_27215,N_26028);
xnor U33798 (N_33798,N_29333,N_29187);
or U33799 (N_33799,N_27308,N_28222);
or U33800 (N_33800,N_29260,N_25837);
nor U33801 (N_33801,N_26874,N_25890);
xnor U33802 (N_33802,N_29135,N_28243);
nor U33803 (N_33803,N_29567,N_26702);
xor U33804 (N_33804,N_26861,N_27702);
or U33805 (N_33805,N_26275,N_29192);
nand U33806 (N_33806,N_28355,N_25374);
and U33807 (N_33807,N_29798,N_27888);
or U33808 (N_33808,N_29921,N_27649);
nor U33809 (N_33809,N_25556,N_26667);
or U33810 (N_33810,N_25402,N_28364);
nand U33811 (N_33811,N_27040,N_29082);
xor U33812 (N_33812,N_29195,N_25942);
and U33813 (N_33813,N_26984,N_25323);
or U33814 (N_33814,N_28586,N_25121);
nor U33815 (N_33815,N_29420,N_25182);
xor U33816 (N_33816,N_27614,N_29096);
or U33817 (N_33817,N_29840,N_28932);
nor U33818 (N_33818,N_26454,N_29997);
or U33819 (N_33819,N_28235,N_27918);
nand U33820 (N_33820,N_28798,N_26905);
xor U33821 (N_33821,N_27909,N_26539);
xor U33822 (N_33822,N_26458,N_29586);
or U33823 (N_33823,N_27070,N_25409);
nand U33824 (N_33824,N_29671,N_26089);
nand U33825 (N_33825,N_25104,N_27529);
xnor U33826 (N_33826,N_28804,N_25807);
xnor U33827 (N_33827,N_27087,N_25500);
or U33828 (N_33828,N_29996,N_27149);
xnor U33829 (N_33829,N_29706,N_28703);
nand U33830 (N_33830,N_29365,N_28141);
nor U33831 (N_33831,N_26466,N_26791);
or U33832 (N_33832,N_26030,N_26477);
and U33833 (N_33833,N_27172,N_26339);
nand U33834 (N_33834,N_29656,N_29052);
and U33835 (N_33835,N_29249,N_29256);
xor U33836 (N_33836,N_26938,N_28232);
or U33837 (N_33837,N_28911,N_25606);
nand U33838 (N_33838,N_29659,N_26371);
and U33839 (N_33839,N_27504,N_26002);
or U33840 (N_33840,N_29839,N_25403);
and U33841 (N_33841,N_28029,N_27983);
or U33842 (N_33842,N_29308,N_29218);
nand U33843 (N_33843,N_29533,N_29949);
xnor U33844 (N_33844,N_25146,N_29091);
xor U33845 (N_33845,N_27588,N_26296);
or U33846 (N_33846,N_26941,N_25161);
or U33847 (N_33847,N_25080,N_29454);
and U33848 (N_33848,N_26471,N_28436);
nor U33849 (N_33849,N_27767,N_27139);
nand U33850 (N_33850,N_29008,N_27896);
and U33851 (N_33851,N_26294,N_27766);
nand U33852 (N_33852,N_25179,N_28038);
nand U33853 (N_33853,N_29697,N_25364);
xnor U33854 (N_33854,N_28006,N_27074);
nor U33855 (N_33855,N_26237,N_25177);
and U33856 (N_33856,N_27234,N_25596);
or U33857 (N_33857,N_27618,N_27693);
and U33858 (N_33858,N_28018,N_27574);
nand U33859 (N_33859,N_27012,N_27441);
xor U33860 (N_33860,N_27163,N_29249);
or U33861 (N_33861,N_25772,N_25450);
nor U33862 (N_33862,N_26044,N_29765);
xor U33863 (N_33863,N_29258,N_25763);
nor U33864 (N_33864,N_25823,N_26356);
xor U33865 (N_33865,N_27812,N_27022);
nand U33866 (N_33866,N_27473,N_26758);
xnor U33867 (N_33867,N_28679,N_29088);
and U33868 (N_33868,N_29158,N_29516);
nand U33869 (N_33869,N_28447,N_26923);
and U33870 (N_33870,N_29894,N_27043);
nand U33871 (N_33871,N_25763,N_26086);
xor U33872 (N_33872,N_29701,N_29908);
nand U33873 (N_33873,N_25900,N_26917);
nor U33874 (N_33874,N_29328,N_27595);
and U33875 (N_33875,N_26469,N_26256);
nor U33876 (N_33876,N_25205,N_25947);
nor U33877 (N_33877,N_27169,N_25957);
nor U33878 (N_33878,N_26334,N_27642);
nor U33879 (N_33879,N_29297,N_27665);
nor U33880 (N_33880,N_25322,N_29924);
and U33881 (N_33881,N_27870,N_25528);
and U33882 (N_33882,N_29771,N_29487);
or U33883 (N_33883,N_27043,N_29477);
or U33884 (N_33884,N_27866,N_26310);
and U33885 (N_33885,N_26702,N_29758);
nor U33886 (N_33886,N_28506,N_26523);
or U33887 (N_33887,N_27293,N_27827);
nor U33888 (N_33888,N_26588,N_27457);
or U33889 (N_33889,N_27602,N_25998);
or U33890 (N_33890,N_26409,N_27967);
nor U33891 (N_33891,N_26776,N_26023);
xor U33892 (N_33892,N_26487,N_29347);
and U33893 (N_33893,N_25319,N_27105);
nor U33894 (N_33894,N_25199,N_29012);
nand U33895 (N_33895,N_25629,N_28677);
and U33896 (N_33896,N_25363,N_28703);
nor U33897 (N_33897,N_28824,N_25005);
nor U33898 (N_33898,N_25386,N_26062);
xnor U33899 (N_33899,N_26428,N_29441);
nor U33900 (N_33900,N_27676,N_29403);
xor U33901 (N_33901,N_28607,N_25474);
xor U33902 (N_33902,N_27705,N_26002);
xor U33903 (N_33903,N_29518,N_29943);
or U33904 (N_33904,N_25396,N_27052);
nand U33905 (N_33905,N_28247,N_27006);
and U33906 (N_33906,N_29000,N_28850);
or U33907 (N_33907,N_28385,N_27467);
nor U33908 (N_33908,N_26232,N_28235);
and U33909 (N_33909,N_25890,N_27828);
nor U33910 (N_33910,N_26570,N_25812);
or U33911 (N_33911,N_28112,N_26263);
nand U33912 (N_33912,N_28609,N_27785);
nor U33913 (N_33913,N_28007,N_28125);
or U33914 (N_33914,N_25610,N_26117);
xor U33915 (N_33915,N_25843,N_26315);
nand U33916 (N_33916,N_25849,N_26270);
or U33917 (N_33917,N_27411,N_26282);
xnor U33918 (N_33918,N_25191,N_25640);
xnor U33919 (N_33919,N_26355,N_28770);
nand U33920 (N_33920,N_26014,N_26078);
xnor U33921 (N_33921,N_25293,N_27008);
and U33922 (N_33922,N_26605,N_27821);
xnor U33923 (N_33923,N_25391,N_28276);
or U33924 (N_33924,N_26577,N_25252);
and U33925 (N_33925,N_28481,N_27014);
and U33926 (N_33926,N_28768,N_29991);
and U33927 (N_33927,N_25035,N_25604);
xnor U33928 (N_33928,N_29335,N_27277);
xor U33929 (N_33929,N_25411,N_25231);
and U33930 (N_33930,N_27745,N_25053);
nand U33931 (N_33931,N_28339,N_29378);
or U33932 (N_33932,N_28825,N_28994);
and U33933 (N_33933,N_28497,N_25796);
and U33934 (N_33934,N_25312,N_25825);
xor U33935 (N_33935,N_29963,N_27200);
xor U33936 (N_33936,N_27747,N_29630);
and U33937 (N_33937,N_26285,N_29434);
nand U33938 (N_33938,N_28972,N_25484);
xnor U33939 (N_33939,N_26737,N_25176);
nor U33940 (N_33940,N_25873,N_25560);
and U33941 (N_33941,N_26268,N_29716);
nand U33942 (N_33942,N_29653,N_27551);
nand U33943 (N_33943,N_25939,N_28676);
and U33944 (N_33944,N_28881,N_27906);
nand U33945 (N_33945,N_29433,N_28080);
or U33946 (N_33946,N_25767,N_26388);
nand U33947 (N_33947,N_27927,N_29228);
nand U33948 (N_33948,N_28104,N_25972);
nor U33949 (N_33949,N_25447,N_28366);
or U33950 (N_33950,N_27032,N_25051);
xor U33951 (N_33951,N_26129,N_25829);
and U33952 (N_33952,N_27135,N_26681);
xnor U33953 (N_33953,N_25263,N_27739);
nand U33954 (N_33954,N_26352,N_29845);
and U33955 (N_33955,N_28677,N_28928);
xor U33956 (N_33956,N_25592,N_28059);
nand U33957 (N_33957,N_27972,N_28379);
and U33958 (N_33958,N_28961,N_25111);
and U33959 (N_33959,N_27169,N_26101);
nor U33960 (N_33960,N_26396,N_28942);
or U33961 (N_33961,N_28077,N_26357);
xnor U33962 (N_33962,N_25018,N_28910);
nand U33963 (N_33963,N_29798,N_27609);
nor U33964 (N_33964,N_26090,N_29024);
xnor U33965 (N_33965,N_25652,N_28887);
or U33966 (N_33966,N_29435,N_25808);
and U33967 (N_33967,N_29646,N_29953);
or U33968 (N_33968,N_27010,N_29619);
nand U33969 (N_33969,N_29006,N_29739);
nor U33970 (N_33970,N_26322,N_28398);
and U33971 (N_33971,N_29506,N_26306);
or U33972 (N_33972,N_28148,N_25296);
nand U33973 (N_33973,N_25337,N_28638);
and U33974 (N_33974,N_29807,N_26667);
nand U33975 (N_33975,N_28806,N_29359);
nand U33976 (N_33976,N_29208,N_28210);
or U33977 (N_33977,N_29716,N_26911);
or U33978 (N_33978,N_25630,N_27323);
xnor U33979 (N_33979,N_28098,N_25105);
xnor U33980 (N_33980,N_25409,N_28193);
or U33981 (N_33981,N_26957,N_25106);
xor U33982 (N_33982,N_27191,N_27506);
xor U33983 (N_33983,N_28535,N_27348);
xnor U33984 (N_33984,N_27960,N_25271);
nor U33985 (N_33985,N_29917,N_27209);
or U33986 (N_33986,N_25825,N_28161);
or U33987 (N_33987,N_28384,N_29571);
nand U33988 (N_33988,N_27219,N_26742);
nor U33989 (N_33989,N_29791,N_25704);
nor U33990 (N_33990,N_28233,N_28166);
and U33991 (N_33991,N_26966,N_25075);
or U33992 (N_33992,N_27300,N_25876);
and U33993 (N_33993,N_29518,N_27743);
and U33994 (N_33994,N_29895,N_26008);
xor U33995 (N_33995,N_27671,N_28492);
or U33996 (N_33996,N_27150,N_26273);
xnor U33997 (N_33997,N_26826,N_28914);
xor U33998 (N_33998,N_29349,N_28671);
xnor U33999 (N_33999,N_28855,N_29185);
nand U34000 (N_34000,N_25969,N_29322);
and U34001 (N_34001,N_29423,N_28720);
xor U34002 (N_34002,N_27243,N_27055);
and U34003 (N_34003,N_26615,N_28715);
and U34004 (N_34004,N_25660,N_27782);
nor U34005 (N_34005,N_29353,N_28583);
and U34006 (N_34006,N_25022,N_27761);
and U34007 (N_34007,N_26813,N_29786);
nand U34008 (N_34008,N_29418,N_28885);
or U34009 (N_34009,N_27901,N_26236);
and U34010 (N_34010,N_25912,N_27558);
and U34011 (N_34011,N_28045,N_29574);
or U34012 (N_34012,N_25984,N_28096);
or U34013 (N_34013,N_28531,N_26826);
and U34014 (N_34014,N_28071,N_29753);
and U34015 (N_34015,N_28101,N_26815);
or U34016 (N_34016,N_26381,N_28059);
nor U34017 (N_34017,N_26065,N_28793);
or U34018 (N_34018,N_26892,N_26204);
nor U34019 (N_34019,N_29164,N_26217);
nand U34020 (N_34020,N_28492,N_28043);
and U34021 (N_34021,N_25049,N_25147);
and U34022 (N_34022,N_29998,N_29102);
and U34023 (N_34023,N_27174,N_27412);
or U34024 (N_34024,N_25615,N_25552);
xor U34025 (N_34025,N_25959,N_26273);
and U34026 (N_34026,N_28143,N_25303);
and U34027 (N_34027,N_29816,N_28308);
xor U34028 (N_34028,N_29827,N_27121);
nand U34029 (N_34029,N_27691,N_28429);
nand U34030 (N_34030,N_27334,N_25252);
xor U34031 (N_34031,N_29664,N_29820);
xor U34032 (N_34032,N_29980,N_25233);
and U34033 (N_34033,N_26957,N_29949);
xnor U34034 (N_34034,N_28937,N_27043);
and U34035 (N_34035,N_26098,N_29100);
nor U34036 (N_34036,N_28475,N_27395);
or U34037 (N_34037,N_25408,N_26551);
xor U34038 (N_34038,N_28609,N_26413);
or U34039 (N_34039,N_26647,N_26936);
or U34040 (N_34040,N_26227,N_29546);
and U34041 (N_34041,N_28167,N_28885);
and U34042 (N_34042,N_26558,N_27096);
xnor U34043 (N_34043,N_25591,N_27409);
xnor U34044 (N_34044,N_27476,N_27536);
nor U34045 (N_34045,N_27635,N_27528);
nand U34046 (N_34046,N_27071,N_27108);
nand U34047 (N_34047,N_27634,N_27291);
xnor U34048 (N_34048,N_28553,N_29908);
nand U34049 (N_34049,N_28884,N_25602);
nand U34050 (N_34050,N_28381,N_26644);
and U34051 (N_34051,N_26027,N_26733);
nor U34052 (N_34052,N_28736,N_25454);
xnor U34053 (N_34053,N_27162,N_27719);
nand U34054 (N_34054,N_25647,N_27289);
or U34055 (N_34055,N_25402,N_26631);
xor U34056 (N_34056,N_27947,N_26449);
xnor U34057 (N_34057,N_27429,N_27466);
or U34058 (N_34058,N_27663,N_27126);
nand U34059 (N_34059,N_28310,N_29926);
xnor U34060 (N_34060,N_27259,N_26743);
nor U34061 (N_34061,N_25109,N_25645);
or U34062 (N_34062,N_25186,N_25056);
and U34063 (N_34063,N_25075,N_26420);
xor U34064 (N_34064,N_27633,N_26504);
nand U34065 (N_34065,N_25063,N_25277);
nor U34066 (N_34066,N_26309,N_26567);
or U34067 (N_34067,N_29769,N_29441);
and U34068 (N_34068,N_29910,N_26960);
nand U34069 (N_34069,N_27096,N_29735);
nand U34070 (N_34070,N_29589,N_27070);
nor U34071 (N_34071,N_27458,N_25851);
xor U34072 (N_34072,N_27629,N_26763);
xnor U34073 (N_34073,N_28735,N_26840);
and U34074 (N_34074,N_28751,N_25470);
nor U34075 (N_34075,N_26154,N_26187);
and U34076 (N_34076,N_27163,N_25845);
nor U34077 (N_34077,N_29326,N_26409);
and U34078 (N_34078,N_28933,N_28401);
nand U34079 (N_34079,N_28935,N_29332);
and U34080 (N_34080,N_29906,N_25122);
nor U34081 (N_34081,N_27052,N_25696);
and U34082 (N_34082,N_25243,N_25050);
and U34083 (N_34083,N_25835,N_29932);
nand U34084 (N_34084,N_25501,N_28163);
and U34085 (N_34085,N_27526,N_26435);
and U34086 (N_34086,N_26138,N_25043);
xor U34087 (N_34087,N_28521,N_28025);
and U34088 (N_34088,N_26988,N_29535);
or U34089 (N_34089,N_29332,N_25577);
nor U34090 (N_34090,N_29958,N_29972);
nor U34091 (N_34091,N_26908,N_25234);
nor U34092 (N_34092,N_29983,N_25866);
and U34093 (N_34093,N_26615,N_28445);
or U34094 (N_34094,N_28046,N_27700);
xnor U34095 (N_34095,N_26550,N_26568);
nor U34096 (N_34096,N_26124,N_29959);
or U34097 (N_34097,N_27034,N_28128);
nor U34098 (N_34098,N_29567,N_25820);
nand U34099 (N_34099,N_27911,N_27939);
or U34100 (N_34100,N_25007,N_25710);
or U34101 (N_34101,N_25922,N_26224);
xor U34102 (N_34102,N_28100,N_29611);
and U34103 (N_34103,N_26796,N_25036);
or U34104 (N_34104,N_28026,N_26350);
and U34105 (N_34105,N_25967,N_27811);
and U34106 (N_34106,N_26432,N_25906);
xor U34107 (N_34107,N_25634,N_26018);
nor U34108 (N_34108,N_28786,N_28639);
xnor U34109 (N_34109,N_28383,N_27583);
xnor U34110 (N_34110,N_27562,N_27244);
nand U34111 (N_34111,N_28123,N_28150);
and U34112 (N_34112,N_29786,N_28041);
nand U34113 (N_34113,N_27483,N_26446);
and U34114 (N_34114,N_25483,N_25805);
or U34115 (N_34115,N_29784,N_26902);
or U34116 (N_34116,N_26954,N_25921);
nor U34117 (N_34117,N_25483,N_28907);
and U34118 (N_34118,N_25149,N_25054);
nor U34119 (N_34119,N_25913,N_29838);
and U34120 (N_34120,N_29784,N_27159);
xnor U34121 (N_34121,N_26256,N_28807);
xnor U34122 (N_34122,N_27737,N_25217);
or U34123 (N_34123,N_25458,N_28336);
nor U34124 (N_34124,N_26158,N_25519);
nor U34125 (N_34125,N_29955,N_29154);
xnor U34126 (N_34126,N_25341,N_26120);
and U34127 (N_34127,N_28117,N_27562);
nand U34128 (N_34128,N_26819,N_27819);
nand U34129 (N_34129,N_28947,N_29132);
nor U34130 (N_34130,N_29579,N_27470);
and U34131 (N_34131,N_27868,N_27451);
xnor U34132 (N_34132,N_25656,N_26703);
or U34133 (N_34133,N_28683,N_26285);
xor U34134 (N_34134,N_28887,N_25072);
nand U34135 (N_34135,N_27106,N_29151);
or U34136 (N_34136,N_25666,N_28785);
and U34137 (N_34137,N_26383,N_28662);
or U34138 (N_34138,N_26985,N_25087);
nor U34139 (N_34139,N_29958,N_26341);
nor U34140 (N_34140,N_26668,N_28554);
nor U34141 (N_34141,N_25974,N_27819);
xor U34142 (N_34142,N_27937,N_25326);
or U34143 (N_34143,N_27772,N_28583);
nand U34144 (N_34144,N_25225,N_26812);
xor U34145 (N_34145,N_28981,N_25189);
or U34146 (N_34146,N_26534,N_27092);
or U34147 (N_34147,N_29624,N_28439);
and U34148 (N_34148,N_27600,N_29522);
nor U34149 (N_34149,N_28637,N_27061);
and U34150 (N_34150,N_29135,N_26854);
or U34151 (N_34151,N_27593,N_28305);
xor U34152 (N_34152,N_25551,N_27354);
or U34153 (N_34153,N_27448,N_27249);
or U34154 (N_34154,N_27432,N_29336);
xor U34155 (N_34155,N_29857,N_27980);
and U34156 (N_34156,N_29972,N_27083);
or U34157 (N_34157,N_28609,N_26229);
xor U34158 (N_34158,N_25302,N_28215);
or U34159 (N_34159,N_29015,N_25964);
nand U34160 (N_34160,N_25266,N_26242);
or U34161 (N_34161,N_26236,N_27582);
xor U34162 (N_34162,N_29269,N_28442);
and U34163 (N_34163,N_29862,N_29259);
or U34164 (N_34164,N_25814,N_28750);
xnor U34165 (N_34165,N_28537,N_29736);
nor U34166 (N_34166,N_26686,N_28788);
nor U34167 (N_34167,N_26554,N_28797);
nand U34168 (N_34168,N_26390,N_28306);
nor U34169 (N_34169,N_27322,N_28000);
or U34170 (N_34170,N_29445,N_29832);
nand U34171 (N_34171,N_26864,N_29115);
nand U34172 (N_34172,N_29786,N_28923);
xor U34173 (N_34173,N_27910,N_26917);
nand U34174 (N_34174,N_25967,N_29685);
or U34175 (N_34175,N_27310,N_29458);
nor U34176 (N_34176,N_25701,N_26964);
xnor U34177 (N_34177,N_26104,N_26857);
and U34178 (N_34178,N_25030,N_25133);
or U34179 (N_34179,N_29283,N_26517);
or U34180 (N_34180,N_28624,N_27489);
or U34181 (N_34181,N_25328,N_27960);
and U34182 (N_34182,N_29031,N_28093);
nor U34183 (N_34183,N_29773,N_29120);
nor U34184 (N_34184,N_25474,N_28309);
nor U34185 (N_34185,N_29890,N_28265);
or U34186 (N_34186,N_27376,N_26433);
and U34187 (N_34187,N_27434,N_26907);
nand U34188 (N_34188,N_28202,N_28534);
xnor U34189 (N_34189,N_28622,N_29176);
nand U34190 (N_34190,N_27313,N_25401);
or U34191 (N_34191,N_28487,N_28514);
and U34192 (N_34192,N_26303,N_28057);
and U34193 (N_34193,N_26146,N_27720);
nor U34194 (N_34194,N_25864,N_28520);
and U34195 (N_34195,N_27075,N_27880);
xor U34196 (N_34196,N_28984,N_28892);
nor U34197 (N_34197,N_25374,N_29572);
nand U34198 (N_34198,N_26104,N_27603);
xor U34199 (N_34199,N_25838,N_25329);
or U34200 (N_34200,N_28366,N_27746);
or U34201 (N_34201,N_28688,N_25114);
nor U34202 (N_34202,N_29313,N_29829);
or U34203 (N_34203,N_29585,N_29430);
and U34204 (N_34204,N_25047,N_25924);
and U34205 (N_34205,N_27383,N_25135);
nand U34206 (N_34206,N_29004,N_28210);
xnor U34207 (N_34207,N_26283,N_26864);
nand U34208 (N_34208,N_29097,N_28408);
and U34209 (N_34209,N_28991,N_29501);
nand U34210 (N_34210,N_26348,N_28163);
nand U34211 (N_34211,N_28753,N_25809);
and U34212 (N_34212,N_28626,N_29306);
nor U34213 (N_34213,N_28964,N_26055);
nor U34214 (N_34214,N_27235,N_25062);
nor U34215 (N_34215,N_29488,N_27933);
xor U34216 (N_34216,N_25903,N_26555);
xnor U34217 (N_34217,N_25032,N_27399);
or U34218 (N_34218,N_28863,N_25542);
and U34219 (N_34219,N_29744,N_25729);
and U34220 (N_34220,N_28872,N_25200);
nand U34221 (N_34221,N_28344,N_26598);
or U34222 (N_34222,N_29875,N_28489);
nor U34223 (N_34223,N_27087,N_27800);
and U34224 (N_34224,N_25279,N_29968);
or U34225 (N_34225,N_29578,N_27466);
or U34226 (N_34226,N_26647,N_27172);
xnor U34227 (N_34227,N_26246,N_25170);
and U34228 (N_34228,N_29223,N_29106);
nand U34229 (N_34229,N_27508,N_28777);
nor U34230 (N_34230,N_29514,N_29214);
nand U34231 (N_34231,N_28503,N_29305);
xor U34232 (N_34232,N_27870,N_27097);
nor U34233 (N_34233,N_28562,N_28478);
or U34234 (N_34234,N_26899,N_29100);
or U34235 (N_34235,N_28167,N_26068);
and U34236 (N_34236,N_26378,N_27008);
or U34237 (N_34237,N_27529,N_28618);
xnor U34238 (N_34238,N_27253,N_27227);
nand U34239 (N_34239,N_25921,N_26201);
or U34240 (N_34240,N_26101,N_27628);
and U34241 (N_34241,N_29270,N_25626);
xnor U34242 (N_34242,N_27786,N_25593);
xnor U34243 (N_34243,N_25740,N_26451);
nand U34244 (N_34244,N_27353,N_28005);
or U34245 (N_34245,N_25929,N_25740);
xor U34246 (N_34246,N_28470,N_29311);
or U34247 (N_34247,N_28150,N_27166);
nand U34248 (N_34248,N_27844,N_26552);
xor U34249 (N_34249,N_29718,N_28575);
and U34250 (N_34250,N_27923,N_26598);
nand U34251 (N_34251,N_28969,N_25246);
nand U34252 (N_34252,N_28803,N_29222);
or U34253 (N_34253,N_27457,N_27470);
and U34254 (N_34254,N_25450,N_26439);
nor U34255 (N_34255,N_27914,N_28320);
and U34256 (N_34256,N_26821,N_27415);
and U34257 (N_34257,N_25724,N_27692);
xor U34258 (N_34258,N_29849,N_28812);
nand U34259 (N_34259,N_26774,N_25445);
nand U34260 (N_34260,N_28102,N_26123);
and U34261 (N_34261,N_27805,N_26170);
and U34262 (N_34262,N_29974,N_26142);
nor U34263 (N_34263,N_29817,N_26498);
nand U34264 (N_34264,N_26782,N_25221);
nand U34265 (N_34265,N_26253,N_26049);
xnor U34266 (N_34266,N_29119,N_26247);
xor U34267 (N_34267,N_29030,N_26736);
and U34268 (N_34268,N_29619,N_26065);
and U34269 (N_34269,N_29033,N_26776);
xnor U34270 (N_34270,N_29216,N_28731);
and U34271 (N_34271,N_26756,N_29283);
xor U34272 (N_34272,N_29908,N_26013);
and U34273 (N_34273,N_25099,N_29389);
xnor U34274 (N_34274,N_29992,N_29433);
nor U34275 (N_34275,N_29363,N_25798);
nor U34276 (N_34276,N_26086,N_26625);
xnor U34277 (N_34277,N_29742,N_26986);
nor U34278 (N_34278,N_29430,N_29148);
xor U34279 (N_34279,N_29636,N_27435);
or U34280 (N_34280,N_29734,N_28437);
xnor U34281 (N_34281,N_27264,N_26591);
nor U34282 (N_34282,N_27920,N_26893);
nand U34283 (N_34283,N_27624,N_29973);
or U34284 (N_34284,N_27024,N_29943);
nand U34285 (N_34285,N_26532,N_26821);
xor U34286 (N_34286,N_27107,N_27150);
xnor U34287 (N_34287,N_25661,N_25679);
or U34288 (N_34288,N_28622,N_25364);
and U34289 (N_34289,N_29846,N_27525);
xnor U34290 (N_34290,N_27774,N_27841);
nor U34291 (N_34291,N_28934,N_26955);
nor U34292 (N_34292,N_29286,N_29328);
nor U34293 (N_34293,N_28137,N_25755);
nor U34294 (N_34294,N_29886,N_26699);
nor U34295 (N_34295,N_29018,N_26059);
xnor U34296 (N_34296,N_29041,N_25773);
nor U34297 (N_34297,N_25905,N_27974);
and U34298 (N_34298,N_25148,N_28157);
or U34299 (N_34299,N_26651,N_27886);
nor U34300 (N_34300,N_29176,N_29757);
or U34301 (N_34301,N_27650,N_26547);
or U34302 (N_34302,N_26444,N_29547);
nand U34303 (N_34303,N_25995,N_28779);
nor U34304 (N_34304,N_27336,N_28252);
nand U34305 (N_34305,N_26709,N_29516);
nand U34306 (N_34306,N_25360,N_27566);
and U34307 (N_34307,N_25597,N_26159);
xnor U34308 (N_34308,N_25183,N_28297);
and U34309 (N_34309,N_26842,N_28887);
xnor U34310 (N_34310,N_29148,N_29974);
xor U34311 (N_34311,N_27532,N_27459);
or U34312 (N_34312,N_25317,N_28663);
and U34313 (N_34313,N_27557,N_27713);
xnor U34314 (N_34314,N_28673,N_25585);
nand U34315 (N_34315,N_25356,N_29718);
nand U34316 (N_34316,N_26375,N_27235);
or U34317 (N_34317,N_28166,N_25834);
and U34318 (N_34318,N_27245,N_27759);
and U34319 (N_34319,N_25062,N_26026);
nand U34320 (N_34320,N_28119,N_27333);
nor U34321 (N_34321,N_28713,N_26411);
and U34322 (N_34322,N_26327,N_26573);
nand U34323 (N_34323,N_28038,N_26135);
and U34324 (N_34324,N_27935,N_28372);
nor U34325 (N_34325,N_25170,N_26674);
and U34326 (N_34326,N_25532,N_25364);
or U34327 (N_34327,N_28167,N_29319);
or U34328 (N_34328,N_29359,N_29688);
or U34329 (N_34329,N_29903,N_29621);
or U34330 (N_34330,N_25445,N_25091);
xnor U34331 (N_34331,N_27031,N_29885);
nor U34332 (N_34332,N_26955,N_29887);
xor U34333 (N_34333,N_27995,N_28615);
and U34334 (N_34334,N_27768,N_28701);
or U34335 (N_34335,N_29131,N_26226);
or U34336 (N_34336,N_27672,N_25542);
xor U34337 (N_34337,N_26835,N_25136);
xnor U34338 (N_34338,N_28263,N_27612);
and U34339 (N_34339,N_27751,N_26883);
nor U34340 (N_34340,N_29179,N_29594);
xnor U34341 (N_34341,N_26529,N_26839);
and U34342 (N_34342,N_25970,N_26138);
nand U34343 (N_34343,N_29835,N_25736);
and U34344 (N_34344,N_26391,N_28900);
and U34345 (N_34345,N_27487,N_25773);
nor U34346 (N_34346,N_26176,N_27189);
nor U34347 (N_34347,N_29488,N_27936);
xor U34348 (N_34348,N_25435,N_27460);
nand U34349 (N_34349,N_25125,N_28496);
nor U34350 (N_34350,N_27630,N_28992);
nand U34351 (N_34351,N_25389,N_27059);
xnor U34352 (N_34352,N_25379,N_28124);
and U34353 (N_34353,N_26042,N_27402);
nand U34354 (N_34354,N_27578,N_25743);
nor U34355 (N_34355,N_26849,N_26683);
nor U34356 (N_34356,N_26436,N_27450);
nand U34357 (N_34357,N_26331,N_29010);
nor U34358 (N_34358,N_29403,N_25240);
nand U34359 (N_34359,N_27688,N_28180);
and U34360 (N_34360,N_29254,N_27713);
or U34361 (N_34361,N_26766,N_27114);
and U34362 (N_34362,N_27977,N_28928);
and U34363 (N_34363,N_27452,N_29367);
and U34364 (N_34364,N_27142,N_27135);
or U34365 (N_34365,N_25490,N_27857);
nand U34366 (N_34366,N_26060,N_25941);
nor U34367 (N_34367,N_27838,N_29202);
and U34368 (N_34368,N_27565,N_29483);
and U34369 (N_34369,N_27060,N_27807);
or U34370 (N_34370,N_26857,N_29732);
nor U34371 (N_34371,N_27909,N_28934);
or U34372 (N_34372,N_26720,N_29677);
nor U34373 (N_34373,N_28300,N_25196);
xor U34374 (N_34374,N_25687,N_25926);
nand U34375 (N_34375,N_29883,N_27511);
xnor U34376 (N_34376,N_25105,N_25209);
nand U34377 (N_34377,N_29461,N_29271);
or U34378 (N_34378,N_25091,N_27734);
nor U34379 (N_34379,N_28673,N_28091);
nor U34380 (N_34380,N_29245,N_27478);
and U34381 (N_34381,N_26053,N_29220);
nand U34382 (N_34382,N_28573,N_27547);
and U34383 (N_34383,N_28441,N_25065);
nor U34384 (N_34384,N_28805,N_25394);
nor U34385 (N_34385,N_25388,N_25663);
or U34386 (N_34386,N_28422,N_27667);
or U34387 (N_34387,N_27397,N_25818);
nand U34388 (N_34388,N_27696,N_26213);
or U34389 (N_34389,N_26494,N_28560);
nand U34390 (N_34390,N_28191,N_29059);
xor U34391 (N_34391,N_26128,N_29552);
xor U34392 (N_34392,N_25851,N_26358);
nand U34393 (N_34393,N_26489,N_26575);
and U34394 (N_34394,N_29967,N_28084);
and U34395 (N_34395,N_26358,N_28125);
and U34396 (N_34396,N_28737,N_28841);
nor U34397 (N_34397,N_28263,N_28898);
nand U34398 (N_34398,N_29638,N_27112);
xnor U34399 (N_34399,N_28591,N_25445);
or U34400 (N_34400,N_25394,N_26911);
nand U34401 (N_34401,N_25160,N_26366);
nor U34402 (N_34402,N_27095,N_28780);
and U34403 (N_34403,N_27063,N_27648);
or U34404 (N_34404,N_28855,N_29628);
or U34405 (N_34405,N_29502,N_28632);
xor U34406 (N_34406,N_27574,N_28799);
and U34407 (N_34407,N_28427,N_26586);
xor U34408 (N_34408,N_28478,N_29548);
and U34409 (N_34409,N_25317,N_29839);
xor U34410 (N_34410,N_29839,N_25418);
xnor U34411 (N_34411,N_25475,N_26331);
nand U34412 (N_34412,N_29053,N_25703);
nor U34413 (N_34413,N_29438,N_28103);
or U34414 (N_34414,N_28023,N_26635);
nor U34415 (N_34415,N_28072,N_25003);
nand U34416 (N_34416,N_28815,N_25790);
and U34417 (N_34417,N_26423,N_26277);
and U34418 (N_34418,N_25416,N_25688);
or U34419 (N_34419,N_26382,N_25294);
and U34420 (N_34420,N_29159,N_26961);
xor U34421 (N_34421,N_29091,N_27061);
nor U34422 (N_34422,N_27452,N_26860);
or U34423 (N_34423,N_27982,N_26831);
nor U34424 (N_34424,N_27549,N_28663);
and U34425 (N_34425,N_25676,N_27735);
nand U34426 (N_34426,N_26698,N_28221);
nor U34427 (N_34427,N_28850,N_29341);
and U34428 (N_34428,N_29454,N_27390);
and U34429 (N_34429,N_29801,N_26052);
or U34430 (N_34430,N_28601,N_29206);
or U34431 (N_34431,N_27555,N_27406);
and U34432 (N_34432,N_28438,N_27300);
xnor U34433 (N_34433,N_27854,N_28678);
nand U34434 (N_34434,N_29518,N_29094);
or U34435 (N_34435,N_26764,N_25485);
xor U34436 (N_34436,N_26803,N_28568);
or U34437 (N_34437,N_28338,N_28475);
or U34438 (N_34438,N_25380,N_28934);
nor U34439 (N_34439,N_28186,N_25546);
and U34440 (N_34440,N_27341,N_27319);
nand U34441 (N_34441,N_28326,N_26331);
nor U34442 (N_34442,N_27188,N_25460);
and U34443 (N_34443,N_25844,N_29956);
nor U34444 (N_34444,N_29308,N_25125);
nor U34445 (N_34445,N_25218,N_26346);
or U34446 (N_34446,N_27806,N_27491);
and U34447 (N_34447,N_26521,N_27307);
xor U34448 (N_34448,N_28192,N_28024);
nand U34449 (N_34449,N_25068,N_26361);
and U34450 (N_34450,N_26518,N_29101);
or U34451 (N_34451,N_26504,N_29401);
and U34452 (N_34452,N_29553,N_25915);
xor U34453 (N_34453,N_28974,N_28103);
xor U34454 (N_34454,N_25854,N_27543);
nor U34455 (N_34455,N_27144,N_27256);
nand U34456 (N_34456,N_26679,N_25939);
and U34457 (N_34457,N_29461,N_26542);
or U34458 (N_34458,N_26407,N_29682);
xnor U34459 (N_34459,N_25917,N_28302);
nand U34460 (N_34460,N_29906,N_26816);
xnor U34461 (N_34461,N_26229,N_28004);
or U34462 (N_34462,N_29754,N_25345);
xor U34463 (N_34463,N_25651,N_27842);
xor U34464 (N_34464,N_28469,N_29799);
and U34465 (N_34465,N_28671,N_28732);
or U34466 (N_34466,N_25132,N_25957);
and U34467 (N_34467,N_25787,N_26465);
nor U34468 (N_34468,N_29013,N_27247);
or U34469 (N_34469,N_29081,N_29266);
xor U34470 (N_34470,N_27158,N_26975);
or U34471 (N_34471,N_28596,N_27010);
or U34472 (N_34472,N_29121,N_26902);
nor U34473 (N_34473,N_28840,N_26820);
xnor U34474 (N_34474,N_25646,N_27442);
or U34475 (N_34475,N_28743,N_28670);
xnor U34476 (N_34476,N_25667,N_28892);
xor U34477 (N_34477,N_25965,N_25715);
nand U34478 (N_34478,N_29325,N_27575);
and U34479 (N_34479,N_28595,N_26989);
xor U34480 (N_34480,N_28275,N_26412);
nand U34481 (N_34481,N_28230,N_29821);
nand U34482 (N_34482,N_27458,N_28745);
nand U34483 (N_34483,N_28774,N_29764);
or U34484 (N_34484,N_26769,N_25603);
nand U34485 (N_34485,N_26546,N_29737);
nand U34486 (N_34486,N_28792,N_27854);
or U34487 (N_34487,N_26135,N_26825);
or U34488 (N_34488,N_28446,N_27317);
or U34489 (N_34489,N_29881,N_27193);
or U34490 (N_34490,N_26257,N_28899);
nor U34491 (N_34491,N_29271,N_28190);
nor U34492 (N_34492,N_28032,N_27492);
nand U34493 (N_34493,N_25013,N_28201);
xor U34494 (N_34494,N_29905,N_29408);
or U34495 (N_34495,N_26946,N_25839);
nand U34496 (N_34496,N_27550,N_29409);
or U34497 (N_34497,N_28195,N_27940);
or U34498 (N_34498,N_25406,N_28663);
nand U34499 (N_34499,N_29780,N_25016);
or U34500 (N_34500,N_25596,N_27986);
xor U34501 (N_34501,N_28384,N_29507);
or U34502 (N_34502,N_29435,N_27738);
nand U34503 (N_34503,N_29878,N_25662);
nand U34504 (N_34504,N_25071,N_26225);
nor U34505 (N_34505,N_28265,N_29282);
nand U34506 (N_34506,N_26611,N_25543);
xnor U34507 (N_34507,N_29196,N_27787);
xnor U34508 (N_34508,N_29135,N_29681);
or U34509 (N_34509,N_26138,N_26346);
xnor U34510 (N_34510,N_25439,N_27394);
xnor U34511 (N_34511,N_25908,N_26967);
or U34512 (N_34512,N_25942,N_27479);
and U34513 (N_34513,N_28821,N_27095);
and U34514 (N_34514,N_25598,N_29789);
or U34515 (N_34515,N_29032,N_26341);
nor U34516 (N_34516,N_27257,N_25947);
or U34517 (N_34517,N_27262,N_29732);
nand U34518 (N_34518,N_27058,N_25410);
nand U34519 (N_34519,N_27825,N_28564);
nand U34520 (N_34520,N_25758,N_27689);
nor U34521 (N_34521,N_26985,N_27166);
xor U34522 (N_34522,N_26302,N_25883);
nor U34523 (N_34523,N_29633,N_26228);
and U34524 (N_34524,N_27062,N_28133);
xor U34525 (N_34525,N_29655,N_27992);
xor U34526 (N_34526,N_28550,N_26281);
or U34527 (N_34527,N_29218,N_28912);
nand U34528 (N_34528,N_25857,N_29134);
nor U34529 (N_34529,N_29890,N_27031);
nor U34530 (N_34530,N_29729,N_29456);
nand U34531 (N_34531,N_29593,N_26055);
xor U34532 (N_34532,N_28150,N_27141);
xnor U34533 (N_34533,N_28961,N_26989);
nor U34534 (N_34534,N_27503,N_27106);
and U34535 (N_34535,N_25853,N_25725);
xnor U34536 (N_34536,N_29290,N_27922);
and U34537 (N_34537,N_28648,N_25875);
and U34538 (N_34538,N_29121,N_26175);
and U34539 (N_34539,N_27195,N_28057);
or U34540 (N_34540,N_29801,N_29710);
and U34541 (N_34541,N_25041,N_25287);
and U34542 (N_34542,N_26906,N_26272);
nand U34543 (N_34543,N_27751,N_27051);
and U34544 (N_34544,N_25023,N_25589);
or U34545 (N_34545,N_26976,N_28028);
nor U34546 (N_34546,N_25932,N_26035);
nor U34547 (N_34547,N_25911,N_28731);
nand U34548 (N_34548,N_29143,N_26269);
nor U34549 (N_34549,N_27439,N_29617);
and U34550 (N_34550,N_25424,N_25929);
nand U34551 (N_34551,N_28816,N_25954);
or U34552 (N_34552,N_28159,N_25915);
nor U34553 (N_34553,N_28836,N_29252);
nand U34554 (N_34554,N_27881,N_29608);
nor U34555 (N_34555,N_25513,N_26733);
or U34556 (N_34556,N_29547,N_25401);
nor U34557 (N_34557,N_28277,N_27343);
and U34558 (N_34558,N_26009,N_25423);
xnor U34559 (N_34559,N_25462,N_28588);
or U34560 (N_34560,N_28905,N_26569);
nor U34561 (N_34561,N_25019,N_28820);
or U34562 (N_34562,N_26469,N_27207);
or U34563 (N_34563,N_25460,N_25644);
or U34564 (N_34564,N_26731,N_25759);
nor U34565 (N_34565,N_29157,N_27653);
nand U34566 (N_34566,N_27818,N_28891);
and U34567 (N_34567,N_27999,N_29395);
or U34568 (N_34568,N_27782,N_25687);
or U34569 (N_34569,N_25334,N_28178);
or U34570 (N_34570,N_27288,N_29218);
and U34571 (N_34571,N_29047,N_25214);
or U34572 (N_34572,N_25246,N_25250);
or U34573 (N_34573,N_28679,N_25018);
nand U34574 (N_34574,N_29406,N_28967);
nor U34575 (N_34575,N_25712,N_29409);
or U34576 (N_34576,N_25983,N_25540);
xnor U34577 (N_34577,N_25401,N_26931);
nand U34578 (N_34578,N_28279,N_26093);
or U34579 (N_34579,N_25723,N_27083);
and U34580 (N_34580,N_27875,N_29069);
and U34581 (N_34581,N_27299,N_29262);
nor U34582 (N_34582,N_27298,N_25318);
and U34583 (N_34583,N_25697,N_25756);
nor U34584 (N_34584,N_25604,N_28989);
nand U34585 (N_34585,N_27186,N_28910);
and U34586 (N_34586,N_29703,N_26802);
xor U34587 (N_34587,N_27422,N_29834);
nor U34588 (N_34588,N_26314,N_29254);
nor U34589 (N_34589,N_27837,N_26650);
nand U34590 (N_34590,N_26914,N_25163);
or U34591 (N_34591,N_28575,N_26691);
or U34592 (N_34592,N_25477,N_28902);
or U34593 (N_34593,N_27082,N_26555);
or U34594 (N_34594,N_28674,N_27450);
xor U34595 (N_34595,N_29161,N_29999);
and U34596 (N_34596,N_29175,N_29849);
nand U34597 (N_34597,N_26836,N_28790);
nor U34598 (N_34598,N_27985,N_28811);
nor U34599 (N_34599,N_29315,N_25344);
nand U34600 (N_34600,N_26105,N_26493);
xnor U34601 (N_34601,N_25381,N_25939);
xor U34602 (N_34602,N_25145,N_28069);
xor U34603 (N_34603,N_29083,N_28110);
nand U34604 (N_34604,N_27162,N_27231);
nor U34605 (N_34605,N_25743,N_28308);
nor U34606 (N_34606,N_25223,N_25222);
or U34607 (N_34607,N_28219,N_29957);
xnor U34608 (N_34608,N_25100,N_26303);
or U34609 (N_34609,N_25537,N_28444);
and U34610 (N_34610,N_26119,N_25010);
or U34611 (N_34611,N_28349,N_29921);
nand U34612 (N_34612,N_26613,N_25720);
nor U34613 (N_34613,N_25350,N_28384);
nor U34614 (N_34614,N_27111,N_27091);
or U34615 (N_34615,N_29106,N_28634);
nor U34616 (N_34616,N_29045,N_27793);
nand U34617 (N_34617,N_29978,N_28816);
nor U34618 (N_34618,N_26621,N_28816);
nor U34619 (N_34619,N_25059,N_25778);
nand U34620 (N_34620,N_28827,N_29876);
and U34621 (N_34621,N_27258,N_25131);
or U34622 (N_34622,N_25690,N_27008);
nand U34623 (N_34623,N_25735,N_27190);
nand U34624 (N_34624,N_28214,N_27371);
and U34625 (N_34625,N_25190,N_29112);
or U34626 (N_34626,N_29111,N_28162);
nor U34627 (N_34627,N_28617,N_27611);
nand U34628 (N_34628,N_25666,N_27543);
and U34629 (N_34629,N_25201,N_26338);
nand U34630 (N_34630,N_28774,N_26678);
and U34631 (N_34631,N_25039,N_25687);
xor U34632 (N_34632,N_28129,N_25102);
and U34633 (N_34633,N_27674,N_27991);
or U34634 (N_34634,N_25516,N_28502);
nor U34635 (N_34635,N_29971,N_25049);
nand U34636 (N_34636,N_25171,N_27238);
nand U34637 (N_34637,N_29551,N_28963);
nor U34638 (N_34638,N_25856,N_29988);
nor U34639 (N_34639,N_27457,N_29238);
and U34640 (N_34640,N_28958,N_29987);
nor U34641 (N_34641,N_26541,N_28035);
xor U34642 (N_34642,N_25811,N_29191);
or U34643 (N_34643,N_27556,N_27476);
or U34644 (N_34644,N_25647,N_28989);
nand U34645 (N_34645,N_25590,N_29863);
nor U34646 (N_34646,N_25229,N_29027);
and U34647 (N_34647,N_25310,N_29497);
xor U34648 (N_34648,N_25143,N_29398);
or U34649 (N_34649,N_26612,N_25265);
nor U34650 (N_34650,N_29868,N_28581);
nor U34651 (N_34651,N_27426,N_29904);
or U34652 (N_34652,N_26810,N_29040);
xnor U34653 (N_34653,N_28519,N_28806);
xor U34654 (N_34654,N_29278,N_27534);
nand U34655 (N_34655,N_28987,N_27690);
or U34656 (N_34656,N_25942,N_28704);
nor U34657 (N_34657,N_26040,N_27621);
nor U34658 (N_34658,N_28805,N_26146);
xnor U34659 (N_34659,N_28651,N_25937);
nand U34660 (N_34660,N_28908,N_25244);
xnor U34661 (N_34661,N_27842,N_26795);
and U34662 (N_34662,N_27980,N_29053);
nand U34663 (N_34663,N_27300,N_28497);
xnor U34664 (N_34664,N_28947,N_29861);
nand U34665 (N_34665,N_25268,N_27833);
or U34666 (N_34666,N_26518,N_27435);
nor U34667 (N_34667,N_28360,N_27635);
xnor U34668 (N_34668,N_29859,N_25668);
and U34669 (N_34669,N_29598,N_26226);
xor U34670 (N_34670,N_28147,N_26295);
xor U34671 (N_34671,N_26672,N_28683);
nand U34672 (N_34672,N_27677,N_29643);
nor U34673 (N_34673,N_29985,N_28159);
xnor U34674 (N_34674,N_29282,N_27369);
xnor U34675 (N_34675,N_28689,N_27311);
and U34676 (N_34676,N_28266,N_26593);
and U34677 (N_34677,N_28936,N_26144);
nand U34678 (N_34678,N_25198,N_26720);
nand U34679 (N_34679,N_26491,N_26826);
xnor U34680 (N_34680,N_26962,N_25704);
nor U34681 (N_34681,N_27729,N_29987);
nand U34682 (N_34682,N_26035,N_26021);
nand U34683 (N_34683,N_28843,N_26155);
nor U34684 (N_34684,N_29390,N_25745);
xor U34685 (N_34685,N_26618,N_27841);
and U34686 (N_34686,N_26468,N_27224);
and U34687 (N_34687,N_29478,N_26719);
nor U34688 (N_34688,N_26322,N_26462);
or U34689 (N_34689,N_25915,N_27790);
or U34690 (N_34690,N_25116,N_28310);
nand U34691 (N_34691,N_27030,N_27386);
or U34692 (N_34692,N_28228,N_25592);
and U34693 (N_34693,N_25353,N_25735);
or U34694 (N_34694,N_28034,N_29709);
nor U34695 (N_34695,N_27983,N_27029);
xnor U34696 (N_34696,N_27092,N_28172);
or U34697 (N_34697,N_27919,N_28213);
nand U34698 (N_34698,N_25155,N_25077);
and U34699 (N_34699,N_25363,N_27506);
xnor U34700 (N_34700,N_28270,N_29885);
or U34701 (N_34701,N_29942,N_25077);
nand U34702 (N_34702,N_25194,N_27068);
nor U34703 (N_34703,N_26875,N_29801);
nor U34704 (N_34704,N_27994,N_29562);
or U34705 (N_34705,N_27626,N_29105);
and U34706 (N_34706,N_26603,N_29460);
nor U34707 (N_34707,N_28386,N_29874);
nor U34708 (N_34708,N_29056,N_29017);
and U34709 (N_34709,N_27670,N_26819);
xor U34710 (N_34710,N_27274,N_27740);
and U34711 (N_34711,N_27112,N_29867);
xnor U34712 (N_34712,N_27129,N_28501);
nand U34713 (N_34713,N_26483,N_29588);
and U34714 (N_34714,N_27944,N_26564);
nand U34715 (N_34715,N_27478,N_26684);
or U34716 (N_34716,N_29342,N_25507);
or U34717 (N_34717,N_28558,N_27532);
nand U34718 (N_34718,N_26839,N_28419);
xor U34719 (N_34719,N_28451,N_29517);
nor U34720 (N_34720,N_25652,N_26571);
nand U34721 (N_34721,N_28121,N_28454);
or U34722 (N_34722,N_29447,N_29718);
nand U34723 (N_34723,N_27931,N_26947);
nor U34724 (N_34724,N_28347,N_28425);
and U34725 (N_34725,N_26830,N_27793);
nor U34726 (N_34726,N_25548,N_29996);
or U34727 (N_34727,N_25291,N_27350);
xor U34728 (N_34728,N_27648,N_29680);
or U34729 (N_34729,N_28635,N_28374);
nor U34730 (N_34730,N_26639,N_29971);
nor U34731 (N_34731,N_28290,N_27369);
xnor U34732 (N_34732,N_25557,N_28907);
xnor U34733 (N_34733,N_28191,N_28222);
nand U34734 (N_34734,N_29773,N_25005);
nand U34735 (N_34735,N_27301,N_26414);
nor U34736 (N_34736,N_25158,N_26223);
nand U34737 (N_34737,N_28145,N_29267);
nor U34738 (N_34738,N_29885,N_26715);
nor U34739 (N_34739,N_29681,N_28848);
or U34740 (N_34740,N_28791,N_27082);
or U34741 (N_34741,N_25425,N_26805);
or U34742 (N_34742,N_26138,N_28068);
xnor U34743 (N_34743,N_25810,N_26044);
nand U34744 (N_34744,N_29362,N_27161);
nor U34745 (N_34745,N_26522,N_25030);
and U34746 (N_34746,N_25641,N_26090);
or U34747 (N_34747,N_28642,N_29822);
and U34748 (N_34748,N_25358,N_25421);
or U34749 (N_34749,N_26088,N_26601);
nor U34750 (N_34750,N_25305,N_28455);
nor U34751 (N_34751,N_28503,N_29659);
or U34752 (N_34752,N_28373,N_26807);
and U34753 (N_34753,N_29604,N_26679);
and U34754 (N_34754,N_25204,N_26650);
nor U34755 (N_34755,N_27128,N_25304);
nor U34756 (N_34756,N_26697,N_25584);
and U34757 (N_34757,N_27194,N_25129);
nand U34758 (N_34758,N_29519,N_25895);
xnor U34759 (N_34759,N_26043,N_27514);
and U34760 (N_34760,N_27866,N_28359);
xor U34761 (N_34761,N_25728,N_27814);
nor U34762 (N_34762,N_29034,N_27045);
or U34763 (N_34763,N_28783,N_29397);
xor U34764 (N_34764,N_28524,N_29589);
xnor U34765 (N_34765,N_29168,N_25336);
xor U34766 (N_34766,N_26335,N_26912);
or U34767 (N_34767,N_26807,N_27235);
xnor U34768 (N_34768,N_25579,N_27336);
or U34769 (N_34769,N_27223,N_28204);
and U34770 (N_34770,N_28867,N_29166);
nor U34771 (N_34771,N_25701,N_29189);
nor U34772 (N_34772,N_25627,N_26260);
nor U34773 (N_34773,N_25787,N_28982);
and U34774 (N_34774,N_29883,N_26160);
nor U34775 (N_34775,N_25765,N_28551);
nor U34776 (N_34776,N_25252,N_27282);
nor U34777 (N_34777,N_29798,N_29441);
or U34778 (N_34778,N_29981,N_25128);
nand U34779 (N_34779,N_26680,N_25365);
xnor U34780 (N_34780,N_28631,N_27922);
or U34781 (N_34781,N_27205,N_26670);
or U34782 (N_34782,N_28414,N_29893);
nand U34783 (N_34783,N_29892,N_29564);
and U34784 (N_34784,N_28100,N_29802);
and U34785 (N_34785,N_27847,N_26943);
or U34786 (N_34786,N_28720,N_29053);
xnor U34787 (N_34787,N_25477,N_28330);
nor U34788 (N_34788,N_29229,N_25950);
nand U34789 (N_34789,N_27748,N_28178);
xor U34790 (N_34790,N_25961,N_25519);
and U34791 (N_34791,N_28315,N_28956);
or U34792 (N_34792,N_29694,N_28770);
and U34793 (N_34793,N_27573,N_26774);
nor U34794 (N_34794,N_28282,N_28419);
and U34795 (N_34795,N_27373,N_28466);
or U34796 (N_34796,N_28358,N_27544);
nor U34797 (N_34797,N_25991,N_25289);
nor U34798 (N_34798,N_29203,N_25501);
nand U34799 (N_34799,N_25835,N_25907);
nand U34800 (N_34800,N_29674,N_28230);
nor U34801 (N_34801,N_26024,N_27279);
xor U34802 (N_34802,N_28436,N_26522);
or U34803 (N_34803,N_25936,N_28151);
or U34804 (N_34804,N_26398,N_25550);
or U34805 (N_34805,N_29287,N_26586);
nor U34806 (N_34806,N_27165,N_26161);
xnor U34807 (N_34807,N_25195,N_26426);
nand U34808 (N_34808,N_25767,N_29169);
xnor U34809 (N_34809,N_29310,N_29952);
nand U34810 (N_34810,N_25191,N_26900);
xnor U34811 (N_34811,N_26308,N_27178);
or U34812 (N_34812,N_28356,N_29221);
or U34813 (N_34813,N_29251,N_26013);
xor U34814 (N_34814,N_29981,N_29967);
and U34815 (N_34815,N_28877,N_26490);
xor U34816 (N_34816,N_25511,N_26300);
nand U34817 (N_34817,N_28084,N_29005);
or U34818 (N_34818,N_25107,N_28657);
nand U34819 (N_34819,N_25763,N_26940);
nor U34820 (N_34820,N_29329,N_26061);
nor U34821 (N_34821,N_27040,N_27933);
nor U34822 (N_34822,N_28578,N_29985);
xnor U34823 (N_34823,N_29702,N_28393);
or U34824 (N_34824,N_29256,N_26036);
or U34825 (N_34825,N_28946,N_25571);
and U34826 (N_34826,N_28967,N_27675);
and U34827 (N_34827,N_27513,N_25746);
or U34828 (N_34828,N_29792,N_27547);
nand U34829 (N_34829,N_27016,N_27680);
and U34830 (N_34830,N_29761,N_27025);
and U34831 (N_34831,N_29418,N_26889);
and U34832 (N_34832,N_27936,N_28322);
nor U34833 (N_34833,N_27846,N_29626);
and U34834 (N_34834,N_25447,N_28609);
nor U34835 (N_34835,N_29955,N_27682);
xnor U34836 (N_34836,N_25832,N_29248);
nand U34837 (N_34837,N_28470,N_29987);
nor U34838 (N_34838,N_25471,N_27113);
or U34839 (N_34839,N_28519,N_27020);
nor U34840 (N_34840,N_27845,N_25014);
nand U34841 (N_34841,N_26681,N_27010);
and U34842 (N_34842,N_25601,N_28578);
nand U34843 (N_34843,N_28482,N_28066);
nand U34844 (N_34844,N_29018,N_27038);
or U34845 (N_34845,N_25973,N_26490);
xor U34846 (N_34846,N_29835,N_27415);
and U34847 (N_34847,N_27374,N_28143);
and U34848 (N_34848,N_29158,N_27477);
xor U34849 (N_34849,N_26299,N_27424);
nor U34850 (N_34850,N_26365,N_27183);
xor U34851 (N_34851,N_29302,N_25554);
nor U34852 (N_34852,N_25681,N_28526);
and U34853 (N_34853,N_28501,N_25290);
and U34854 (N_34854,N_25928,N_28137);
or U34855 (N_34855,N_28659,N_25503);
nand U34856 (N_34856,N_26372,N_27163);
and U34857 (N_34857,N_29390,N_26991);
or U34858 (N_34858,N_25320,N_26053);
or U34859 (N_34859,N_25543,N_28189);
xnor U34860 (N_34860,N_25084,N_29286);
nor U34861 (N_34861,N_25111,N_27168);
xnor U34862 (N_34862,N_26269,N_26400);
nand U34863 (N_34863,N_26691,N_26643);
xor U34864 (N_34864,N_28515,N_28847);
xor U34865 (N_34865,N_25683,N_29310);
and U34866 (N_34866,N_26777,N_27474);
nor U34867 (N_34867,N_29140,N_27192);
nand U34868 (N_34868,N_25090,N_27196);
nor U34869 (N_34869,N_25741,N_26017);
and U34870 (N_34870,N_27636,N_26155);
xor U34871 (N_34871,N_29548,N_26810);
xor U34872 (N_34872,N_27114,N_27807);
nand U34873 (N_34873,N_25611,N_26510);
and U34874 (N_34874,N_28260,N_29207);
or U34875 (N_34875,N_28595,N_25552);
nand U34876 (N_34876,N_28267,N_28942);
and U34877 (N_34877,N_29635,N_28149);
nand U34878 (N_34878,N_29798,N_27317);
or U34879 (N_34879,N_26253,N_25839);
xor U34880 (N_34880,N_28216,N_25845);
nor U34881 (N_34881,N_26655,N_26047);
xnor U34882 (N_34882,N_25427,N_29646);
xor U34883 (N_34883,N_26636,N_27602);
or U34884 (N_34884,N_26362,N_28137);
xor U34885 (N_34885,N_26799,N_25753);
nand U34886 (N_34886,N_25829,N_26695);
nor U34887 (N_34887,N_26370,N_28993);
nand U34888 (N_34888,N_28943,N_26316);
xnor U34889 (N_34889,N_27310,N_28804);
nor U34890 (N_34890,N_26747,N_29441);
and U34891 (N_34891,N_26817,N_26234);
nand U34892 (N_34892,N_25206,N_25063);
nor U34893 (N_34893,N_26195,N_29524);
nor U34894 (N_34894,N_26722,N_26129);
nor U34895 (N_34895,N_25589,N_26872);
nand U34896 (N_34896,N_28561,N_29945);
nor U34897 (N_34897,N_26589,N_29404);
xor U34898 (N_34898,N_26904,N_25411);
nand U34899 (N_34899,N_25346,N_27011);
and U34900 (N_34900,N_29491,N_28888);
nand U34901 (N_34901,N_27754,N_25109);
xnor U34902 (N_34902,N_25747,N_29854);
and U34903 (N_34903,N_26421,N_28679);
nand U34904 (N_34904,N_26939,N_25716);
nor U34905 (N_34905,N_29716,N_29031);
and U34906 (N_34906,N_26848,N_29822);
xnor U34907 (N_34907,N_27020,N_26171);
xnor U34908 (N_34908,N_27550,N_29774);
or U34909 (N_34909,N_27955,N_28111);
xor U34910 (N_34910,N_28102,N_27074);
and U34911 (N_34911,N_25624,N_26264);
xnor U34912 (N_34912,N_27422,N_29873);
xor U34913 (N_34913,N_29589,N_28957);
nand U34914 (N_34914,N_25368,N_29589);
or U34915 (N_34915,N_25002,N_29946);
or U34916 (N_34916,N_25038,N_26041);
or U34917 (N_34917,N_25339,N_29738);
nor U34918 (N_34918,N_25637,N_28501);
xnor U34919 (N_34919,N_25302,N_27256);
xnor U34920 (N_34920,N_25655,N_29560);
nor U34921 (N_34921,N_28445,N_28654);
xnor U34922 (N_34922,N_25161,N_27868);
nand U34923 (N_34923,N_29761,N_26524);
nand U34924 (N_34924,N_27968,N_28712);
xnor U34925 (N_34925,N_25442,N_29742);
nand U34926 (N_34926,N_27533,N_26545);
or U34927 (N_34927,N_29874,N_27223);
xnor U34928 (N_34928,N_25585,N_28456);
nor U34929 (N_34929,N_26601,N_28513);
xnor U34930 (N_34930,N_25651,N_28730);
or U34931 (N_34931,N_29565,N_27920);
nor U34932 (N_34932,N_26631,N_29896);
nand U34933 (N_34933,N_29558,N_28298);
xor U34934 (N_34934,N_29726,N_28847);
or U34935 (N_34935,N_29549,N_28729);
nor U34936 (N_34936,N_26185,N_26976);
nand U34937 (N_34937,N_25018,N_28123);
nand U34938 (N_34938,N_26338,N_27556);
or U34939 (N_34939,N_28244,N_26537);
or U34940 (N_34940,N_28050,N_26221);
nand U34941 (N_34941,N_25985,N_29068);
nand U34942 (N_34942,N_28334,N_29765);
nor U34943 (N_34943,N_25314,N_27707);
and U34944 (N_34944,N_29837,N_26295);
xor U34945 (N_34945,N_25589,N_26635);
nor U34946 (N_34946,N_29173,N_28635);
xor U34947 (N_34947,N_27283,N_27204);
nand U34948 (N_34948,N_28768,N_29787);
nor U34949 (N_34949,N_29863,N_28593);
nor U34950 (N_34950,N_28258,N_27809);
xnor U34951 (N_34951,N_26638,N_27784);
and U34952 (N_34952,N_27570,N_27732);
or U34953 (N_34953,N_27536,N_28044);
nor U34954 (N_34954,N_27812,N_26571);
and U34955 (N_34955,N_28069,N_28356);
and U34956 (N_34956,N_25305,N_28850);
and U34957 (N_34957,N_27884,N_29284);
and U34958 (N_34958,N_25832,N_28921);
xor U34959 (N_34959,N_26646,N_29074);
or U34960 (N_34960,N_26633,N_28202);
nor U34961 (N_34961,N_26582,N_28507);
nand U34962 (N_34962,N_25884,N_29607);
nor U34963 (N_34963,N_25060,N_25577);
and U34964 (N_34964,N_26802,N_28371);
xnor U34965 (N_34965,N_29799,N_28119);
or U34966 (N_34966,N_27077,N_28615);
nand U34967 (N_34967,N_25393,N_28820);
nand U34968 (N_34968,N_26041,N_28854);
nor U34969 (N_34969,N_28650,N_27370);
nor U34970 (N_34970,N_29132,N_28041);
or U34971 (N_34971,N_27792,N_27237);
or U34972 (N_34972,N_25414,N_29219);
nand U34973 (N_34973,N_27536,N_26922);
xor U34974 (N_34974,N_28945,N_29394);
nand U34975 (N_34975,N_28790,N_27183);
nand U34976 (N_34976,N_28128,N_25233);
and U34977 (N_34977,N_25568,N_25687);
and U34978 (N_34978,N_29544,N_26542);
and U34979 (N_34979,N_26655,N_27365);
nand U34980 (N_34980,N_28936,N_27313);
or U34981 (N_34981,N_28763,N_27177);
nand U34982 (N_34982,N_25205,N_29422);
nor U34983 (N_34983,N_29338,N_28355);
nand U34984 (N_34984,N_29209,N_27121);
nand U34985 (N_34985,N_25688,N_28252);
or U34986 (N_34986,N_25016,N_27015);
or U34987 (N_34987,N_29476,N_29004);
nor U34988 (N_34988,N_27254,N_25812);
nor U34989 (N_34989,N_28218,N_27783);
xor U34990 (N_34990,N_25578,N_27035);
nand U34991 (N_34991,N_28970,N_26127);
nor U34992 (N_34992,N_26395,N_27482);
and U34993 (N_34993,N_26180,N_26023);
xnor U34994 (N_34994,N_26208,N_26508);
xor U34995 (N_34995,N_29093,N_25096);
nor U34996 (N_34996,N_28875,N_28916);
nor U34997 (N_34997,N_25430,N_29341);
nand U34998 (N_34998,N_26166,N_25796);
xnor U34999 (N_34999,N_28383,N_29580);
nand U35000 (N_35000,N_34538,N_34036);
nand U35001 (N_35001,N_32431,N_31031);
nand U35002 (N_35002,N_31251,N_32067);
nor U35003 (N_35003,N_32268,N_34549);
nand U35004 (N_35004,N_30840,N_32908);
or U35005 (N_35005,N_33393,N_33497);
and U35006 (N_35006,N_33560,N_33549);
nor U35007 (N_35007,N_32889,N_31219);
nor U35008 (N_35008,N_33421,N_33412);
nand U35009 (N_35009,N_30688,N_30525);
and U35010 (N_35010,N_34791,N_30985);
nand U35011 (N_35011,N_32633,N_30966);
and U35012 (N_35012,N_31874,N_33568);
or U35013 (N_35013,N_34199,N_31741);
nor U35014 (N_35014,N_31752,N_32440);
nand U35015 (N_35015,N_32789,N_32470);
and U35016 (N_35016,N_34304,N_31249);
and U35017 (N_35017,N_32746,N_30786);
nand U35018 (N_35018,N_31570,N_33191);
or U35019 (N_35019,N_32629,N_30078);
and U35020 (N_35020,N_34873,N_34546);
nand U35021 (N_35021,N_32326,N_31533);
or U35022 (N_35022,N_33755,N_33288);
or U35023 (N_35023,N_31764,N_34466);
nor U35024 (N_35024,N_34092,N_33611);
and U35025 (N_35025,N_31236,N_31212);
or U35026 (N_35026,N_34990,N_32142);
xnor U35027 (N_35027,N_30658,N_34240);
and U35028 (N_35028,N_32356,N_34554);
nor U35029 (N_35029,N_30946,N_34817);
nor U35030 (N_35030,N_34797,N_32744);
xnor U35031 (N_35031,N_31282,N_32305);
nand U35032 (N_35032,N_31609,N_34456);
and U35033 (N_35033,N_32137,N_30549);
and U35034 (N_35034,N_32288,N_32405);
xnor U35035 (N_35035,N_32188,N_31837);
and U35036 (N_35036,N_31319,N_31182);
nor U35037 (N_35037,N_30811,N_33380);
nand U35038 (N_35038,N_32297,N_32684);
or U35039 (N_35039,N_32892,N_31008);
nand U35040 (N_35040,N_30652,N_32290);
xor U35041 (N_35041,N_32542,N_31929);
nand U35042 (N_35042,N_34056,N_33167);
nor U35043 (N_35043,N_33116,N_34155);
or U35044 (N_35044,N_30064,N_32500);
or U35045 (N_35045,N_31353,N_31638);
xor U35046 (N_35046,N_34094,N_31035);
nand U35047 (N_35047,N_32360,N_34574);
xor U35048 (N_35048,N_31542,N_31107);
nand U35049 (N_35049,N_33088,N_30940);
nand U35050 (N_35050,N_30687,N_33702);
xor U35051 (N_35051,N_33881,N_31198);
and U35052 (N_35052,N_30018,N_34945);
xnor U35053 (N_35053,N_31015,N_30794);
and U35054 (N_35054,N_32639,N_34951);
xnor U35055 (N_35055,N_32795,N_34750);
nand U35056 (N_35056,N_33573,N_30858);
or U35057 (N_35057,N_30425,N_32947);
or U35058 (N_35058,N_33169,N_30548);
nand U35059 (N_35059,N_33907,N_32233);
xnor U35060 (N_35060,N_30554,N_31655);
and U35061 (N_35061,N_34484,N_30350);
nor U35062 (N_35062,N_34086,N_34698);
nand U35063 (N_35063,N_33661,N_32589);
xnor U35064 (N_35064,N_34046,N_30187);
and U35065 (N_35065,N_34408,N_33496);
and U35066 (N_35066,N_32257,N_32365);
or U35067 (N_35067,N_32077,N_34838);
nand U35068 (N_35068,N_33632,N_33769);
and U35069 (N_35069,N_33397,N_33452);
and U35070 (N_35070,N_32557,N_30233);
xnor U35071 (N_35071,N_32753,N_32362);
xor U35072 (N_35072,N_32095,N_31998);
nor U35073 (N_35073,N_31750,N_31535);
nand U35074 (N_35074,N_31481,N_33679);
or U35075 (N_35075,N_33969,N_31339);
and U35076 (N_35076,N_30952,N_31322);
nand U35077 (N_35077,N_34650,N_33998);
or U35078 (N_35078,N_33882,N_32767);
or U35079 (N_35079,N_33043,N_34610);
nor U35080 (N_35080,N_32839,N_32541);
and U35081 (N_35081,N_33562,N_33791);
nand U35082 (N_35082,N_32818,N_34100);
nand U35083 (N_35083,N_33592,N_32309);
nand U35084 (N_35084,N_32285,N_32748);
and U35085 (N_35085,N_30844,N_34831);
nor U35086 (N_35086,N_34050,N_30628);
or U35087 (N_35087,N_31624,N_30224);
or U35088 (N_35088,N_30632,N_32241);
or U35089 (N_35089,N_31875,N_31746);
xor U35090 (N_35090,N_31981,N_31788);
xor U35091 (N_35091,N_31038,N_34804);
or U35092 (N_35092,N_31711,N_34087);
nand U35093 (N_35093,N_32112,N_31231);
and U35094 (N_35094,N_34453,N_31157);
nand U35095 (N_35095,N_34489,N_30085);
or U35096 (N_35096,N_33555,N_31414);
xor U35097 (N_35097,N_34236,N_33871);
or U35098 (N_35098,N_34904,N_31019);
nor U35099 (N_35099,N_34935,N_30958);
nor U35100 (N_35100,N_30755,N_33261);
xor U35101 (N_35101,N_34544,N_32458);
xor U35102 (N_35102,N_32595,N_31190);
nand U35103 (N_35103,N_30981,N_31923);
xor U35104 (N_35104,N_31623,N_32729);
nand U35105 (N_35105,N_31745,N_32199);
nor U35106 (N_35106,N_32336,N_31590);
nor U35107 (N_35107,N_31964,N_31857);
nor U35108 (N_35108,N_34064,N_34523);
xnor U35109 (N_35109,N_33122,N_31021);
nand U35110 (N_35110,N_33321,N_34424);
and U35111 (N_35111,N_32837,N_32054);
and U35112 (N_35112,N_31680,N_32177);
xor U35113 (N_35113,N_31861,N_31519);
or U35114 (N_35114,N_34387,N_30633);
and U35115 (N_35115,N_31254,N_32087);
nor U35116 (N_35116,N_34077,N_30691);
nor U35117 (N_35117,N_31354,N_31170);
xor U35118 (N_35118,N_34073,N_32606);
xor U35119 (N_35119,N_32946,N_32669);
nand U35120 (N_35120,N_31876,N_32190);
nand U35121 (N_35121,N_30039,N_34220);
nor U35122 (N_35122,N_34451,N_33461);
and U35123 (N_35123,N_32006,N_32666);
nand U35124 (N_35124,N_32555,N_30759);
xor U35125 (N_35125,N_34899,N_30196);
nor U35126 (N_35126,N_34914,N_33268);
or U35127 (N_35127,N_32221,N_30556);
nand U35128 (N_35128,N_33761,N_30870);
nand U35129 (N_35129,N_34105,N_30474);
and U35130 (N_35130,N_32307,N_34430);
and U35131 (N_35131,N_33964,N_32016);
xor U35132 (N_35132,N_32192,N_31303);
nand U35133 (N_35133,N_34250,N_30733);
and U35134 (N_35134,N_30322,N_32625);
nand U35135 (N_35135,N_33920,N_30345);
or U35136 (N_35136,N_33922,N_33509);
or U35137 (N_35137,N_32600,N_34004);
nor U35138 (N_35138,N_31869,N_33246);
nor U35139 (N_35139,N_34340,N_33439);
and U35140 (N_35140,N_33061,N_32989);
or U35141 (N_35141,N_32149,N_31499);
or U35142 (N_35142,N_31438,N_34009);
xnor U35143 (N_35143,N_32623,N_31286);
and U35144 (N_35144,N_32264,N_32978);
nand U35145 (N_35145,N_31677,N_30585);
and U35146 (N_35146,N_32870,N_30390);
or U35147 (N_35147,N_33996,N_33831);
xor U35148 (N_35148,N_30401,N_31900);
and U35149 (N_35149,N_31824,N_34291);
or U35150 (N_35150,N_32782,N_30243);
nand U35151 (N_35151,N_34630,N_33241);
nor U35152 (N_35152,N_32184,N_31662);
xnor U35153 (N_35153,N_30026,N_32621);
and U35154 (N_35154,N_34496,N_31281);
or U35155 (N_35155,N_34389,N_34794);
xnor U35156 (N_35156,N_30222,N_30572);
or U35157 (N_35157,N_33574,N_30800);
and U35158 (N_35158,N_33958,N_30129);
xnor U35159 (N_35159,N_33128,N_34908);
nand U35160 (N_35160,N_31531,N_34853);
nor U35161 (N_35161,N_30262,N_31435);
and U35162 (N_35162,N_34511,N_32531);
xnor U35163 (N_35163,N_30290,N_31132);
nor U35164 (N_35164,N_34798,N_34980);
or U35165 (N_35165,N_31980,N_30355);
nand U35166 (N_35166,N_33571,N_30827);
nor U35167 (N_35167,N_31368,N_30792);
nor U35168 (N_35168,N_30143,N_31300);
xnor U35169 (N_35169,N_30208,N_30573);
nand U35170 (N_35170,N_34720,N_30410);
xnor U35171 (N_35171,N_31790,N_34499);
and U35172 (N_35172,N_30889,N_32921);
xor U35173 (N_35173,N_30854,N_31886);
xor U35174 (N_35174,N_34557,N_31881);
or U35175 (N_35175,N_32056,N_33876);
nand U35176 (N_35176,N_31241,N_31243);
and U35177 (N_35177,N_33586,N_32240);
or U35178 (N_35178,N_33142,N_34471);
and U35179 (N_35179,N_30877,N_33019);
nand U35180 (N_35180,N_34618,N_30689);
or U35181 (N_35181,N_34502,N_34763);
xor U35182 (N_35182,N_34742,N_34918);
nor U35183 (N_35183,N_33857,N_30588);
and U35184 (N_35184,N_30875,N_31738);
or U35185 (N_35185,N_30964,N_34427);
and U35186 (N_35186,N_30957,N_33943);
and U35187 (N_35187,N_34171,N_31203);
nand U35188 (N_35188,N_33726,N_31871);
xnor U35189 (N_35189,N_33327,N_33029);
or U35190 (N_35190,N_30824,N_33223);
xnor U35191 (N_35191,N_34076,N_33620);
or U35192 (N_35192,N_32652,N_33607);
nor U35193 (N_35193,N_33753,N_30686);
and U35194 (N_35194,N_32964,N_31919);
and U35195 (N_35195,N_31997,N_30570);
nand U35196 (N_35196,N_31625,N_34774);
and U35197 (N_35197,N_32965,N_31124);
and U35198 (N_35198,N_30641,N_34604);
xnor U35199 (N_35199,N_31852,N_30988);
or U35200 (N_35200,N_31513,N_30301);
nor U35201 (N_35201,N_32327,N_31859);
or U35202 (N_35202,N_33877,N_32717);
and U35203 (N_35203,N_30145,N_34813);
nand U35204 (N_35204,N_32357,N_33704);
or U35205 (N_35205,N_31493,N_32770);
xnor U35206 (N_35206,N_33427,N_32738);
or U35207 (N_35207,N_31768,N_30168);
or U35208 (N_35208,N_34120,N_30151);
xnor U35209 (N_35209,N_32715,N_34870);
nor U35210 (N_35210,N_33060,N_32074);
or U35211 (N_35211,N_31393,N_31547);
or U35212 (N_35212,N_32665,N_30458);
or U35213 (N_35213,N_32133,N_34925);
and U35214 (N_35214,N_33546,N_33801);
nand U35215 (N_35215,N_33101,N_32413);
or U35216 (N_35216,N_34677,N_30447);
or U35217 (N_35217,N_34378,N_32752);
and U35218 (N_35218,N_34308,N_30690);
nor U35219 (N_35219,N_34059,N_31460);
nor U35220 (N_35220,N_33936,N_30341);
or U35221 (N_35221,N_31194,N_33294);
and U35222 (N_35222,N_32803,N_30919);
or U35223 (N_35223,N_32654,N_32857);
nand U35224 (N_35224,N_33822,N_34590);
or U35225 (N_35225,N_30561,N_30300);
nor U35226 (N_35226,N_31462,N_32788);
or U35227 (N_35227,N_33262,N_33697);
or U35228 (N_35228,N_31934,N_31659);
or U35229 (N_35229,N_33733,N_34216);
xnor U35230 (N_35230,N_34629,N_33691);
and U35231 (N_35231,N_34653,N_31598);
and U35232 (N_35232,N_34493,N_33621);
nand U35233 (N_35233,N_31708,N_34930);
or U35234 (N_35234,N_32914,N_33619);
and U35235 (N_35235,N_32804,N_32676);
xnor U35236 (N_35236,N_34124,N_31005);
or U35237 (N_35237,N_32709,N_32312);
xor U35238 (N_35238,N_31851,N_32143);
nor U35239 (N_35239,N_31806,N_34293);
nand U35240 (N_35240,N_33038,N_31895);
or U35241 (N_35241,N_31574,N_32529);
nand U35242 (N_35242,N_31388,N_34117);
or U35243 (N_35243,N_34419,N_34837);
xor U35244 (N_35244,N_33398,N_33593);
xnor U35245 (N_35245,N_34331,N_34102);
nor U35246 (N_35246,N_31389,N_33940);
xor U35247 (N_35247,N_34839,N_33935);
or U35248 (N_35248,N_30935,N_32934);
nor U35249 (N_35249,N_33174,N_32952);
nand U35250 (N_35250,N_31780,N_32945);
and U35251 (N_35251,N_31826,N_33501);
nor U35252 (N_35252,N_34369,N_32012);
nor U35253 (N_35253,N_33915,N_31080);
xor U35254 (N_35254,N_33768,N_31817);
and U35255 (N_35255,N_33670,N_33325);
xor U35256 (N_35256,N_30160,N_32527);
or U35257 (N_35257,N_34234,N_33222);
xnor U35258 (N_35258,N_34128,N_33135);
nand U35259 (N_35259,N_31293,N_34697);
nor U35260 (N_35260,N_30193,N_33519);
nand U35261 (N_35261,N_32602,N_30539);
nor U35262 (N_35262,N_32960,N_32929);
xnor U35263 (N_35263,N_33087,N_33422);
and U35264 (N_35264,N_34858,N_30834);
or U35265 (N_35265,N_34141,N_34101);
and U35266 (N_35266,N_32483,N_34846);
and U35267 (N_35267,N_34472,N_33093);
xnor U35268 (N_35268,N_30865,N_34452);
and U35269 (N_35269,N_31577,N_31762);
xor U35270 (N_35270,N_32535,N_30389);
and U35271 (N_35271,N_31222,N_32662);
or U35272 (N_35272,N_31619,N_31543);
or U35273 (N_35273,N_31647,N_32951);
or U35274 (N_35274,N_34907,N_33471);
and U35275 (N_35275,N_34663,N_32745);
xnor U35276 (N_35276,N_30154,N_33486);
xor U35277 (N_35277,N_30394,N_34354);
xnor U35278 (N_35278,N_33503,N_33291);
and U35279 (N_35279,N_32941,N_30882);
or U35280 (N_35280,N_30065,N_30926);
nand U35281 (N_35281,N_30663,N_30318);
nor U35282 (N_35282,N_30014,N_34151);
nor U35283 (N_35283,N_31694,N_31425);
and U35284 (N_35284,N_34473,N_33376);
nand U35285 (N_35285,N_32501,N_34396);
xnor U35286 (N_35286,N_30538,N_34275);
and U35287 (N_35287,N_30745,N_33508);
nand U35288 (N_35288,N_30651,N_33187);
xnor U35289 (N_35289,N_34140,N_33090);
and U35290 (N_35290,N_31306,N_34126);
and U35291 (N_35291,N_32522,N_31471);
nand U35292 (N_35292,N_32024,N_34806);
xnor U35293 (N_35293,N_31413,N_32512);
nor U35294 (N_35294,N_32497,N_31759);
nand U35295 (N_35295,N_30540,N_31226);
xor U35296 (N_35296,N_32502,N_31360);
xor U35297 (N_35297,N_31349,N_30897);
and U35298 (N_35298,N_32273,N_34208);
nand U35299 (N_35299,N_31630,N_30427);
and U35300 (N_35300,N_31473,N_34821);
or U35301 (N_35301,N_30010,N_34045);
and U35302 (N_35302,N_30264,N_30866);
xnor U35303 (N_35303,N_30861,N_30161);
nor U35304 (N_35304,N_34707,N_33548);
nand U35305 (N_35305,N_32217,N_30325);
or U35306 (N_35306,N_31576,N_30051);
nor U35307 (N_35307,N_32815,N_33602);
and U35308 (N_35308,N_32106,N_32841);
nand U35309 (N_35309,N_34439,N_30031);
or U35310 (N_35310,N_31893,N_34416);
and U35311 (N_35311,N_33027,N_33572);
and U35312 (N_35312,N_34764,N_31915);
or U35313 (N_35313,N_33228,N_32831);
or U35314 (N_35314,N_33933,N_30584);
xnor U35315 (N_35315,N_32656,N_30320);
nand U35316 (N_35316,N_30909,N_30209);
nor U35317 (N_35317,N_32569,N_32301);
nor U35318 (N_35318,N_33971,N_34558);
nor U35319 (N_35319,N_34048,N_31928);
nor U35320 (N_35320,N_33338,N_30551);
xnor U35321 (N_35321,N_30265,N_30750);
and U35322 (N_35322,N_30781,N_30612);
xnor U35323 (N_35323,N_30176,N_31100);
or U35324 (N_35324,N_31366,N_34668);
xnor U35325 (N_35325,N_30435,N_34719);
xor U35326 (N_35326,N_30197,N_33848);
nand U35327 (N_35327,N_30312,N_32830);
or U35328 (N_35328,N_34789,N_31468);
or U35329 (N_35329,N_30052,N_34700);
xor U35330 (N_35330,N_30823,N_31395);
xnor U35331 (N_35331,N_33561,N_32671);
nand U35332 (N_35332,N_33792,N_31283);
or U35333 (N_35333,N_33874,N_31514);
nand U35334 (N_35334,N_32775,N_31744);
nor U35335 (N_35335,N_32537,N_33221);
and U35336 (N_35336,N_32222,N_32247);
xnor U35337 (N_35337,N_30229,N_31309);
and U35338 (N_35338,N_32781,N_30841);
or U35339 (N_35339,N_33622,N_32597);
nand U35340 (N_35340,N_33146,N_34034);
nand U35341 (N_35341,N_30920,N_30250);
or U35342 (N_35342,N_33094,N_32287);
or U35343 (N_35343,N_30395,N_34039);
and U35344 (N_35344,N_32088,N_32879);
nor U35345 (N_35345,N_30146,N_33742);
nor U35346 (N_35346,N_32904,N_32319);
and U35347 (N_35347,N_31996,N_30796);
nor U35348 (N_35348,N_30880,N_31469);
nand U35349 (N_35349,N_32797,N_31010);
xnor U35350 (N_35350,N_34127,N_31736);
or U35351 (N_35351,N_31727,N_31036);
nor U35352 (N_35352,N_31795,N_30158);
xnor U35353 (N_35353,N_34560,N_33759);
nor U35354 (N_35354,N_30657,N_34768);
or U35355 (N_35355,N_32371,N_30313);
nand U35356 (N_35356,N_32253,N_32577);
nor U35357 (N_35357,N_30507,N_32099);
xor U35358 (N_35358,N_32072,N_32456);
or U35359 (N_35359,N_34884,N_34758);
nor U35360 (N_35360,N_31688,N_31179);
xor U35361 (N_35361,N_31451,N_33516);
nor U35362 (N_35362,N_32918,N_31020);
nor U35363 (N_35363,N_34682,N_30440);
nand U35364 (N_35364,N_33207,N_31160);
nand U35365 (N_35365,N_31683,N_30040);
xor U35366 (N_35366,N_32286,N_30953);
xor U35367 (N_35367,N_34204,N_33131);
nor U35368 (N_35368,N_33968,N_33558);
xnor U35369 (N_35369,N_32768,N_34706);
nand U35370 (N_35370,N_34344,N_31865);
or U35371 (N_35371,N_31705,N_32705);
nand U35372 (N_35372,N_31457,N_30816);
nor U35373 (N_35373,N_33069,N_32386);
nor U35374 (N_35374,N_30675,N_31568);
xor U35375 (N_35375,N_33766,N_30741);
nand U35376 (N_35376,N_33749,N_32708);
or U35377 (N_35377,N_32103,N_30429);
or U35378 (N_35378,N_30121,N_32341);
and U35379 (N_35379,N_32675,N_33247);
xor U35380 (N_35380,N_30375,N_32591);
xor U35381 (N_35381,N_30439,N_30363);
nor U35382 (N_35382,N_34476,N_34944);
or U35383 (N_35383,N_32911,N_30407);
or U35384 (N_35384,N_34031,N_32592);
nor U35385 (N_35385,N_30057,N_34891);
xor U35386 (N_35386,N_33036,N_31532);
and U35387 (N_35387,N_30452,N_33419);
and U35388 (N_35388,N_30600,N_30084);
and U35389 (N_35389,N_32802,N_32552);
and U35390 (N_35390,N_32491,N_32179);
and U35391 (N_35391,N_32399,N_30291);
and U35392 (N_35392,N_30522,N_34169);
xor U35393 (N_35393,N_31489,N_33667);
and U35394 (N_35394,N_32495,N_34982);
nand U35395 (N_35395,N_30106,N_30177);
xnor U35396 (N_35396,N_33790,N_31108);
xnor U35397 (N_35397,N_31995,N_33827);
and U35398 (N_35398,N_34157,N_34395);
or U35399 (N_35399,N_31025,N_34805);
and U35400 (N_35400,N_34449,N_33377);
xnor U35401 (N_35401,N_30028,N_34620);
and U35402 (N_35402,N_33627,N_31687);
or U35403 (N_35403,N_32648,N_30483);
or U35404 (N_35404,N_31663,N_32865);
and U35405 (N_35405,N_34265,N_32953);
nand U35406 (N_35406,N_34294,N_31954);
nand U35407 (N_35407,N_33719,N_34403);
nand U35408 (N_35408,N_30183,N_33804);
nand U35409 (N_35409,N_34210,N_32875);
xnor U35410 (N_35410,N_32463,N_32031);
xor U35411 (N_35411,N_34368,N_30102);
nor U35412 (N_35412,N_33298,N_31410);
xor U35413 (N_35413,N_32146,N_34961);
nand U35414 (N_35414,N_30062,N_30459);
xor U35415 (N_35415,N_33066,N_30284);
or U35416 (N_35416,N_30785,N_32342);
and U35417 (N_35417,N_33028,N_31152);
or U35418 (N_35418,N_30500,N_31097);
xor U35419 (N_35419,N_31841,N_31063);
and U35420 (N_35420,N_31678,N_30068);
xor U35421 (N_35421,N_31320,N_30139);
xnor U35422 (N_35422,N_33476,N_30075);
nor U35423 (N_35423,N_33757,N_30122);
or U35424 (N_35424,N_30697,N_30047);
or U35425 (N_35425,N_32955,N_30192);
or U35426 (N_35426,N_32814,N_33152);
nand U35427 (N_35427,N_33724,N_31866);
or U35428 (N_35428,N_33316,N_31175);
and U35429 (N_35429,N_33104,N_32044);
nor U35430 (N_35430,N_32182,N_31753);
and U35431 (N_35431,N_31381,N_33151);
xnor U35432 (N_35432,N_32355,N_32211);
nor U35433 (N_35433,N_32777,N_32741);
or U35434 (N_35434,N_33711,N_32271);
or U35435 (N_35435,N_34874,N_30608);
nand U35436 (N_35436,N_32765,N_32895);
nor U35437 (N_35437,N_30970,N_31940);
xor U35438 (N_35438,N_32393,N_32073);
nor U35439 (N_35439,N_32695,N_32065);
and U35440 (N_35440,N_30267,N_31094);
nor U35441 (N_35441,N_30782,N_30069);
nand U35442 (N_35442,N_31700,N_33656);
nand U35443 (N_35443,N_34184,N_34233);
or U35444 (N_35444,N_32736,N_30828);
or U35445 (N_35445,N_31073,N_30636);
nand U35446 (N_35446,N_33973,N_31208);
nor U35447 (N_35447,N_31653,N_33125);
xor U35448 (N_35448,N_33367,N_33331);
nor U35449 (N_35449,N_30488,N_31636);
xnor U35450 (N_35450,N_32565,N_31661);
xnor U35451 (N_35451,N_33363,N_30232);
nand U35452 (N_35452,N_33547,N_30076);
xnor U35453 (N_35453,N_34252,N_33959);
or U35454 (N_35454,N_31279,N_33781);
xnor U35455 (N_35455,N_34296,N_32873);
or U35456 (N_35456,N_34090,N_32219);
xnor U35457 (N_35457,N_34959,N_31023);
xnor U35458 (N_35458,N_30117,N_32332);
and U35459 (N_35459,N_34588,N_34415);
nor U35460 (N_35460,N_31846,N_33353);
xor U35461 (N_35461,N_34801,N_31390);
and U35462 (N_35462,N_31441,N_30976);
and U35463 (N_35463,N_32813,N_33771);
or U35464 (N_35464,N_30058,N_33931);
xnor U35465 (N_35465,N_32859,N_30619);
and U35466 (N_35466,N_34775,N_33689);
xnor U35467 (N_35467,N_32427,N_31838);
or U35468 (N_35468,N_30761,N_31452);
nor U35469 (N_35469,N_30236,N_32367);
nand U35470 (N_35470,N_34379,N_33946);
xnor U35471 (N_35471,N_31739,N_34053);
and U35472 (N_35472,N_30676,N_34316);
and U35473 (N_35473,N_33832,N_30293);
nand U35474 (N_35474,N_31580,N_34788);
or U35475 (N_35475,N_31141,N_31467);
and U35476 (N_35476,N_31692,N_32673);
and U35477 (N_35477,N_32350,N_30937);
xor U35478 (N_35478,N_30510,N_30030);
nand U35479 (N_35479,N_34080,N_33278);
nor U35480 (N_35480,N_33015,N_32683);
or U35481 (N_35481,N_34219,N_33039);
nor U35482 (N_35482,N_34373,N_30769);
or U35483 (N_35483,N_32966,N_32215);
and U35484 (N_35484,N_30529,N_30904);
xnor U35485 (N_35485,N_32269,N_32718);
and U35486 (N_35486,N_31784,N_34310);
xor U35487 (N_35487,N_30569,N_34782);
xor U35488 (N_35488,N_34382,N_30627);
xor U35489 (N_35489,N_32213,N_30990);
or U35490 (N_35490,N_30172,N_33609);
nor U35491 (N_35491,N_30077,N_33576);
or U35492 (N_35492,N_32825,N_32050);
nand U35493 (N_35493,N_30346,N_34109);
nand U35494 (N_35494,N_32267,N_32205);
nand U35495 (N_35495,N_32218,N_32171);
xor U35496 (N_35496,N_30837,N_33559);
nor U35497 (N_35497,N_30516,N_34149);
or U35498 (N_35498,N_34751,N_30083);
nor U35499 (N_35499,N_32335,N_30526);
nor U35500 (N_35500,N_31767,N_30616);
or U35501 (N_35501,N_34760,N_34063);
xor U35502 (N_35502,N_32270,N_32200);
or U35503 (N_35503,N_30441,N_33282);
nor U35504 (N_35504,N_34085,N_31536);
nor U35505 (N_35505,N_31658,N_34563);
or U35506 (N_35506,N_34865,N_32144);
and U35507 (N_35507,N_31382,N_32863);
or U35508 (N_35508,N_30005,N_32384);
nor U35509 (N_35509,N_34409,N_33355);
and U35510 (N_35510,N_32339,N_30002);
or U35511 (N_35511,N_34435,N_34723);
xnor U35512 (N_35512,N_30148,N_33156);
nor U35513 (N_35513,N_34400,N_32689);
xnor U35514 (N_35514,N_34417,N_34598);
nand U35515 (N_35515,N_32272,N_30024);
nor U35516 (N_35516,N_34327,N_34477);
xor U35517 (N_35517,N_33009,N_34299);
nor U35518 (N_35518,N_32315,N_32576);
nand U35519 (N_35519,N_31949,N_32869);
nor U35520 (N_35520,N_31966,N_31029);
nor U35521 (N_35521,N_33944,N_34426);
or U35522 (N_35522,N_31362,N_30324);
nand U35523 (N_35523,N_31255,N_32607);
or U35524 (N_35524,N_32148,N_30757);
nand U35525 (N_35525,N_34625,N_32560);
and U35526 (N_35526,N_30023,N_30557);
and U35527 (N_35527,N_34407,N_34665);
or U35528 (N_35528,N_31402,N_32845);
xor U35529 (N_35529,N_31823,N_34061);
and U35530 (N_35530,N_33690,N_30261);
nand U35531 (N_35531,N_32450,N_30927);
and U35532 (N_35532,N_32351,N_30822);
xor U35533 (N_35533,N_30163,N_33447);
or U35534 (N_35534,N_30931,N_32796);
xor U35535 (N_35535,N_32062,N_30144);
nor U35536 (N_35536,N_34676,N_30432);
nor U35537 (N_35537,N_32739,N_32994);
nand U35538 (N_35538,N_30285,N_32354);
xor U35539 (N_35539,N_32283,N_33880);
and U35540 (N_35540,N_32868,N_33924);
or U35541 (N_35541,N_33939,N_32277);
or U35542 (N_35542,N_34238,N_33491);
xnor U35543 (N_35543,N_32145,N_32370);
xor U35544 (N_35544,N_34114,N_33368);
or U35545 (N_35545,N_34834,N_34121);
or U35546 (N_35546,N_33214,N_30918);
xnor U35547 (N_35547,N_30704,N_31186);
and U35548 (N_35548,N_34527,N_31990);
nor U35549 (N_35549,N_30836,N_34529);
nor U35550 (N_35550,N_33623,N_30544);
or U35551 (N_35551,N_30956,N_30430);
nor U35552 (N_35552,N_34547,N_34679);
or U35553 (N_35553,N_33974,N_34249);
or U35554 (N_35554,N_33898,N_33437);
nor U35555 (N_35555,N_33820,N_31800);
xnor U35556 (N_35556,N_30977,N_30063);
and U35557 (N_35557,N_32838,N_33403);
or U35558 (N_35558,N_34615,N_34281);
or U35559 (N_35559,N_34507,N_32015);
or U35560 (N_35560,N_30524,N_30535);
xor U35561 (N_35561,N_31804,N_32020);
and U35562 (N_35562,N_33722,N_31524);
and U35563 (N_35563,N_31131,N_34991);
or U35564 (N_35564,N_33232,N_33853);
xor U35565 (N_35565,N_33815,N_31703);
nand U35566 (N_35566,N_32025,N_33414);
or U35567 (N_35567,N_30211,N_33587);
nor U35568 (N_35568,N_32396,N_31510);
xor U35569 (N_35569,N_33340,N_34418);
xor U35570 (N_35570,N_34569,N_30118);
or U35571 (N_35571,N_30595,N_33890);
and U35572 (N_35572,N_34552,N_30716);
nand U35573 (N_35573,N_32798,N_30424);
and U35574 (N_35574,N_34186,N_30624);
and U35575 (N_35575,N_30819,N_33057);
and U35576 (N_35576,N_34649,N_34548);
nor U35577 (N_35577,N_33919,N_33052);
or U35578 (N_35578,N_31047,N_31554);
nand U35579 (N_35579,N_31067,N_30127);
and U35580 (N_35580,N_31373,N_32189);
xnor U35581 (N_35581,N_32476,N_31747);
or U35582 (N_35582,N_34460,N_30520);
nor U35583 (N_35583,N_34670,N_32094);
or U35584 (N_35584,N_30388,N_31466);
nand U35585 (N_35585,N_33731,N_34543);
nor U35586 (N_35586,N_34277,N_31879);
nand U35587 (N_35587,N_34584,N_31994);
or U35588 (N_35588,N_32936,N_33710);
nand U35589 (N_35589,N_34158,N_33810);
and U35590 (N_35590,N_30356,N_33798);
and U35591 (N_35591,N_32670,N_33337);
nand U35592 (N_35592,N_34886,N_30577);
and U35593 (N_35593,N_30917,N_32254);
and U35594 (N_35594,N_30936,N_33530);
xor U35595 (N_35595,N_32419,N_33451);
xor U35596 (N_35596,N_31975,N_34479);
nand U35597 (N_35597,N_32039,N_33195);
nor U35598 (N_35598,N_32259,N_30692);
xor U35599 (N_35599,N_34332,N_30041);
xor U35600 (N_35600,N_34033,N_31465);
and U35601 (N_35601,N_34088,N_33784);
nor U35602 (N_35602,N_32840,N_34857);
or U35603 (N_35603,N_31220,N_32348);
nor U35604 (N_35604,N_31614,N_30302);
or U35605 (N_35605,N_34498,N_34897);
nand U35606 (N_35606,N_34261,N_33653);
nand U35607 (N_35607,N_30820,N_34826);
nand U35608 (N_35608,N_32195,N_34330);
and U35609 (N_35609,N_34492,N_32400);
or U35610 (N_35610,N_32722,N_31830);
and U35611 (N_35611,N_33588,N_32210);
nand U35612 (N_35612,N_31384,N_34026);
nand U35613 (N_35613,N_30174,N_31258);
nor U35614 (N_35614,N_33114,N_34165);
xnor U35615 (N_35615,N_34083,N_30428);
and U35616 (N_35616,N_33999,N_34889);
or U35617 (N_35617,N_31461,N_33952);
or U35618 (N_35618,N_31316,N_31211);
xor U35619 (N_35619,N_31724,N_33124);
nand U35620 (N_35620,N_33031,N_30805);
or U35621 (N_35621,N_31626,N_32426);
or U35622 (N_35622,N_34885,N_32225);
nand U35623 (N_35623,N_33362,N_32997);
or U35624 (N_35624,N_31145,N_32853);
xor U35625 (N_35625,N_32429,N_31178);
nand U35626 (N_35626,N_34132,N_31403);
and U35627 (N_35627,N_34565,N_33188);
xnor U35628 (N_35628,N_32248,N_33349);
or U35629 (N_35629,N_32762,N_31550);
nor U35630 (N_35630,N_31938,N_34328);
nand U35631 (N_35631,N_34346,N_31297);
xnor U35632 (N_35632,N_30715,N_30082);
nor U35633 (N_35633,N_31561,N_32246);
nor U35634 (N_35634,N_33049,N_32848);
or U35635 (N_35635,N_31668,N_30242);
and U35636 (N_35636,N_30306,N_30448);
xnor U35637 (N_35637,N_30737,N_33425);
or U35638 (N_35638,N_33237,N_32972);
and U35639 (N_35639,N_32122,N_34792);
or U35640 (N_35640,N_31261,N_30973);
xnor U35641 (N_35641,N_30027,N_33194);
nand U35642 (N_35642,N_33828,N_33307);
nand U35643 (N_35643,N_34860,N_33258);
nand U35644 (N_35644,N_32570,N_34280);
nor U35645 (N_35645,N_33443,N_34254);
nand U35646 (N_35646,N_30862,N_33903);
xnor U35647 (N_35647,N_30699,N_34580);
or U35648 (N_35648,N_34799,N_33252);
nand U35649 (N_35649,N_31599,N_33747);
xor U35650 (N_35650,N_31552,N_34749);
or U35651 (N_35651,N_31086,N_32151);
or U35652 (N_35652,N_30517,N_32826);
nor U35653 (N_35653,N_33489,N_31237);
xnor U35654 (N_35654,N_33721,N_32161);
xor U35655 (N_35655,N_30481,N_34264);
nand U35656 (N_35656,N_31715,N_30289);
or U35657 (N_35657,N_30565,N_32956);
and U35658 (N_35658,N_30848,N_32323);
xor U35659 (N_35659,N_32091,N_33779);
nand U35660 (N_35660,N_34242,N_33170);
xnor U35661 (N_35661,N_32982,N_31936);
and U35662 (N_35662,N_33430,N_34965);
and U35663 (N_35663,N_34709,N_31726);
nor U35664 (N_35664,N_31137,N_31257);
xnor U35665 (N_35665,N_32503,N_34223);
xnor U35666 (N_35666,N_33647,N_31517);
nand U35667 (N_35667,N_32703,N_34992);
or U35668 (N_35668,N_31154,N_30170);
or U35669 (N_35669,N_32694,N_34779);
nand U35670 (N_35670,N_32661,N_31357);
nand U35671 (N_35671,N_32078,N_34075);
and U35672 (N_35672,N_34830,N_34913);
nand U35673 (N_35673,N_30592,N_32209);
xor U35674 (N_35674,N_33440,N_32991);
nor U35675 (N_35675,N_32810,N_34600);
nor U35676 (N_35676,N_31246,N_30227);
or U35677 (N_35677,N_33844,N_31099);
and U35678 (N_35678,N_33041,N_33841);
or U35679 (N_35679,N_33020,N_32174);
xnor U35680 (N_35680,N_33963,N_34783);
or U35681 (N_35681,N_34772,N_31487);
nand U35682 (N_35682,N_33692,N_33554);
nand U35683 (N_35683,N_31645,N_32156);
or U35684 (N_35684,N_31486,N_30408);
nand U35685 (N_35685,N_32478,N_34425);
or U35686 (N_35686,N_34936,N_30932);
nand U35687 (N_35687,N_32707,N_33660);
nor U35688 (N_35688,N_30392,N_31399);
xnor U35689 (N_35689,N_34634,N_31809);
xnor U35690 (N_35690,N_33078,N_30668);
and U35691 (N_35691,N_32706,N_34734);
and U35692 (N_35692,N_34360,N_30705);
xnor U35693 (N_35693,N_33364,N_32017);
and U35694 (N_35694,N_33986,N_31159);
or U35695 (N_35695,N_34333,N_33780);
xor U35696 (N_35696,N_32725,N_32163);
xor U35697 (N_35697,N_31690,N_31840);
nor U35698 (N_35698,N_33400,N_33409);
or U35699 (N_35699,N_34465,N_31167);
nor U35700 (N_35700,N_31165,N_30167);
or U35701 (N_35701,N_33255,N_34659);
xnor U35702 (N_35702,N_33677,N_33396);
xor U35703 (N_35703,N_30270,N_34729);
xor U35704 (N_35704,N_30329,N_34652);
or U35705 (N_35705,N_31347,N_33825);
and U35706 (N_35706,N_33916,N_30527);
and U35707 (N_35707,N_34248,N_32959);
xnor U35708 (N_35708,N_30029,N_33674);
xor U35709 (N_35709,N_34535,N_32420);
xor U35710 (N_35710,N_33138,N_32053);
or U35711 (N_35711,N_32764,N_34043);
or U35712 (N_35712,N_30879,N_31555);
xnor U35713 (N_35713,N_33240,N_31456);
and U35714 (N_35714,N_32776,N_34947);
xor U35715 (N_35715,N_32435,N_32925);
xor U35716 (N_35716,N_34747,N_32720);
xor U35717 (N_35717,N_32410,N_30249);
nor U35718 (N_35718,N_34269,N_33299);
or U35719 (N_35719,N_30316,N_30693);
xnor U35720 (N_35720,N_34695,N_32422);
nor U35721 (N_35721,N_32833,N_34509);
xnor U35722 (N_35722,N_32646,N_34581);
nand U35723 (N_35723,N_33625,N_33004);
xor U35724 (N_35724,N_32505,N_33468);
nor U35725 (N_35725,N_30043,N_33648);
nand U35726 (N_35726,N_33345,N_30983);
xor U35727 (N_35727,N_33663,N_31204);
xnor U35728 (N_35728,N_33068,N_33531);
and U35729 (N_35729,N_30776,N_34638);
and U35730 (N_35730,N_30808,N_32906);
or U35731 (N_35731,N_34404,N_30466);
nor U35732 (N_35732,N_31868,N_30764);
nor U35733 (N_35733,N_34325,N_30241);
nor U35734 (N_35734,N_32134,N_32526);
nand U35735 (N_35735,N_34470,N_32856);
and U35736 (N_35736,N_32444,N_33339);
nor U35737 (N_35737,N_33525,N_33474);
xor U35738 (N_35738,N_33106,N_34006);
or U35739 (N_35739,N_31558,N_30700);
or U35740 (N_35740,N_31829,N_33517);
xor U35741 (N_35741,N_33109,N_31247);
and U35742 (N_35742,N_34674,N_31062);
nand U35743 (N_35743,N_33809,N_32383);
xnor U35744 (N_35744,N_30116,N_32004);
nor U35745 (N_35745,N_32058,N_32749);
xnor U35746 (N_35746,N_33161,N_32519);
and U35747 (N_35747,N_30560,N_33048);
and U35748 (N_35748,N_33313,N_31172);
or U35749 (N_35749,N_32252,N_32084);
xor U35750 (N_35750,N_31722,N_33723);
nand U35751 (N_35751,N_34585,N_33287);
nor U35752 (N_35752,N_34855,N_32786);
or U35753 (N_35753,N_33144,N_31464);
nand U35754 (N_35754,N_33867,N_34434);
or U35755 (N_35755,N_31064,N_32185);
nor U35756 (N_35756,N_33285,N_32548);
xnor U35757 (N_35757,N_30226,N_33650);
xnor U35758 (N_35758,N_34969,N_33712);
and U35759 (N_35759,N_31960,N_31057);
nor U35760 (N_35760,N_33025,N_32640);
nand U35761 (N_35761,N_34137,N_32352);
and U35762 (N_35762,N_34012,N_33834);
or U35763 (N_35763,N_32872,N_34463);
or U35764 (N_35764,N_31916,N_34079);
xnor U35765 (N_35765,N_30537,N_31839);
or U35766 (N_35766,N_33030,N_33098);
or U35767 (N_35767,N_30453,N_30980);
xnor U35768 (N_35768,N_34741,N_30634);
and U35769 (N_35769,N_34540,N_30485);
and U35770 (N_35770,N_30072,N_31491);
or U35771 (N_35771,N_34376,N_33595);
nand U35772 (N_35772,N_32414,N_33213);
and U35773 (N_35773,N_31470,N_32877);
and U35774 (N_35774,N_33870,N_33359);
xor U35775 (N_35775,N_31440,N_30442);
or U35776 (N_35776,N_34450,N_31386);
xnor U35777 (N_35777,N_31449,N_31921);
or U35778 (N_35778,N_33118,N_30799);
nor U35779 (N_35779,N_34622,N_33005);
or U35780 (N_35780,N_32465,N_32381);
and U35781 (N_35781,N_34097,N_33628);
xnor U35782 (N_35782,N_30812,N_33688);
xnor U35783 (N_35783,N_30279,N_33190);
xnor U35784 (N_35784,N_32582,N_30685);
or U35785 (N_35785,N_31484,N_33159);
and U35786 (N_35786,N_33072,N_34038);
and U35787 (N_35787,N_33800,N_33817);
nand U35788 (N_35788,N_32645,N_32643);
nor U35789 (N_35789,N_30189,N_30383);
or U35790 (N_35790,N_30006,N_30762);
nor U35791 (N_35791,N_30922,N_31991);
or U35792 (N_35792,N_31660,N_32580);
xnor U35793 (N_35793,N_33694,N_33035);
xnor U35794 (N_35794,N_32318,N_30421);
xnor U35795 (N_35795,N_30613,N_34481);
or U35796 (N_35796,N_33344,N_32398);
or U35797 (N_35797,N_34769,N_34883);
nand U35798 (N_35798,N_34894,N_31071);
nand U35799 (N_35799,N_31052,N_33381);
nor U35800 (N_35800,N_33754,N_30670);
xor U35801 (N_35801,N_31351,N_34550);
or U35802 (N_35802,N_34671,N_30914);
xor U35803 (N_35803,N_32878,N_34461);
and U35804 (N_35804,N_32510,N_31214);
and U35805 (N_35805,N_32011,N_34909);
nand U35806 (N_35806,N_33310,N_32329);
or U35807 (N_35807,N_32130,N_30943);
nand U35808 (N_35808,N_31301,N_31843);
xor U35809 (N_35809,N_32170,N_33434);
nor U35810 (N_35810,N_30860,N_33387);
nor U35811 (N_35811,N_31967,N_34974);
nand U35812 (N_35812,N_31122,N_32711);
nor U35813 (N_35813,N_31259,N_32913);
nand U35814 (N_35814,N_34374,N_31693);
or U35815 (N_35815,N_34895,N_30337);
nand U35816 (N_35816,N_34448,N_33487);
or U35817 (N_35817,N_31447,N_32926);
xnor U35818 (N_35818,N_30090,N_31608);
nand U35819 (N_35819,N_31507,N_31883);
nand U35820 (N_35820,N_34669,N_33323);
xor U35821 (N_35821,N_30022,N_32035);
and U35822 (N_35822,N_32667,N_34644);
nand U35823 (N_35823,N_33193,N_31618);
xnor U35824 (N_35824,N_31006,N_33073);
nand U35825 (N_35825,N_34521,N_32766);
or U35826 (N_35826,N_31268,N_31430);
or U35827 (N_35827,N_31078,N_30353);
and U35828 (N_35828,N_33488,N_32887);
xnor U35829 (N_35829,N_30961,N_33895);
or U35830 (N_35830,N_32896,N_34051);
nand U35831 (N_35831,N_32461,N_32256);
and U35832 (N_35832,N_33365,N_32567);
nor U35833 (N_35833,N_32829,N_33407);
nor U35834 (N_35834,N_33472,N_34422);
nand U35835 (N_35835,N_33886,N_32983);
and U35836 (N_35836,N_33492,N_33204);
xnor U35837 (N_35837,N_31567,N_32971);
nand U35838 (N_35838,N_30607,N_31889);
and U35839 (N_35839,N_34807,N_31898);
nor U35840 (N_35840,N_32561,N_32617);
nor U35841 (N_35841,N_30276,N_32479);
and U35842 (N_35842,N_33604,N_30277);
or U35843 (N_35843,N_34251,N_30112);
xnor U35844 (N_35844,N_33914,N_32518);
and U35845 (N_35845,N_32702,N_32801);
xor U35846 (N_35846,N_33987,N_33811);
nand U35847 (N_35847,N_33417,N_34297);
nand U35848 (N_35848,N_31116,N_34429);
or U35849 (N_35849,N_32847,N_32598);
and U35850 (N_35850,N_31287,N_31920);
nand U35851 (N_35851,N_30414,N_33217);
xor U35852 (N_35852,N_34703,N_30469);
nor U35853 (N_35853,N_33937,N_33989);
nand U35854 (N_35854,N_32821,N_30225);
nand U35855 (N_35855,N_31405,N_32849);
or U35856 (N_35856,N_33037,N_30609);
or U35857 (N_35857,N_33957,N_30594);
and U35858 (N_35858,N_31695,N_33645);
xnor U35859 (N_35859,N_30644,N_32785);
and U35860 (N_35860,N_32284,N_30944);
nand U35861 (N_35861,N_30708,N_30945);
nor U35862 (N_35862,N_30296,N_32509);
nand U35863 (N_35863,N_31091,N_32604);
nor U35864 (N_35864,N_30868,N_33108);
and U35865 (N_35865,N_34993,N_33736);
nand U35866 (N_35866,N_34028,N_32037);
nand U35867 (N_35867,N_33875,N_33175);
and U35868 (N_35868,N_33714,N_33921);
or U35869 (N_35869,N_34728,N_32737);
nand U35870 (N_35870,N_31559,N_31833);
xnor U35871 (N_35871,N_33231,N_31406);
and U35872 (N_35872,N_31371,N_31401);
xnor U35873 (N_35873,N_31359,N_34551);
xnor U35874 (N_35874,N_31537,N_32274);
xor U35875 (N_35875,N_31022,N_30159);
nor U35876 (N_35876,N_32530,N_31761);
xor U35877 (N_35877,N_31093,N_32790);
nor U35878 (N_35878,N_34999,N_32726);
or U35879 (N_35879,N_30825,N_31267);
nand U35880 (N_35880,N_32637,N_33543);
nor U35881 (N_35881,N_32340,N_34320);
or U35882 (N_35882,N_33390,N_34878);
nand U35883 (N_35883,N_30604,N_30258);
xnor U35884 (N_35884,N_34603,N_34645);
nor U35885 (N_35885,N_30991,N_30107);
or U35886 (N_35886,N_32610,N_33007);
or U35887 (N_35887,N_32235,N_31478);
nand U35888 (N_35888,N_32232,N_30271);
nand U35889 (N_35889,N_31607,N_34825);
nand U35890 (N_35890,N_31704,N_31947);
xor U35891 (N_35891,N_34490,N_32359);
and U35892 (N_35892,N_34892,N_31757);
and U35893 (N_35893,N_33885,N_32186);
nor U35894 (N_35894,N_31437,N_34657);
nand U35895 (N_35895,N_32320,N_30778);
nor U35896 (N_35896,N_31540,N_32893);
or U35897 (N_35897,N_30842,N_32477);
and U35898 (N_35898,N_31217,N_34202);
and U35899 (N_35899,N_30259,N_34491);
and U35900 (N_35900,N_30237,N_31977);
or U35901 (N_35901,N_30984,N_32158);
nor U35902 (N_35902,N_31411,N_30743);
nand U35903 (N_35903,N_33977,N_31557);
nand U35904 (N_35904,N_32314,N_30801);
and U35905 (N_35905,N_32636,N_34273);
nand U35906 (N_35906,N_32172,N_32558);
nor U35907 (N_35907,N_33685,N_31586);
nand U35908 (N_35908,N_33833,N_34049);
xnor U35909 (N_35909,N_33157,N_30767);
or U35910 (N_35910,N_30153,N_30263);
xor U35911 (N_35911,N_30310,N_32533);
xnor U35912 (N_35912,N_32412,N_31126);
and U35913 (N_35913,N_34533,N_32931);
nor U35914 (N_35914,N_34687,N_32346);
nand U35915 (N_35915,N_34289,N_34940);
or U35916 (N_35916,N_30110,N_32772);
nand U35917 (N_35917,N_34849,N_34568);
nand U35918 (N_35918,N_32583,N_34932);
nor U35919 (N_35919,N_30770,N_31195);
xor U35920 (N_35920,N_30864,N_30340);
xor U35921 (N_35921,N_34385,N_31476);
nand U35922 (N_35922,N_32915,N_31164);
xor U35923 (N_35923,N_33201,N_30454);
and U35924 (N_35924,N_31017,N_30587);
and U35925 (N_35925,N_34530,N_34694);
and U35926 (N_35926,N_34337,N_31370);
xor U35927 (N_35927,N_30821,N_32430);
xor U35928 (N_35928,N_30286,N_30484);
xnor U35929 (N_35929,N_31667,N_32942);
or U35930 (N_35930,N_31814,N_33145);
or U35931 (N_35931,N_31290,N_34156);
or U35932 (N_35932,N_33236,N_32442);
nor U35933 (N_35933,N_33123,N_30996);
nor U35934 (N_35934,N_31825,N_30379);
nand U35935 (N_35935,N_30297,N_32051);
xnor U35936 (N_35936,N_34954,N_33438);
xor U35937 (N_35937,N_34276,N_31787);
or U35938 (N_35938,N_30257,N_34745);
nor U35939 (N_35939,N_33606,N_32009);
or U35940 (N_35940,N_33816,N_30832);
or U35941 (N_35941,N_30220,N_33413);
nand U35942 (N_35942,N_31400,N_30790);
and U35943 (N_35943,N_31740,N_31490);
and U35944 (N_35944,N_31065,N_32928);
nand U35945 (N_35945,N_30221,N_31959);
xor U35946 (N_35946,N_32076,N_33470);
and U35947 (N_35947,N_31174,N_30740);
or U35948 (N_35948,N_31951,N_33954);
nand U35949 (N_35949,N_31163,N_32173);
or U35950 (N_35950,N_31941,N_33673);
and U35951 (N_35951,N_33750,N_33311);
nor U35952 (N_35952,N_33613,N_30777);
and U35953 (N_35953,N_32380,N_30532);
nor U35954 (N_35954,N_30660,N_33348);
xor U35955 (N_35955,N_33752,N_31153);
nor U35956 (N_35956,N_32401,N_33082);
and U35957 (N_35957,N_32998,N_31066);
and U35958 (N_35958,N_31189,N_31818);
or U35959 (N_35959,N_33675,N_31272);
xnor U35960 (N_35960,N_32668,N_30491);
and U35961 (N_35961,N_34302,N_33658);
nand U35962 (N_35962,N_31993,N_31387);
and U35963 (N_35963,N_34989,N_34113);
xnor U35964 (N_35964,N_30032,N_33389);
and U35965 (N_35965,N_30004,N_34893);
and U35966 (N_35966,N_30783,N_32373);
and U35967 (N_35967,N_31495,N_30712);
xor U35968 (N_35968,N_30119,N_33120);
nor U35969 (N_35969,N_34710,N_31556);
nand U35970 (N_35970,N_33900,N_34288);
xor U35971 (N_35971,N_33636,N_30212);
nor U35972 (N_35972,N_30579,N_31127);
nor U35973 (N_35973,N_34744,N_32933);
nand U35974 (N_35974,N_33358,N_34303);
or U35975 (N_35975,N_33051,N_30201);
and U35976 (N_35976,N_34911,N_31146);
nand U35977 (N_35977,N_33659,N_34214);
nor U35978 (N_35978,N_31068,N_33245);
or U35979 (N_35979,N_34739,N_34110);
or U35980 (N_35980,N_32337,N_32899);
nor U35981 (N_35981,N_31836,N_30434);
and U35982 (N_35982,N_31075,N_34570);
and U35983 (N_35983,N_34027,N_30698);
nor U35984 (N_35984,N_32407,N_34879);
or U35985 (N_35985,N_33725,N_33283);
xnor U35986 (N_35986,N_30661,N_34060);
or U35987 (N_35987,N_31248,N_32980);
nand U35988 (N_35988,N_33640,N_34562);
or U35989 (N_35989,N_31506,N_34666);
nand U35990 (N_35990,N_34812,N_31791);
and U35991 (N_35991,N_34247,N_33843);
and U35992 (N_35992,N_32492,N_34194);
and U35993 (N_35993,N_32724,N_30589);
and U35994 (N_35994,N_33557,N_33113);
nor U35995 (N_35995,N_33990,N_33322);
or U35996 (N_35996,N_32379,N_34985);
and U35997 (N_35997,N_34457,N_30969);
and U35998 (N_35998,N_32366,N_30019);
nor U35999 (N_35999,N_33859,N_34468);
nand U36000 (N_36000,N_34357,N_33010);
nor U36001 (N_36001,N_31924,N_31294);
nand U36002 (N_36002,N_30273,N_33858);
nor U36003 (N_36003,N_34129,N_32939);
or U36004 (N_36004,N_33079,N_34052);
nor U36005 (N_36005,N_30511,N_32026);
and U36006 (N_36006,N_34654,N_33888);
nor U36007 (N_36007,N_33256,N_31742);
xnor U36008 (N_36008,N_33328,N_32927);
nor U36009 (N_36009,N_32079,N_34661);
and U36010 (N_36010,N_31847,N_32816);
nor U36011 (N_36011,N_33680,N_31045);
nor U36012 (N_36012,N_32860,N_34420);
xnor U36013 (N_36013,N_31862,N_34777);
nor U36014 (N_36014,N_34957,N_32187);
and U36015 (N_36015,N_30734,N_30294);
nor U36016 (N_36016,N_34833,N_33192);
nor U36017 (N_36017,N_31657,N_31545);
and U36018 (N_36018,N_32375,N_33894);
or U36019 (N_36019,N_34197,N_33394);
nor U36020 (N_36020,N_33239,N_33506);
xnor U36021 (N_36021,N_34081,N_30411);
nor U36022 (N_36022,N_34721,N_31908);
or U36023 (N_36023,N_33671,N_30642);
nor U36024 (N_36024,N_31758,N_30863);
nand U36025 (N_36025,N_33789,N_30646);
or U36026 (N_36026,N_31424,N_30165);
nand U36027 (N_36027,N_31429,N_34987);
nand U36028 (N_36028,N_33951,N_30999);
nor U36029 (N_36029,N_34014,N_32275);
nand U36030 (N_36030,N_30826,N_31138);
nor U36031 (N_36031,N_32292,N_30468);
xnor U36032 (N_36032,N_30519,N_31546);
xor U36033 (N_36033,N_30563,N_30338);
and U36034 (N_36034,N_31773,N_31206);
xor U36035 (N_36035,N_30482,N_32000);
nor U36036 (N_36036,N_34480,N_31044);
nor U36037 (N_36037,N_33695,N_30810);
nor U36038 (N_36038,N_31974,N_30552);
or U36039 (N_36039,N_32207,N_31376);
nor U36040 (N_36040,N_34245,N_32353);
xnor U36041 (N_36041,N_34506,N_33301);
nand U36042 (N_36042,N_33084,N_34370);
nand U36043 (N_36043,N_33405,N_30347);
nand U36044 (N_36044,N_34266,N_31213);
or U36045 (N_36045,N_31229,N_34790);
or U36046 (N_36046,N_33099,N_34556);
and U36047 (N_36047,N_34716,N_31291);
or U36048 (N_36048,N_31482,N_33873);
or U36049 (N_36049,N_34537,N_30571);
nor U36050 (N_36050,N_33184,N_34229);
nand U36051 (N_36051,N_32150,N_32674);
and U36052 (N_36052,N_32228,N_34931);
nor U36053 (N_36053,N_30130,N_32508);
nor U36054 (N_36054,N_34253,N_31055);
xnor U36055 (N_36055,N_34752,N_30094);
and U36056 (N_36056,N_34759,N_32310);
nand U36057 (N_36057,N_33378,N_34108);
nand U36058 (N_36058,N_30706,N_32663);
or U36059 (N_36059,N_32719,N_31342);
nand U36060 (N_36060,N_32063,N_31450);
or U36061 (N_36061,N_33566,N_30833);
and U36062 (N_36062,N_34428,N_31685);
xnor U36063 (N_36063,N_33823,N_34841);
and U36064 (N_36064,N_31142,N_32474);
nor U36065 (N_36065,N_32507,N_34054);
nand U36066 (N_36066,N_33652,N_31539);
or U36067 (N_36067,N_34306,N_34257);
and U36068 (N_36068,N_34942,N_30815);
or U36069 (N_36069,N_30443,N_33705);
or U36070 (N_36070,N_34915,N_32962);
nand U36071 (N_36071,N_33696,N_33267);
or U36072 (N_36072,N_31612,N_31600);
and U36073 (N_36073,N_33788,N_30558);
or U36074 (N_36074,N_34082,N_31813);
xnor U36075 (N_36075,N_32279,N_31786);
nor U36076 (N_36076,N_34692,N_33601);
or U36077 (N_36077,N_31032,N_34364);
nand U36078 (N_36078,N_30012,N_32014);
and U36079 (N_36079,N_31305,N_34827);
nand U36080 (N_36080,N_31573,N_32443);
and U36081 (N_36081,N_34997,N_33735);
or U36082 (N_36082,N_33693,N_34188);
xor U36083 (N_36083,N_33179,N_32198);
nand U36084 (N_36084,N_33580,N_31815);
or U36085 (N_36085,N_30659,N_33250);
nand U36086 (N_36086,N_30911,N_31584);
and U36087 (N_36087,N_34903,N_34948);
and U36088 (N_36088,N_34290,N_30629);
nand U36089 (N_36089,N_34740,N_33026);
or U36090 (N_36090,N_33545,N_33681);
nor U36091 (N_36091,N_31803,N_33186);
xor U36092 (N_36092,N_33366,N_31180);
xor U36093 (N_36093,N_30445,N_33289);
nand U36094 (N_36094,N_31596,N_31404);
nand U36095 (N_36095,N_33202,N_32686);
xor U36096 (N_36096,N_30317,N_31380);
and U36097 (N_36097,N_33799,N_31326);
xor U36098 (N_36098,N_33347,N_31642);
xnor U36099 (N_36099,N_34756,N_30493);
nand U36100 (N_36100,N_32075,N_33083);
or U36101 (N_36101,N_32974,N_34875);
nand U36102 (N_36102,N_32001,N_34068);
and U36103 (N_36103,N_33149,N_34596);
xor U36104 (N_36104,N_32963,N_32249);
nor U36105 (N_36105,N_31459,N_34513);
nand U36106 (N_36106,N_34341,N_33295);
nor U36107 (N_36107,N_33356,N_30288);
xor U36108 (N_36108,N_32787,N_30818);
or U36109 (N_36109,N_31930,N_33166);
or U36110 (N_36110,N_34164,N_32572);
xnor U36111 (N_36111,N_31631,N_33455);
xor U36112 (N_36112,N_30336,N_34057);
nand U36113 (N_36113,N_30240,N_30169);
nand U36114 (N_36114,N_31882,N_30404);
nand U36115 (N_36115,N_32135,N_33458);
nand U36116 (N_36116,N_30382,N_31148);
xor U36117 (N_36117,N_31569,N_32242);
nor U36118 (N_36118,N_34977,N_31777);
nor U36119 (N_36119,N_34522,N_31329);
nand U36120 (N_36120,N_32255,N_34362);
or U36121 (N_36121,N_34962,N_31117);
nor U36122 (N_36122,N_31216,N_33129);
nor U36123 (N_36123,N_33901,N_33738);
nor U36124 (N_36124,N_30011,N_34138);
and U36125 (N_36125,N_34474,N_32042);
nand U36126 (N_36126,N_30748,N_31615);
nor U36127 (N_36127,N_30732,N_31168);
xnor U36128 (N_36128,N_32261,N_30721);
or U36129 (N_36129,N_30528,N_34803);
and U36130 (N_36130,N_32657,N_34375);
nor U36131 (N_36131,N_33532,N_30036);
or U36132 (N_36132,N_31083,N_34335);
nor U36133 (N_36133,N_33281,N_31252);
nand U36134 (N_36134,N_31053,N_34844);
or U36135 (N_36135,N_34771,N_30583);
and U36136 (N_36136,N_33334,N_34847);
and U36137 (N_36137,N_32033,N_34125);
nor U36138 (N_36138,N_31385,N_31521);
or U36139 (N_36139,N_30747,N_33806);
and U36140 (N_36140,N_32432,N_31106);
or U36141 (N_36141,N_30274,N_34258);
nand U36142 (N_36142,N_30681,N_33276);
and U36143 (N_36143,N_31096,N_32109);
nand U36144 (N_36144,N_32057,N_31644);
xnor U36145 (N_36145,N_34268,N_33699);
or U36146 (N_36146,N_34691,N_30021);
and U36147 (N_36147,N_34401,N_31743);
or U36148 (N_36148,N_31505,N_32389);
nor U36149 (N_36149,N_30061,N_33080);
and U36150 (N_36150,N_31419,N_33585);
nor U36151 (N_36151,N_32969,N_32013);
nand U36152 (N_36152,N_34816,N_33598);
and U36153 (N_36153,N_31069,N_33993);
and U36154 (N_36154,N_31523,N_31765);
nand U36155 (N_36155,N_30971,N_31398);
xnor U36156 (N_36156,N_33401,N_31943);
xnor U36157 (N_36157,N_31903,N_31613);
and U36158 (N_36158,N_33432,N_31674);
xnor U36159 (N_36159,N_32759,N_34017);
nor U36160 (N_36160,N_30942,N_30384);
or U36161 (N_36161,N_33091,N_32363);
nor U36162 (N_36162,N_30103,N_30091);
nand U36163 (N_36163,N_33199,N_31014);
nand U36164 (N_36164,N_34019,N_30109);
nor U36165 (N_36165,N_30625,N_34662);
nor U36166 (N_36166,N_32687,N_30674);
xor U36167 (N_36167,N_31088,N_30218);
nand U36168 (N_36168,N_34811,N_31679);
xor U36169 (N_36169,N_32052,N_33617);
and U36170 (N_36170,N_31651,N_33495);
and U36171 (N_36171,N_33100,N_30887);
xnor U36172 (N_36172,N_32635,N_34820);
xnor U36173 (N_36173,N_33869,N_32119);
xnor U36174 (N_36174,N_31910,N_31332);
or U36175 (N_36175,N_32237,N_33826);
and U36176 (N_36176,N_33046,N_33225);
and U36177 (N_36177,N_31723,N_33164);
or U36178 (N_36178,N_31110,N_32475);
and U36179 (N_36179,N_32032,N_30035);
or U36180 (N_36180,N_30883,N_30393);
nor U36181 (N_36181,N_31606,N_32783);
or U36182 (N_36182,N_33821,N_32364);
or U36183 (N_36183,N_32160,N_32626);
nand U36184 (N_36184,N_33515,N_34591);
and U36185 (N_36185,N_31264,N_34766);
and U36186 (N_36186,N_34753,N_34345);
nand U36187 (N_36187,N_31832,N_30731);
nand U36188 (N_36188,N_34518,N_30309);
xnor U36189 (N_36189,N_34748,N_31113);
and U36190 (N_36190,N_34953,N_33785);
or U36191 (N_36191,N_33635,N_30376);
nand U36192 (N_36192,N_31292,N_33955);
and U36193 (N_36193,N_31760,N_32611);
or U36194 (N_36194,N_33158,N_34244);
or U36195 (N_36195,N_31751,N_34864);
nand U36196 (N_36196,N_30846,N_31565);
or U36197 (N_36197,N_30667,N_32957);
nor U36198 (N_36198,N_32609,N_30568);
nand U36199 (N_36199,N_30803,N_33866);
and U36200 (N_36200,N_32328,N_31896);
xnor U36201 (N_36201,N_32751,N_30147);
and U36202 (N_36202,N_31714,N_32603);
xnor U36203 (N_36203,N_32343,N_32018);
nand U36204 (N_36204,N_32763,N_32846);
xnor U36205 (N_36205,N_30649,N_32943);
nor U36206 (N_36206,N_32449,N_31805);
or U36207 (N_36207,N_30003,N_31643);
and U36208 (N_36208,N_32950,N_33463);
nor U36209 (N_36209,N_30728,N_32549);
and U36210 (N_36210,N_34020,N_33861);
xor U36211 (N_36211,N_30843,N_31365);
nor U36212 (N_36212,N_33460,N_32514);
xnor U36213 (N_36213,N_31207,N_31770);
nor U36214 (N_36214,N_31344,N_32977);
nand U36215 (N_36215,N_31394,N_33300);
nor U36216 (N_36216,N_34636,N_31616);
or U36217 (N_36217,N_34626,N_34614);
and U36218 (N_36218,N_30155,N_33059);
nor U36219 (N_36219,N_32448,N_33845);
nand U36220 (N_36220,N_31578,N_30974);
or U36221 (N_36221,N_34553,N_30412);
and U36222 (N_36222,N_34624,N_33814);
nand U36223 (N_36223,N_32528,N_33505);
or U36224 (N_36224,N_31639,N_32126);
or U36225 (N_36225,N_32791,N_34193);
or U36226 (N_36226,N_30081,N_34278);
and U36227 (N_36227,N_31077,N_30253);
nand U36228 (N_36228,N_31051,N_33141);
nand U36229 (N_36229,N_33284,N_30166);
nand U36230 (N_36230,N_34516,N_33727);
or U36231 (N_36231,N_33119,N_34003);
nand U36232 (N_36232,N_30915,N_31635);
nand U36233 (N_36233,N_33103,N_30418);
or U36234 (N_36234,N_30142,N_32049);
nor U36235 (N_36235,N_30847,N_32434);
or U36236 (N_36236,N_32325,N_31433);
nand U36237 (N_36237,N_34693,N_32534);
and U36238 (N_36238,N_30446,N_30779);
or U36239 (N_36239,N_31684,N_33643);
nor U36240 (N_36240,N_32905,N_30907);
nand U36241 (N_36241,N_33909,N_34421);
xor U36242 (N_36242,N_31628,N_32300);
xnor U36243 (N_36243,N_32655,N_32466);
nor U36244 (N_36244,N_34796,N_32113);
nand U36245 (N_36245,N_31622,N_33795);
or U36246 (N_36246,N_30694,N_33860);
and U36247 (N_36247,N_31318,N_33306);
or U36248 (N_36248,N_30647,N_30321);
and U36249 (N_36249,N_30954,N_32515);
and U36250 (N_36250,N_31942,N_30037);
and U36251 (N_36251,N_34305,N_32152);
or U36252 (N_36252,N_30219,N_33829);
or U36253 (N_36253,N_33478,N_34809);
or U36254 (N_36254,N_31177,N_32324);
nor U36255 (N_36255,N_34338,N_33942);
or U36256 (N_36256,N_33303,N_31796);
and U36257 (N_36257,N_31927,N_30982);
nor U36258 (N_36258,N_34314,N_30080);
and U36259 (N_36259,N_31706,N_30615);
nor U36260 (N_36260,N_31748,N_32023);
and U36261 (N_36261,N_30774,N_34433);
xnor U36262 (N_36262,N_33196,N_33666);
nand U36263 (N_36263,N_31582,N_32333);
nand U36264 (N_36264,N_33490,N_34613);
nor U36265 (N_36265,N_34696,N_31571);
or U36266 (N_36266,N_30397,N_32658);
or U36267 (N_36267,N_32524,N_31511);
nor U36268 (N_36268,N_34454,N_31295);
and U36269 (N_36269,N_34123,N_34952);
xnor U36270 (N_36270,N_33741,N_33210);
nand U36271 (N_36271,N_33763,N_34432);
or U36272 (N_36272,N_32334,N_32516);
nand U36273 (N_36273,N_33384,N_31850);
nor U36274 (N_36274,N_32901,N_32543);
xor U36275 (N_36275,N_30042,N_32330);
xor U36276 (N_36276,N_34755,N_30962);
and U36277 (N_36277,N_31939,N_31485);
and U36278 (N_36278,N_30120,N_31030);
xor U36279 (N_36279,N_34397,N_34840);
xor U36280 (N_36280,N_31230,N_33314);
or U36281 (N_36281,N_34225,N_32117);
or U36282 (N_36282,N_31961,N_30182);
xor U36283 (N_36283,N_30281,N_34872);
or U36284 (N_36284,N_34519,N_32086);
nand U36285 (N_36285,N_33233,N_34501);
nor U36286 (N_36286,N_33259,N_33406);
nand U36287 (N_36287,N_34013,N_32459);
or U36288 (N_36288,N_34656,N_33399);
xor U36289 (N_36289,N_32919,N_30292);
and U36290 (N_36290,N_32055,N_32226);
nor U36291 (N_36291,N_31043,N_30478);
xnor U36292 (N_36292,N_31059,N_32154);
nor U36293 (N_36293,N_30986,N_31946);
nand U36294 (N_36294,N_31420,N_31266);
xor U36295 (N_36295,N_34182,N_33324);
and U36296 (N_36296,N_32944,N_31633);
nand U36297 (N_36297,N_30280,N_34173);
and U36298 (N_36298,N_33535,N_34133);
and U36299 (N_36299,N_34515,N_31092);
or U36300 (N_36300,N_30930,N_33441);
xor U36301 (N_36301,N_31335,N_34189);
and U36302 (N_36302,N_30000,N_33756);
xnor U36303 (N_36303,N_31494,N_30342);
nand U36304 (N_36304,N_33180,N_34607);
nor U36305 (N_36305,N_32376,N_30780);
or U36306 (N_36306,N_33270,N_30874);
xnor U36307 (N_36307,N_31497,N_34780);
or U36308 (N_36308,N_34469,N_34298);
nand U36309 (N_36309,N_30244,N_32756);
nand U36310 (N_36310,N_32984,N_33249);
and U36311 (N_36311,N_31912,N_33293);
and U36312 (N_36312,N_34062,N_31675);
nand U36313 (N_36313,N_33524,N_30610);
xor U36314 (N_36314,N_30473,N_32303);
nand U36315 (N_36315,N_33850,N_34822);
nand U36316 (N_36316,N_30807,N_34994);
nor U36317 (N_36317,N_33341,N_34047);
nand U36318 (N_36318,N_30096,N_31525);
xnor U36319 (N_36319,N_32294,N_30839);
or U36320 (N_36320,N_30640,N_30791);
and U36321 (N_36321,N_30895,N_32750);
or U36322 (N_36322,N_31503,N_33534);
nand U36323 (N_36323,N_30213,N_31891);
nor U36324 (N_36324,N_31196,N_31827);
nor U36325 (N_36325,N_30157,N_31058);
nand U36326 (N_36326,N_32935,N_32114);
nor U36327 (N_36327,N_30593,N_33248);
or U36328 (N_36328,N_33279,N_33134);
nand U36329 (N_36329,N_30489,N_30829);
nor U36330 (N_36330,N_32691,N_30993);
or U36331 (N_36331,N_33126,N_32421);
and U36332 (N_36332,N_31444,N_32281);
nand U36333 (N_36333,N_30352,N_33235);
or U36334 (N_36334,N_34786,N_33382);
nor U36335 (N_36335,N_32344,N_31718);
and U36336 (N_36336,N_33319,N_34738);
xor U36337 (N_36337,N_33758,N_34776);
and U36338 (N_36338,N_33975,N_33429);
and U36339 (N_36339,N_34154,N_31789);
nand U36340 (N_36340,N_33021,N_34285);
or U36341 (N_36341,N_33715,N_30599);
and U36342 (N_36342,N_34196,N_32403);
nor U36343 (N_36343,N_32374,N_34967);
xor U36344 (N_36344,N_31421,N_34170);
or U36345 (N_36345,N_32852,N_31771);
xor U36346 (N_36346,N_30965,N_33074);
or U36347 (N_36347,N_33045,N_33578);
and U36348 (N_36348,N_34828,N_32278);
or U36349 (N_36349,N_30377,N_30308);
nand U36350 (N_36350,N_30928,N_31367);
nor U36351 (N_36351,N_34002,N_31808);
or U36352 (N_36352,N_30426,N_34814);
nor U36353 (N_36353,N_33424,N_34317);
nor U36354 (N_36354,N_31445,N_30204);
nor U36355 (N_36355,N_30115,N_32488);
xor U36356 (N_36356,N_34178,N_34413);
or U36357 (N_36357,N_33357,N_33056);
nand U36358 (N_36358,N_34423,N_31793);
xor U36359 (N_36359,N_30381,N_31710);
xor U36360 (N_36360,N_32800,N_32082);
or U36361 (N_36361,N_30327,N_34406);
nand U36362 (N_36362,N_34681,N_32116);
nor U36363 (N_36363,N_32096,N_33849);
and U36364 (N_36364,N_31950,N_32506);
and U36365 (N_36365,N_33132,N_32224);
nor U36366 (N_36366,N_33375,N_34215);
xnor U36367 (N_36367,N_32489,N_31828);
xor U36368 (N_36368,N_31166,N_32605);
nor U36369 (N_36369,N_30141,N_34655);
or U36370 (N_36370,N_32423,N_33541);
and U36371 (N_36371,N_32289,N_34084);
nor U36372 (N_36372,N_30680,N_33966);
nand U36373 (N_36373,N_31298,N_30357);
or U36374 (N_36374,N_34390,N_34532);
nand U36375 (N_36375,N_34508,N_33896);
xor U36376 (N_36376,N_34070,N_30717);
or U36377 (N_36377,N_33431,N_34445);
or U36378 (N_36378,N_33637,N_30742);
and U36379 (N_36379,N_31274,N_32807);
and U36380 (N_36380,N_34673,N_32981);
and U36381 (N_36381,N_32194,N_31604);
and U36382 (N_36382,N_32559,N_31520);
xnor U36383 (N_36383,N_31095,N_34672);
or U36384 (N_36384,N_31144,N_31056);
and U36385 (N_36385,N_32627,N_30016);
and U36386 (N_36386,N_30886,N_31004);
nor U36387 (N_36387,N_33840,N_33182);
and U36388 (N_36388,N_30804,N_34160);
nand U36389 (N_36389,N_30247,N_33564);
or U36390 (N_36390,N_30621,N_33513);
nor U36391 (N_36391,N_32819,N_32299);
nand U36392 (N_36392,N_33570,N_31119);
or U36393 (N_36393,N_31269,N_31007);
nor U36394 (N_36394,N_32391,N_34227);
and U36395 (N_36395,N_33638,N_32047);
xor U36396 (N_36396,N_33678,N_32880);
nand U36397 (N_36397,N_30872,N_34143);
nand U36398 (N_36398,N_32263,N_31820);
nor U36399 (N_36399,N_31984,N_30503);
or U36400 (N_36400,N_34964,N_30180);
or U36401 (N_36401,N_31192,N_32993);
nor U36402 (N_36402,N_30916,N_32551);
nor U36403 (N_36403,N_31587,N_30191);
xor U36404 (N_36404,N_32132,N_33631);
nand U36405 (N_36405,N_34561,N_31583);
and U36406 (N_36406,N_34534,N_33507);
or U36407 (N_36407,N_32409,N_33787);
and U36408 (N_36408,N_31669,N_32940);
xor U36409 (N_36409,N_30097,N_32550);
and U36410 (N_36410,N_31105,N_31074);
xnor U36411 (N_36411,N_31225,N_32641);
or U36412 (N_36412,N_33739,N_31215);
nor U36413 (N_36413,N_33897,N_31877);
and U36414 (N_36414,N_31887,N_33624);
and U36415 (N_36415,N_31121,N_34851);
xnor U36416 (N_36416,N_30251,N_33855);
xor U36417 (N_36417,N_33552,N_34309);
or U36418 (N_36418,N_30044,N_34981);
nand U36419 (N_36419,N_34919,N_30903);
nor U36420 (N_36420,N_32002,N_33446);
xor U36421 (N_36421,N_33796,N_33482);
nor U36422 (N_36422,N_31454,N_34366);
or U36423 (N_36423,N_31120,N_31037);
nand U36424 (N_36424,N_31139,N_31581);
nand U36425 (N_36425,N_30409,N_31181);
nor U36426 (N_36426,N_30278,N_32547);
or U36427 (N_36427,N_33493,N_33536);
nor U36428 (N_36428,N_30260,N_34313);
nor U36429 (N_36429,N_31989,N_34579);
nand U36430 (N_36430,N_31327,N_34001);
nor U36431 (N_36431,N_32111,N_33544);
nor U36432 (N_36432,N_34069,N_34572);
nand U36433 (N_36433,N_30200,N_32714);
xor U36434 (N_36434,N_34605,N_32302);
and U36435 (N_36435,N_33494,N_30216);
and U36436 (N_36436,N_34386,N_30575);
xor U36437 (N_36437,N_31448,N_30578);
and U36438 (N_36438,N_30333,N_32036);
nand U36439 (N_36439,N_34916,N_31799);
or U36440 (N_36440,N_30501,N_33105);
nor U36441 (N_36441,N_31089,N_34567);
or U36442 (N_36442,N_32306,N_32613);
xnor U36443 (N_36443,N_33315,N_30857);
xor U36444 (N_36444,N_32882,N_31592);
and U36445 (N_36445,N_34365,N_31529);
xnor U36446 (N_36446,N_34181,N_31654);
nand U36447 (N_36447,N_30724,N_31090);
nor U36448 (N_36448,N_33556,N_31262);
xnor U36449 (N_36449,N_30521,N_32139);
nor U36450 (N_36450,N_31244,N_32584);
nor U36451 (N_36451,N_33350,N_32811);
xnor U36452 (N_36452,N_33686,N_31453);
and U36453 (N_36453,N_34986,N_34648);
xor U36454 (N_36454,N_30695,N_33136);
nor U36455 (N_36455,N_31104,N_32779);
nor U36456 (N_36456,N_33014,N_33150);
or U36457 (N_36457,N_33997,N_31769);
nand U36458 (N_36458,N_31885,N_32581);
nand U36459 (N_36459,N_34230,N_34689);
nand U36460 (N_36460,N_32216,N_33706);
nand U36461 (N_36461,N_34627,N_32616);
xnor U36462 (N_36462,N_33070,N_30275);
nand U36463 (N_36463,N_31024,N_32520);
xor U36464 (N_36464,N_31548,N_30314);
nand U36465 (N_36465,N_31781,N_30606);
nor U36466 (N_36466,N_34393,N_31201);
nand U36467 (N_36467,N_34958,N_33805);
nand U36468 (N_36468,N_32243,N_30531);
nand U36469 (N_36469,N_30464,N_33889);
nand U36470 (N_36470,N_31336,N_30402);
and U36471 (N_36471,N_33483,N_33729);
or U36472 (N_36472,N_30164,N_30735);
nand U36473 (N_36473,N_30248,N_32699);
xnor U36474 (N_36474,N_34176,N_33537);
xnor U36475 (N_36475,N_30775,N_33698);
nor U36476 (N_36476,N_33523,N_32792);
and U36477 (N_36477,N_31311,N_33081);
xor U36478 (N_36478,N_30967,N_33062);
nor U36479 (N_36479,N_30763,N_33342);
nor U36480 (N_36480,N_34025,N_31171);
xor U36481 (N_36481,N_33465,N_32822);
or U36482 (N_36482,N_30859,N_33642);
nand U36483 (N_36483,N_31082,N_34905);
nor U36484 (N_36484,N_31816,N_32385);
xnor U36485 (N_36485,N_30462,N_34972);
and U36486 (N_36486,N_31656,N_33392);
nand U36487 (N_36487,N_30477,N_34348);
and U36488 (N_36488,N_31634,N_34023);
nand U36489 (N_36489,N_34343,N_30351);
nor U36490 (N_36490,N_33388,N_31143);
nand U36491 (N_36491,N_31713,N_34392);
nand U36492 (N_36492,N_31873,N_33603);
xor U36493 (N_36493,N_32438,N_33740);
and U36494 (N_36494,N_32754,N_30602);
xor U36495 (N_36495,N_30678,N_33522);
xor U36496 (N_36496,N_34483,N_33189);
and U36497 (N_36497,N_31988,N_33893);
or U36498 (N_36498,N_30088,N_33011);
xnor U36499 (N_36499,N_34441,N_30972);
xor U36500 (N_36500,N_33006,N_34725);
and U36501 (N_36501,N_30509,N_32019);
or U36502 (N_36502,N_30190,N_34007);
nand U36503 (N_36503,N_31909,N_32843);
and U36504 (N_36504,N_34044,N_33863);
xnor U36505 (N_36505,N_30726,N_33717);
and U36506 (N_36506,N_33569,N_31965);
nand U36507 (N_36507,N_33305,N_31324);
nor U36508 (N_36508,N_32030,N_32387);
nor U36509 (N_36509,N_34399,N_34440);
and U36510 (N_36510,N_32930,N_30053);
nor U36511 (N_36511,N_33423,N_34267);
nor U36512 (N_36512,N_31118,N_31610);
xnor U36513 (N_36513,N_30656,N_30497);
or U36514 (N_36514,N_34232,N_32730);
xnor U36515 (N_36515,N_30545,N_31566);
and U36516 (N_36516,N_32098,N_30787);
and U36517 (N_36517,N_32987,N_32614);
nand U36518 (N_36518,N_33962,N_33980);
nor U36519 (N_36519,N_34447,N_30754);
nor U36520 (N_36520,N_31968,N_33177);
or U36521 (N_36521,N_30086,N_32571);
or U36522 (N_36522,N_31835,N_31265);
and U36523 (N_36523,N_31632,N_30722);
nand U36524 (N_36524,N_30095,N_33662);
or U36525 (N_36525,N_34628,N_31101);
nand U36526 (N_36526,N_32979,N_34767);
xnor U36527 (N_36527,N_30711,N_30795);
nor U36528 (N_36528,N_31169,N_34147);
xor U36529 (N_36529,N_31436,N_34733);
nor U36530 (N_36530,N_30884,N_32451);
nor U36531 (N_36531,N_31512,N_34793);
or U36532 (N_36532,N_34573,N_33865);
nand U36533 (N_36533,N_31970,N_30515);
xor U36534 (N_36534,N_33514,N_30056);
nand U36535 (N_36535,N_32428,N_34359);
and U36536 (N_36536,N_30562,N_32436);
or U36537 (N_36537,N_32388,N_34322);
xor U36538 (N_36538,N_34646,N_34235);
or U36539 (N_36539,N_33500,N_34205);
and U36540 (N_36540,N_32203,N_34398);
or U36541 (N_36541,N_32060,N_31340);
nor U36542 (N_36542,N_34583,N_30079);
and U36543 (N_36543,N_33055,N_34287);
or U36544 (N_36544,N_33336,N_32912);
and U36545 (N_36545,N_31374,N_34207);
xor U36546 (N_36546,N_30400,N_32713);
xnor U36547 (N_36547,N_31018,N_34890);
and U36548 (N_36548,N_30431,N_34021);
or U36549 (N_36549,N_30888,N_32437);
nor U36550 (N_36550,N_34955,N_33457);
nand U36551 (N_36551,N_30753,N_30576);
xnor U36552 (N_36552,N_31026,N_32183);
and U36553 (N_36553,N_30703,N_31697);
and U36554 (N_36554,N_31202,N_33905);
and U36555 (N_36555,N_31979,N_33242);
and U36556 (N_36556,N_32854,N_30099);
nor U36557 (N_36557,N_30178,N_31958);
or U36558 (N_36558,N_31774,N_30929);
or U36559 (N_36559,N_34159,N_31671);
nor U36560 (N_36560,N_30017,N_30152);
nand U36561 (N_36561,N_34119,N_32556);
or U36562 (N_36562,N_33732,N_33426);
nor U36563 (N_36563,N_34150,N_34576);
or U36564 (N_36564,N_34148,N_34525);
nor U36565 (N_36565,N_31689,N_34611);
or U36566 (N_36566,N_32204,N_34274);
xnor U36567 (N_36567,N_34520,N_30460);
and U36568 (N_36568,N_30344,N_32731);
nor U36569 (N_36569,N_31049,N_34526);
xnor U36570 (N_36570,N_32778,N_33263);
xnor U36571 (N_36571,N_32457,N_31572);
xnor U36572 (N_36572,N_32773,N_34939);
and U36573 (N_36573,N_31188,N_33212);
nor U36574 (N_36574,N_31239,N_33130);
nor U36575 (N_36575,N_34712,N_30506);
or U36576 (N_36576,N_30495,N_32932);
nand U36577 (N_36577,N_30372,N_30637);
or U36578 (N_36578,N_30045,N_34018);
and U36579 (N_36579,N_30101,N_31831);
or U36580 (N_36580,N_33260,N_34381);
xnor U36581 (N_36581,N_30547,N_34361);
or U36582 (N_36582,N_32685,N_34660);
and U36583 (N_36583,N_34819,N_34979);
or U36584 (N_36584,N_34111,N_33326);
xor U36585 (N_36585,N_30650,N_31084);
xnor U36586 (N_36586,N_32191,N_33605);
and U36587 (N_36587,N_32231,N_31897);
and U36588 (N_36588,N_31591,N_34191);
xnor U36589 (N_36589,N_31377,N_31858);
nor U36590 (N_36590,N_31779,N_31235);
or U36591 (N_36591,N_30789,N_32871);
nand U36592 (N_36592,N_33994,N_34035);
nor U36593 (N_36593,N_30673,N_30677);
nand U36594 (N_36594,N_32884,N_32107);
xor U36595 (N_36595,N_30852,N_31735);
and U36596 (N_36596,N_34988,N_30643);
nand U36597 (N_36597,N_32280,N_30727);
nand U36598 (N_36598,N_32368,N_32539);
nand U36599 (N_36599,N_31728,N_32532);
nand U36600 (N_36600,N_31844,N_32080);
or U36601 (N_36601,N_32916,N_31999);
or U36602 (N_36602,N_31890,N_31492);
xnor U36603 (N_36603,N_34717,N_31502);
or U36604 (N_36604,N_32369,N_31953);
nand U36605 (N_36605,N_31242,N_33716);
xnor U36606 (N_36606,N_33502,N_34494);
xor U36607 (N_36607,N_33526,N_32647);
xor U36608 (N_36608,N_30008,N_34835);
nand U36609 (N_36609,N_34286,N_31140);
or U36610 (N_36610,N_31867,N_33253);
and U36611 (N_36611,N_33979,N_31048);
and U36612 (N_36612,N_30921,N_31001);
and U36613 (N_36613,N_30758,N_30136);
or U36614 (N_36614,N_31115,N_33140);
or U36615 (N_36615,N_32780,N_30701);
xor U36616 (N_36616,N_30746,N_32361);
nor U36617 (N_36617,N_30751,N_31328);
and U36618 (N_36618,N_33280,N_32885);
nor U36619 (N_36619,N_33208,N_33917);
or U36620 (N_36620,N_33418,N_30245);
nand U36621 (N_36621,N_33374,N_34868);
nor U36622 (N_36622,N_32562,N_33462);
nand U36623 (N_36623,N_30149,N_32311);
nor U36624 (N_36624,N_34071,N_31794);
nor U36625 (N_36625,N_30188,N_32040);
and U36626 (N_36626,N_30546,N_30900);
xor U36627 (N_36627,N_34072,N_34342);
xnor U36628 (N_36628,N_34929,N_33676);
nand U36629 (N_36629,N_34089,N_34270);
and U36630 (N_36630,N_31431,N_32937);
and U36631 (N_36631,N_32866,N_34927);
nand U36632 (N_36632,N_31296,N_32417);
or U36633 (N_36633,N_34139,N_34116);
nor U36634 (N_36634,N_31811,N_33856);
or U36635 (N_36635,N_33017,N_34355);
and U36636 (N_36636,N_32693,N_31807);
or U36637 (N_36637,N_32651,N_30574);
nor U36638 (N_36638,N_31696,N_33296);
or U36639 (N_36639,N_30639,N_32108);
and U36640 (N_36640,N_30814,N_33459);
xnor U36641 (N_36641,N_33846,N_32262);
nand U36642 (N_36642,N_31992,N_32624);
and U36643 (N_36643,N_33147,N_31334);
nor U36644 (N_36644,N_31270,N_32672);
xor U36645 (N_36645,N_33251,N_34802);
and U36646 (N_36646,N_31925,N_31937);
nand U36647 (N_36647,N_30326,N_30105);
and U36648 (N_36648,N_30369,N_30361);
nand U36649 (N_36649,N_32446,N_32938);
or U36650 (N_36650,N_33930,N_33163);
nand U36651 (N_36651,N_34810,N_34363);
nand U36652 (N_36652,N_30682,N_33133);
nor U36653 (N_36653,N_31285,N_30020);
and U36654 (N_36654,N_32631,N_30311);
nand U36655 (N_36655,N_32101,N_34861);
nor U36656 (N_36656,N_33824,N_33230);
nand U36657 (N_36657,N_33976,N_34495);
xor U36658 (N_36658,N_34260,N_33591);
nor U36659 (N_36659,N_30359,N_30138);
or U36660 (N_36660,N_30893,N_31597);
and U36661 (N_36661,N_31649,N_32090);
and U36662 (N_36662,N_33703,N_31396);
xnor U36663 (N_36663,N_34263,N_31355);
xnor U36664 (N_36664,N_31480,N_32282);
nand U36665 (N_36665,N_31914,N_33264);
nor U36666 (N_36666,N_34601,N_32521);
nor U36667 (N_36667,N_33211,N_34351);
xnor U36668 (N_36668,N_32948,N_33369);
nand U36669 (N_36669,N_34845,N_30793);
or U36670 (N_36670,N_31500,N_34876);
xor U36671 (N_36671,N_32523,N_33590);
nand U36672 (N_36672,N_30111,N_31538);
and U36673 (N_36673,N_34172,N_31855);
nand U36674 (N_36674,N_34651,N_31755);
xor U36675 (N_36675,N_31983,N_30797);
and U36676 (N_36676,N_33778,N_34545);
and U36677 (N_36677,N_32728,N_30765);
xor U36678 (N_36678,N_33599,N_33600);
or U36679 (N_36679,N_32727,N_30156);
or U36680 (N_36680,N_34910,N_33589);
nor U36681 (N_36681,N_31210,N_33485);
and U36682 (N_36682,N_32593,N_30060);
or U36683 (N_36683,N_31477,N_30366);
xnor U36684 (N_36684,N_31588,N_30534);
or U36685 (N_36685,N_31917,N_31238);
nor U36686 (N_36686,N_32761,N_30239);
or U36687 (N_36687,N_32677,N_32794);
nand U36688 (N_36688,N_33102,N_33641);
nand U36689 (N_36689,N_30181,N_32291);
and U36690 (N_36690,N_32085,N_32129);
and U36691 (N_36691,N_34528,N_32615);
xor U36692 (N_36692,N_30617,N_32317);
xor U36693 (N_36693,N_33830,N_34920);
nor U36694 (N_36694,N_32377,N_34497);
or U36695 (N_36695,N_30514,N_31717);
nand U36696 (N_36696,N_30567,N_33983);
nand U36697 (N_36697,N_33610,N_33707);
or U36698 (N_36698,N_34869,N_31356);
or U36699 (N_36699,N_31000,N_30150);
xor U36700 (N_36700,N_30662,N_32525);
xor U36701 (N_36701,N_30496,N_32620);
xor U36702 (N_36702,N_34850,N_31904);
nor U36703 (N_36703,N_34640,N_34938);
nand U36704 (N_36704,N_30214,N_30948);
nor U36705 (N_36705,N_31849,N_31423);
and U36706 (N_36706,N_31629,N_34037);
and U36707 (N_36707,N_31205,N_30683);
or U36708 (N_36708,N_33511,N_33371);
or U36709 (N_36709,N_31948,N_32970);
xor U36710 (N_36710,N_34737,N_31081);
nor U36711 (N_36711,N_30104,N_30335);
or U36712 (N_36712,N_32201,N_31854);
nor U36713 (N_36713,N_30541,N_34201);
or U36714 (N_36714,N_31346,N_34459);
xnor U36715 (N_36715,N_30597,N_32812);
and U36716 (N_36716,N_32622,N_34736);
nand U36717 (N_36717,N_32734,N_30403);
and U36718 (N_36718,N_33911,N_34272);
or U36719 (N_36719,N_31664,N_34279);
nand U36720 (N_36720,N_30266,N_34996);
xnor U36721 (N_36721,N_30461,N_33629);
nand U36722 (N_36722,N_32486,N_31228);
nand U36723 (N_36723,N_33402,N_30601);
nor U36724 (N_36724,N_32511,N_31834);
xnor U36725 (N_36725,N_34318,N_30234);
and U36726 (N_36726,N_33540,N_32358);
nand U36727 (N_36727,N_32378,N_32513);
and U36728 (N_36728,N_34971,N_33127);
and U36729 (N_36729,N_33539,N_34241);
and U36730 (N_36730,N_33577,N_34675);
nor U36731 (N_36731,N_32659,N_32540);
nor U36732 (N_36732,N_32599,N_30979);
xnor U36733 (N_36733,N_30654,N_32902);
nor U36734 (N_36734,N_30463,N_31041);
nor U36735 (N_36735,N_34637,N_34218);
nand U36736 (N_36736,N_33086,N_31046);
xor U36737 (N_36737,N_31341,N_33553);
nor U36738 (N_36738,N_30738,N_30283);
and U36739 (N_36739,N_34301,N_34485);
nand U36740 (N_36740,N_34198,N_31918);
nand U36741 (N_36741,N_32757,N_31732);
and U36742 (N_36742,N_34730,N_31737);
or U36743 (N_36743,N_33596,N_32850);
nand U36744 (N_36744,N_33360,N_30913);
nor U36745 (N_36745,N_32642,N_33033);
xor U36746 (N_36746,N_32471,N_31488);
xnor U36747 (N_36747,N_32851,N_33745);
xnor U36748 (N_36748,N_33504,N_30230);
xor U36749 (N_36749,N_31331,N_33330);
nor U36750 (N_36750,N_34212,N_34336);
xor U36751 (N_36751,N_34726,N_34104);
and U36752 (N_36752,N_33616,N_34231);
xor U36753 (N_36753,N_30472,N_33772);
nor U36754 (N_36754,N_33420,N_30391);
and U36755 (N_36755,N_33197,N_31102);
nor U36756 (N_36756,N_30938,N_33408);
and U36757 (N_36757,N_33329,N_34829);
nand U36758 (N_36758,N_31158,N_31358);
xnor U36759 (N_36759,N_30475,N_33110);
xnor U36760 (N_36760,N_31627,N_34510);
or U36761 (N_36761,N_33229,N_31428);
and U36762 (N_36762,N_33477,N_30533);
or U36763 (N_36763,N_33835,N_34524);
nor U36764 (N_36764,N_32563,N_32212);
nand U36765 (N_36765,N_33008,N_33762);
xor U36766 (N_36766,N_32630,N_33902);
xor U36767 (N_36767,N_33286,N_31240);
xnor U36768 (N_36768,N_34621,N_34467);
nand U36769 (N_36769,N_31072,N_30254);
nand U36770 (N_36770,N_32634,N_30374);
nand U36771 (N_36771,N_31969,N_31701);
xnor U36772 (N_36772,N_32517,N_34055);
xor U36773 (N_36773,N_33456,N_34112);
nor U36774 (N_36774,N_33290,N_34024);
or U36775 (N_36775,N_34008,N_31952);
nand U36776 (N_36776,N_34578,N_34787);
and U36777 (N_36777,N_33978,N_30071);
or U36778 (N_36778,N_30885,N_33464);
nand U36779 (N_36779,N_34667,N_31128);
nor U36780 (N_36780,N_34566,N_32236);
and U36781 (N_36781,N_33618,N_30255);
or U36782 (N_36782,N_33720,N_33904);
and U36783 (N_36783,N_30162,N_33352);
and U36784 (N_36784,N_33178,N_31463);
and U36785 (N_36785,N_30367,N_33945);
nor U36786 (N_36786,N_30555,N_33238);
xnor U36787 (N_36787,N_31307,N_34941);
and U36788 (N_36788,N_34185,N_30508);
and U36789 (N_36789,N_32349,N_31227);
nor U36790 (N_36790,N_30339,N_31534);
xor U36791 (N_36791,N_34166,N_30140);
nor U36792 (N_36792,N_33302,N_31372);
xor U36793 (N_36793,N_32296,N_31562);
nor U36794 (N_36794,N_33949,N_33972);
xor U36795 (N_36795,N_34922,N_32124);
and U36796 (N_36796,N_33092,N_32774);
nor U36797 (N_36797,N_31528,N_32331);
nor U36798 (N_36798,N_30630,N_31944);
or U36799 (N_36799,N_30749,N_31666);
nand U36800 (N_36800,N_33528,N_33453);
nor U36801 (N_36801,N_31027,N_32147);
or U36802 (N_36802,N_34852,N_30179);
xnor U36803 (N_36803,N_34367,N_31775);
nand U36804 (N_36804,N_30334,N_34848);
xor U36805 (N_36805,N_31853,N_30596);
nor U36806 (N_36806,N_32723,N_31763);
xnor U36807 (N_36807,N_32664,N_32864);
or U36808 (N_36808,N_34394,N_33646);
xor U36809 (N_36809,N_34917,N_31819);
xor U36810 (N_36810,N_34724,N_31317);
nand U36811 (N_36811,N_30089,N_31504);
and U36812 (N_36812,N_34658,N_32083);
xnor U36813 (N_36813,N_33205,N_34347);
and U36814 (N_36814,N_34718,N_33234);
nor U36815 (N_36815,N_34011,N_34761);
nor U36816 (N_36816,N_33063,N_33521);
nor U36817 (N_36817,N_32907,N_33992);
or U36818 (N_36818,N_34239,N_32202);
or U36819 (N_36819,N_33498,N_31233);
nor U36820 (N_36820,N_34443,N_34255);
and U36821 (N_36821,N_32590,N_33277);
nand U36822 (N_36822,N_31973,N_30498);
or U36823 (N_36823,N_34192,N_34823);
nor U36824 (N_36824,N_30416,N_32996);
or U36825 (N_36825,N_32842,N_32234);
xnor U36826 (N_36826,N_31913,N_34067);
nor U36827 (N_36827,N_33510,N_33575);
xor U36828 (N_36828,N_30502,N_33934);
xor U36829 (N_36829,N_33415,N_32897);
and U36830 (N_36830,N_34356,N_34686);
xnor U36831 (N_36831,N_31221,N_33373);
nor U36832 (N_36832,N_31733,N_34107);
nor U36833 (N_36833,N_33836,N_32999);
nand U36834 (N_36834,N_31987,N_33775);
nand U36835 (N_36835,N_34863,N_31527);
and U36836 (N_36836,N_30523,N_33700);
xnor U36837 (N_36837,N_33173,N_31343);
xnor U36838 (N_36838,N_34391,N_34319);
nand U36839 (N_36839,N_34203,N_34608);
nand U36840 (N_36840,N_34887,N_32481);
and U36841 (N_36841,N_32392,N_32827);
nor U36842 (N_36842,N_30305,N_33563);
nor U36843 (N_36843,N_31016,N_34800);
nor U36844 (N_36844,N_31409,N_30744);
nand U36845 (N_36845,N_30343,N_33433);
or U36846 (N_36846,N_34284,N_33058);
xor U36847 (N_36847,N_30331,N_33818);
xnor U36848 (N_36848,N_34380,N_30238);
nand U36849 (N_36849,N_31682,N_32682);
nor U36850 (N_36850,N_31412,N_34949);
nand U36851 (N_36851,N_30709,N_31509);
xnor U36852 (N_36852,N_33542,N_33054);
or U36853 (N_36853,N_31348,N_34115);
and U36854 (N_36854,N_34881,N_32568);
or U36855 (N_36855,N_32922,N_32828);
or U36856 (N_36856,N_31363,N_33770);
and U36857 (N_36857,N_33984,N_31042);
and U36858 (N_36858,N_34431,N_30892);
or U36859 (N_36859,N_31407,N_31734);
nand U36860 (N_36860,N_34597,N_30007);
and U36861 (N_36861,N_32093,N_33274);
and U36862 (N_36862,N_34542,N_30125);
nand U36863 (N_36863,N_34200,N_32482);
xor U36864 (N_36864,N_31676,N_30941);
nand U36865 (N_36865,N_31114,N_32544);
nand U36866 (N_36866,N_34504,N_30386);
and U36867 (N_36867,N_32644,N_32618);
nand U36868 (N_36868,N_30471,N_33379);
nand U36869 (N_36869,N_30499,N_32418);
and U36870 (N_36870,N_33892,N_31549);
xnor U36871 (N_36871,N_32454,N_32923);
nand U36872 (N_36872,N_34963,N_32546);
nor U36873 (N_36873,N_32799,N_33435);
xnor U36874 (N_36874,N_32573,N_30126);
nand U36875 (N_36875,N_33155,N_33469);
xnor U36876 (N_36876,N_30679,N_33967);
nand U36877 (N_36877,N_31673,N_34711);
nand U36878 (N_36878,N_33803,N_34616);
nand U36879 (N_36879,N_33634,N_30171);
and U36880 (N_36880,N_32027,N_30513);
or U36881 (N_36881,N_33923,N_32678);
or U36882 (N_36882,N_33273,N_32976);
nor U36883 (N_36883,N_33292,N_33947);
or U36884 (N_36884,N_32992,N_34599);
xor U36885 (N_36885,N_33912,N_33777);
nand U36886 (N_36886,N_31870,N_31070);
and U36887 (N_36887,N_34934,N_30635);
xor U36888 (N_36888,N_31778,N_33395);
or U36889 (N_36889,N_30505,N_33002);
nor U36890 (N_36890,N_32164,N_30405);
or U36891 (N_36891,N_34438,N_32041);
xnor U36892 (N_36892,N_33076,N_32596);
nand U36893 (N_36893,N_33985,N_30906);
nand U36894 (N_36894,N_30856,N_34880);
xnor U36895 (N_36895,N_34444,N_30215);
xnor U36896 (N_36896,N_30671,N_32632);
nor U36897 (N_36897,N_34808,N_32587);
and U36898 (N_36898,N_31193,N_32159);
nand U36899 (N_36899,N_34300,N_33797);
and U36900 (N_36900,N_33794,N_33473);
and U36901 (N_36901,N_30873,N_33097);
or U36902 (N_36902,N_30132,N_34818);
and U36903 (N_36903,N_33938,N_34862);
xnor U36904 (N_36904,N_33713,N_31872);
nor U36905 (N_36905,N_30348,N_32227);
and U36906 (N_36906,N_32784,N_33682);
nor U36907 (N_36907,N_31391,N_34832);
or U36908 (N_36908,N_31079,N_34702);
xnor U36909 (N_36909,N_34924,N_32069);
nor U36910 (N_36910,N_31323,N_33567);
and U36911 (N_36911,N_31234,N_32861);
nand U36912 (N_36912,N_33346,N_32910);
and U36913 (N_36913,N_31416,N_32742);
or U36914 (N_36914,N_31801,N_34078);
nor U36915 (N_36915,N_30295,N_33819);
nor U36916 (N_36916,N_34683,N_30304);
nand U36917 (N_36917,N_31721,N_30902);
or U36918 (N_36918,N_33411,N_34968);
xnor U36919 (N_36919,N_33529,N_33480);
nand U36920 (N_36920,N_30055,N_33584);
nor U36921 (N_36921,N_33404,N_30878);
or U36922 (N_36922,N_32836,N_31640);
nor U36923 (N_36923,N_33883,N_30713);
nand U36924 (N_36924,N_31563,N_30752);
nor U36925 (N_36925,N_33948,N_34592);
xnor U36926 (N_36926,N_32883,N_31798);
or U36927 (N_36927,N_30137,N_33001);
xnor U36928 (N_36928,N_34315,N_32102);
or U36929 (N_36929,N_31185,N_34978);
and U36930 (N_36930,N_32416,N_32100);
nor U36931 (N_36931,N_31156,N_30899);
nand U36932 (N_36932,N_33746,N_30282);
or U36933 (N_36933,N_33018,N_34577);
nand U36934 (N_36934,N_33594,N_30933);
and U36935 (N_36935,N_30924,N_30559);
and U36936 (N_36936,N_31276,N_30330);
or U36937 (N_36937,N_30580,N_30490);
and U36938 (N_36938,N_34016,N_32167);
nor U36939 (N_36939,N_30582,N_30655);
or U36940 (N_36940,N_33837,N_32898);
nor U36941 (N_36941,N_32008,N_31472);
or U36942 (N_36942,N_33851,N_34350);
or U36943 (N_36943,N_34282,N_33807);
nor U36944 (N_36944,N_33802,N_32045);
or U36945 (N_36945,N_31223,N_32251);
xor U36946 (N_36946,N_30206,N_30067);
and U36947 (N_36947,N_31962,N_34593);
xnor U36948 (N_36948,N_31129,N_30013);
or U36949 (N_36949,N_32769,N_33484);
or U36950 (N_36950,N_32579,N_33884);
nor U36951 (N_36951,N_31756,N_30665);
or U36952 (N_36952,N_30373,N_34984);
or U36953 (N_36953,N_33764,N_31439);
xnor U36954 (N_36954,N_32022,N_34921);
or U36955 (N_36955,N_31061,N_32425);
xor U36956 (N_36956,N_32097,N_32585);
xnor U36957 (N_36957,N_32048,N_31931);
nor U36958 (N_36958,N_30645,N_34995);
nand U36959 (N_36959,N_31802,N_31621);
and U36960 (N_36960,N_32735,N_34478);
nor U36961 (N_36961,N_32293,N_34902);
or U36962 (N_36962,N_34701,N_34746);
and U36963 (N_36963,N_33878,N_34096);
or U36964 (N_36964,N_30025,N_31134);
nand U36965 (N_36965,N_31731,N_32404);
and U36966 (N_36966,N_31446,N_31350);
or U36967 (N_36967,N_34323,N_34442);
nand U36968 (N_36968,N_34217,N_34937);
and U36969 (N_36969,N_31458,N_32588);
nand U36970 (N_36970,N_31455,N_33203);
nor U36971 (N_36971,N_34512,N_32382);
or U36972 (N_36972,N_33067,N_31076);
xor U36973 (N_36973,N_34353,N_34871);
or U36974 (N_36974,N_30987,N_34098);
and U36975 (N_36975,N_34487,N_31432);
nor U36976 (N_36976,N_31209,N_30050);
nor U36977 (N_36977,N_31515,N_34713);
xnor U36978 (N_36978,N_34405,N_33776);
and U36979 (N_36979,N_33852,N_32295);
nor U36980 (N_36980,N_30894,N_31498);
and U36981 (N_36981,N_33220,N_34032);
and U36982 (N_36982,N_32153,N_32844);
or U36983 (N_36983,N_33908,N_30975);
xnor U36984 (N_36984,N_33654,N_31860);
or U36985 (N_36985,N_33928,N_32110);
or U36986 (N_36986,N_30710,N_30960);
and U36987 (N_36987,N_30838,N_34928);
nor U36988 (N_36988,N_32468,N_32066);
nor U36989 (N_36989,N_33003,N_33927);
and U36990 (N_36990,N_32961,N_33391);
or U36991 (N_36991,N_34586,N_32649);
nor U36992 (N_36992,N_32176,N_32397);
xor U36993 (N_36993,N_33932,N_32487);
nand U36994 (N_36994,N_31766,N_32990);
nand U36995 (N_36995,N_30672,N_32891);
nor U36996 (N_36996,N_30653,N_34856);
xnor U36997 (N_36997,N_32081,N_31040);
or U36998 (N_36998,N_31034,N_31012);
xnor U36999 (N_36999,N_33137,N_30959);
nand U37000 (N_37000,N_32601,N_33649);
xnor U37001 (N_37001,N_30358,N_31352);
or U37002 (N_37002,N_32806,N_33728);
and U37003 (N_37003,N_34602,N_32061);
or U37004 (N_37004,N_32698,N_31273);
and U37005 (N_37005,N_30867,N_33168);
nor U37006 (N_37006,N_32165,N_32986);
and U37007 (N_37007,N_30387,N_34795);
nor U37008 (N_37008,N_31161,N_33960);
nor U37009 (N_37009,N_33445,N_31957);
and U37010 (N_37010,N_34619,N_34770);
or U37011 (N_37011,N_34898,N_32338);
nand U37012 (N_37012,N_33838,N_34015);
and U37013 (N_37013,N_32586,N_31085);
nand U37014 (N_37014,N_33970,N_32028);
xor U37015 (N_37015,N_30365,N_30830);
and U37016 (N_37016,N_30194,N_30813);
or U37017 (N_37017,N_32740,N_32138);
nand U37018 (N_37018,N_30768,N_34690);
or U37019 (N_37019,N_34785,N_31670);
xnor U37020 (N_37020,N_31526,N_33887);
xor U37021 (N_37021,N_30203,N_32157);
xor U37022 (N_37022,N_34091,N_33272);
nor U37023 (N_37023,N_31288,N_31028);
xor U37024 (N_37024,N_33879,N_31111);
or U37025 (N_37025,N_31922,N_34180);
nand U37026 (N_37026,N_31901,N_31650);
and U37027 (N_37027,N_33095,N_30210);
nor U37028 (N_37028,N_30413,N_31483);
nand U37029 (N_37029,N_30951,N_31709);
nand U37030 (N_37030,N_34896,N_32071);
xnor U37031 (N_37031,N_31646,N_30423);
and U37032 (N_37032,N_33065,N_33176);
xnor U37033 (N_37033,N_33748,N_32452);
or U37034 (N_37034,N_31691,N_34966);
nor U37035 (N_37035,N_32494,N_33096);
nand U37036 (N_37036,N_30853,N_30049);
nand U37037 (N_37037,N_33995,N_30947);
nand U37038 (N_37038,N_33016,N_32638);
nor U37039 (N_37039,N_34042,N_34635);
and U37040 (N_37040,N_31971,N_31544);
nand U37041 (N_37041,N_32136,N_30784);
or U37042 (N_37042,N_32168,N_33644);
nand U37043 (N_37043,N_34531,N_32855);
or U37044 (N_37044,N_34541,N_32876);
nand U37045 (N_37045,N_32988,N_30591);
nor U37046 (N_37046,N_33034,N_31103);
or U37047 (N_37047,N_32408,N_32313);
xnor U37048 (N_37048,N_31720,N_31184);
or U37049 (N_37049,N_34183,N_33744);
and U37050 (N_37050,N_31797,N_32127);
and U37051 (N_37051,N_33615,N_31594);
xor U37052 (N_37052,N_32688,N_34224);
nor U37053 (N_37053,N_30070,N_32701);
nor U37054 (N_37054,N_32196,N_30100);
or U37055 (N_37055,N_32574,N_30256);
nor U37056 (N_37056,N_32823,N_34029);
and U37057 (N_37057,N_30845,N_30451);
or U37058 (N_37058,N_33783,N_34175);
nor U37059 (N_37059,N_34135,N_30714);
nand U37060 (N_37060,N_34312,N_30487);
nand U37061 (N_37061,N_33085,N_32692);
nand U37062 (N_37062,N_32345,N_34762);
nor U37063 (N_37063,N_34536,N_33981);
and U37064 (N_37064,N_32308,N_34836);
or U37065 (N_37065,N_34482,N_33436);
or U37066 (N_37066,N_34246,N_32566);
xnor U37067 (N_37067,N_30098,N_34680);
xnor U37068 (N_37068,N_30184,N_31253);
nand U37069 (N_37069,N_33925,N_34010);
or U37070 (N_37070,N_33154,N_31474);
nand U37071 (N_37071,N_31725,N_34093);
nor U37072 (N_37072,N_30354,N_32175);
or U37073 (N_37073,N_33612,N_31313);
nor U37074 (N_37074,N_32469,N_31136);
or U37075 (N_37075,N_34781,N_31783);
and U37076 (N_37076,N_34410,N_30398);
or U37077 (N_37077,N_32499,N_33385);
nor U37078 (N_37078,N_32834,N_34956);
and U37079 (N_37079,N_31250,N_30033);
nand U37080 (N_37080,N_33143,N_31050);
or U37081 (N_37081,N_32007,N_32743);
nor U37082 (N_37082,N_31284,N_34732);
nor U37083 (N_37083,N_32862,N_31899);
xnor U37084 (N_37084,N_31945,N_31199);
xor U37085 (N_37085,N_31729,N_32619);
nor U37086 (N_37086,N_30756,N_34187);
nand U37087 (N_37087,N_31856,N_34715);
and U37088 (N_37088,N_31601,N_31982);
or U37089 (N_37089,N_31098,N_33669);
xor U37090 (N_37090,N_30467,N_31906);
nor U37091 (N_37091,N_34623,N_34388);
and U37092 (N_37092,N_30684,N_32473);
nor U37093 (N_37093,N_32244,N_33597);
nor U37094 (N_37094,N_34946,N_32697);
and U37095 (N_37095,N_31821,N_31637);
nor U37096 (N_37096,N_32564,N_31427);
or U37097 (N_37097,N_32128,N_33918);
xor U37098 (N_37098,N_33012,N_31888);
or U37099 (N_37099,N_32760,N_34209);
or U37100 (N_37100,N_34161,N_32835);
xnor U37101 (N_37101,N_31672,N_30912);
xnor U37102 (N_37102,N_34145,N_34177);
or U37103 (N_37103,N_30963,N_30319);
and U37104 (N_37104,N_31585,N_33383);
nand U37105 (N_37105,N_31935,N_30855);
xor U37106 (N_37106,N_33988,N_34488);
nand U37107 (N_37107,N_31299,N_32321);
nand U37108 (N_37108,N_31369,N_32472);
or U37109 (N_37109,N_30798,N_30202);
xnor U37110 (N_37110,N_31516,N_30059);
nand U37111 (N_37111,N_32858,N_31956);
xnor U37112 (N_37112,N_33183,N_34901);
xor U37113 (N_37113,N_30622,N_34866);
or U37114 (N_37114,N_30199,N_30923);
nor U37115 (N_37115,N_34058,N_33709);
nand U37116 (N_37116,N_31130,N_31719);
nand U37117 (N_37117,N_30420,N_33813);
and U37118 (N_37118,N_33354,N_33165);
xor U37119 (N_37119,N_31620,N_31932);
and U37120 (N_37120,N_31589,N_32220);
or U37121 (N_37121,N_31772,N_34339);
nor U37122 (N_37122,N_33518,N_32029);
or U37123 (N_37123,N_32808,N_34765);
and U37124 (N_37124,N_30092,N_33481);
nand U37125 (N_37125,N_34722,N_31289);
or U37126 (N_37126,N_30901,N_34975);
xor U37127 (N_37127,N_30908,N_32490);
xor U37128 (N_37128,N_34259,N_30719);
and U37129 (N_37129,N_31955,N_30614);
or U37130 (N_37130,N_30399,N_31310);
nand U37131 (N_37131,N_34595,N_32696);
xor U37132 (N_37132,N_34455,N_32545);
nor U37133 (N_37133,N_31681,N_34144);
nand U37134 (N_37134,N_33064,N_32206);
nand U37135 (N_37135,N_32462,N_34555);
and U37136 (N_37136,N_32260,N_33773);
nand U37137 (N_37137,N_32178,N_30736);
xor U37138 (N_37138,N_31200,N_31333);
or U37139 (N_37139,N_33416,N_30720);
xnor U37140 (N_37140,N_33581,N_33765);
and U37141 (N_37141,N_30185,N_31575);
or U37142 (N_37142,N_33047,N_31308);
nor U37143 (N_37143,N_31151,N_32123);
nor U37144 (N_37144,N_32653,N_32690);
nand U37145 (N_37145,N_34539,N_32721);
and U37146 (N_37146,N_33442,N_33000);
and U37147 (N_37147,N_33044,N_33718);
nor U37148 (N_37148,N_33198,N_34486);
nor U37149 (N_37149,N_33864,N_33153);
nand U37150 (N_37150,N_34973,N_33847);
nand U37151 (N_37151,N_30046,N_32092);
nor U37152 (N_37152,N_31330,N_34162);
nand U37153 (N_37153,N_30205,N_34384);
nand U37154 (N_37154,N_34324,N_33121);
or U37155 (N_37155,N_30898,N_32347);
and U37156 (N_37156,N_30038,N_31039);
xor U37157 (N_37157,N_33982,N_30195);
nor U37158 (N_37158,N_31011,N_32394);
xnor U37159 (N_37159,N_30437,N_30881);
xnor U37160 (N_37160,N_32424,N_34517);
or U37161 (N_37161,N_30235,N_34699);
nor U37162 (N_37162,N_33614,N_33320);
and U37163 (N_37163,N_34983,N_31894);
xor U37164 (N_37164,N_30470,N_33024);
nor U37165 (N_37165,N_32755,N_31776);
nor U37166 (N_37166,N_34867,N_34349);
and U37167 (N_37167,N_34334,N_33215);
nand U37168 (N_37168,N_32239,N_34168);
nand U37169 (N_37169,N_34134,N_30406);
and U37170 (N_37170,N_32258,N_32166);
nand U37171 (N_37171,N_32372,N_34589);
nand U37172 (N_37172,N_30998,N_30207);
and U37173 (N_37173,N_32141,N_31665);
nor U37174 (N_37174,N_34685,N_33899);
nor U37175 (N_37175,N_34022,N_32214);
xnor U37176 (N_37176,N_31087,N_30332);
and U37177 (N_37177,N_30444,N_31147);
or U37178 (N_37178,N_32732,N_34933);
and U37179 (N_37179,N_31135,N_33961);
xor U37180 (N_37180,N_30536,N_31224);
nor U37181 (N_37181,N_32229,N_31810);
nand U37182 (N_37182,N_34854,N_34642);
and U37183 (N_37183,N_33941,N_32298);
nand U37184 (N_37184,N_34131,N_34237);
and U37185 (N_37185,N_30504,N_30246);
nand U37186 (N_37186,N_30869,N_32553);
xnor U37187 (N_37187,N_33608,N_33538);
or U37188 (N_37188,N_34122,N_32612);
or U37189 (N_37189,N_30349,N_31595);
nand U37190 (N_37190,N_34163,N_31422);
xor U37191 (N_37191,N_32070,N_30417);
nand U37192 (N_37192,N_31149,N_31060);
or U37193 (N_37193,N_31716,N_31508);
or U37194 (N_37194,N_31325,N_33760);
and U37195 (N_37195,N_32208,N_30198);
xor U37196 (N_37196,N_30802,N_33913);
nand U37197 (N_37197,N_34271,N_30950);
xor U37198 (N_37198,N_31686,N_32975);
nand U37199 (N_37199,N_34295,N_30543);
nand U37200 (N_37200,N_31418,N_34708);
nor U37201 (N_37201,N_31417,N_31501);
nor U37202 (N_37202,N_32820,N_31972);
or U37203 (N_37203,N_32903,N_30131);
xnor U37204 (N_37204,N_33450,N_31155);
nand U37205 (N_37205,N_32276,N_33687);
or U37206 (N_37206,N_31749,N_34371);
nand U37207 (N_37207,N_30992,N_31985);
and U37208 (N_37208,N_31187,N_33148);
or U37209 (N_37209,N_33312,N_33200);
nand U37210 (N_37210,N_30486,N_33171);
and U37211 (N_37211,N_31863,N_30896);
nor U37212 (N_37212,N_31564,N_31338);
xnor U37213 (N_37213,N_30457,N_34912);
xnor U37214 (N_37214,N_33361,N_33444);
xnor U37215 (N_37215,N_33672,N_34475);
or U37216 (N_37216,N_34226,N_30723);
or U37217 (N_37217,N_33664,N_32131);
and U37218 (N_37218,N_33162,N_33040);
or U37219 (N_37219,N_31397,N_34773);
and U37220 (N_37220,N_31518,N_33297);
nor U37221 (N_37221,N_33665,N_32712);
and U37222 (N_37222,N_33265,N_33343);
xnor U37223 (N_37223,N_32973,N_32193);
nor U37224 (N_37224,N_31880,N_33209);
or U37225 (N_37225,N_33318,N_30093);
and U37226 (N_37226,N_34704,N_33767);
xor U37227 (N_37227,N_32949,N_32484);
nand U37228 (N_37228,N_34976,N_32104);
and U37229 (N_37229,N_34103,N_30586);
and U37230 (N_37230,N_30542,N_34383);
nor U37231 (N_37231,N_31754,N_34688);
or U37232 (N_37232,N_30378,N_31605);
nor U37233 (N_37233,N_32115,N_33372);
xnor U37234 (N_37234,N_33266,N_31442);
xnor U37235 (N_37235,N_30905,N_30512);
or U37236 (N_37236,N_30370,N_32181);
nand U37237 (N_37237,N_31218,N_34000);
xor U37238 (N_37238,N_30766,N_34612);
nand U37239 (N_37239,N_33639,N_31530);
xor U37240 (N_37240,N_31009,N_32068);
nor U37241 (N_37241,N_30217,N_30272);
nor U37242 (N_37242,N_33751,N_33965);
or U37243 (N_37243,N_30648,N_34136);
nor U37244 (N_37244,N_34358,N_33579);
or U37245 (N_37245,N_34436,N_31551);
nand U37246 (N_37246,N_33910,N_34571);
nor U37247 (N_37247,N_31933,N_32480);
nor U37248 (N_37248,N_34179,N_32455);
or U37249 (N_37249,N_32886,N_34352);
or U37250 (N_37250,N_30968,N_32395);
or U37251 (N_37251,N_31337,N_34641);
nor U37252 (N_37252,N_34843,N_34213);
or U37253 (N_37253,N_34735,N_33467);
xor U37254 (N_37254,N_32140,N_30328);
xnor U37255 (N_37255,N_31475,N_30530);
nor U37256 (N_37256,N_34074,N_33630);
and U37257 (N_37257,N_33071,N_34414);
xnor U37258 (N_37258,N_30605,N_33050);
xnor U37259 (N_37259,N_30123,N_33479);
xor U37260 (N_37260,N_30307,N_31579);
nand U37261 (N_37261,N_30298,N_32710);
xor U37262 (N_37262,N_30995,N_33023);
or U37263 (N_37263,N_31321,N_31884);
xnor U37264 (N_37264,N_32554,N_30303);
nor U37265 (N_37265,N_32920,N_31848);
or U37266 (N_37266,N_31652,N_33032);
xnor U37267 (N_37267,N_33269,N_34643);
nor U37268 (N_37268,N_30175,N_33743);
nand U37269 (N_37269,N_31277,N_30564);
xor U37270 (N_37270,N_31443,N_30380);
and U37271 (N_37271,N_34142,N_31792);
and U37272 (N_37272,N_34743,N_30371);
and U37273 (N_37273,N_30480,N_33730);
xor U37274 (N_37274,N_30494,N_31712);
xnor U37275 (N_37275,N_32046,N_34307);
nor U37276 (N_37276,N_30994,N_33386);
or U37277 (N_37277,N_33111,N_31698);
and U37278 (N_37278,N_33657,N_30455);
nand U37279 (N_37279,N_32704,N_34754);
or U37280 (N_37280,N_31986,N_32594);
nand U37281 (N_37281,N_34877,N_30871);
and U37282 (N_37282,N_32266,N_33475);
nand U37283 (N_37283,N_30997,N_31911);
nor U37284 (N_37284,N_30730,N_30450);
nand U37285 (N_37285,N_34559,N_33512);
and U37286 (N_37286,N_34190,N_31648);
and U37287 (N_37287,N_30465,N_30664);
xor U37288 (N_37288,N_34998,N_31109);
nand U37289 (N_37289,N_33651,N_33906);
nand U37290 (N_37290,N_34647,N_33428);
or U37291 (N_37291,N_32650,N_32758);
or U37292 (N_37292,N_33533,N_34206);
or U37293 (N_37293,N_33582,N_34130);
and U37294 (N_37294,N_33370,N_30955);
nand U37295 (N_37295,N_34462,N_32445);
or U37296 (N_37296,N_30518,N_32155);
xor U37297 (N_37297,N_32493,N_30252);
xor U37298 (N_37298,N_30809,N_33466);
xnor U37299 (N_37299,N_32105,N_34970);
nor U37300 (N_37300,N_33499,N_31123);
nand U37301 (N_37301,N_30073,N_31976);
nand U37302 (N_37302,N_33077,N_31785);
xnor U37303 (N_37303,N_33075,N_34065);
nor U37304 (N_37304,N_32245,N_32824);
and U37305 (N_37305,N_33782,N_34311);
or U37306 (N_37306,N_30788,N_31408);
xnor U37307 (N_37307,N_31263,N_34464);
nor U37308 (N_37308,N_32439,N_34582);
nor U37309 (N_37309,N_30581,N_32498);
nand U37310 (N_37310,N_34377,N_31963);
nand U37311 (N_37311,N_31112,N_33117);
xnor U37312 (N_37312,N_34118,N_33872);
and U37313 (N_37313,N_34960,N_30456);
or U37314 (N_37314,N_34678,N_32805);
nand U37315 (N_37315,N_31641,N_31415);
nand U37316 (N_37316,N_32162,N_34503);
nor U37317 (N_37317,N_34040,N_34784);
xnor U37318 (N_37318,N_31617,N_34099);
and U37319 (N_37319,N_33089,N_33839);
and U37320 (N_37320,N_34714,N_33053);
and U37321 (N_37321,N_31812,N_34664);
nand U37322 (N_37322,N_32680,N_32832);
nor U37323 (N_37323,N_30806,N_30128);
or U37324 (N_37324,N_32003,N_34292);
or U37325 (N_37325,N_31280,N_33550);
and U37326 (N_37326,N_30476,N_32059);
or U37327 (N_37327,N_33551,N_34005);
nand U37328 (N_37328,N_33991,N_34609);
nand U37329 (N_37329,N_34505,N_33668);
or U37330 (N_37330,N_30135,N_31378);
or U37331 (N_37331,N_33275,N_32660);
xnor U37332 (N_37332,N_33950,N_34575);
and U37333 (N_37333,N_30817,N_31173);
and U37334 (N_37334,N_33737,N_31603);
and U37335 (N_37335,N_33107,N_30419);
and U37336 (N_37336,N_32995,N_34594);
xnor U37337 (N_37337,N_34243,N_34402);
or U37338 (N_37338,N_31707,N_32197);
xnor U37339 (N_37339,N_30696,N_34152);
nor U37340 (N_37340,N_30362,N_33655);
nor U37341 (N_37341,N_32496,N_32034);
or U37342 (N_37342,N_34222,N_32467);
nand U37343 (N_37343,N_32406,N_31902);
nor U37344 (N_37344,N_31730,N_31013);
and U37345 (N_37345,N_32021,N_33226);
or U37346 (N_37346,N_30015,N_31315);
or U37347 (N_37347,N_34221,N_30739);
nand U37348 (N_37348,N_32900,N_33410);
xor U37349 (N_37349,N_30989,N_34174);
or U37350 (N_37350,N_34458,N_31150);
xnor U37351 (N_37351,N_34950,N_31560);
nor U37352 (N_37352,N_32010,N_30702);
nand U37353 (N_37353,N_30760,N_31302);
or U37354 (N_37354,N_32968,N_30299);
nand U37355 (N_37355,N_34842,N_34326);
nor U37356 (N_37356,N_32453,N_31003);
or U37357 (N_37357,N_31379,N_34437);
and U37358 (N_37358,N_30550,N_34095);
xor U37359 (N_37359,N_31383,N_30074);
or U37360 (N_37360,N_33956,N_32909);
nor U37361 (N_37361,N_32223,N_34778);
nor U37362 (N_37362,N_32238,N_33172);
nand U37363 (N_37363,N_30433,N_30771);
nand U37364 (N_37364,N_31842,N_31864);
nand U37365 (N_37365,N_31191,N_30009);
or U37366 (N_37366,N_31304,N_32265);
xnor U37367 (N_37367,N_31176,N_30910);
nand U37368 (N_37368,N_34926,N_30626);
xor U37369 (N_37369,N_31602,N_34211);
nor U37370 (N_37370,N_32250,N_31271);
xnor U37371 (N_37371,N_30669,N_32485);
and U37372 (N_37372,N_32169,N_30134);
and U37373 (N_37373,N_32578,N_31907);
nor U37374 (N_37374,N_33219,N_34684);
and U37375 (N_37375,N_31033,N_32038);
nor U37376 (N_37376,N_30849,N_33351);
nor U37377 (N_37377,N_32043,N_33042);
nor U37378 (N_37378,N_30108,N_30133);
or U37379 (N_37379,N_33317,N_32230);
or U37380 (N_37380,N_30934,N_30087);
xnor U37381 (N_37381,N_34500,N_30269);
and U37382 (N_37382,N_32120,N_33583);
nand U37383 (N_37383,N_31892,N_33185);
or U37384 (N_37384,N_32700,N_30034);
and U37385 (N_37385,N_34606,N_30603);
nor U37386 (N_37386,N_31392,N_31553);
and U37387 (N_37387,N_34705,N_34283);
and U37388 (N_37388,N_33774,N_34815);
and U37389 (N_37389,N_32809,N_31162);
xnor U37390 (N_37390,N_32679,N_34631);
xnor U37391 (N_37391,N_32390,N_32441);
or U37392 (N_37392,N_32958,N_31245);
or U37393 (N_37393,N_30891,N_34859);
or U37394 (N_37394,N_33734,N_30287);
nor U37395 (N_37395,N_34066,N_33926);
and U37396 (N_37396,N_33565,N_30666);
or U37397 (N_37397,N_33842,N_30385);
xnor U37398 (N_37398,N_31699,N_34882);
xnor U37399 (N_37399,N_31314,N_33868);
and U37400 (N_37400,N_34256,N_32118);
xor U37401 (N_37401,N_32888,N_32415);
or U37402 (N_37402,N_31183,N_34030);
nand U37403 (N_37403,N_34146,N_31702);
nor U37404 (N_37404,N_33527,N_30422);
nand U37405 (N_37405,N_34900,N_34329);
xor U37406 (N_37406,N_30492,N_30590);
nor U37407 (N_37407,N_30638,N_34888);
nor U37408 (N_37408,N_30001,N_33633);
and U37409 (N_37409,N_31364,N_33013);
nor U37410 (N_37410,N_30368,N_32125);
nor U37411 (N_37411,N_30315,N_33335);
or U37412 (N_37412,N_32874,N_33449);
nand U37413 (N_37413,N_33206,N_32867);
xnor U37414 (N_37414,N_30436,N_31426);
nand U37415 (N_37415,N_33243,N_32447);
xor U37416 (N_37416,N_33333,N_31260);
nor U37417 (N_37417,N_33224,N_30360);
and U37418 (N_37418,N_34167,N_32575);
or U37419 (N_37419,N_31345,N_30725);
nand U37420 (N_37420,N_30835,N_33454);
nand U37421 (N_37421,N_30364,N_31434);
nor U37422 (N_37422,N_30623,N_30566);
and U37423 (N_37423,N_32628,N_31125);
nand U37424 (N_37424,N_31541,N_30231);
nor U37425 (N_37425,N_33862,N_31479);
xor U37426 (N_37426,N_32924,N_34632);
and U37427 (N_37427,N_30718,N_30773);
xnor U37428 (N_37428,N_32747,N_30925);
and U37429 (N_37429,N_32538,N_34195);
or U37430 (N_37430,N_32881,N_33308);
xor U37431 (N_37431,N_30729,N_32316);
nor U37432 (N_37432,N_33115,N_31611);
or U37433 (N_37433,N_33309,N_34633);
nand U37434 (N_37434,N_33520,N_30978);
nor U37435 (N_37435,N_34153,N_30228);
nor U37436 (N_37436,N_30707,N_30851);
nand U37437 (N_37437,N_31278,N_31232);
xnor U37438 (N_37438,N_30949,N_30186);
and U37439 (N_37439,N_31978,N_30048);
nor U37440 (N_37440,N_31522,N_33257);
and U37441 (N_37441,N_30876,N_32890);
nand U37442 (N_37442,N_30772,N_30223);
nor U37443 (N_37443,N_33626,N_34041);
nor U37444 (N_37444,N_31197,N_34923);
nand U37445 (N_37445,N_34262,N_34106);
nand U37446 (N_37446,N_34943,N_31256);
nor U37447 (N_37447,N_32402,N_33891);
or U37448 (N_37448,N_31275,N_30620);
nor U37449 (N_37449,N_30449,N_30939);
nor U37450 (N_37450,N_33953,N_32504);
or U37451 (N_37451,N_32536,N_32121);
nor U37452 (N_37452,N_31822,N_33304);
or U37453 (N_37453,N_32608,N_34617);
nor U37454 (N_37454,N_31593,N_30415);
xnor U37455 (N_37455,N_34412,N_32180);
nand U37456 (N_37456,N_31133,N_30113);
or U37457 (N_37457,N_31878,N_33139);
nor U37458 (N_37458,N_32433,N_32411);
or U37459 (N_37459,N_34639,N_33684);
or U37460 (N_37460,N_30831,N_32733);
and U37461 (N_37461,N_33227,N_32322);
xnor U37462 (N_37462,N_33271,N_32716);
or U37463 (N_37463,N_32817,N_34514);
nand U37464 (N_37464,N_33218,N_31375);
nand U37465 (N_37465,N_34587,N_30479);
and U37466 (N_37466,N_31905,N_31926);
nor U37467 (N_37467,N_33244,N_30611);
or U37468 (N_37468,N_30323,N_30438);
xnor U37469 (N_37469,N_31782,N_33854);
nand U37470 (N_37470,N_30553,N_33793);
nor U37471 (N_37471,N_31054,N_34321);
nand U37472 (N_37472,N_34564,N_32967);
xor U37473 (N_37473,N_32894,N_33254);
nor U37474 (N_37474,N_30066,N_34411);
nand U37475 (N_37475,N_32089,N_30124);
xor U37476 (N_37476,N_33216,N_32005);
and U37477 (N_37477,N_33708,N_32681);
nor U37478 (N_37478,N_33683,N_30054);
nand U37479 (N_37479,N_32917,N_34731);
or U37480 (N_37480,N_31496,N_31845);
nor U37481 (N_37481,N_34906,N_32954);
and U37482 (N_37482,N_33808,N_32985);
nand U37483 (N_37483,N_34446,N_34228);
nand U37484 (N_37484,N_32064,N_32793);
or U37485 (N_37485,N_32304,N_34757);
nand U37486 (N_37486,N_30114,N_33812);
xnor U37487 (N_37487,N_33448,N_30631);
and U37488 (N_37488,N_30268,N_33701);
and U37489 (N_37489,N_33786,N_34824);
nand U37490 (N_37490,N_34727,N_30890);
nand U37491 (N_37491,N_33929,N_33181);
or U37492 (N_37492,N_34372,N_30850);
or U37493 (N_37493,N_33160,N_33332);
and U37494 (N_37494,N_30618,N_32771);
or U37495 (N_37495,N_31312,N_30598);
or U37496 (N_37496,N_33112,N_30173);
nand U37497 (N_37497,N_32464,N_30396);
xnor U37498 (N_37498,N_33022,N_31002);
or U37499 (N_37499,N_32460,N_31361);
and U37500 (N_37500,N_30188,N_32833);
and U37501 (N_37501,N_33788,N_32148);
or U37502 (N_37502,N_31846,N_33705);
nand U37503 (N_37503,N_30183,N_31093);
or U37504 (N_37504,N_31616,N_33287);
nand U37505 (N_37505,N_34558,N_30585);
nand U37506 (N_37506,N_33248,N_33776);
nand U37507 (N_37507,N_34575,N_30222);
xnor U37508 (N_37508,N_31023,N_33588);
xnor U37509 (N_37509,N_34465,N_33020);
and U37510 (N_37510,N_34149,N_32666);
xor U37511 (N_37511,N_34251,N_34926);
nor U37512 (N_37512,N_31394,N_31547);
or U37513 (N_37513,N_31873,N_30198);
nor U37514 (N_37514,N_31777,N_32801);
xor U37515 (N_37515,N_30246,N_33001);
nand U37516 (N_37516,N_32638,N_33697);
or U37517 (N_37517,N_31112,N_34905);
xor U37518 (N_37518,N_33319,N_34119);
nor U37519 (N_37519,N_33899,N_33288);
nor U37520 (N_37520,N_34583,N_33572);
xor U37521 (N_37521,N_34352,N_32363);
nand U37522 (N_37522,N_32772,N_33721);
and U37523 (N_37523,N_30730,N_32336);
xnor U37524 (N_37524,N_33085,N_34909);
and U37525 (N_37525,N_33585,N_31017);
and U37526 (N_37526,N_32979,N_34086);
nand U37527 (N_37527,N_32690,N_31923);
nand U37528 (N_37528,N_33317,N_33664);
and U37529 (N_37529,N_34797,N_34170);
or U37530 (N_37530,N_32403,N_31970);
nor U37531 (N_37531,N_33685,N_34397);
nor U37532 (N_37532,N_31210,N_30816);
nand U37533 (N_37533,N_31589,N_34356);
and U37534 (N_37534,N_31398,N_33627);
nand U37535 (N_37535,N_31782,N_31074);
nor U37536 (N_37536,N_32261,N_33215);
or U37537 (N_37537,N_30607,N_32237);
xor U37538 (N_37538,N_30976,N_32586);
and U37539 (N_37539,N_33498,N_34964);
nand U37540 (N_37540,N_33434,N_32868);
or U37541 (N_37541,N_32084,N_31135);
xor U37542 (N_37542,N_30696,N_34827);
and U37543 (N_37543,N_33468,N_33727);
nand U37544 (N_37544,N_30549,N_32465);
nand U37545 (N_37545,N_30701,N_34694);
and U37546 (N_37546,N_32302,N_33365);
nor U37547 (N_37547,N_31913,N_30686);
and U37548 (N_37548,N_30664,N_33967);
xnor U37549 (N_37549,N_32886,N_33668);
xor U37550 (N_37550,N_30447,N_32155);
nor U37551 (N_37551,N_31507,N_31333);
or U37552 (N_37552,N_34127,N_33175);
nor U37553 (N_37553,N_32645,N_32614);
nand U37554 (N_37554,N_32900,N_32205);
nor U37555 (N_37555,N_30334,N_33954);
nand U37556 (N_37556,N_34105,N_31084);
nor U37557 (N_37557,N_34274,N_33182);
or U37558 (N_37558,N_32499,N_31865);
or U37559 (N_37559,N_33776,N_32891);
nor U37560 (N_37560,N_31251,N_30128);
and U37561 (N_37561,N_31663,N_33991);
nor U37562 (N_37562,N_34263,N_34509);
nor U37563 (N_37563,N_34556,N_33580);
xor U37564 (N_37564,N_30670,N_34742);
and U37565 (N_37565,N_32813,N_34930);
xnor U37566 (N_37566,N_30052,N_33057);
xor U37567 (N_37567,N_33723,N_34027);
nand U37568 (N_37568,N_33559,N_32661);
nor U37569 (N_37569,N_30465,N_30507);
or U37570 (N_37570,N_33365,N_33039);
and U37571 (N_37571,N_33652,N_30514);
xnor U37572 (N_37572,N_32071,N_30053);
xor U37573 (N_37573,N_34524,N_30980);
xor U37574 (N_37574,N_31701,N_30457);
nor U37575 (N_37575,N_32089,N_31056);
xnor U37576 (N_37576,N_31075,N_30819);
or U37577 (N_37577,N_31149,N_31382);
xnor U37578 (N_37578,N_33614,N_31902);
nor U37579 (N_37579,N_33642,N_32192);
nor U37580 (N_37580,N_32167,N_34721);
and U37581 (N_37581,N_34117,N_30392);
nand U37582 (N_37582,N_34770,N_32764);
or U37583 (N_37583,N_31719,N_31472);
nor U37584 (N_37584,N_34970,N_34909);
nand U37585 (N_37585,N_31521,N_33220);
nand U37586 (N_37586,N_31738,N_34729);
nand U37587 (N_37587,N_33846,N_34398);
nand U37588 (N_37588,N_33217,N_33279);
nor U37589 (N_37589,N_31572,N_30629);
xor U37590 (N_37590,N_31357,N_32829);
or U37591 (N_37591,N_34237,N_33042);
xor U37592 (N_37592,N_34492,N_34902);
and U37593 (N_37593,N_30534,N_33404);
xor U37594 (N_37594,N_34528,N_33336);
nor U37595 (N_37595,N_31579,N_33053);
and U37596 (N_37596,N_31889,N_32714);
or U37597 (N_37597,N_30033,N_34067);
and U37598 (N_37598,N_32774,N_32070);
and U37599 (N_37599,N_34946,N_31381);
nand U37600 (N_37600,N_31108,N_33712);
xnor U37601 (N_37601,N_33342,N_30018);
and U37602 (N_37602,N_32384,N_34618);
xor U37603 (N_37603,N_31780,N_33204);
or U37604 (N_37604,N_31320,N_34409);
nand U37605 (N_37605,N_32062,N_31378);
nor U37606 (N_37606,N_33454,N_33769);
nor U37607 (N_37607,N_32673,N_30184);
and U37608 (N_37608,N_34354,N_30189);
or U37609 (N_37609,N_32846,N_31052);
nand U37610 (N_37610,N_34209,N_33719);
and U37611 (N_37611,N_31764,N_30181);
and U37612 (N_37612,N_33295,N_32949);
or U37613 (N_37613,N_34493,N_33596);
xnor U37614 (N_37614,N_33155,N_30728);
nor U37615 (N_37615,N_34112,N_30990);
nor U37616 (N_37616,N_34762,N_34777);
xor U37617 (N_37617,N_32573,N_32662);
xor U37618 (N_37618,N_32490,N_32520);
and U37619 (N_37619,N_34410,N_31945);
xnor U37620 (N_37620,N_31324,N_31063);
nand U37621 (N_37621,N_34025,N_30243);
xor U37622 (N_37622,N_33814,N_33195);
and U37623 (N_37623,N_32213,N_30958);
or U37624 (N_37624,N_31753,N_30206);
xnor U37625 (N_37625,N_32637,N_34226);
nor U37626 (N_37626,N_34472,N_33915);
and U37627 (N_37627,N_33402,N_30688);
nand U37628 (N_37628,N_31284,N_30603);
and U37629 (N_37629,N_30139,N_30602);
and U37630 (N_37630,N_34518,N_32390);
xor U37631 (N_37631,N_32828,N_32939);
xnor U37632 (N_37632,N_32681,N_30686);
nor U37633 (N_37633,N_32743,N_30287);
nand U37634 (N_37634,N_32189,N_33688);
and U37635 (N_37635,N_34187,N_30408);
xor U37636 (N_37636,N_30090,N_34589);
nor U37637 (N_37637,N_31904,N_30496);
xnor U37638 (N_37638,N_32954,N_34353);
or U37639 (N_37639,N_34420,N_31283);
nand U37640 (N_37640,N_32087,N_33800);
or U37641 (N_37641,N_31547,N_33235);
nor U37642 (N_37642,N_34769,N_33838);
xor U37643 (N_37643,N_32784,N_33070);
or U37644 (N_37644,N_33313,N_31101);
nor U37645 (N_37645,N_32458,N_30282);
nand U37646 (N_37646,N_32950,N_33722);
xnor U37647 (N_37647,N_32527,N_30304);
nand U37648 (N_37648,N_31608,N_30048);
nand U37649 (N_37649,N_30464,N_31733);
xor U37650 (N_37650,N_34751,N_34388);
nor U37651 (N_37651,N_33391,N_32240);
and U37652 (N_37652,N_30786,N_31256);
nor U37653 (N_37653,N_30995,N_33942);
xor U37654 (N_37654,N_31344,N_31379);
xnor U37655 (N_37655,N_33983,N_33609);
xnor U37656 (N_37656,N_32106,N_32299);
nand U37657 (N_37657,N_30452,N_30785);
and U37658 (N_37658,N_32781,N_30755);
nand U37659 (N_37659,N_34427,N_34869);
nor U37660 (N_37660,N_33411,N_32360);
or U37661 (N_37661,N_33854,N_32970);
xnor U37662 (N_37662,N_31924,N_30612);
xnor U37663 (N_37663,N_30842,N_33743);
xnor U37664 (N_37664,N_34250,N_32558);
or U37665 (N_37665,N_32804,N_34876);
xor U37666 (N_37666,N_32192,N_30802);
nor U37667 (N_37667,N_32957,N_34315);
and U37668 (N_37668,N_30097,N_33420);
nand U37669 (N_37669,N_33417,N_32108);
and U37670 (N_37670,N_31838,N_31130);
or U37671 (N_37671,N_31580,N_32696);
xor U37672 (N_37672,N_30571,N_31804);
nand U37673 (N_37673,N_30025,N_33210);
nand U37674 (N_37674,N_34428,N_31238);
xor U37675 (N_37675,N_30468,N_33222);
nor U37676 (N_37676,N_32808,N_34414);
or U37677 (N_37677,N_31966,N_32214);
nor U37678 (N_37678,N_30319,N_34282);
nand U37679 (N_37679,N_34931,N_31278);
nor U37680 (N_37680,N_34693,N_33094);
xnor U37681 (N_37681,N_34250,N_31037);
nand U37682 (N_37682,N_32531,N_33765);
nand U37683 (N_37683,N_34526,N_34495);
nand U37684 (N_37684,N_31068,N_30554);
xor U37685 (N_37685,N_34885,N_33198);
nor U37686 (N_37686,N_32870,N_34663);
and U37687 (N_37687,N_34057,N_32276);
xnor U37688 (N_37688,N_33418,N_31343);
and U37689 (N_37689,N_33888,N_33301);
nor U37690 (N_37690,N_34682,N_32600);
and U37691 (N_37691,N_30394,N_34726);
nand U37692 (N_37692,N_31837,N_31294);
xor U37693 (N_37693,N_31105,N_33952);
nand U37694 (N_37694,N_31030,N_34380);
xor U37695 (N_37695,N_30238,N_31474);
nor U37696 (N_37696,N_34069,N_34312);
xor U37697 (N_37697,N_33209,N_34232);
nor U37698 (N_37698,N_30919,N_30312);
and U37699 (N_37699,N_33899,N_30361);
nor U37700 (N_37700,N_31760,N_33398);
xnor U37701 (N_37701,N_32073,N_34778);
and U37702 (N_37702,N_31404,N_34981);
or U37703 (N_37703,N_32458,N_33376);
nor U37704 (N_37704,N_30203,N_34080);
xnor U37705 (N_37705,N_34052,N_32872);
xnor U37706 (N_37706,N_31655,N_30633);
nor U37707 (N_37707,N_34270,N_31801);
nand U37708 (N_37708,N_33775,N_30651);
or U37709 (N_37709,N_31904,N_31942);
nor U37710 (N_37710,N_32684,N_32317);
nand U37711 (N_37711,N_31970,N_34190);
or U37712 (N_37712,N_31036,N_30316);
and U37713 (N_37713,N_33691,N_30917);
and U37714 (N_37714,N_32789,N_31241);
and U37715 (N_37715,N_31550,N_30828);
xnor U37716 (N_37716,N_31860,N_31214);
xnor U37717 (N_37717,N_32011,N_30030);
nor U37718 (N_37718,N_30718,N_34150);
and U37719 (N_37719,N_31649,N_34035);
and U37720 (N_37720,N_33849,N_34033);
or U37721 (N_37721,N_32640,N_34757);
or U37722 (N_37722,N_30772,N_32040);
nand U37723 (N_37723,N_34953,N_33245);
nor U37724 (N_37724,N_32716,N_33251);
xor U37725 (N_37725,N_33335,N_34139);
nor U37726 (N_37726,N_30928,N_30098);
nand U37727 (N_37727,N_30751,N_34193);
xnor U37728 (N_37728,N_33696,N_30546);
or U37729 (N_37729,N_31377,N_32961);
and U37730 (N_37730,N_31633,N_32572);
nand U37731 (N_37731,N_30377,N_31705);
xnor U37732 (N_37732,N_32391,N_30460);
nor U37733 (N_37733,N_30418,N_31040);
nand U37734 (N_37734,N_30469,N_34879);
nand U37735 (N_37735,N_31544,N_33906);
nor U37736 (N_37736,N_33860,N_32340);
or U37737 (N_37737,N_33325,N_30203);
nand U37738 (N_37738,N_30878,N_32707);
and U37739 (N_37739,N_33204,N_30681);
nor U37740 (N_37740,N_31265,N_30421);
nor U37741 (N_37741,N_34463,N_32931);
or U37742 (N_37742,N_30158,N_32958);
nor U37743 (N_37743,N_32788,N_33445);
xor U37744 (N_37744,N_31709,N_30594);
nor U37745 (N_37745,N_31313,N_31809);
nor U37746 (N_37746,N_34385,N_30277);
or U37747 (N_37747,N_31749,N_32756);
nand U37748 (N_37748,N_30111,N_30576);
and U37749 (N_37749,N_30809,N_32785);
nand U37750 (N_37750,N_34858,N_30808);
nor U37751 (N_37751,N_31929,N_34015);
or U37752 (N_37752,N_34909,N_32708);
and U37753 (N_37753,N_33417,N_33051);
or U37754 (N_37754,N_31095,N_30687);
and U37755 (N_37755,N_34757,N_32576);
or U37756 (N_37756,N_31718,N_30595);
nor U37757 (N_37757,N_32621,N_33567);
nand U37758 (N_37758,N_31119,N_30881);
xnor U37759 (N_37759,N_33089,N_32637);
nand U37760 (N_37760,N_34490,N_33602);
nor U37761 (N_37761,N_30662,N_31417);
nor U37762 (N_37762,N_30996,N_32134);
xor U37763 (N_37763,N_32465,N_30259);
xor U37764 (N_37764,N_31457,N_32012);
nor U37765 (N_37765,N_31151,N_34106);
or U37766 (N_37766,N_31882,N_34765);
nand U37767 (N_37767,N_32153,N_30299);
nor U37768 (N_37768,N_32068,N_34569);
or U37769 (N_37769,N_31477,N_32542);
xor U37770 (N_37770,N_32558,N_33275);
nand U37771 (N_37771,N_34945,N_30603);
and U37772 (N_37772,N_30623,N_31204);
xor U37773 (N_37773,N_31467,N_31638);
nand U37774 (N_37774,N_34868,N_31723);
and U37775 (N_37775,N_33722,N_33770);
xnor U37776 (N_37776,N_34361,N_33912);
or U37777 (N_37777,N_34152,N_33722);
nand U37778 (N_37778,N_30682,N_31624);
nand U37779 (N_37779,N_30552,N_30812);
and U37780 (N_37780,N_31915,N_30343);
and U37781 (N_37781,N_34140,N_31327);
and U37782 (N_37782,N_30765,N_31871);
xor U37783 (N_37783,N_33756,N_34198);
and U37784 (N_37784,N_32433,N_30519);
xor U37785 (N_37785,N_31378,N_34945);
and U37786 (N_37786,N_34196,N_34741);
xor U37787 (N_37787,N_31349,N_31339);
and U37788 (N_37788,N_32361,N_34166);
xor U37789 (N_37789,N_30479,N_31321);
nand U37790 (N_37790,N_30857,N_33085);
xnor U37791 (N_37791,N_32560,N_34224);
or U37792 (N_37792,N_30377,N_31580);
nor U37793 (N_37793,N_33519,N_30551);
nand U37794 (N_37794,N_34202,N_30120);
nand U37795 (N_37795,N_30309,N_33020);
nor U37796 (N_37796,N_33261,N_33238);
nand U37797 (N_37797,N_33851,N_33323);
nor U37798 (N_37798,N_30627,N_30801);
nand U37799 (N_37799,N_33486,N_33693);
xnor U37800 (N_37800,N_31008,N_32414);
and U37801 (N_37801,N_34633,N_34040);
xor U37802 (N_37802,N_30593,N_33317);
and U37803 (N_37803,N_31178,N_32141);
and U37804 (N_37804,N_30354,N_31838);
and U37805 (N_37805,N_31485,N_31724);
or U37806 (N_37806,N_30919,N_33578);
and U37807 (N_37807,N_30452,N_34179);
xnor U37808 (N_37808,N_34280,N_31762);
xnor U37809 (N_37809,N_30698,N_32929);
or U37810 (N_37810,N_32444,N_34945);
xor U37811 (N_37811,N_32793,N_34250);
or U37812 (N_37812,N_30483,N_34207);
nand U37813 (N_37813,N_34435,N_32375);
and U37814 (N_37814,N_31672,N_30246);
and U37815 (N_37815,N_33541,N_32481);
nand U37816 (N_37816,N_30172,N_32895);
and U37817 (N_37817,N_34374,N_30362);
and U37818 (N_37818,N_33518,N_31309);
and U37819 (N_37819,N_34377,N_32398);
and U37820 (N_37820,N_30464,N_33727);
nor U37821 (N_37821,N_32745,N_34495);
or U37822 (N_37822,N_34309,N_32000);
nand U37823 (N_37823,N_33130,N_31299);
or U37824 (N_37824,N_30552,N_31076);
xnor U37825 (N_37825,N_30088,N_32834);
nor U37826 (N_37826,N_34407,N_31896);
nor U37827 (N_37827,N_34252,N_32127);
nor U37828 (N_37828,N_31257,N_34547);
and U37829 (N_37829,N_31567,N_31643);
or U37830 (N_37830,N_30334,N_33398);
or U37831 (N_37831,N_30618,N_34716);
nor U37832 (N_37832,N_32234,N_32548);
xnor U37833 (N_37833,N_31031,N_33108);
nand U37834 (N_37834,N_31769,N_31838);
nor U37835 (N_37835,N_33005,N_33566);
xor U37836 (N_37836,N_30951,N_31800);
or U37837 (N_37837,N_33965,N_30534);
or U37838 (N_37838,N_34620,N_30577);
and U37839 (N_37839,N_34512,N_34375);
and U37840 (N_37840,N_31814,N_34347);
nor U37841 (N_37841,N_34737,N_34281);
and U37842 (N_37842,N_31440,N_30251);
and U37843 (N_37843,N_30118,N_30704);
nor U37844 (N_37844,N_30306,N_30641);
nand U37845 (N_37845,N_33249,N_30256);
and U37846 (N_37846,N_31306,N_31175);
nand U37847 (N_37847,N_30591,N_34786);
nand U37848 (N_37848,N_33831,N_31008);
xnor U37849 (N_37849,N_33373,N_31871);
or U37850 (N_37850,N_32764,N_33503);
and U37851 (N_37851,N_32944,N_30006);
xnor U37852 (N_37852,N_30329,N_33910);
xnor U37853 (N_37853,N_30631,N_30948);
xor U37854 (N_37854,N_30890,N_32039);
nor U37855 (N_37855,N_34894,N_31066);
nor U37856 (N_37856,N_30472,N_32278);
or U37857 (N_37857,N_33645,N_34341);
and U37858 (N_37858,N_31302,N_30776);
xor U37859 (N_37859,N_30514,N_33581);
nand U37860 (N_37860,N_34667,N_34714);
xnor U37861 (N_37861,N_30876,N_33720);
and U37862 (N_37862,N_30654,N_33003);
nand U37863 (N_37863,N_34378,N_33449);
nor U37864 (N_37864,N_31549,N_31281);
or U37865 (N_37865,N_33443,N_30858);
and U37866 (N_37866,N_34910,N_33440);
and U37867 (N_37867,N_33331,N_34778);
and U37868 (N_37868,N_32862,N_30773);
and U37869 (N_37869,N_31250,N_33144);
nand U37870 (N_37870,N_32285,N_33588);
nor U37871 (N_37871,N_31554,N_31059);
xor U37872 (N_37872,N_33670,N_31029);
nor U37873 (N_37873,N_32198,N_34382);
nor U37874 (N_37874,N_30411,N_30471);
nand U37875 (N_37875,N_30254,N_32954);
nand U37876 (N_37876,N_31425,N_30633);
nor U37877 (N_37877,N_33349,N_34268);
and U37878 (N_37878,N_30767,N_32855);
nor U37879 (N_37879,N_30876,N_32766);
or U37880 (N_37880,N_33068,N_31196);
nand U37881 (N_37881,N_31670,N_34677);
nor U37882 (N_37882,N_31286,N_32526);
and U37883 (N_37883,N_33986,N_32666);
or U37884 (N_37884,N_33037,N_34416);
nand U37885 (N_37885,N_34803,N_32306);
and U37886 (N_37886,N_32899,N_31109);
nand U37887 (N_37887,N_33115,N_30199);
or U37888 (N_37888,N_30154,N_32242);
and U37889 (N_37889,N_34968,N_31619);
nor U37890 (N_37890,N_34508,N_33710);
xnor U37891 (N_37891,N_32242,N_32199);
nand U37892 (N_37892,N_34186,N_30605);
xor U37893 (N_37893,N_30671,N_34607);
nor U37894 (N_37894,N_31896,N_34819);
or U37895 (N_37895,N_33925,N_32850);
nand U37896 (N_37896,N_30184,N_33689);
nand U37897 (N_37897,N_32027,N_31749);
xnor U37898 (N_37898,N_32415,N_33341);
nand U37899 (N_37899,N_34534,N_32724);
and U37900 (N_37900,N_32640,N_31383);
nand U37901 (N_37901,N_33720,N_33721);
nand U37902 (N_37902,N_33952,N_30259);
xnor U37903 (N_37903,N_31539,N_31120);
nand U37904 (N_37904,N_33451,N_31349);
nor U37905 (N_37905,N_30284,N_30936);
xnor U37906 (N_37906,N_33835,N_31549);
xnor U37907 (N_37907,N_32432,N_34127);
and U37908 (N_37908,N_34727,N_34025);
xor U37909 (N_37909,N_32602,N_33310);
and U37910 (N_37910,N_32162,N_31833);
xor U37911 (N_37911,N_34603,N_30585);
or U37912 (N_37912,N_33531,N_33247);
nand U37913 (N_37913,N_30661,N_30804);
nand U37914 (N_37914,N_34801,N_33767);
or U37915 (N_37915,N_34208,N_33833);
xor U37916 (N_37916,N_30874,N_31109);
xor U37917 (N_37917,N_30084,N_32971);
and U37918 (N_37918,N_33529,N_30867);
or U37919 (N_37919,N_30603,N_30839);
nand U37920 (N_37920,N_31950,N_34634);
nand U37921 (N_37921,N_32012,N_33979);
or U37922 (N_37922,N_31129,N_33205);
xor U37923 (N_37923,N_30692,N_34974);
nor U37924 (N_37924,N_33448,N_30485);
or U37925 (N_37925,N_30958,N_30340);
nand U37926 (N_37926,N_30941,N_34668);
nor U37927 (N_37927,N_33216,N_30169);
nand U37928 (N_37928,N_30927,N_31231);
and U37929 (N_37929,N_34671,N_31918);
nand U37930 (N_37930,N_31505,N_30343);
nand U37931 (N_37931,N_30216,N_34527);
nor U37932 (N_37932,N_33958,N_30309);
or U37933 (N_37933,N_32316,N_33833);
nor U37934 (N_37934,N_33301,N_32102);
nor U37935 (N_37935,N_31317,N_33785);
nand U37936 (N_37936,N_31837,N_34106);
nand U37937 (N_37937,N_32740,N_31922);
or U37938 (N_37938,N_33243,N_31962);
or U37939 (N_37939,N_33589,N_32445);
nor U37940 (N_37940,N_33204,N_34952);
or U37941 (N_37941,N_30448,N_34838);
nor U37942 (N_37942,N_32885,N_32101);
nor U37943 (N_37943,N_33269,N_31196);
nand U37944 (N_37944,N_32649,N_32769);
xor U37945 (N_37945,N_30456,N_32238);
xnor U37946 (N_37946,N_33877,N_31394);
xnor U37947 (N_37947,N_30724,N_31726);
nor U37948 (N_37948,N_32575,N_34169);
and U37949 (N_37949,N_34639,N_31952);
xor U37950 (N_37950,N_32124,N_31440);
and U37951 (N_37951,N_33475,N_32108);
xnor U37952 (N_37952,N_30610,N_33967);
xnor U37953 (N_37953,N_32763,N_33791);
nand U37954 (N_37954,N_31002,N_34178);
nand U37955 (N_37955,N_32298,N_33881);
and U37956 (N_37956,N_31742,N_32532);
nor U37957 (N_37957,N_34730,N_34504);
or U37958 (N_37958,N_31348,N_33948);
nor U37959 (N_37959,N_33926,N_33436);
nand U37960 (N_37960,N_32522,N_33723);
nor U37961 (N_37961,N_33124,N_31895);
xnor U37962 (N_37962,N_32030,N_34642);
and U37963 (N_37963,N_30398,N_34940);
nor U37964 (N_37964,N_33945,N_33792);
and U37965 (N_37965,N_31940,N_32198);
nor U37966 (N_37966,N_30785,N_30579);
and U37967 (N_37967,N_30916,N_30360);
nor U37968 (N_37968,N_30337,N_30221);
nand U37969 (N_37969,N_33277,N_32721);
xor U37970 (N_37970,N_30857,N_31399);
nand U37971 (N_37971,N_31980,N_33296);
or U37972 (N_37972,N_30198,N_34232);
nand U37973 (N_37973,N_33069,N_32146);
and U37974 (N_37974,N_31997,N_31347);
xnor U37975 (N_37975,N_33736,N_33988);
nand U37976 (N_37976,N_30876,N_33364);
and U37977 (N_37977,N_32198,N_33424);
xor U37978 (N_37978,N_30498,N_30550);
and U37979 (N_37979,N_34877,N_30542);
xnor U37980 (N_37980,N_32816,N_34608);
nor U37981 (N_37981,N_32139,N_32043);
xor U37982 (N_37982,N_33247,N_30469);
xor U37983 (N_37983,N_30585,N_31578);
xnor U37984 (N_37984,N_33120,N_32624);
or U37985 (N_37985,N_33171,N_31347);
and U37986 (N_37986,N_33124,N_30693);
and U37987 (N_37987,N_34542,N_30297);
nand U37988 (N_37988,N_31239,N_32021);
xnor U37989 (N_37989,N_34714,N_30384);
nand U37990 (N_37990,N_33581,N_34599);
xnor U37991 (N_37991,N_32471,N_33748);
xnor U37992 (N_37992,N_31271,N_33260);
nand U37993 (N_37993,N_30347,N_31725);
xor U37994 (N_37994,N_34425,N_33723);
and U37995 (N_37995,N_32369,N_31174);
or U37996 (N_37996,N_31852,N_31052);
nor U37997 (N_37997,N_33629,N_31809);
xnor U37998 (N_37998,N_32258,N_33460);
or U37999 (N_37999,N_34380,N_31234);
xor U38000 (N_38000,N_31355,N_31974);
xor U38001 (N_38001,N_32114,N_30590);
xor U38002 (N_38002,N_33416,N_34045);
xnor U38003 (N_38003,N_32651,N_34339);
and U38004 (N_38004,N_30196,N_30881);
or U38005 (N_38005,N_33470,N_31306);
and U38006 (N_38006,N_31714,N_34007);
and U38007 (N_38007,N_33962,N_34048);
or U38008 (N_38008,N_30296,N_33309);
xnor U38009 (N_38009,N_30009,N_34677);
or U38010 (N_38010,N_30336,N_31813);
or U38011 (N_38011,N_30767,N_34181);
and U38012 (N_38012,N_33009,N_30711);
xnor U38013 (N_38013,N_33729,N_30014);
xor U38014 (N_38014,N_31042,N_34599);
xnor U38015 (N_38015,N_34616,N_31329);
xor U38016 (N_38016,N_32686,N_30693);
xor U38017 (N_38017,N_32726,N_33665);
xnor U38018 (N_38018,N_33223,N_33579);
xnor U38019 (N_38019,N_31557,N_30125);
and U38020 (N_38020,N_34551,N_32226);
or U38021 (N_38021,N_30558,N_34725);
xnor U38022 (N_38022,N_30003,N_31355);
and U38023 (N_38023,N_30373,N_32856);
xor U38024 (N_38024,N_32352,N_32042);
nor U38025 (N_38025,N_31565,N_32259);
xnor U38026 (N_38026,N_34823,N_34556);
and U38027 (N_38027,N_30605,N_30254);
and U38028 (N_38028,N_30955,N_30959);
nand U38029 (N_38029,N_31909,N_31095);
or U38030 (N_38030,N_33659,N_30121);
or U38031 (N_38031,N_30953,N_32419);
or U38032 (N_38032,N_33355,N_30793);
nand U38033 (N_38033,N_30928,N_30410);
or U38034 (N_38034,N_32649,N_34193);
and U38035 (N_38035,N_32622,N_34545);
nand U38036 (N_38036,N_33900,N_30541);
xor U38037 (N_38037,N_34419,N_30719);
nor U38038 (N_38038,N_30652,N_31597);
nand U38039 (N_38039,N_30987,N_32561);
or U38040 (N_38040,N_30414,N_31163);
xnor U38041 (N_38041,N_34691,N_31277);
nor U38042 (N_38042,N_33662,N_33162);
nand U38043 (N_38043,N_34513,N_30736);
and U38044 (N_38044,N_30734,N_34883);
xnor U38045 (N_38045,N_30161,N_34912);
nor U38046 (N_38046,N_30133,N_32338);
xnor U38047 (N_38047,N_30983,N_31106);
nor U38048 (N_38048,N_33603,N_32024);
nand U38049 (N_38049,N_33232,N_32473);
nand U38050 (N_38050,N_31229,N_30889);
xor U38051 (N_38051,N_31987,N_33026);
nor U38052 (N_38052,N_32848,N_34986);
nand U38053 (N_38053,N_31629,N_32223);
nand U38054 (N_38054,N_34276,N_31433);
nand U38055 (N_38055,N_33387,N_30431);
nor U38056 (N_38056,N_33799,N_32295);
xnor U38057 (N_38057,N_34034,N_33173);
xnor U38058 (N_38058,N_31620,N_31748);
or U38059 (N_38059,N_31757,N_33710);
nand U38060 (N_38060,N_33371,N_34480);
and U38061 (N_38061,N_33412,N_30462);
or U38062 (N_38062,N_32493,N_34982);
or U38063 (N_38063,N_31905,N_33554);
and U38064 (N_38064,N_30346,N_30612);
or U38065 (N_38065,N_33838,N_32355);
xor U38066 (N_38066,N_34017,N_31229);
and U38067 (N_38067,N_31287,N_32413);
nor U38068 (N_38068,N_32225,N_30512);
nand U38069 (N_38069,N_34676,N_30486);
and U38070 (N_38070,N_34038,N_30372);
xnor U38071 (N_38071,N_30909,N_34917);
nand U38072 (N_38072,N_33403,N_33303);
nand U38073 (N_38073,N_34422,N_31878);
nand U38074 (N_38074,N_31401,N_30109);
nor U38075 (N_38075,N_32908,N_33820);
xnor U38076 (N_38076,N_30696,N_31703);
and U38077 (N_38077,N_33744,N_34654);
nor U38078 (N_38078,N_32644,N_31941);
and U38079 (N_38079,N_33173,N_34701);
nor U38080 (N_38080,N_34239,N_34257);
xor U38081 (N_38081,N_30266,N_34056);
nor U38082 (N_38082,N_30215,N_30159);
nand U38083 (N_38083,N_32159,N_31066);
nor U38084 (N_38084,N_33399,N_32238);
nand U38085 (N_38085,N_33558,N_33889);
or U38086 (N_38086,N_33307,N_31161);
nand U38087 (N_38087,N_34004,N_34390);
and U38088 (N_38088,N_33386,N_34465);
or U38089 (N_38089,N_30533,N_30492);
and U38090 (N_38090,N_30582,N_34536);
or U38091 (N_38091,N_34752,N_33344);
nand U38092 (N_38092,N_34445,N_30103);
and U38093 (N_38093,N_31101,N_30573);
xor U38094 (N_38094,N_34100,N_32365);
or U38095 (N_38095,N_30396,N_32924);
or U38096 (N_38096,N_31786,N_34992);
or U38097 (N_38097,N_34238,N_30062);
and U38098 (N_38098,N_33318,N_33483);
or U38099 (N_38099,N_30113,N_30543);
xnor U38100 (N_38100,N_32804,N_34764);
nand U38101 (N_38101,N_30451,N_32491);
or U38102 (N_38102,N_32436,N_30315);
and U38103 (N_38103,N_32908,N_32995);
and U38104 (N_38104,N_32688,N_32645);
xor U38105 (N_38105,N_31259,N_33590);
and U38106 (N_38106,N_34460,N_30083);
nor U38107 (N_38107,N_30512,N_31584);
xor U38108 (N_38108,N_31652,N_33880);
or U38109 (N_38109,N_31862,N_30151);
xnor U38110 (N_38110,N_34316,N_33943);
nor U38111 (N_38111,N_32665,N_31477);
xnor U38112 (N_38112,N_33517,N_30761);
or U38113 (N_38113,N_32153,N_34230);
nor U38114 (N_38114,N_30666,N_33026);
xnor U38115 (N_38115,N_30175,N_30783);
nor U38116 (N_38116,N_33592,N_33265);
xnor U38117 (N_38117,N_30997,N_33076);
xnor U38118 (N_38118,N_30493,N_34929);
nor U38119 (N_38119,N_31490,N_31062);
nand U38120 (N_38120,N_30406,N_31784);
nand U38121 (N_38121,N_31263,N_33009);
or U38122 (N_38122,N_31784,N_31167);
or U38123 (N_38123,N_31435,N_34619);
nand U38124 (N_38124,N_30231,N_33177);
xor U38125 (N_38125,N_34342,N_31680);
or U38126 (N_38126,N_34199,N_34354);
nor U38127 (N_38127,N_31320,N_32312);
nor U38128 (N_38128,N_33775,N_31641);
nand U38129 (N_38129,N_30535,N_33031);
nand U38130 (N_38130,N_30279,N_33210);
nand U38131 (N_38131,N_32728,N_30538);
xor U38132 (N_38132,N_32434,N_33359);
xor U38133 (N_38133,N_30459,N_32196);
or U38134 (N_38134,N_34154,N_32977);
or U38135 (N_38135,N_30152,N_31612);
nor U38136 (N_38136,N_30234,N_34146);
nand U38137 (N_38137,N_34951,N_34447);
nand U38138 (N_38138,N_31553,N_34107);
nor U38139 (N_38139,N_32836,N_33670);
nand U38140 (N_38140,N_31622,N_30299);
nand U38141 (N_38141,N_34219,N_33578);
xor U38142 (N_38142,N_34016,N_30413);
nor U38143 (N_38143,N_30441,N_34202);
or U38144 (N_38144,N_33015,N_30725);
xor U38145 (N_38145,N_32988,N_32759);
nor U38146 (N_38146,N_33623,N_33576);
nor U38147 (N_38147,N_33517,N_31724);
nor U38148 (N_38148,N_34413,N_32878);
or U38149 (N_38149,N_34535,N_33584);
nor U38150 (N_38150,N_31997,N_30760);
xor U38151 (N_38151,N_33516,N_30732);
nor U38152 (N_38152,N_33617,N_30184);
xnor U38153 (N_38153,N_31087,N_33746);
xor U38154 (N_38154,N_33642,N_30572);
and U38155 (N_38155,N_33697,N_34708);
nor U38156 (N_38156,N_30765,N_34352);
xor U38157 (N_38157,N_32715,N_33931);
or U38158 (N_38158,N_31973,N_30326);
xor U38159 (N_38159,N_32967,N_34373);
and U38160 (N_38160,N_31897,N_30171);
or U38161 (N_38161,N_30920,N_30681);
xnor U38162 (N_38162,N_34593,N_33586);
xnor U38163 (N_38163,N_33060,N_32443);
and U38164 (N_38164,N_32260,N_33549);
and U38165 (N_38165,N_33468,N_32054);
or U38166 (N_38166,N_33841,N_30363);
xnor U38167 (N_38167,N_31774,N_33724);
or U38168 (N_38168,N_31988,N_34735);
xor U38169 (N_38169,N_34033,N_33048);
or U38170 (N_38170,N_32036,N_34854);
and U38171 (N_38171,N_33696,N_33225);
nor U38172 (N_38172,N_30307,N_33090);
and U38173 (N_38173,N_31443,N_34683);
nor U38174 (N_38174,N_31084,N_30699);
nor U38175 (N_38175,N_31389,N_32094);
xor U38176 (N_38176,N_34254,N_31612);
and U38177 (N_38177,N_31583,N_30141);
nor U38178 (N_38178,N_32473,N_33817);
nand U38179 (N_38179,N_31412,N_33762);
and U38180 (N_38180,N_32240,N_31513);
or U38181 (N_38181,N_34604,N_34299);
nor U38182 (N_38182,N_31940,N_32956);
xnor U38183 (N_38183,N_34662,N_34504);
or U38184 (N_38184,N_33724,N_34083);
and U38185 (N_38185,N_31890,N_31936);
xor U38186 (N_38186,N_33038,N_32487);
xor U38187 (N_38187,N_32236,N_31286);
nor U38188 (N_38188,N_33109,N_33647);
and U38189 (N_38189,N_32178,N_33466);
xor U38190 (N_38190,N_33992,N_32693);
or U38191 (N_38191,N_30746,N_32374);
or U38192 (N_38192,N_32485,N_33008);
nand U38193 (N_38193,N_32382,N_34020);
or U38194 (N_38194,N_30051,N_33056);
or U38195 (N_38195,N_32787,N_31543);
nor U38196 (N_38196,N_34953,N_33884);
nand U38197 (N_38197,N_31287,N_33930);
nor U38198 (N_38198,N_33207,N_33098);
and U38199 (N_38199,N_33424,N_31685);
xor U38200 (N_38200,N_34100,N_30999);
or U38201 (N_38201,N_31559,N_34318);
nor U38202 (N_38202,N_30473,N_30073);
and U38203 (N_38203,N_34875,N_32573);
nor U38204 (N_38204,N_31797,N_32244);
or U38205 (N_38205,N_30646,N_33301);
nor U38206 (N_38206,N_34939,N_33761);
nor U38207 (N_38207,N_34982,N_31775);
nand U38208 (N_38208,N_32939,N_32457);
and U38209 (N_38209,N_30271,N_33037);
nand U38210 (N_38210,N_33829,N_34124);
and U38211 (N_38211,N_30913,N_33864);
nor U38212 (N_38212,N_32664,N_30264);
nor U38213 (N_38213,N_32220,N_32016);
and U38214 (N_38214,N_34050,N_33250);
and U38215 (N_38215,N_30100,N_34146);
xor U38216 (N_38216,N_34492,N_32905);
nand U38217 (N_38217,N_34927,N_30382);
nand U38218 (N_38218,N_34776,N_33104);
or U38219 (N_38219,N_33890,N_34699);
or U38220 (N_38220,N_32174,N_33925);
xnor U38221 (N_38221,N_32371,N_34093);
nor U38222 (N_38222,N_30271,N_31199);
and U38223 (N_38223,N_32924,N_33674);
and U38224 (N_38224,N_34524,N_33042);
or U38225 (N_38225,N_31328,N_32109);
nor U38226 (N_38226,N_30661,N_34080);
or U38227 (N_38227,N_34007,N_34794);
or U38228 (N_38228,N_34227,N_30949);
nor U38229 (N_38229,N_31194,N_33927);
and U38230 (N_38230,N_32190,N_30323);
xor U38231 (N_38231,N_33028,N_30580);
or U38232 (N_38232,N_33259,N_33272);
nor U38233 (N_38233,N_34824,N_33205);
nand U38234 (N_38234,N_34366,N_34684);
nand U38235 (N_38235,N_32102,N_33336);
xor U38236 (N_38236,N_31059,N_33993);
nor U38237 (N_38237,N_31109,N_30266);
and U38238 (N_38238,N_32898,N_33342);
and U38239 (N_38239,N_33894,N_32614);
and U38240 (N_38240,N_31852,N_34243);
and U38241 (N_38241,N_30382,N_32926);
xor U38242 (N_38242,N_34325,N_30273);
or U38243 (N_38243,N_34186,N_31208);
xnor U38244 (N_38244,N_33013,N_32883);
or U38245 (N_38245,N_33627,N_31697);
nor U38246 (N_38246,N_30515,N_34155);
xor U38247 (N_38247,N_34988,N_34066);
or U38248 (N_38248,N_31567,N_31162);
nand U38249 (N_38249,N_32682,N_32392);
nor U38250 (N_38250,N_31796,N_30642);
and U38251 (N_38251,N_34967,N_33209);
or U38252 (N_38252,N_34083,N_32000);
and U38253 (N_38253,N_33845,N_31530);
or U38254 (N_38254,N_30023,N_30764);
nor U38255 (N_38255,N_31439,N_33207);
nor U38256 (N_38256,N_31134,N_32070);
and U38257 (N_38257,N_34777,N_32798);
xnor U38258 (N_38258,N_34296,N_30035);
or U38259 (N_38259,N_33810,N_32448);
and U38260 (N_38260,N_33451,N_30120);
and U38261 (N_38261,N_32232,N_34168);
nand U38262 (N_38262,N_32575,N_33296);
or U38263 (N_38263,N_30983,N_30064);
xor U38264 (N_38264,N_32444,N_31961);
and U38265 (N_38265,N_33890,N_30462);
xnor U38266 (N_38266,N_34507,N_30298);
or U38267 (N_38267,N_30224,N_32132);
and U38268 (N_38268,N_33323,N_31907);
nand U38269 (N_38269,N_31490,N_32790);
xnor U38270 (N_38270,N_34599,N_31892);
and U38271 (N_38271,N_30042,N_33762);
nand U38272 (N_38272,N_31219,N_30112);
nand U38273 (N_38273,N_30275,N_30715);
nor U38274 (N_38274,N_31488,N_32395);
and U38275 (N_38275,N_31027,N_34483);
nor U38276 (N_38276,N_31332,N_30674);
and U38277 (N_38277,N_33480,N_34107);
or U38278 (N_38278,N_33570,N_30241);
or U38279 (N_38279,N_32391,N_31796);
and U38280 (N_38280,N_34208,N_30382);
nand U38281 (N_38281,N_32559,N_33293);
and U38282 (N_38282,N_33123,N_33274);
or U38283 (N_38283,N_33270,N_31553);
xnor U38284 (N_38284,N_33527,N_34882);
xnor U38285 (N_38285,N_33177,N_34113);
and U38286 (N_38286,N_32433,N_34463);
nor U38287 (N_38287,N_33547,N_32802);
and U38288 (N_38288,N_33445,N_31012);
or U38289 (N_38289,N_30867,N_34805);
or U38290 (N_38290,N_31360,N_33619);
xnor U38291 (N_38291,N_33478,N_30046);
nor U38292 (N_38292,N_32024,N_34598);
and U38293 (N_38293,N_32820,N_34407);
nor U38294 (N_38294,N_31762,N_32036);
or U38295 (N_38295,N_32649,N_30855);
nor U38296 (N_38296,N_30973,N_34685);
xnor U38297 (N_38297,N_34451,N_34148);
nor U38298 (N_38298,N_34909,N_33132);
and U38299 (N_38299,N_34591,N_30537);
xor U38300 (N_38300,N_32311,N_33410);
nor U38301 (N_38301,N_33937,N_32008);
nand U38302 (N_38302,N_33875,N_32288);
xor U38303 (N_38303,N_33536,N_34873);
xor U38304 (N_38304,N_31646,N_34801);
nand U38305 (N_38305,N_31684,N_30430);
xor U38306 (N_38306,N_32370,N_30658);
nor U38307 (N_38307,N_34081,N_30829);
and U38308 (N_38308,N_33742,N_32702);
and U38309 (N_38309,N_31059,N_34486);
and U38310 (N_38310,N_31680,N_30527);
or U38311 (N_38311,N_32711,N_33065);
nand U38312 (N_38312,N_30568,N_30899);
and U38313 (N_38313,N_32463,N_34354);
nand U38314 (N_38314,N_33363,N_32554);
xor U38315 (N_38315,N_30035,N_34221);
nand U38316 (N_38316,N_30321,N_32147);
nand U38317 (N_38317,N_32022,N_32119);
nand U38318 (N_38318,N_31475,N_30353);
or U38319 (N_38319,N_33687,N_34820);
nand U38320 (N_38320,N_30366,N_34686);
xnor U38321 (N_38321,N_30981,N_33140);
or U38322 (N_38322,N_32521,N_31347);
nor U38323 (N_38323,N_32398,N_33587);
and U38324 (N_38324,N_34878,N_30433);
nand U38325 (N_38325,N_32279,N_33875);
or U38326 (N_38326,N_31646,N_31419);
nand U38327 (N_38327,N_34157,N_34110);
nand U38328 (N_38328,N_32423,N_31813);
nand U38329 (N_38329,N_33421,N_30923);
nor U38330 (N_38330,N_31470,N_31935);
xor U38331 (N_38331,N_30038,N_33148);
xor U38332 (N_38332,N_33752,N_31578);
and U38333 (N_38333,N_30691,N_32164);
and U38334 (N_38334,N_30950,N_33916);
xnor U38335 (N_38335,N_30825,N_32091);
or U38336 (N_38336,N_32367,N_33724);
and U38337 (N_38337,N_34073,N_32953);
xor U38338 (N_38338,N_30715,N_31530);
and U38339 (N_38339,N_30052,N_30049);
or U38340 (N_38340,N_34210,N_30050);
nor U38341 (N_38341,N_33276,N_32801);
xnor U38342 (N_38342,N_32930,N_34266);
xor U38343 (N_38343,N_34735,N_34176);
or U38344 (N_38344,N_32899,N_33023);
nand U38345 (N_38345,N_30228,N_30369);
xor U38346 (N_38346,N_33879,N_33572);
xnor U38347 (N_38347,N_34487,N_32361);
or U38348 (N_38348,N_33133,N_33125);
or U38349 (N_38349,N_31605,N_33770);
nor U38350 (N_38350,N_33848,N_31117);
nand U38351 (N_38351,N_34462,N_34416);
nand U38352 (N_38352,N_33651,N_34723);
xnor U38353 (N_38353,N_30198,N_34969);
and U38354 (N_38354,N_33848,N_30909);
or U38355 (N_38355,N_31263,N_34548);
nor U38356 (N_38356,N_34533,N_33163);
nand U38357 (N_38357,N_31716,N_33163);
and U38358 (N_38358,N_32135,N_33590);
or U38359 (N_38359,N_34615,N_33717);
nor U38360 (N_38360,N_34390,N_30102);
nand U38361 (N_38361,N_33011,N_30272);
or U38362 (N_38362,N_31579,N_32146);
xnor U38363 (N_38363,N_32098,N_34073);
nand U38364 (N_38364,N_33463,N_34786);
and U38365 (N_38365,N_32099,N_32011);
or U38366 (N_38366,N_30584,N_30087);
or U38367 (N_38367,N_34950,N_31080);
nand U38368 (N_38368,N_33466,N_33225);
xor U38369 (N_38369,N_34404,N_33792);
nand U38370 (N_38370,N_30331,N_34968);
nand U38371 (N_38371,N_32125,N_33079);
and U38372 (N_38372,N_33832,N_34812);
xor U38373 (N_38373,N_33524,N_30899);
nand U38374 (N_38374,N_32146,N_31165);
nand U38375 (N_38375,N_33613,N_31156);
nand U38376 (N_38376,N_34111,N_33682);
or U38377 (N_38377,N_31649,N_31073);
or U38378 (N_38378,N_34265,N_30511);
nand U38379 (N_38379,N_31299,N_31611);
nand U38380 (N_38380,N_31140,N_30545);
xor U38381 (N_38381,N_34138,N_31834);
nor U38382 (N_38382,N_34688,N_33894);
xor U38383 (N_38383,N_32959,N_32669);
and U38384 (N_38384,N_30640,N_34594);
xnor U38385 (N_38385,N_32940,N_30136);
xnor U38386 (N_38386,N_33542,N_34399);
or U38387 (N_38387,N_31715,N_33798);
nand U38388 (N_38388,N_32590,N_30449);
nor U38389 (N_38389,N_31009,N_32715);
xor U38390 (N_38390,N_31553,N_32970);
nand U38391 (N_38391,N_32786,N_34091);
nand U38392 (N_38392,N_31003,N_33962);
nor U38393 (N_38393,N_34291,N_30380);
xnor U38394 (N_38394,N_32604,N_32385);
and U38395 (N_38395,N_34247,N_34192);
nor U38396 (N_38396,N_34549,N_31789);
and U38397 (N_38397,N_34592,N_33274);
nor U38398 (N_38398,N_33741,N_32204);
xnor U38399 (N_38399,N_34468,N_34435);
and U38400 (N_38400,N_33137,N_30355);
nand U38401 (N_38401,N_33788,N_33266);
nor U38402 (N_38402,N_34217,N_31680);
xnor U38403 (N_38403,N_31792,N_34007);
nor U38404 (N_38404,N_34199,N_30497);
nor U38405 (N_38405,N_33721,N_34534);
xor U38406 (N_38406,N_33343,N_33912);
and U38407 (N_38407,N_30502,N_34788);
and U38408 (N_38408,N_34099,N_30063);
xnor U38409 (N_38409,N_32211,N_34158);
and U38410 (N_38410,N_33046,N_31663);
and U38411 (N_38411,N_33615,N_33482);
nor U38412 (N_38412,N_33230,N_32409);
xor U38413 (N_38413,N_30612,N_34836);
xor U38414 (N_38414,N_30555,N_34542);
nor U38415 (N_38415,N_34043,N_32755);
and U38416 (N_38416,N_33097,N_33431);
or U38417 (N_38417,N_33787,N_30441);
nor U38418 (N_38418,N_30333,N_30972);
xor U38419 (N_38419,N_31089,N_30340);
or U38420 (N_38420,N_31738,N_31906);
and U38421 (N_38421,N_32384,N_34521);
and U38422 (N_38422,N_30056,N_31591);
nor U38423 (N_38423,N_32941,N_31142);
xnor U38424 (N_38424,N_31224,N_30882);
xor U38425 (N_38425,N_30540,N_31804);
nand U38426 (N_38426,N_32982,N_33749);
or U38427 (N_38427,N_30401,N_30584);
and U38428 (N_38428,N_30478,N_31165);
or U38429 (N_38429,N_32506,N_34775);
and U38430 (N_38430,N_31577,N_31626);
xnor U38431 (N_38431,N_32089,N_34043);
and U38432 (N_38432,N_32793,N_30722);
nor U38433 (N_38433,N_34123,N_31556);
and U38434 (N_38434,N_34597,N_34882);
or U38435 (N_38435,N_34941,N_34235);
nor U38436 (N_38436,N_32604,N_30461);
or U38437 (N_38437,N_34280,N_31091);
nand U38438 (N_38438,N_33354,N_30283);
nand U38439 (N_38439,N_34193,N_33331);
and U38440 (N_38440,N_32599,N_32281);
and U38441 (N_38441,N_34135,N_32495);
nand U38442 (N_38442,N_31403,N_32952);
or U38443 (N_38443,N_33280,N_32685);
or U38444 (N_38444,N_34955,N_30426);
nor U38445 (N_38445,N_30039,N_33561);
or U38446 (N_38446,N_31243,N_30805);
or U38447 (N_38447,N_33530,N_30945);
nand U38448 (N_38448,N_31553,N_30105);
and U38449 (N_38449,N_32724,N_34564);
nand U38450 (N_38450,N_30316,N_33498);
and U38451 (N_38451,N_34335,N_31634);
xnor U38452 (N_38452,N_33917,N_34316);
xnor U38453 (N_38453,N_32686,N_32612);
and U38454 (N_38454,N_32034,N_31070);
nand U38455 (N_38455,N_33930,N_34511);
nand U38456 (N_38456,N_31981,N_30987);
or U38457 (N_38457,N_33246,N_33788);
and U38458 (N_38458,N_31772,N_33810);
xnor U38459 (N_38459,N_31215,N_33175);
or U38460 (N_38460,N_34732,N_34583);
nor U38461 (N_38461,N_34308,N_33687);
nor U38462 (N_38462,N_30438,N_32283);
nor U38463 (N_38463,N_30106,N_32608);
nor U38464 (N_38464,N_32564,N_31484);
xor U38465 (N_38465,N_31457,N_30102);
or U38466 (N_38466,N_34612,N_33568);
nand U38467 (N_38467,N_32903,N_34074);
or U38468 (N_38468,N_33636,N_34707);
nor U38469 (N_38469,N_34992,N_32129);
nand U38470 (N_38470,N_33961,N_32873);
xor U38471 (N_38471,N_31710,N_31097);
nand U38472 (N_38472,N_31349,N_31249);
xnor U38473 (N_38473,N_32245,N_30383);
nand U38474 (N_38474,N_34082,N_32728);
nor U38475 (N_38475,N_30222,N_33772);
nand U38476 (N_38476,N_32630,N_33096);
and U38477 (N_38477,N_32349,N_32257);
nor U38478 (N_38478,N_34950,N_30432);
or U38479 (N_38479,N_34932,N_30224);
xor U38480 (N_38480,N_33269,N_32792);
and U38481 (N_38481,N_32486,N_33026);
and U38482 (N_38482,N_33648,N_33348);
xnor U38483 (N_38483,N_34807,N_33663);
or U38484 (N_38484,N_32520,N_32908);
nand U38485 (N_38485,N_32040,N_32082);
nand U38486 (N_38486,N_34084,N_30724);
and U38487 (N_38487,N_30677,N_30520);
xor U38488 (N_38488,N_31683,N_34905);
nand U38489 (N_38489,N_34498,N_31822);
nand U38490 (N_38490,N_32360,N_30409);
or U38491 (N_38491,N_33832,N_31554);
and U38492 (N_38492,N_33321,N_34053);
nand U38493 (N_38493,N_32385,N_33201);
nor U38494 (N_38494,N_34603,N_30540);
or U38495 (N_38495,N_31871,N_32104);
nand U38496 (N_38496,N_31652,N_30363);
nor U38497 (N_38497,N_33715,N_30014);
xnor U38498 (N_38498,N_31154,N_32246);
nor U38499 (N_38499,N_34542,N_31668);
xnor U38500 (N_38500,N_33864,N_31946);
nor U38501 (N_38501,N_33850,N_33442);
or U38502 (N_38502,N_34926,N_31368);
nand U38503 (N_38503,N_32871,N_33216);
xnor U38504 (N_38504,N_34855,N_32298);
nor U38505 (N_38505,N_31659,N_34564);
or U38506 (N_38506,N_34763,N_33695);
nor U38507 (N_38507,N_33067,N_30787);
nor U38508 (N_38508,N_34691,N_31582);
nand U38509 (N_38509,N_30885,N_30575);
and U38510 (N_38510,N_33242,N_30585);
nor U38511 (N_38511,N_31262,N_33427);
xor U38512 (N_38512,N_31006,N_34209);
and U38513 (N_38513,N_31470,N_33388);
xor U38514 (N_38514,N_34747,N_32852);
xor U38515 (N_38515,N_33523,N_31565);
xor U38516 (N_38516,N_34200,N_34802);
nand U38517 (N_38517,N_32103,N_32681);
and U38518 (N_38518,N_34652,N_34697);
xnor U38519 (N_38519,N_33034,N_34285);
nand U38520 (N_38520,N_33260,N_31677);
xnor U38521 (N_38521,N_33201,N_30114);
nand U38522 (N_38522,N_31225,N_34015);
nor U38523 (N_38523,N_33574,N_32212);
nor U38524 (N_38524,N_31277,N_32739);
nor U38525 (N_38525,N_33953,N_31016);
or U38526 (N_38526,N_34780,N_32372);
nor U38527 (N_38527,N_34683,N_30058);
or U38528 (N_38528,N_32852,N_30670);
or U38529 (N_38529,N_34502,N_30918);
or U38530 (N_38530,N_33725,N_32244);
nand U38531 (N_38531,N_34337,N_33880);
nand U38532 (N_38532,N_33676,N_34376);
nand U38533 (N_38533,N_32830,N_30494);
and U38534 (N_38534,N_33417,N_31551);
and U38535 (N_38535,N_32875,N_34000);
or U38536 (N_38536,N_30198,N_30980);
nand U38537 (N_38537,N_33749,N_31213);
xor U38538 (N_38538,N_33999,N_33745);
and U38539 (N_38539,N_34914,N_31120);
nor U38540 (N_38540,N_32582,N_31747);
and U38541 (N_38541,N_34435,N_33492);
and U38542 (N_38542,N_31494,N_31273);
nand U38543 (N_38543,N_32226,N_31481);
and U38544 (N_38544,N_32821,N_32968);
xor U38545 (N_38545,N_31052,N_32747);
and U38546 (N_38546,N_34749,N_31515);
nor U38547 (N_38547,N_30732,N_32443);
and U38548 (N_38548,N_30367,N_34852);
nand U38549 (N_38549,N_31223,N_31719);
nor U38550 (N_38550,N_31747,N_31816);
or U38551 (N_38551,N_31118,N_30115);
or U38552 (N_38552,N_30980,N_32565);
xnor U38553 (N_38553,N_34601,N_32388);
xnor U38554 (N_38554,N_33710,N_32364);
and U38555 (N_38555,N_32715,N_30953);
nand U38556 (N_38556,N_32561,N_30318);
or U38557 (N_38557,N_30612,N_34591);
nand U38558 (N_38558,N_31884,N_32013);
xnor U38559 (N_38559,N_32259,N_34740);
xor U38560 (N_38560,N_31158,N_31551);
nand U38561 (N_38561,N_30956,N_33311);
nand U38562 (N_38562,N_33069,N_32227);
nand U38563 (N_38563,N_32375,N_33145);
and U38564 (N_38564,N_34133,N_30172);
nand U38565 (N_38565,N_33244,N_34397);
xnor U38566 (N_38566,N_34226,N_32909);
and U38567 (N_38567,N_31444,N_34637);
xor U38568 (N_38568,N_33006,N_30758);
or U38569 (N_38569,N_33670,N_31104);
and U38570 (N_38570,N_33510,N_34957);
or U38571 (N_38571,N_33978,N_33732);
or U38572 (N_38572,N_30075,N_33818);
and U38573 (N_38573,N_34008,N_34930);
nor U38574 (N_38574,N_31050,N_33154);
or U38575 (N_38575,N_32359,N_34136);
nand U38576 (N_38576,N_30324,N_30975);
or U38577 (N_38577,N_32713,N_33837);
and U38578 (N_38578,N_31452,N_34223);
and U38579 (N_38579,N_32748,N_32431);
nand U38580 (N_38580,N_34319,N_30512);
or U38581 (N_38581,N_31530,N_32343);
or U38582 (N_38582,N_32707,N_33571);
xor U38583 (N_38583,N_31487,N_34133);
or U38584 (N_38584,N_34244,N_32860);
and U38585 (N_38585,N_30745,N_33369);
nor U38586 (N_38586,N_31964,N_32704);
or U38587 (N_38587,N_34531,N_31701);
xor U38588 (N_38588,N_34089,N_31188);
or U38589 (N_38589,N_31897,N_34875);
and U38590 (N_38590,N_32491,N_31520);
nor U38591 (N_38591,N_31841,N_31053);
or U38592 (N_38592,N_30274,N_31141);
and U38593 (N_38593,N_33382,N_31244);
and U38594 (N_38594,N_33246,N_33811);
nor U38595 (N_38595,N_32768,N_31274);
or U38596 (N_38596,N_33947,N_32796);
nor U38597 (N_38597,N_33183,N_30721);
xor U38598 (N_38598,N_30281,N_31729);
xor U38599 (N_38599,N_33651,N_31427);
and U38600 (N_38600,N_30843,N_30391);
and U38601 (N_38601,N_30041,N_31835);
nand U38602 (N_38602,N_31205,N_33320);
xor U38603 (N_38603,N_34870,N_34919);
nor U38604 (N_38604,N_34736,N_30616);
or U38605 (N_38605,N_33570,N_33774);
and U38606 (N_38606,N_32157,N_30710);
and U38607 (N_38607,N_34637,N_30360);
nand U38608 (N_38608,N_34390,N_30407);
or U38609 (N_38609,N_30089,N_30536);
xor U38610 (N_38610,N_34544,N_33560);
or U38611 (N_38611,N_31102,N_30378);
nor U38612 (N_38612,N_31677,N_34195);
xnor U38613 (N_38613,N_32240,N_34666);
xnor U38614 (N_38614,N_32853,N_31201);
and U38615 (N_38615,N_32496,N_32137);
and U38616 (N_38616,N_33666,N_33513);
nand U38617 (N_38617,N_33836,N_34474);
or U38618 (N_38618,N_33574,N_33961);
xor U38619 (N_38619,N_34171,N_32092);
or U38620 (N_38620,N_33462,N_34279);
and U38621 (N_38621,N_30766,N_33219);
and U38622 (N_38622,N_33922,N_31607);
nand U38623 (N_38623,N_32578,N_33719);
and U38624 (N_38624,N_33828,N_33969);
or U38625 (N_38625,N_31645,N_30813);
and U38626 (N_38626,N_31684,N_34634);
xnor U38627 (N_38627,N_34789,N_34821);
or U38628 (N_38628,N_33570,N_34888);
or U38629 (N_38629,N_33146,N_30081);
nor U38630 (N_38630,N_32224,N_34836);
nand U38631 (N_38631,N_30873,N_32539);
or U38632 (N_38632,N_30472,N_34449);
and U38633 (N_38633,N_33135,N_34844);
nand U38634 (N_38634,N_34552,N_33817);
or U38635 (N_38635,N_31322,N_30714);
nor U38636 (N_38636,N_33475,N_32333);
nor U38637 (N_38637,N_34862,N_34010);
nand U38638 (N_38638,N_32260,N_30959);
xor U38639 (N_38639,N_31986,N_32091);
nor U38640 (N_38640,N_30444,N_30453);
nor U38641 (N_38641,N_31510,N_33582);
nor U38642 (N_38642,N_33708,N_30019);
xnor U38643 (N_38643,N_30637,N_33431);
and U38644 (N_38644,N_30925,N_32948);
xor U38645 (N_38645,N_30271,N_30803);
and U38646 (N_38646,N_31777,N_34760);
or U38647 (N_38647,N_31958,N_31892);
xor U38648 (N_38648,N_33676,N_32580);
nand U38649 (N_38649,N_34786,N_32685);
xor U38650 (N_38650,N_32301,N_33807);
or U38651 (N_38651,N_34698,N_33425);
nand U38652 (N_38652,N_31342,N_34904);
nor U38653 (N_38653,N_30952,N_30727);
or U38654 (N_38654,N_34865,N_31161);
and U38655 (N_38655,N_32271,N_34267);
nand U38656 (N_38656,N_32950,N_32914);
xor U38657 (N_38657,N_34650,N_32407);
xnor U38658 (N_38658,N_30804,N_30499);
or U38659 (N_38659,N_34388,N_31211);
xnor U38660 (N_38660,N_31628,N_34833);
xnor U38661 (N_38661,N_32888,N_30010);
nor U38662 (N_38662,N_33113,N_31067);
or U38663 (N_38663,N_33442,N_32262);
and U38664 (N_38664,N_33552,N_33992);
nor U38665 (N_38665,N_31564,N_30421);
and U38666 (N_38666,N_30873,N_31415);
nor U38667 (N_38667,N_33547,N_32860);
xnor U38668 (N_38668,N_31655,N_32547);
xnor U38669 (N_38669,N_33400,N_33628);
or U38670 (N_38670,N_33519,N_33207);
xor U38671 (N_38671,N_34733,N_33864);
nor U38672 (N_38672,N_31666,N_34161);
and U38673 (N_38673,N_32860,N_31153);
or U38674 (N_38674,N_30704,N_33830);
or U38675 (N_38675,N_32274,N_30531);
and U38676 (N_38676,N_30033,N_32987);
nand U38677 (N_38677,N_31198,N_32602);
and U38678 (N_38678,N_32949,N_32306);
nor U38679 (N_38679,N_34176,N_34466);
nor U38680 (N_38680,N_32967,N_33788);
or U38681 (N_38681,N_31391,N_32065);
and U38682 (N_38682,N_34768,N_33226);
or U38683 (N_38683,N_34696,N_32117);
nor U38684 (N_38684,N_32310,N_31998);
nand U38685 (N_38685,N_33373,N_31924);
xor U38686 (N_38686,N_30604,N_31362);
or U38687 (N_38687,N_32725,N_33344);
xor U38688 (N_38688,N_32558,N_33607);
nor U38689 (N_38689,N_31453,N_33423);
and U38690 (N_38690,N_31000,N_31738);
nor U38691 (N_38691,N_31607,N_31504);
nor U38692 (N_38692,N_33100,N_34160);
or U38693 (N_38693,N_34628,N_30201);
nand U38694 (N_38694,N_33167,N_34891);
xor U38695 (N_38695,N_32710,N_32111);
nand U38696 (N_38696,N_34808,N_34273);
xor U38697 (N_38697,N_32144,N_31279);
nand U38698 (N_38698,N_31040,N_31566);
or U38699 (N_38699,N_31915,N_33129);
nor U38700 (N_38700,N_34073,N_30376);
and U38701 (N_38701,N_31145,N_31405);
xor U38702 (N_38702,N_34204,N_34955);
nor U38703 (N_38703,N_32236,N_33138);
nand U38704 (N_38704,N_34100,N_30288);
nand U38705 (N_38705,N_30108,N_34484);
or U38706 (N_38706,N_31440,N_31930);
nand U38707 (N_38707,N_33885,N_33221);
nand U38708 (N_38708,N_34788,N_32946);
and U38709 (N_38709,N_31423,N_30975);
nor U38710 (N_38710,N_31981,N_31397);
or U38711 (N_38711,N_33106,N_33432);
or U38712 (N_38712,N_33960,N_33424);
nand U38713 (N_38713,N_30891,N_30112);
nor U38714 (N_38714,N_34829,N_31390);
xnor U38715 (N_38715,N_34030,N_31447);
xnor U38716 (N_38716,N_32189,N_33876);
nand U38717 (N_38717,N_30633,N_33294);
xnor U38718 (N_38718,N_31708,N_30569);
or U38719 (N_38719,N_33345,N_31786);
nand U38720 (N_38720,N_33743,N_31875);
nand U38721 (N_38721,N_33903,N_30727);
or U38722 (N_38722,N_31388,N_33285);
nor U38723 (N_38723,N_33575,N_32998);
or U38724 (N_38724,N_31023,N_30466);
nor U38725 (N_38725,N_30630,N_34797);
nor U38726 (N_38726,N_33621,N_31000);
or U38727 (N_38727,N_31111,N_31998);
or U38728 (N_38728,N_30398,N_33105);
nor U38729 (N_38729,N_33172,N_33097);
or U38730 (N_38730,N_32533,N_30623);
xor U38731 (N_38731,N_32506,N_32962);
or U38732 (N_38732,N_32812,N_30784);
xnor U38733 (N_38733,N_31023,N_31306);
xnor U38734 (N_38734,N_31395,N_31286);
nor U38735 (N_38735,N_31031,N_33131);
or U38736 (N_38736,N_33662,N_34225);
xnor U38737 (N_38737,N_34429,N_30116);
and U38738 (N_38738,N_32060,N_33754);
or U38739 (N_38739,N_30224,N_33491);
nand U38740 (N_38740,N_34552,N_32865);
or U38741 (N_38741,N_30688,N_31495);
or U38742 (N_38742,N_30781,N_33152);
xnor U38743 (N_38743,N_33743,N_33407);
nand U38744 (N_38744,N_33479,N_33492);
or U38745 (N_38745,N_31323,N_31338);
nor U38746 (N_38746,N_33947,N_32412);
xnor U38747 (N_38747,N_30228,N_31466);
nor U38748 (N_38748,N_30259,N_33433);
and U38749 (N_38749,N_32143,N_34882);
or U38750 (N_38750,N_32759,N_32293);
nor U38751 (N_38751,N_30695,N_31546);
or U38752 (N_38752,N_33779,N_30642);
or U38753 (N_38753,N_33022,N_33157);
nand U38754 (N_38754,N_32862,N_33411);
nand U38755 (N_38755,N_34845,N_34374);
nand U38756 (N_38756,N_30396,N_32546);
xor U38757 (N_38757,N_34610,N_31258);
nand U38758 (N_38758,N_31325,N_33159);
nand U38759 (N_38759,N_33894,N_30234);
or U38760 (N_38760,N_30015,N_33666);
nand U38761 (N_38761,N_32164,N_30564);
and U38762 (N_38762,N_30061,N_33051);
and U38763 (N_38763,N_34700,N_34272);
and U38764 (N_38764,N_30674,N_34469);
and U38765 (N_38765,N_33427,N_33980);
nor U38766 (N_38766,N_33660,N_32349);
xnor U38767 (N_38767,N_31577,N_34394);
nand U38768 (N_38768,N_30761,N_33083);
nand U38769 (N_38769,N_34852,N_31584);
xor U38770 (N_38770,N_31536,N_33153);
xor U38771 (N_38771,N_31222,N_33003);
xnor U38772 (N_38772,N_30112,N_30340);
xor U38773 (N_38773,N_31036,N_34310);
xor U38774 (N_38774,N_33874,N_32074);
or U38775 (N_38775,N_31299,N_31834);
xor U38776 (N_38776,N_30367,N_32517);
nor U38777 (N_38777,N_34760,N_33342);
or U38778 (N_38778,N_30037,N_33844);
nand U38779 (N_38779,N_33686,N_32257);
nor U38780 (N_38780,N_30040,N_31438);
nor U38781 (N_38781,N_31859,N_31348);
and U38782 (N_38782,N_33369,N_30307);
and U38783 (N_38783,N_31885,N_33232);
xor U38784 (N_38784,N_34732,N_33858);
or U38785 (N_38785,N_33465,N_30488);
or U38786 (N_38786,N_34804,N_31922);
nor U38787 (N_38787,N_31436,N_33598);
or U38788 (N_38788,N_33661,N_31616);
nand U38789 (N_38789,N_31756,N_34931);
nor U38790 (N_38790,N_31331,N_30448);
nand U38791 (N_38791,N_30628,N_31358);
xnor U38792 (N_38792,N_32383,N_33024);
nor U38793 (N_38793,N_33024,N_34257);
and U38794 (N_38794,N_34972,N_32090);
or U38795 (N_38795,N_34030,N_33161);
nor U38796 (N_38796,N_31150,N_30750);
or U38797 (N_38797,N_33388,N_30872);
xnor U38798 (N_38798,N_31102,N_34875);
and U38799 (N_38799,N_34746,N_30323);
or U38800 (N_38800,N_31870,N_31217);
and U38801 (N_38801,N_30934,N_34656);
and U38802 (N_38802,N_32144,N_32381);
nand U38803 (N_38803,N_34634,N_32709);
nor U38804 (N_38804,N_34881,N_30609);
nand U38805 (N_38805,N_32988,N_31524);
or U38806 (N_38806,N_33683,N_32406);
and U38807 (N_38807,N_30862,N_33752);
nor U38808 (N_38808,N_31671,N_30804);
and U38809 (N_38809,N_34542,N_30481);
nand U38810 (N_38810,N_33701,N_33222);
or U38811 (N_38811,N_30224,N_32615);
nor U38812 (N_38812,N_32170,N_34457);
xnor U38813 (N_38813,N_32672,N_34382);
nand U38814 (N_38814,N_30917,N_34718);
or U38815 (N_38815,N_34040,N_34780);
nor U38816 (N_38816,N_31596,N_32676);
and U38817 (N_38817,N_30318,N_30441);
and U38818 (N_38818,N_34332,N_32812);
nand U38819 (N_38819,N_32093,N_32198);
and U38820 (N_38820,N_32904,N_31453);
xor U38821 (N_38821,N_34627,N_34624);
nand U38822 (N_38822,N_32965,N_32669);
nand U38823 (N_38823,N_32445,N_30824);
xnor U38824 (N_38824,N_30788,N_34730);
or U38825 (N_38825,N_30852,N_32334);
nand U38826 (N_38826,N_32920,N_34999);
or U38827 (N_38827,N_30005,N_32802);
xor U38828 (N_38828,N_30626,N_32667);
and U38829 (N_38829,N_33750,N_31178);
and U38830 (N_38830,N_33297,N_31783);
or U38831 (N_38831,N_33995,N_34192);
nor U38832 (N_38832,N_32105,N_32276);
or U38833 (N_38833,N_34020,N_31909);
and U38834 (N_38834,N_31683,N_32738);
nor U38835 (N_38835,N_31961,N_33491);
or U38836 (N_38836,N_30845,N_31061);
nor U38837 (N_38837,N_31800,N_32504);
nand U38838 (N_38838,N_33460,N_34174);
and U38839 (N_38839,N_31014,N_32545);
or U38840 (N_38840,N_33201,N_30079);
nand U38841 (N_38841,N_31178,N_32781);
nor U38842 (N_38842,N_33466,N_30296);
and U38843 (N_38843,N_32244,N_30899);
xor U38844 (N_38844,N_31387,N_33844);
nor U38845 (N_38845,N_32071,N_33502);
nor U38846 (N_38846,N_30482,N_33455);
or U38847 (N_38847,N_31338,N_30932);
nand U38848 (N_38848,N_32431,N_32055);
nand U38849 (N_38849,N_34432,N_31986);
or U38850 (N_38850,N_30600,N_31381);
or U38851 (N_38851,N_30122,N_33269);
or U38852 (N_38852,N_34871,N_33122);
and U38853 (N_38853,N_30389,N_31319);
nand U38854 (N_38854,N_31618,N_31240);
nor U38855 (N_38855,N_33958,N_34378);
nand U38856 (N_38856,N_34637,N_31282);
nor U38857 (N_38857,N_31751,N_34181);
nand U38858 (N_38858,N_34000,N_33815);
or U38859 (N_38859,N_34956,N_34313);
xor U38860 (N_38860,N_31704,N_32399);
nor U38861 (N_38861,N_33168,N_32766);
nand U38862 (N_38862,N_32018,N_33945);
and U38863 (N_38863,N_31180,N_32736);
xnor U38864 (N_38864,N_30877,N_30114);
xnor U38865 (N_38865,N_32952,N_34331);
and U38866 (N_38866,N_32330,N_33573);
or U38867 (N_38867,N_34365,N_30845);
nor U38868 (N_38868,N_30053,N_30769);
nand U38869 (N_38869,N_30094,N_32126);
xor U38870 (N_38870,N_34481,N_34465);
nand U38871 (N_38871,N_31232,N_31085);
and U38872 (N_38872,N_31142,N_31836);
or U38873 (N_38873,N_34119,N_34031);
nand U38874 (N_38874,N_33120,N_31630);
or U38875 (N_38875,N_34775,N_34175);
nor U38876 (N_38876,N_33446,N_30402);
xnor U38877 (N_38877,N_32524,N_34604);
xnor U38878 (N_38878,N_33822,N_33071);
xnor U38879 (N_38879,N_31994,N_30013);
xnor U38880 (N_38880,N_32014,N_31455);
and U38881 (N_38881,N_33230,N_30243);
xor U38882 (N_38882,N_34560,N_30223);
nor U38883 (N_38883,N_33511,N_34964);
and U38884 (N_38884,N_33258,N_30059);
nand U38885 (N_38885,N_34143,N_31829);
nor U38886 (N_38886,N_34363,N_32058);
or U38887 (N_38887,N_32548,N_31289);
xnor U38888 (N_38888,N_32642,N_32416);
and U38889 (N_38889,N_34420,N_31565);
and U38890 (N_38890,N_30403,N_33069);
xnor U38891 (N_38891,N_34274,N_30733);
or U38892 (N_38892,N_34876,N_32026);
nand U38893 (N_38893,N_30149,N_31972);
nand U38894 (N_38894,N_32519,N_34741);
nor U38895 (N_38895,N_31567,N_33785);
nand U38896 (N_38896,N_34657,N_32124);
and U38897 (N_38897,N_32017,N_33013);
and U38898 (N_38898,N_33176,N_34539);
or U38899 (N_38899,N_34971,N_31245);
and U38900 (N_38900,N_31993,N_34858);
xor U38901 (N_38901,N_32697,N_34171);
nand U38902 (N_38902,N_32842,N_34198);
or U38903 (N_38903,N_30375,N_32507);
xnor U38904 (N_38904,N_30240,N_30806);
xnor U38905 (N_38905,N_30236,N_33673);
nor U38906 (N_38906,N_34174,N_32714);
and U38907 (N_38907,N_33854,N_30843);
nand U38908 (N_38908,N_30303,N_30559);
and U38909 (N_38909,N_34285,N_32933);
nand U38910 (N_38910,N_33763,N_34113);
or U38911 (N_38911,N_34485,N_34701);
nor U38912 (N_38912,N_30241,N_34118);
xnor U38913 (N_38913,N_31869,N_30594);
or U38914 (N_38914,N_33791,N_30222);
and U38915 (N_38915,N_34201,N_30408);
nand U38916 (N_38916,N_34909,N_34725);
nor U38917 (N_38917,N_33429,N_34318);
and U38918 (N_38918,N_30290,N_30727);
xor U38919 (N_38919,N_31828,N_33241);
nand U38920 (N_38920,N_31414,N_33340);
xnor U38921 (N_38921,N_31605,N_30573);
or U38922 (N_38922,N_30743,N_34115);
nand U38923 (N_38923,N_33350,N_31301);
or U38924 (N_38924,N_31032,N_31502);
nand U38925 (N_38925,N_30938,N_33558);
xnor U38926 (N_38926,N_31583,N_33994);
nand U38927 (N_38927,N_34648,N_30859);
nand U38928 (N_38928,N_33009,N_30691);
xor U38929 (N_38929,N_32872,N_30291);
nor U38930 (N_38930,N_33861,N_30241);
or U38931 (N_38931,N_30175,N_30409);
or U38932 (N_38932,N_32002,N_32850);
nand U38933 (N_38933,N_31158,N_33868);
nand U38934 (N_38934,N_31578,N_31114);
and U38935 (N_38935,N_33031,N_30796);
nand U38936 (N_38936,N_33664,N_30858);
and U38937 (N_38937,N_30202,N_32628);
xor U38938 (N_38938,N_34606,N_31786);
or U38939 (N_38939,N_30047,N_32973);
nor U38940 (N_38940,N_34598,N_32429);
or U38941 (N_38941,N_30191,N_32905);
and U38942 (N_38942,N_33556,N_31637);
and U38943 (N_38943,N_32898,N_34899);
and U38944 (N_38944,N_34547,N_31107);
nand U38945 (N_38945,N_32742,N_31143);
or U38946 (N_38946,N_32418,N_33710);
nand U38947 (N_38947,N_30327,N_33160);
or U38948 (N_38948,N_30214,N_33935);
xor U38949 (N_38949,N_31091,N_32214);
nand U38950 (N_38950,N_32608,N_34312);
nor U38951 (N_38951,N_32964,N_31177);
nand U38952 (N_38952,N_34384,N_34661);
and U38953 (N_38953,N_30488,N_30353);
nand U38954 (N_38954,N_32500,N_33851);
nor U38955 (N_38955,N_30580,N_33312);
or U38956 (N_38956,N_31287,N_34635);
nand U38957 (N_38957,N_34103,N_30490);
nor U38958 (N_38958,N_30054,N_30805);
nand U38959 (N_38959,N_31761,N_33864);
nand U38960 (N_38960,N_31423,N_32407);
nor U38961 (N_38961,N_31191,N_30690);
xnor U38962 (N_38962,N_32434,N_32407);
nand U38963 (N_38963,N_32499,N_34471);
and U38964 (N_38964,N_31929,N_33015);
or U38965 (N_38965,N_34582,N_32440);
or U38966 (N_38966,N_32461,N_31866);
and U38967 (N_38967,N_32123,N_30202);
or U38968 (N_38968,N_32749,N_33142);
xor U38969 (N_38969,N_33533,N_32351);
nand U38970 (N_38970,N_33346,N_31848);
or U38971 (N_38971,N_34999,N_34614);
nor U38972 (N_38972,N_34437,N_32981);
and U38973 (N_38973,N_32718,N_31734);
or U38974 (N_38974,N_30817,N_34883);
or U38975 (N_38975,N_32270,N_31847);
nor U38976 (N_38976,N_33578,N_30904);
and U38977 (N_38977,N_31587,N_30610);
and U38978 (N_38978,N_31889,N_31605);
or U38979 (N_38979,N_34556,N_33173);
xor U38980 (N_38980,N_30367,N_32450);
or U38981 (N_38981,N_32445,N_32631);
nand U38982 (N_38982,N_32065,N_32570);
nor U38983 (N_38983,N_31167,N_31251);
xor U38984 (N_38984,N_30272,N_33493);
nor U38985 (N_38985,N_31159,N_34200);
nor U38986 (N_38986,N_30123,N_33931);
or U38987 (N_38987,N_30438,N_32410);
or U38988 (N_38988,N_30693,N_32766);
and U38989 (N_38989,N_33147,N_31835);
or U38990 (N_38990,N_32336,N_32760);
nand U38991 (N_38991,N_31312,N_33733);
and U38992 (N_38992,N_31526,N_30906);
nor U38993 (N_38993,N_31711,N_31108);
nand U38994 (N_38994,N_33961,N_30776);
nor U38995 (N_38995,N_31952,N_30453);
nor U38996 (N_38996,N_32738,N_30874);
or U38997 (N_38997,N_31028,N_32636);
nor U38998 (N_38998,N_32787,N_33502);
nand U38999 (N_38999,N_33400,N_31201);
xor U39000 (N_39000,N_34010,N_30159);
nor U39001 (N_39001,N_32193,N_30272);
nor U39002 (N_39002,N_32390,N_34656);
nand U39003 (N_39003,N_31466,N_34976);
xnor U39004 (N_39004,N_31799,N_34372);
nand U39005 (N_39005,N_31134,N_32357);
nor U39006 (N_39006,N_32399,N_33314);
or U39007 (N_39007,N_33605,N_33158);
nand U39008 (N_39008,N_31346,N_33689);
or U39009 (N_39009,N_33660,N_31130);
or U39010 (N_39010,N_33319,N_33110);
nor U39011 (N_39011,N_34269,N_30039);
nand U39012 (N_39012,N_32015,N_32394);
xor U39013 (N_39013,N_33258,N_34734);
and U39014 (N_39014,N_34936,N_32488);
and U39015 (N_39015,N_31793,N_34153);
xor U39016 (N_39016,N_34040,N_30249);
nand U39017 (N_39017,N_34268,N_34192);
nor U39018 (N_39018,N_33072,N_31742);
or U39019 (N_39019,N_32896,N_34721);
and U39020 (N_39020,N_31761,N_33117);
xnor U39021 (N_39021,N_34365,N_31854);
nor U39022 (N_39022,N_31560,N_33189);
xor U39023 (N_39023,N_34373,N_32494);
and U39024 (N_39024,N_33569,N_33539);
nor U39025 (N_39025,N_30783,N_33036);
or U39026 (N_39026,N_34484,N_32926);
nand U39027 (N_39027,N_31405,N_30733);
or U39028 (N_39028,N_31322,N_32136);
or U39029 (N_39029,N_32102,N_31025);
or U39030 (N_39030,N_31009,N_32109);
and U39031 (N_39031,N_30953,N_34377);
nand U39032 (N_39032,N_31152,N_34609);
and U39033 (N_39033,N_34516,N_33479);
xor U39034 (N_39034,N_31857,N_30249);
or U39035 (N_39035,N_33317,N_33704);
and U39036 (N_39036,N_34801,N_34930);
nand U39037 (N_39037,N_30389,N_31232);
or U39038 (N_39038,N_33525,N_33614);
nor U39039 (N_39039,N_31355,N_31277);
nand U39040 (N_39040,N_34754,N_34580);
or U39041 (N_39041,N_32835,N_34415);
or U39042 (N_39042,N_30097,N_34889);
nor U39043 (N_39043,N_33915,N_31569);
or U39044 (N_39044,N_31446,N_34113);
and U39045 (N_39045,N_34580,N_30987);
nor U39046 (N_39046,N_31032,N_34999);
nor U39047 (N_39047,N_30206,N_31726);
nand U39048 (N_39048,N_33249,N_30794);
nand U39049 (N_39049,N_32579,N_30865);
and U39050 (N_39050,N_34744,N_30865);
and U39051 (N_39051,N_33389,N_32013);
nor U39052 (N_39052,N_34320,N_32813);
nand U39053 (N_39053,N_31109,N_34916);
nor U39054 (N_39054,N_33092,N_32048);
nor U39055 (N_39055,N_32984,N_33875);
and U39056 (N_39056,N_32188,N_31582);
or U39057 (N_39057,N_30526,N_31869);
xor U39058 (N_39058,N_34565,N_34100);
or U39059 (N_39059,N_30472,N_33448);
and U39060 (N_39060,N_33781,N_30074);
nor U39061 (N_39061,N_34446,N_34221);
xor U39062 (N_39062,N_33001,N_32110);
nor U39063 (N_39063,N_30803,N_34688);
nand U39064 (N_39064,N_32970,N_31074);
nor U39065 (N_39065,N_34708,N_30375);
or U39066 (N_39066,N_33595,N_30599);
and U39067 (N_39067,N_33131,N_31849);
xor U39068 (N_39068,N_33738,N_31088);
and U39069 (N_39069,N_32329,N_30504);
nand U39070 (N_39070,N_30727,N_31218);
and U39071 (N_39071,N_33996,N_31552);
and U39072 (N_39072,N_34358,N_31397);
xnor U39073 (N_39073,N_30518,N_30962);
or U39074 (N_39074,N_31085,N_33013);
nor U39075 (N_39075,N_31716,N_33412);
or U39076 (N_39076,N_31790,N_34115);
or U39077 (N_39077,N_30446,N_32021);
nand U39078 (N_39078,N_34637,N_34959);
and U39079 (N_39079,N_33038,N_32067);
nor U39080 (N_39080,N_30752,N_32974);
or U39081 (N_39081,N_32567,N_31066);
and U39082 (N_39082,N_34430,N_32773);
nor U39083 (N_39083,N_31002,N_31893);
nand U39084 (N_39084,N_31541,N_34405);
and U39085 (N_39085,N_31244,N_32298);
nand U39086 (N_39086,N_31907,N_30464);
or U39087 (N_39087,N_31180,N_34040);
and U39088 (N_39088,N_33149,N_31009);
xnor U39089 (N_39089,N_32611,N_30131);
or U39090 (N_39090,N_34716,N_34758);
xnor U39091 (N_39091,N_31784,N_33676);
and U39092 (N_39092,N_33686,N_31860);
and U39093 (N_39093,N_32023,N_31907);
xor U39094 (N_39094,N_30788,N_33768);
nand U39095 (N_39095,N_34604,N_31540);
nor U39096 (N_39096,N_34371,N_32409);
and U39097 (N_39097,N_32471,N_30460);
or U39098 (N_39098,N_31048,N_30739);
nor U39099 (N_39099,N_30648,N_34729);
xor U39100 (N_39100,N_34781,N_32751);
nor U39101 (N_39101,N_32782,N_32616);
or U39102 (N_39102,N_32080,N_33133);
nor U39103 (N_39103,N_30730,N_32230);
nor U39104 (N_39104,N_34444,N_32473);
nor U39105 (N_39105,N_31921,N_33137);
nand U39106 (N_39106,N_33133,N_30926);
xor U39107 (N_39107,N_34264,N_30471);
nand U39108 (N_39108,N_30902,N_33004);
nand U39109 (N_39109,N_30080,N_33635);
and U39110 (N_39110,N_32186,N_33108);
nand U39111 (N_39111,N_32208,N_31350);
or U39112 (N_39112,N_34820,N_31124);
nor U39113 (N_39113,N_30025,N_32051);
nand U39114 (N_39114,N_30039,N_30959);
xor U39115 (N_39115,N_33739,N_32542);
nand U39116 (N_39116,N_30474,N_33679);
xnor U39117 (N_39117,N_31028,N_30696);
nand U39118 (N_39118,N_34333,N_30864);
xnor U39119 (N_39119,N_34254,N_32038);
nand U39120 (N_39120,N_31820,N_34604);
nor U39121 (N_39121,N_30495,N_34786);
nand U39122 (N_39122,N_32871,N_33726);
or U39123 (N_39123,N_33931,N_31562);
xor U39124 (N_39124,N_34022,N_30952);
nor U39125 (N_39125,N_30119,N_31650);
and U39126 (N_39126,N_34110,N_31245);
nand U39127 (N_39127,N_30200,N_34309);
or U39128 (N_39128,N_32958,N_33414);
nand U39129 (N_39129,N_30268,N_30610);
nor U39130 (N_39130,N_33001,N_32864);
nand U39131 (N_39131,N_32749,N_34364);
or U39132 (N_39132,N_30371,N_34977);
xor U39133 (N_39133,N_30432,N_33577);
and U39134 (N_39134,N_30223,N_30822);
and U39135 (N_39135,N_33485,N_34623);
nor U39136 (N_39136,N_31888,N_30549);
nand U39137 (N_39137,N_30264,N_32632);
nor U39138 (N_39138,N_33455,N_30125);
nand U39139 (N_39139,N_31025,N_34036);
and U39140 (N_39140,N_32743,N_34413);
nor U39141 (N_39141,N_31485,N_33666);
nand U39142 (N_39142,N_30496,N_34922);
and U39143 (N_39143,N_31629,N_32490);
and U39144 (N_39144,N_33976,N_32574);
and U39145 (N_39145,N_30599,N_32252);
nor U39146 (N_39146,N_31279,N_31644);
xor U39147 (N_39147,N_30791,N_30903);
nor U39148 (N_39148,N_34785,N_32190);
nand U39149 (N_39149,N_31794,N_30092);
or U39150 (N_39150,N_32186,N_33356);
xnor U39151 (N_39151,N_34352,N_31814);
or U39152 (N_39152,N_32045,N_33970);
and U39153 (N_39153,N_33619,N_30795);
and U39154 (N_39154,N_31729,N_30383);
and U39155 (N_39155,N_30340,N_33922);
nand U39156 (N_39156,N_33026,N_32911);
and U39157 (N_39157,N_33417,N_31557);
nor U39158 (N_39158,N_30662,N_33747);
or U39159 (N_39159,N_34406,N_30917);
xnor U39160 (N_39160,N_34349,N_32100);
and U39161 (N_39161,N_32402,N_31461);
nand U39162 (N_39162,N_32378,N_30370);
or U39163 (N_39163,N_33748,N_31770);
xor U39164 (N_39164,N_33990,N_32916);
nand U39165 (N_39165,N_31906,N_32735);
or U39166 (N_39166,N_34784,N_30968);
nor U39167 (N_39167,N_34483,N_33099);
or U39168 (N_39168,N_31863,N_34440);
or U39169 (N_39169,N_33913,N_33725);
nor U39170 (N_39170,N_30122,N_30397);
or U39171 (N_39171,N_34874,N_30363);
nand U39172 (N_39172,N_33998,N_34983);
nand U39173 (N_39173,N_30299,N_34776);
nand U39174 (N_39174,N_32815,N_30065);
nand U39175 (N_39175,N_34163,N_34783);
xnor U39176 (N_39176,N_30187,N_34568);
and U39177 (N_39177,N_33629,N_33525);
or U39178 (N_39178,N_33524,N_32296);
xnor U39179 (N_39179,N_30700,N_30447);
or U39180 (N_39180,N_32258,N_31315);
nand U39181 (N_39181,N_33413,N_32322);
nand U39182 (N_39182,N_34230,N_33008);
or U39183 (N_39183,N_33156,N_33487);
nor U39184 (N_39184,N_31472,N_34394);
nor U39185 (N_39185,N_30428,N_32683);
nor U39186 (N_39186,N_30980,N_34773);
xnor U39187 (N_39187,N_32280,N_32276);
and U39188 (N_39188,N_32048,N_34098);
nor U39189 (N_39189,N_33968,N_34447);
nor U39190 (N_39190,N_32340,N_34286);
nand U39191 (N_39191,N_34672,N_30038);
and U39192 (N_39192,N_33136,N_30627);
and U39193 (N_39193,N_32036,N_34203);
nand U39194 (N_39194,N_33861,N_34052);
nor U39195 (N_39195,N_33657,N_31224);
and U39196 (N_39196,N_34582,N_30207);
xnor U39197 (N_39197,N_34217,N_32533);
and U39198 (N_39198,N_31015,N_33154);
nand U39199 (N_39199,N_34451,N_34089);
nand U39200 (N_39200,N_32904,N_32490);
xor U39201 (N_39201,N_30488,N_31957);
nand U39202 (N_39202,N_32877,N_30837);
xnor U39203 (N_39203,N_33397,N_32915);
or U39204 (N_39204,N_30492,N_32932);
xnor U39205 (N_39205,N_34720,N_31600);
and U39206 (N_39206,N_33324,N_31821);
nor U39207 (N_39207,N_32401,N_34843);
nor U39208 (N_39208,N_30903,N_33806);
nand U39209 (N_39209,N_31611,N_33928);
or U39210 (N_39210,N_32132,N_34472);
or U39211 (N_39211,N_30044,N_30969);
nand U39212 (N_39212,N_30806,N_31633);
or U39213 (N_39213,N_30863,N_31219);
xor U39214 (N_39214,N_30225,N_31822);
or U39215 (N_39215,N_32502,N_31718);
xnor U39216 (N_39216,N_32859,N_33836);
nor U39217 (N_39217,N_30979,N_33392);
nor U39218 (N_39218,N_33805,N_33108);
or U39219 (N_39219,N_31421,N_30627);
or U39220 (N_39220,N_31868,N_30558);
or U39221 (N_39221,N_32965,N_32925);
xnor U39222 (N_39222,N_31565,N_33052);
nand U39223 (N_39223,N_33971,N_32632);
or U39224 (N_39224,N_30443,N_31814);
or U39225 (N_39225,N_31961,N_33674);
nand U39226 (N_39226,N_34111,N_34151);
xor U39227 (N_39227,N_31834,N_33497);
xnor U39228 (N_39228,N_30435,N_31175);
and U39229 (N_39229,N_30789,N_31965);
or U39230 (N_39230,N_30920,N_30304);
xnor U39231 (N_39231,N_34265,N_31323);
nor U39232 (N_39232,N_33028,N_34210);
nand U39233 (N_39233,N_31427,N_34443);
and U39234 (N_39234,N_32989,N_30294);
nor U39235 (N_39235,N_33830,N_31393);
xnor U39236 (N_39236,N_34531,N_32519);
nand U39237 (N_39237,N_31351,N_31541);
or U39238 (N_39238,N_33109,N_30086);
nor U39239 (N_39239,N_34973,N_34806);
nor U39240 (N_39240,N_31832,N_32026);
xor U39241 (N_39241,N_32520,N_31991);
xor U39242 (N_39242,N_34483,N_34855);
and U39243 (N_39243,N_34624,N_30670);
nand U39244 (N_39244,N_32775,N_31249);
and U39245 (N_39245,N_34770,N_31650);
and U39246 (N_39246,N_30554,N_31503);
and U39247 (N_39247,N_32119,N_33725);
and U39248 (N_39248,N_33689,N_31281);
xor U39249 (N_39249,N_33837,N_34343);
nor U39250 (N_39250,N_33992,N_34336);
xor U39251 (N_39251,N_32554,N_31891);
and U39252 (N_39252,N_31619,N_34180);
or U39253 (N_39253,N_32176,N_31177);
nand U39254 (N_39254,N_30515,N_34900);
or U39255 (N_39255,N_30830,N_31422);
xor U39256 (N_39256,N_31910,N_30301);
nand U39257 (N_39257,N_31437,N_30095);
and U39258 (N_39258,N_30416,N_31010);
or U39259 (N_39259,N_32425,N_30679);
or U39260 (N_39260,N_32395,N_30807);
nand U39261 (N_39261,N_30452,N_33315);
xor U39262 (N_39262,N_32709,N_32780);
nand U39263 (N_39263,N_30803,N_31579);
or U39264 (N_39264,N_32306,N_31517);
nand U39265 (N_39265,N_33549,N_32650);
and U39266 (N_39266,N_34680,N_31801);
xnor U39267 (N_39267,N_33338,N_31155);
or U39268 (N_39268,N_31086,N_31533);
nor U39269 (N_39269,N_33952,N_33041);
nand U39270 (N_39270,N_33892,N_34254);
and U39271 (N_39271,N_31690,N_32089);
and U39272 (N_39272,N_34609,N_34269);
xor U39273 (N_39273,N_34039,N_33270);
and U39274 (N_39274,N_32753,N_33988);
nor U39275 (N_39275,N_34779,N_32103);
nand U39276 (N_39276,N_33546,N_30819);
xnor U39277 (N_39277,N_32275,N_33267);
or U39278 (N_39278,N_31162,N_33078);
nor U39279 (N_39279,N_31137,N_34122);
and U39280 (N_39280,N_30873,N_31262);
and U39281 (N_39281,N_34390,N_31224);
or U39282 (N_39282,N_31240,N_33069);
and U39283 (N_39283,N_33675,N_31669);
nand U39284 (N_39284,N_34415,N_33584);
nand U39285 (N_39285,N_33348,N_31087);
or U39286 (N_39286,N_34354,N_32330);
nand U39287 (N_39287,N_30987,N_30615);
nand U39288 (N_39288,N_32772,N_32800);
nand U39289 (N_39289,N_31149,N_34563);
or U39290 (N_39290,N_32526,N_32587);
or U39291 (N_39291,N_30115,N_30896);
or U39292 (N_39292,N_30685,N_34074);
and U39293 (N_39293,N_32339,N_33470);
xnor U39294 (N_39294,N_31312,N_30997);
and U39295 (N_39295,N_32883,N_33358);
or U39296 (N_39296,N_34911,N_34889);
or U39297 (N_39297,N_33203,N_34548);
nor U39298 (N_39298,N_34251,N_31454);
and U39299 (N_39299,N_32922,N_32554);
nor U39300 (N_39300,N_32825,N_33498);
nand U39301 (N_39301,N_33956,N_34205);
nand U39302 (N_39302,N_31767,N_31618);
and U39303 (N_39303,N_32003,N_33936);
nand U39304 (N_39304,N_30609,N_33505);
nor U39305 (N_39305,N_30189,N_33810);
and U39306 (N_39306,N_33751,N_34663);
and U39307 (N_39307,N_34660,N_32617);
xor U39308 (N_39308,N_31235,N_33505);
or U39309 (N_39309,N_34184,N_32034);
and U39310 (N_39310,N_34359,N_32388);
and U39311 (N_39311,N_32871,N_31515);
nand U39312 (N_39312,N_30388,N_30569);
or U39313 (N_39313,N_30897,N_31227);
nand U39314 (N_39314,N_33877,N_33023);
nor U39315 (N_39315,N_31992,N_32351);
xor U39316 (N_39316,N_30171,N_31061);
nand U39317 (N_39317,N_33660,N_32929);
xor U39318 (N_39318,N_33399,N_31296);
nor U39319 (N_39319,N_32098,N_33572);
or U39320 (N_39320,N_31633,N_31517);
nand U39321 (N_39321,N_32359,N_32134);
nand U39322 (N_39322,N_33818,N_31439);
and U39323 (N_39323,N_32502,N_34003);
or U39324 (N_39324,N_31327,N_34123);
nand U39325 (N_39325,N_30136,N_30054);
xor U39326 (N_39326,N_30960,N_30316);
xnor U39327 (N_39327,N_30702,N_30120);
nor U39328 (N_39328,N_33225,N_31310);
xnor U39329 (N_39329,N_31366,N_30631);
nand U39330 (N_39330,N_33186,N_30804);
or U39331 (N_39331,N_33295,N_34949);
or U39332 (N_39332,N_31022,N_34011);
nand U39333 (N_39333,N_30553,N_31115);
xnor U39334 (N_39334,N_33653,N_30305);
and U39335 (N_39335,N_30947,N_30666);
xor U39336 (N_39336,N_33863,N_30319);
or U39337 (N_39337,N_32566,N_31931);
nand U39338 (N_39338,N_34880,N_34729);
nand U39339 (N_39339,N_30127,N_34823);
and U39340 (N_39340,N_31123,N_32352);
xnor U39341 (N_39341,N_30739,N_34540);
nand U39342 (N_39342,N_31273,N_32020);
or U39343 (N_39343,N_30439,N_33205);
nand U39344 (N_39344,N_30668,N_32145);
or U39345 (N_39345,N_30103,N_32403);
and U39346 (N_39346,N_33729,N_30547);
or U39347 (N_39347,N_31939,N_31497);
and U39348 (N_39348,N_30823,N_33168);
or U39349 (N_39349,N_34298,N_34160);
or U39350 (N_39350,N_33786,N_33286);
xor U39351 (N_39351,N_33732,N_33924);
or U39352 (N_39352,N_31540,N_32286);
and U39353 (N_39353,N_31200,N_30132);
nor U39354 (N_39354,N_32092,N_32742);
or U39355 (N_39355,N_31342,N_30810);
and U39356 (N_39356,N_33078,N_30473);
nand U39357 (N_39357,N_32338,N_34653);
xnor U39358 (N_39358,N_30942,N_32450);
and U39359 (N_39359,N_31749,N_33325);
nand U39360 (N_39360,N_34639,N_33878);
nand U39361 (N_39361,N_33836,N_31702);
nand U39362 (N_39362,N_34212,N_31788);
nor U39363 (N_39363,N_32813,N_32056);
xor U39364 (N_39364,N_34323,N_30579);
nor U39365 (N_39365,N_30389,N_30934);
nand U39366 (N_39366,N_32781,N_32940);
nor U39367 (N_39367,N_31719,N_30536);
nor U39368 (N_39368,N_32762,N_34152);
nor U39369 (N_39369,N_31524,N_30650);
xor U39370 (N_39370,N_30057,N_31941);
xor U39371 (N_39371,N_34795,N_32983);
xnor U39372 (N_39372,N_34120,N_33240);
nor U39373 (N_39373,N_30954,N_31821);
and U39374 (N_39374,N_34164,N_34376);
and U39375 (N_39375,N_34556,N_33725);
xnor U39376 (N_39376,N_31005,N_33109);
nor U39377 (N_39377,N_31574,N_33502);
nand U39378 (N_39378,N_32871,N_32999);
or U39379 (N_39379,N_34141,N_31942);
xnor U39380 (N_39380,N_33566,N_34330);
and U39381 (N_39381,N_31799,N_31844);
nand U39382 (N_39382,N_31185,N_33142);
or U39383 (N_39383,N_31065,N_32763);
xnor U39384 (N_39384,N_30828,N_32278);
or U39385 (N_39385,N_31307,N_30123);
xor U39386 (N_39386,N_34549,N_33463);
and U39387 (N_39387,N_33691,N_30937);
nand U39388 (N_39388,N_30499,N_33266);
xor U39389 (N_39389,N_31211,N_31314);
or U39390 (N_39390,N_32991,N_30541);
nand U39391 (N_39391,N_31768,N_31488);
nand U39392 (N_39392,N_30654,N_31023);
nor U39393 (N_39393,N_30152,N_33416);
and U39394 (N_39394,N_34979,N_30682);
or U39395 (N_39395,N_34229,N_34801);
nand U39396 (N_39396,N_33560,N_32605);
and U39397 (N_39397,N_31129,N_31328);
or U39398 (N_39398,N_34653,N_33736);
nor U39399 (N_39399,N_34651,N_30444);
xnor U39400 (N_39400,N_30330,N_30948);
nand U39401 (N_39401,N_31809,N_32980);
xnor U39402 (N_39402,N_33272,N_30609);
nor U39403 (N_39403,N_31744,N_31070);
xnor U39404 (N_39404,N_34718,N_33691);
nor U39405 (N_39405,N_31665,N_31530);
nand U39406 (N_39406,N_33444,N_30588);
xnor U39407 (N_39407,N_31070,N_32393);
xnor U39408 (N_39408,N_33761,N_31841);
and U39409 (N_39409,N_33412,N_30641);
nand U39410 (N_39410,N_31504,N_32412);
and U39411 (N_39411,N_31234,N_33593);
nor U39412 (N_39412,N_30063,N_32945);
and U39413 (N_39413,N_33636,N_31230);
or U39414 (N_39414,N_34286,N_32039);
nand U39415 (N_39415,N_31473,N_34281);
and U39416 (N_39416,N_30042,N_31897);
nand U39417 (N_39417,N_33956,N_32994);
nand U39418 (N_39418,N_34049,N_30829);
xor U39419 (N_39419,N_32647,N_31362);
and U39420 (N_39420,N_34391,N_33054);
nand U39421 (N_39421,N_34412,N_31673);
xor U39422 (N_39422,N_30591,N_33115);
and U39423 (N_39423,N_32667,N_32453);
or U39424 (N_39424,N_32704,N_32421);
nor U39425 (N_39425,N_30508,N_31399);
nor U39426 (N_39426,N_31074,N_34171);
or U39427 (N_39427,N_30563,N_31142);
and U39428 (N_39428,N_33710,N_34224);
nor U39429 (N_39429,N_31265,N_34312);
or U39430 (N_39430,N_31117,N_34912);
nor U39431 (N_39431,N_34874,N_33761);
xnor U39432 (N_39432,N_33630,N_34288);
and U39433 (N_39433,N_30385,N_30691);
and U39434 (N_39434,N_32570,N_34395);
and U39435 (N_39435,N_33925,N_31843);
xor U39436 (N_39436,N_32538,N_34831);
nor U39437 (N_39437,N_31614,N_31637);
and U39438 (N_39438,N_31675,N_30148);
and U39439 (N_39439,N_30484,N_33953);
nand U39440 (N_39440,N_32276,N_30325);
nor U39441 (N_39441,N_30658,N_32244);
xor U39442 (N_39442,N_33205,N_32479);
nor U39443 (N_39443,N_30910,N_32369);
nor U39444 (N_39444,N_31766,N_30055);
or U39445 (N_39445,N_31828,N_32277);
and U39446 (N_39446,N_32367,N_32739);
and U39447 (N_39447,N_33963,N_31232);
nand U39448 (N_39448,N_32230,N_32408);
xor U39449 (N_39449,N_30493,N_33563);
xnor U39450 (N_39450,N_33911,N_33873);
nor U39451 (N_39451,N_32019,N_31802);
nor U39452 (N_39452,N_34811,N_31326);
nor U39453 (N_39453,N_31365,N_31448);
nor U39454 (N_39454,N_33911,N_30637);
or U39455 (N_39455,N_31561,N_32961);
nand U39456 (N_39456,N_31862,N_31269);
nor U39457 (N_39457,N_34147,N_30648);
and U39458 (N_39458,N_30683,N_33541);
nand U39459 (N_39459,N_33372,N_34937);
and U39460 (N_39460,N_33090,N_32904);
nor U39461 (N_39461,N_34293,N_34694);
nor U39462 (N_39462,N_32539,N_31473);
or U39463 (N_39463,N_32886,N_31181);
nor U39464 (N_39464,N_31528,N_32003);
and U39465 (N_39465,N_31301,N_30212);
nor U39466 (N_39466,N_30161,N_33607);
and U39467 (N_39467,N_34630,N_31781);
nand U39468 (N_39468,N_33259,N_30135);
and U39469 (N_39469,N_30080,N_33817);
xor U39470 (N_39470,N_34300,N_34015);
and U39471 (N_39471,N_33036,N_30695);
nand U39472 (N_39472,N_33441,N_30159);
or U39473 (N_39473,N_31379,N_32130);
or U39474 (N_39474,N_31309,N_31720);
nand U39475 (N_39475,N_33615,N_31011);
nor U39476 (N_39476,N_34842,N_30886);
nor U39477 (N_39477,N_30119,N_32096);
or U39478 (N_39478,N_32035,N_30495);
xnor U39479 (N_39479,N_33104,N_33768);
nand U39480 (N_39480,N_30266,N_30789);
and U39481 (N_39481,N_30888,N_31405);
or U39482 (N_39482,N_31940,N_33180);
nor U39483 (N_39483,N_32917,N_34351);
or U39484 (N_39484,N_33331,N_31207);
nand U39485 (N_39485,N_34532,N_31993);
nand U39486 (N_39486,N_30027,N_33700);
xor U39487 (N_39487,N_34926,N_32868);
and U39488 (N_39488,N_32370,N_33380);
nor U39489 (N_39489,N_31310,N_32086);
nor U39490 (N_39490,N_31645,N_34104);
and U39491 (N_39491,N_31970,N_30983);
nor U39492 (N_39492,N_30019,N_32209);
or U39493 (N_39493,N_33141,N_34321);
xor U39494 (N_39494,N_34662,N_32260);
nor U39495 (N_39495,N_31610,N_33257);
and U39496 (N_39496,N_33626,N_31320);
xnor U39497 (N_39497,N_33223,N_32136);
nor U39498 (N_39498,N_30835,N_33712);
xor U39499 (N_39499,N_31994,N_31181);
nor U39500 (N_39500,N_31615,N_30594);
and U39501 (N_39501,N_30460,N_33090);
or U39502 (N_39502,N_33895,N_32470);
xor U39503 (N_39503,N_32626,N_34882);
nor U39504 (N_39504,N_33273,N_34633);
nor U39505 (N_39505,N_32222,N_33855);
nand U39506 (N_39506,N_32632,N_34806);
nand U39507 (N_39507,N_32866,N_32216);
xnor U39508 (N_39508,N_34515,N_31903);
xor U39509 (N_39509,N_33379,N_32779);
and U39510 (N_39510,N_33367,N_34851);
and U39511 (N_39511,N_31687,N_34774);
xnor U39512 (N_39512,N_30695,N_32936);
or U39513 (N_39513,N_34175,N_32069);
nand U39514 (N_39514,N_32707,N_30117);
nand U39515 (N_39515,N_31124,N_30405);
or U39516 (N_39516,N_33465,N_32378);
and U39517 (N_39517,N_33419,N_30548);
nand U39518 (N_39518,N_33929,N_31526);
nand U39519 (N_39519,N_33007,N_31313);
and U39520 (N_39520,N_32824,N_31368);
nand U39521 (N_39521,N_34258,N_34937);
and U39522 (N_39522,N_32792,N_32166);
and U39523 (N_39523,N_33110,N_30311);
or U39524 (N_39524,N_31753,N_34988);
or U39525 (N_39525,N_32430,N_30238);
xor U39526 (N_39526,N_30943,N_30374);
xor U39527 (N_39527,N_32816,N_31860);
xnor U39528 (N_39528,N_33127,N_33532);
or U39529 (N_39529,N_30146,N_30580);
xnor U39530 (N_39530,N_30044,N_33501);
or U39531 (N_39531,N_31046,N_30897);
or U39532 (N_39532,N_34591,N_30646);
xnor U39533 (N_39533,N_31600,N_32659);
or U39534 (N_39534,N_32936,N_34478);
nand U39535 (N_39535,N_31966,N_33122);
nand U39536 (N_39536,N_32739,N_34141);
xnor U39537 (N_39537,N_32394,N_31489);
and U39538 (N_39538,N_31055,N_34752);
or U39539 (N_39539,N_31957,N_31244);
and U39540 (N_39540,N_30245,N_32914);
and U39541 (N_39541,N_32796,N_33321);
xnor U39542 (N_39542,N_34808,N_32717);
nand U39543 (N_39543,N_31376,N_30762);
and U39544 (N_39544,N_31780,N_34891);
nor U39545 (N_39545,N_34960,N_30959);
nor U39546 (N_39546,N_34608,N_31219);
and U39547 (N_39547,N_34812,N_30417);
and U39548 (N_39548,N_31417,N_32253);
nor U39549 (N_39549,N_33690,N_33921);
xor U39550 (N_39550,N_30765,N_33847);
nand U39551 (N_39551,N_32214,N_33358);
xor U39552 (N_39552,N_32585,N_30160);
and U39553 (N_39553,N_34174,N_30854);
nand U39554 (N_39554,N_33623,N_31579);
nor U39555 (N_39555,N_34162,N_30247);
and U39556 (N_39556,N_34325,N_34011);
nor U39557 (N_39557,N_32007,N_32894);
nor U39558 (N_39558,N_33895,N_30608);
nand U39559 (N_39559,N_30494,N_33987);
xnor U39560 (N_39560,N_31969,N_32387);
xor U39561 (N_39561,N_31648,N_34481);
nand U39562 (N_39562,N_33278,N_31925);
and U39563 (N_39563,N_30625,N_34235);
nand U39564 (N_39564,N_33493,N_34890);
nand U39565 (N_39565,N_31434,N_33773);
xnor U39566 (N_39566,N_34838,N_34686);
and U39567 (N_39567,N_33022,N_31151);
or U39568 (N_39568,N_34313,N_33184);
nand U39569 (N_39569,N_31533,N_33710);
nor U39570 (N_39570,N_33300,N_34522);
xnor U39571 (N_39571,N_30649,N_30424);
nor U39572 (N_39572,N_34668,N_32747);
and U39573 (N_39573,N_33608,N_30315);
xnor U39574 (N_39574,N_34988,N_31940);
nor U39575 (N_39575,N_32680,N_33546);
or U39576 (N_39576,N_34502,N_32919);
xnor U39577 (N_39577,N_32716,N_34720);
nor U39578 (N_39578,N_30786,N_31967);
or U39579 (N_39579,N_33494,N_31153);
and U39580 (N_39580,N_31389,N_32303);
xnor U39581 (N_39581,N_30740,N_30781);
xnor U39582 (N_39582,N_30282,N_30640);
and U39583 (N_39583,N_33479,N_33956);
and U39584 (N_39584,N_32551,N_33203);
xor U39585 (N_39585,N_34850,N_30255);
nor U39586 (N_39586,N_32856,N_32931);
xnor U39587 (N_39587,N_30920,N_31287);
nand U39588 (N_39588,N_33773,N_31056);
nand U39589 (N_39589,N_31438,N_34586);
nor U39590 (N_39590,N_33953,N_33170);
or U39591 (N_39591,N_30454,N_34670);
xnor U39592 (N_39592,N_31354,N_33168);
nor U39593 (N_39593,N_31762,N_33844);
xnor U39594 (N_39594,N_30517,N_30924);
nand U39595 (N_39595,N_33924,N_32504);
or U39596 (N_39596,N_33629,N_31993);
nor U39597 (N_39597,N_32258,N_32981);
and U39598 (N_39598,N_31664,N_34619);
nand U39599 (N_39599,N_33126,N_30066);
nor U39600 (N_39600,N_31016,N_30517);
nor U39601 (N_39601,N_32997,N_33518);
or U39602 (N_39602,N_34271,N_34200);
or U39603 (N_39603,N_33938,N_31929);
nand U39604 (N_39604,N_33107,N_32185);
nand U39605 (N_39605,N_30967,N_32118);
nor U39606 (N_39606,N_34051,N_32129);
nor U39607 (N_39607,N_34778,N_32447);
or U39608 (N_39608,N_32543,N_34526);
xor U39609 (N_39609,N_30901,N_33088);
nand U39610 (N_39610,N_33122,N_30071);
nor U39611 (N_39611,N_33810,N_31430);
xor U39612 (N_39612,N_32284,N_31067);
xnor U39613 (N_39613,N_31560,N_34088);
xor U39614 (N_39614,N_32095,N_32150);
nand U39615 (N_39615,N_32444,N_30727);
nand U39616 (N_39616,N_30585,N_33279);
nand U39617 (N_39617,N_34759,N_30623);
and U39618 (N_39618,N_32419,N_32596);
nand U39619 (N_39619,N_34940,N_31329);
or U39620 (N_39620,N_34313,N_31614);
xnor U39621 (N_39621,N_30371,N_32082);
or U39622 (N_39622,N_31292,N_34137);
nand U39623 (N_39623,N_32263,N_33900);
xor U39624 (N_39624,N_31362,N_32555);
or U39625 (N_39625,N_32659,N_34966);
nand U39626 (N_39626,N_31174,N_33256);
nand U39627 (N_39627,N_31572,N_30786);
and U39628 (N_39628,N_32875,N_31198);
and U39629 (N_39629,N_30074,N_33608);
nand U39630 (N_39630,N_30306,N_31545);
and U39631 (N_39631,N_31214,N_34243);
or U39632 (N_39632,N_30819,N_34952);
xor U39633 (N_39633,N_34895,N_32805);
nor U39634 (N_39634,N_33955,N_30058);
nor U39635 (N_39635,N_31054,N_31257);
nor U39636 (N_39636,N_31205,N_30209);
or U39637 (N_39637,N_32797,N_30919);
or U39638 (N_39638,N_32047,N_31167);
nor U39639 (N_39639,N_31418,N_33461);
or U39640 (N_39640,N_34397,N_34767);
and U39641 (N_39641,N_33956,N_33419);
xor U39642 (N_39642,N_33561,N_33661);
xnor U39643 (N_39643,N_32800,N_34559);
nor U39644 (N_39644,N_32069,N_32786);
or U39645 (N_39645,N_33817,N_31509);
and U39646 (N_39646,N_30001,N_33837);
or U39647 (N_39647,N_33133,N_33401);
nand U39648 (N_39648,N_30740,N_33850);
nor U39649 (N_39649,N_30822,N_31478);
and U39650 (N_39650,N_30737,N_33690);
and U39651 (N_39651,N_33301,N_33106);
nand U39652 (N_39652,N_33068,N_32188);
nand U39653 (N_39653,N_32735,N_33288);
and U39654 (N_39654,N_34766,N_33028);
and U39655 (N_39655,N_34138,N_34829);
and U39656 (N_39656,N_32969,N_33746);
and U39657 (N_39657,N_34904,N_32492);
and U39658 (N_39658,N_30740,N_33648);
and U39659 (N_39659,N_30975,N_31049);
and U39660 (N_39660,N_30497,N_32463);
xnor U39661 (N_39661,N_34152,N_32032);
nor U39662 (N_39662,N_32602,N_33825);
xor U39663 (N_39663,N_31615,N_32483);
xnor U39664 (N_39664,N_32391,N_31915);
xnor U39665 (N_39665,N_33587,N_34629);
nand U39666 (N_39666,N_32268,N_30160);
nand U39667 (N_39667,N_33144,N_34887);
xnor U39668 (N_39668,N_32110,N_34392);
or U39669 (N_39669,N_32999,N_31986);
nor U39670 (N_39670,N_32114,N_33242);
and U39671 (N_39671,N_32195,N_31488);
nor U39672 (N_39672,N_34435,N_33762);
and U39673 (N_39673,N_34689,N_30387);
nor U39674 (N_39674,N_30887,N_31523);
xnor U39675 (N_39675,N_33688,N_31879);
xor U39676 (N_39676,N_32640,N_34230);
and U39677 (N_39677,N_30562,N_34014);
nor U39678 (N_39678,N_33301,N_31687);
and U39679 (N_39679,N_34182,N_30372);
and U39680 (N_39680,N_33478,N_34536);
nor U39681 (N_39681,N_31463,N_31694);
and U39682 (N_39682,N_32409,N_31298);
and U39683 (N_39683,N_33712,N_31302);
or U39684 (N_39684,N_34171,N_34934);
or U39685 (N_39685,N_33107,N_31125);
and U39686 (N_39686,N_33499,N_33286);
nand U39687 (N_39687,N_33418,N_33210);
or U39688 (N_39688,N_33542,N_34374);
and U39689 (N_39689,N_31331,N_31309);
nand U39690 (N_39690,N_30920,N_32844);
or U39691 (N_39691,N_31934,N_34165);
xnor U39692 (N_39692,N_30865,N_32854);
or U39693 (N_39693,N_32214,N_31834);
and U39694 (N_39694,N_30001,N_30789);
nor U39695 (N_39695,N_31066,N_31071);
xor U39696 (N_39696,N_30251,N_34510);
nand U39697 (N_39697,N_31663,N_32727);
or U39698 (N_39698,N_33561,N_33221);
and U39699 (N_39699,N_33041,N_30176);
nand U39700 (N_39700,N_32388,N_34857);
nor U39701 (N_39701,N_34187,N_33388);
and U39702 (N_39702,N_31243,N_34851);
nor U39703 (N_39703,N_33186,N_31890);
nand U39704 (N_39704,N_33809,N_34995);
xor U39705 (N_39705,N_30037,N_30517);
nand U39706 (N_39706,N_31331,N_34337);
xnor U39707 (N_39707,N_34505,N_30760);
xnor U39708 (N_39708,N_32268,N_30563);
xor U39709 (N_39709,N_33458,N_32922);
or U39710 (N_39710,N_33433,N_33040);
nor U39711 (N_39711,N_30627,N_33970);
and U39712 (N_39712,N_34114,N_33246);
or U39713 (N_39713,N_30914,N_33323);
and U39714 (N_39714,N_33017,N_34552);
and U39715 (N_39715,N_33416,N_31387);
and U39716 (N_39716,N_31688,N_32265);
nor U39717 (N_39717,N_32569,N_31755);
xnor U39718 (N_39718,N_34903,N_32555);
nor U39719 (N_39719,N_34949,N_31761);
nor U39720 (N_39720,N_34068,N_33587);
xnor U39721 (N_39721,N_30617,N_33050);
and U39722 (N_39722,N_33305,N_30952);
or U39723 (N_39723,N_33290,N_33831);
and U39724 (N_39724,N_32010,N_32750);
or U39725 (N_39725,N_33597,N_32646);
nor U39726 (N_39726,N_30407,N_32816);
xnor U39727 (N_39727,N_30188,N_34203);
or U39728 (N_39728,N_34215,N_31632);
nand U39729 (N_39729,N_31400,N_30518);
nand U39730 (N_39730,N_31096,N_33762);
or U39731 (N_39731,N_31332,N_33475);
nand U39732 (N_39732,N_30573,N_30463);
or U39733 (N_39733,N_31588,N_34099);
nor U39734 (N_39734,N_33139,N_33959);
and U39735 (N_39735,N_31432,N_32644);
nand U39736 (N_39736,N_31825,N_31490);
and U39737 (N_39737,N_33903,N_30807);
nor U39738 (N_39738,N_31403,N_33593);
nand U39739 (N_39739,N_34209,N_32544);
and U39740 (N_39740,N_30258,N_30721);
or U39741 (N_39741,N_32991,N_32229);
nand U39742 (N_39742,N_33790,N_34331);
or U39743 (N_39743,N_33682,N_34397);
nand U39744 (N_39744,N_33783,N_32887);
nand U39745 (N_39745,N_32679,N_30486);
nor U39746 (N_39746,N_31378,N_30969);
nand U39747 (N_39747,N_30650,N_33684);
xor U39748 (N_39748,N_30181,N_33497);
xnor U39749 (N_39749,N_32167,N_32546);
or U39750 (N_39750,N_31348,N_31929);
xor U39751 (N_39751,N_33450,N_31901);
nor U39752 (N_39752,N_32034,N_30731);
nand U39753 (N_39753,N_32823,N_34578);
xnor U39754 (N_39754,N_33806,N_30720);
or U39755 (N_39755,N_30764,N_32030);
xor U39756 (N_39756,N_34351,N_32821);
or U39757 (N_39757,N_34269,N_33402);
nand U39758 (N_39758,N_33328,N_33628);
or U39759 (N_39759,N_30495,N_34308);
nand U39760 (N_39760,N_31921,N_30478);
and U39761 (N_39761,N_34499,N_31387);
and U39762 (N_39762,N_34304,N_32168);
and U39763 (N_39763,N_30418,N_32341);
nor U39764 (N_39764,N_30546,N_30754);
nand U39765 (N_39765,N_30816,N_30669);
xor U39766 (N_39766,N_30439,N_31521);
nand U39767 (N_39767,N_31264,N_32320);
nor U39768 (N_39768,N_31393,N_30979);
and U39769 (N_39769,N_31416,N_33035);
nor U39770 (N_39770,N_32448,N_31709);
nor U39771 (N_39771,N_31224,N_30851);
or U39772 (N_39772,N_34585,N_33607);
and U39773 (N_39773,N_31771,N_32247);
nand U39774 (N_39774,N_31910,N_34961);
or U39775 (N_39775,N_31150,N_31621);
nor U39776 (N_39776,N_33092,N_32750);
or U39777 (N_39777,N_31911,N_30556);
or U39778 (N_39778,N_34829,N_34836);
or U39779 (N_39779,N_31760,N_33796);
xnor U39780 (N_39780,N_33504,N_34292);
xor U39781 (N_39781,N_30657,N_30541);
nor U39782 (N_39782,N_31321,N_32460);
xor U39783 (N_39783,N_31219,N_34464);
xnor U39784 (N_39784,N_34335,N_31004);
xor U39785 (N_39785,N_30532,N_30888);
and U39786 (N_39786,N_33458,N_33653);
nor U39787 (N_39787,N_30721,N_30185);
nand U39788 (N_39788,N_34058,N_32313);
nor U39789 (N_39789,N_34200,N_34845);
or U39790 (N_39790,N_33309,N_31516);
xnor U39791 (N_39791,N_30267,N_33967);
nand U39792 (N_39792,N_34551,N_33610);
xor U39793 (N_39793,N_34355,N_33543);
or U39794 (N_39794,N_32985,N_31584);
nand U39795 (N_39795,N_31103,N_31393);
or U39796 (N_39796,N_32254,N_33222);
and U39797 (N_39797,N_32804,N_30828);
and U39798 (N_39798,N_30550,N_30078);
or U39799 (N_39799,N_33096,N_33756);
nand U39800 (N_39800,N_34436,N_34014);
xor U39801 (N_39801,N_33975,N_31630);
and U39802 (N_39802,N_34245,N_31150);
nand U39803 (N_39803,N_31819,N_31281);
nand U39804 (N_39804,N_33431,N_31931);
nor U39805 (N_39805,N_34037,N_33865);
xnor U39806 (N_39806,N_30392,N_31943);
nand U39807 (N_39807,N_32205,N_34196);
or U39808 (N_39808,N_31049,N_33586);
nor U39809 (N_39809,N_34378,N_31552);
nor U39810 (N_39810,N_33202,N_32061);
or U39811 (N_39811,N_33727,N_33227);
nor U39812 (N_39812,N_34386,N_34121);
and U39813 (N_39813,N_31693,N_33726);
xnor U39814 (N_39814,N_30583,N_31864);
and U39815 (N_39815,N_32443,N_32955);
nand U39816 (N_39816,N_34364,N_32226);
or U39817 (N_39817,N_30315,N_32374);
and U39818 (N_39818,N_33415,N_33360);
and U39819 (N_39819,N_31723,N_33104);
nand U39820 (N_39820,N_34129,N_34248);
xnor U39821 (N_39821,N_32818,N_33830);
xnor U39822 (N_39822,N_33303,N_34467);
nand U39823 (N_39823,N_32468,N_32747);
xor U39824 (N_39824,N_30028,N_32061);
nand U39825 (N_39825,N_32613,N_32414);
nor U39826 (N_39826,N_31308,N_30174);
nand U39827 (N_39827,N_32225,N_32910);
nand U39828 (N_39828,N_32010,N_34067);
or U39829 (N_39829,N_34858,N_31227);
xnor U39830 (N_39830,N_34055,N_30149);
nor U39831 (N_39831,N_34792,N_33834);
nand U39832 (N_39832,N_32139,N_30613);
and U39833 (N_39833,N_31917,N_34553);
nand U39834 (N_39834,N_33022,N_32089);
nand U39835 (N_39835,N_33003,N_34106);
xnor U39836 (N_39836,N_34721,N_32333);
or U39837 (N_39837,N_32305,N_30906);
or U39838 (N_39838,N_31102,N_32446);
xor U39839 (N_39839,N_34602,N_32035);
xnor U39840 (N_39840,N_32199,N_33599);
nand U39841 (N_39841,N_30658,N_31202);
nor U39842 (N_39842,N_34693,N_33491);
nand U39843 (N_39843,N_30650,N_31762);
nand U39844 (N_39844,N_30692,N_31551);
nand U39845 (N_39845,N_31832,N_33819);
xnor U39846 (N_39846,N_31004,N_33525);
nor U39847 (N_39847,N_30307,N_33314);
and U39848 (N_39848,N_30253,N_32631);
nor U39849 (N_39849,N_34965,N_33919);
and U39850 (N_39850,N_34222,N_33191);
or U39851 (N_39851,N_31629,N_30598);
xor U39852 (N_39852,N_31121,N_32096);
nand U39853 (N_39853,N_33411,N_31011);
nand U39854 (N_39854,N_31322,N_33185);
and U39855 (N_39855,N_31591,N_30796);
and U39856 (N_39856,N_30679,N_34426);
or U39857 (N_39857,N_31158,N_30851);
and U39858 (N_39858,N_33724,N_32982);
xnor U39859 (N_39859,N_30935,N_31383);
xnor U39860 (N_39860,N_31666,N_30273);
nor U39861 (N_39861,N_32676,N_32191);
nor U39862 (N_39862,N_33700,N_34396);
and U39863 (N_39863,N_32306,N_31612);
xor U39864 (N_39864,N_30506,N_32234);
and U39865 (N_39865,N_34598,N_32251);
nor U39866 (N_39866,N_33650,N_32871);
xor U39867 (N_39867,N_32462,N_34475);
xnor U39868 (N_39868,N_32502,N_33152);
and U39869 (N_39869,N_30161,N_30957);
or U39870 (N_39870,N_33655,N_31442);
xnor U39871 (N_39871,N_31702,N_32437);
nor U39872 (N_39872,N_32502,N_34344);
nor U39873 (N_39873,N_34466,N_30328);
nor U39874 (N_39874,N_31802,N_33453);
nor U39875 (N_39875,N_33720,N_33244);
nor U39876 (N_39876,N_31754,N_34552);
nand U39877 (N_39877,N_33336,N_34327);
and U39878 (N_39878,N_33078,N_30040);
xnor U39879 (N_39879,N_34682,N_31973);
nor U39880 (N_39880,N_31522,N_34138);
nor U39881 (N_39881,N_30569,N_33349);
xor U39882 (N_39882,N_32344,N_30027);
nand U39883 (N_39883,N_34952,N_33733);
nor U39884 (N_39884,N_34332,N_32574);
nand U39885 (N_39885,N_31689,N_34440);
nor U39886 (N_39886,N_31992,N_30005);
and U39887 (N_39887,N_34838,N_30346);
nor U39888 (N_39888,N_33795,N_30611);
nor U39889 (N_39889,N_33680,N_32105);
xor U39890 (N_39890,N_34234,N_34143);
xor U39891 (N_39891,N_31734,N_33038);
nand U39892 (N_39892,N_34815,N_34712);
or U39893 (N_39893,N_34407,N_31914);
xor U39894 (N_39894,N_33877,N_31536);
nor U39895 (N_39895,N_31109,N_30812);
nand U39896 (N_39896,N_31700,N_32996);
nor U39897 (N_39897,N_30951,N_33804);
nand U39898 (N_39898,N_31422,N_33353);
nand U39899 (N_39899,N_32557,N_32830);
xnor U39900 (N_39900,N_33447,N_30474);
xor U39901 (N_39901,N_30654,N_30981);
xnor U39902 (N_39902,N_31376,N_34227);
and U39903 (N_39903,N_31165,N_31342);
nor U39904 (N_39904,N_34954,N_32281);
or U39905 (N_39905,N_31546,N_32885);
nand U39906 (N_39906,N_34152,N_31085);
nand U39907 (N_39907,N_34967,N_30935);
xnor U39908 (N_39908,N_30029,N_31800);
nand U39909 (N_39909,N_31991,N_30317);
nand U39910 (N_39910,N_32879,N_30060);
nand U39911 (N_39911,N_30765,N_30496);
nor U39912 (N_39912,N_30929,N_32870);
or U39913 (N_39913,N_32157,N_31265);
nor U39914 (N_39914,N_30845,N_31226);
or U39915 (N_39915,N_32111,N_32007);
or U39916 (N_39916,N_31924,N_34804);
nor U39917 (N_39917,N_33508,N_32810);
nand U39918 (N_39918,N_31143,N_32393);
and U39919 (N_39919,N_30997,N_33168);
nand U39920 (N_39920,N_33020,N_32252);
and U39921 (N_39921,N_31244,N_33895);
or U39922 (N_39922,N_32524,N_32673);
or U39923 (N_39923,N_31289,N_31324);
nor U39924 (N_39924,N_30320,N_34655);
or U39925 (N_39925,N_30341,N_34124);
and U39926 (N_39926,N_30847,N_32829);
nor U39927 (N_39927,N_30838,N_33775);
nand U39928 (N_39928,N_31846,N_34602);
nand U39929 (N_39929,N_31899,N_32063);
nand U39930 (N_39930,N_34971,N_30928);
nand U39931 (N_39931,N_31467,N_34882);
nand U39932 (N_39932,N_31877,N_31828);
xor U39933 (N_39933,N_30669,N_30471);
and U39934 (N_39934,N_34489,N_33362);
nor U39935 (N_39935,N_34248,N_32013);
xnor U39936 (N_39936,N_32197,N_31408);
and U39937 (N_39937,N_34103,N_31517);
and U39938 (N_39938,N_31573,N_33624);
or U39939 (N_39939,N_32277,N_31354);
nand U39940 (N_39940,N_34763,N_31506);
and U39941 (N_39941,N_34771,N_34556);
or U39942 (N_39942,N_34097,N_31373);
or U39943 (N_39943,N_32622,N_33814);
xor U39944 (N_39944,N_34091,N_34276);
or U39945 (N_39945,N_31839,N_34531);
nor U39946 (N_39946,N_34314,N_32137);
or U39947 (N_39947,N_34954,N_33476);
nand U39948 (N_39948,N_30480,N_31967);
or U39949 (N_39949,N_32332,N_31544);
and U39950 (N_39950,N_33734,N_31454);
nand U39951 (N_39951,N_34761,N_34013);
nor U39952 (N_39952,N_32771,N_33625);
nor U39953 (N_39953,N_31693,N_31487);
nor U39954 (N_39954,N_33974,N_32222);
nand U39955 (N_39955,N_33304,N_31324);
nor U39956 (N_39956,N_31365,N_32939);
xnor U39957 (N_39957,N_32949,N_31199);
nor U39958 (N_39958,N_30202,N_34758);
xor U39959 (N_39959,N_30832,N_30545);
nor U39960 (N_39960,N_34832,N_31214);
or U39961 (N_39961,N_33710,N_32511);
xnor U39962 (N_39962,N_32797,N_32326);
nor U39963 (N_39963,N_30397,N_32320);
or U39964 (N_39964,N_33454,N_31521);
xor U39965 (N_39965,N_33559,N_34547);
nand U39966 (N_39966,N_31633,N_34991);
nand U39967 (N_39967,N_32078,N_32444);
nand U39968 (N_39968,N_33706,N_32622);
xor U39969 (N_39969,N_33829,N_32681);
nand U39970 (N_39970,N_33664,N_33750);
or U39971 (N_39971,N_34196,N_30805);
nand U39972 (N_39972,N_33526,N_33459);
and U39973 (N_39973,N_34409,N_33989);
and U39974 (N_39974,N_33572,N_34745);
xnor U39975 (N_39975,N_32869,N_33094);
xnor U39976 (N_39976,N_34889,N_32532);
xnor U39977 (N_39977,N_31595,N_33929);
and U39978 (N_39978,N_34375,N_31777);
and U39979 (N_39979,N_31605,N_30175);
nand U39980 (N_39980,N_32778,N_33631);
and U39981 (N_39981,N_33936,N_30618);
or U39982 (N_39982,N_34673,N_32360);
nand U39983 (N_39983,N_34350,N_34704);
and U39984 (N_39984,N_30406,N_31040);
and U39985 (N_39985,N_31855,N_30869);
or U39986 (N_39986,N_31965,N_34987);
nor U39987 (N_39987,N_32883,N_30918);
nor U39988 (N_39988,N_33077,N_34387);
or U39989 (N_39989,N_33819,N_32524);
or U39990 (N_39990,N_30137,N_33535);
or U39991 (N_39991,N_32269,N_33631);
nor U39992 (N_39992,N_32290,N_32456);
xor U39993 (N_39993,N_34607,N_30314);
or U39994 (N_39994,N_31350,N_33225);
or U39995 (N_39995,N_32072,N_32594);
or U39996 (N_39996,N_31436,N_34911);
or U39997 (N_39997,N_33119,N_30736);
and U39998 (N_39998,N_30259,N_34152);
and U39999 (N_39999,N_32841,N_32995);
xnor U40000 (N_40000,N_36603,N_37389);
or U40001 (N_40001,N_38488,N_37893);
xnor U40002 (N_40002,N_38539,N_38319);
nor U40003 (N_40003,N_36222,N_38869);
nor U40004 (N_40004,N_38544,N_35032);
nor U40005 (N_40005,N_38413,N_36054);
and U40006 (N_40006,N_39977,N_38937);
or U40007 (N_40007,N_37248,N_36423);
and U40008 (N_40008,N_35970,N_39909);
nand U40009 (N_40009,N_38829,N_37836);
nand U40010 (N_40010,N_39594,N_36400);
and U40011 (N_40011,N_37977,N_37864);
or U40012 (N_40012,N_37286,N_38681);
and U40013 (N_40013,N_36030,N_36316);
or U40014 (N_40014,N_37386,N_39466);
and U40015 (N_40015,N_37014,N_36043);
xnor U40016 (N_40016,N_38577,N_38325);
xor U40017 (N_40017,N_35479,N_37591);
or U40018 (N_40018,N_39046,N_39770);
or U40019 (N_40019,N_36154,N_35303);
nand U40020 (N_40020,N_37867,N_36348);
nand U40021 (N_40021,N_35268,N_37353);
nor U40022 (N_40022,N_35209,N_39652);
nand U40023 (N_40023,N_39571,N_36701);
nor U40024 (N_40024,N_37122,N_38884);
nor U40025 (N_40025,N_39035,N_39173);
nand U40026 (N_40026,N_37880,N_36172);
and U40027 (N_40027,N_37720,N_39147);
nand U40028 (N_40028,N_35779,N_38445);
or U40029 (N_40029,N_36979,N_35146);
and U40030 (N_40030,N_37242,N_37993);
or U40031 (N_40031,N_37297,N_37770);
nand U40032 (N_40032,N_37070,N_39142);
nand U40033 (N_40033,N_35556,N_35871);
xor U40034 (N_40034,N_38055,N_39056);
nand U40035 (N_40035,N_39239,N_36507);
xnor U40036 (N_40036,N_38099,N_39815);
xor U40037 (N_40037,N_36343,N_39792);
and U40038 (N_40038,N_38134,N_37903);
and U40039 (N_40039,N_36394,N_37978);
nand U40040 (N_40040,N_39442,N_36063);
or U40041 (N_40041,N_38020,N_39771);
xor U40042 (N_40042,N_37200,N_38284);
and U40043 (N_40043,N_38012,N_39537);
or U40044 (N_40044,N_35222,N_37898);
and U40045 (N_40045,N_35802,N_39673);
nor U40046 (N_40046,N_37011,N_36415);
nand U40047 (N_40047,N_36015,N_39775);
and U40048 (N_40048,N_39163,N_35287);
nand U40049 (N_40049,N_36688,N_39176);
xor U40050 (N_40050,N_39181,N_38062);
and U40051 (N_40051,N_35201,N_39472);
or U40052 (N_40052,N_39004,N_37722);
xnor U40053 (N_40053,N_36721,N_36941);
xor U40054 (N_40054,N_38542,N_39689);
and U40055 (N_40055,N_39152,N_37562);
or U40056 (N_40056,N_35772,N_35811);
xor U40057 (N_40057,N_36028,N_39658);
nor U40058 (N_40058,N_37422,N_36782);
nor U40059 (N_40059,N_39477,N_39108);
or U40060 (N_40060,N_37377,N_35440);
nand U40061 (N_40061,N_36821,N_35696);
and U40062 (N_40062,N_36545,N_39078);
and U40063 (N_40063,N_36712,N_35463);
nand U40064 (N_40064,N_37910,N_37401);
xor U40065 (N_40065,N_38934,N_37037);
or U40066 (N_40066,N_35043,N_38187);
and U40067 (N_40067,N_35776,N_37282);
nand U40068 (N_40068,N_35049,N_36196);
xnor U40069 (N_40069,N_37698,N_39855);
xor U40070 (N_40070,N_37628,N_36909);
xnor U40071 (N_40071,N_36745,N_35788);
or U40072 (N_40072,N_37211,N_36053);
or U40073 (N_40073,N_37511,N_36337);
and U40074 (N_40074,N_38212,N_38905);
and U40075 (N_40075,N_37696,N_36977);
nand U40076 (N_40076,N_35053,N_37808);
nand U40077 (N_40077,N_38311,N_37520);
nor U40078 (N_40078,N_35832,N_39077);
nor U40079 (N_40079,N_37428,N_37912);
or U40080 (N_40080,N_36068,N_39647);
nor U40081 (N_40081,N_39653,N_38589);
nor U40082 (N_40082,N_39259,N_37429);
or U40083 (N_40083,N_39710,N_36528);
and U40084 (N_40084,N_35985,N_39500);
xnor U40085 (N_40085,N_38135,N_38971);
xnor U40086 (N_40086,N_37356,N_38595);
and U40087 (N_40087,N_38504,N_39878);
nor U40088 (N_40088,N_38685,N_38691);
xor U40089 (N_40089,N_35159,N_35390);
nand U40090 (N_40090,N_36322,N_35600);
nor U40091 (N_40091,N_39356,N_38633);
xnor U40092 (N_40092,N_39481,N_35228);
xor U40093 (N_40093,N_35437,N_39742);
nand U40094 (N_40094,N_35286,N_35660);
and U40095 (N_40095,N_38973,N_39225);
or U40096 (N_40096,N_36881,N_35766);
nand U40097 (N_40097,N_36574,N_35745);
nor U40098 (N_40098,N_35509,N_38551);
and U40099 (N_40099,N_36864,N_38947);
xor U40100 (N_40100,N_35328,N_35547);
nand U40101 (N_40101,N_36862,N_37071);
xnor U40102 (N_40102,N_36890,N_39404);
xnor U40103 (N_40103,N_35719,N_39797);
and U40104 (N_40104,N_35502,N_38571);
nor U40105 (N_40105,N_35526,N_38716);
nand U40106 (N_40106,N_38080,N_36263);
nor U40107 (N_40107,N_39799,N_35410);
xnor U40108 (N_40108,N_35572,N_37460);
nand U40109 (N_40109,N_38793,N_35536);
xnor U40110 (N_40110,N_37941,N_38735);
nor U40111 (N_40111,N_36406,N_36946);
xnor U40112 (N_40112,N_39055,N_37534);
nand U40113 (N_40113,N_37443,N_36796);
and U40114 (N_40114,N_36808,N_37485);
nand U40115 (N_40115,N_38151,N_39819);
or U40116 (N_40116,N_36611,N_37212);
and U40117 (N_40117,N_37156,N_35177);
and U40118 (N_40118,N_35761,N_39458);
nor U40119 (N_40119,N_39629,N_35105);
or U40120 (N_40120,N_37889,N_35198);
nand U40121 (N_40121,N_37635,N_36131);
nand U40122 (N_40122,N_37495,N_37195);
xnor U40123 (N_40123,N_39730,N_37043);
nor U40124 (N_40124,N_35363,N_37819);
or U40125 (N_40125,N_35578,N_39119);
xor U40126 (N_40126,N_35817,N_39268);
nand U40127 (N_40127,N_35601,N_38082);
and U40128 (N_40128,N_37087,N_35293);
xor U40129 (N_40129,N_38465,N_36670);
xnor U40130 (N_40130,N_37247,N_35013);
and U40131 (N_40131,N_39403,N_35521);
nand U40132 (N_40132,N_37782,N_36535);
or U40133 (N_40133,N_38895,N_35839);
xnor U40134 (N_40134,N_35940,N_36328);
xnor U40135 (N_40135,N_36044,N_38297);
xor U40136 (N_40136,N_39635,N_37791);
nand U40137 (N_40137,N_38576,N_39414);
xor U40138 (N_40138,N_38052,N_39378);
xnor U40139 (N_40139,N_36693,N_38156);
nor U40140 (N_40140,N_39503,N_39619);
or U40141 (N_40141,N_37330,N_39674);
xor U40142 (N_40142,N_35626,N_37250);
and U40143 (N_40143,N_38513,N_39428);
nand U40144 (N_40144,N_36565,N_38254);
nand U40145 (N_40145,N_36359,N_36181);
xor U40146 (N_40146,N_39047,N_39830);
or U40147 (N_40147,N_36681,N_39185);
nor U40148 (N_40148,N_38514,N_37610);
nor U40149 (N_40149,N_39218,N_36967);
nor U40150 (N_40150,N_35001,N_36876);
nor U40151 (N_40151,N_38825,N_38060);
and U40152 (N_40152,N_38555,N_36934);
xor U40153 (N_40153,N_39029,N_38653);
or U40154 (N_40154,N_37291,N_37254);
nor U40155 (N_40155,N_38105,N_39501);
xor U40156 (N_40156,N_35525,N_36998);
or U40157 (N_40157,N_35492,N_37338);
nand U40158 (N_40158,N_37293,N_36445);
xnor U40159 (N_40159,N_39256,N_35330);
nor U40160 (N_40160,N_37048,N_38567);
or U40161 (N_40161,N_37750,N_36072);
and U40162 (N_40162,N_37568,N_35487);
xnor U40163 (N_40163,N_37036,N_35425);
or U40164 (N_40164,N_38473,N_35948);
xor U40165 (N_40165,N_36041,N_39849);
xor U40166 (N_40166,N_38705,N_38597);
nand U40167 (N_40167,N_36293,N_38910);
or U40168 (N_40168,N_37380,N_39339);
nor U40169 (N_40169,N_35755,N_38215);
and U40170 (N_40170,N_37243,N_38774);
or U40171 (N_40171,N_37308,N_37040);
and U40172 (N_40172,N_37502,N_38260);
nor U40173 (N_40173,N_36382,N_38987);
xor U40174 (N_40174,N_39470,N_35362);
or U40175 (N_40175,N_36246,N_38783);
xor U40176 (N_40176,N_38833,N_35831);
or U40177 (N_40177,N_37968,N_35971);
nand U40178 (N_40178,N_36674,N_35978);
or U40179 (N_40179,N_35067,N_35099);
and U40180 (N_40180,N_38917,N_36676);
and U40181 (N_40181,N_35218,N_38250);
or U40182 (N_40182,N_35684,N_35106);
nor U40183 (N_40183,N_39872,N_38725);
nor U40184 (N_40184,N_37285,N_37833);
xnor U40185 (N_40185,N_36793,N_39267);
or U40186 (N_40186,N_35200,N_35383);
and U40187 (N_40187,N_37795,N_38933);
or U40188 (N_40188,N_38913,N_38265);
and U40189 (N_40189,N_35242,N_37283);
or U40190 (N_40190,N_38185,N_38647);
xnor U40191 (N_40191,N_38394,N_37999);
nor U40192 (N_40192,N_35493,N_35511);
or U40193 (N_40193,N_38509,N_35056);
nand U40194 (N_40194,N_35789,N_38815);
and U40195 (N_40195,N_35651,N_37112);
nand U40196 (N_40196,N_38130,N_36970);
or U40197 (N_40197,N_35281,N_35878);
or U40198 (N_40198,N_38481,N_37376);
xor U40199 (N_40199,N_35954,N_36464);
or U40200 (N_40200,N_38040,N_36550);
and U40201 (N_40201,N_36219,N_35340);
nor U40202 (N_40202,N_35091,N_38415);
or U40203 (N_40203,N_37986,N_35849);
nor U40204 (N_40204,N_35720,N_36612);
xnor U40205 (N_40205,N_38333,N_36245);
nand U40206 (N_40206,N_38124,N_38512);
or U40207 (N_40207,N_37202,N_35296);
or U40208 (N_40208,N_36650,N_37224);
xnor U40209 (N_40209,N_37671,N_37328);
nand U40210 (N_40210,N_37663,N_36857);
nand U40211 (N_40211,N_37094,N_37454);
or U40212 (N_40212,N_37571,N_35711);
nand U40213 (N_40213,N_39111,N_35958);
or U40214 (N_40214,N_36945,N_37585);
xnor U40215 (N_40215,N_36476,N_39827);
xnor U40216 (N_40216,N_35939,N_36547);
and U40217 (N_40217,N_37597,N_38898);
nand U40218 (N_40218,N_37371,N_38469);
xnor U40219 (N_40219,N_35313,N_36931);
xor U40220 (N_40220,N_39332,N_35285);
and U40221 (N_40221,N_37452,N_39129);
and U40222 (N_40222,N_35927,N_36659);
xnor U40223 (N_40223,N_37827,N_39490);
xnor U40224 (N_40224,N_38457,N_38068);
or U40225 (N_40225,N_35609,N_38952);
nor U40226 (N_40226,N_36960,N_39755);
nor U40227 (N_40227,N_39014,N_36278);
xor U40228 (N_40228,N_37095,N_36018);
and U40229 (N_40229,N_36695,N_35284);
nor U40230 (N_40230,N_35797,N_37113);
and U40231 (N_40231,N_38063,N_35171);
nor U40232 (N_40232,N_39419,N_36040);
nand U40233 (N_40233,N_35860,N_37575);
nand U40234 (N_40234,N_35596,N_39602);
or U40235 (N_40235,N_35499,N_39237);
nand U40236 (N_40236,N_37260,N_39675);
nor U40237 (N_40237,N_38820,N_37984);
nand U40238 (N_40238,N_35644,N_35851);
or U40239 (N_40239,N_38516,N_36839);
xor U40240 (N_40240,N_37801,N_39936);
nor U40241 (N_40241,N_39456,N_38744);
or U40242 (N_40242,N_37375,N_36236);
or U40243 (N_40243,N_39604,N_35768);
or U40244 (N_40244,N_39308,N_39130);
nand U40245 (N_40245,N_36904,N_39822);
nand U40246 (N_40246,N_38304,N_39449);
and U40247 (N_40247,N_39717,N_36552);
xor U40248 (N_40248,N_39930,N_38550);
nand U40249 (N_40249,N_36664,N_35522);
and U40250 (N_40250,N_38092,N_35709);
nand U40251 (N_40251,N_38339,N_37574);
xor U40252 (N_40252,N_39128,N_38949);
and U40253 (N_40253,N_35305,N_37305);
xor U40254 (N_40254,N_35504,N_36927);
nor U40255 (N_40255,N_39778,N_38464);
or U40256 (N_40256,N_38618,N_38975);
nand U40257 (N_40257,N_37336,N_38030);
nor U40258 (N_40258,N_38125,N_35167);
and U40259 (N_40259,N_37431,N_36867);
and U40260 (N_40260,N_39915,N_36773);
or U40261 (N_40261,N_38919,N_38310);
xnor U40262 (N_40262,N_38948,N_36250);
nor U40263 (N_40263,N_38792,N_39609);
xor U40264 (N_40264,N_35678,N_39985);
xnor U40265 (N_40265,N_37455,N_35751);
nor U40266 (N_40266,N_39581,N_39338);
and U40267 (N_40267,N_38737,N_37398);
and U40268 (N_40268,N_35844,N_37588);
and U40269 (N_40269,N_38538,N_36972);
nand U40270 (N_40270,N_38643,N_39499);
or U40271 (N_40271,N_36296,N_39840);
or U40272 (N_40272,N_36694,N_39281);
and U40273 (N_40273,N_37846,N_36461);
or U40274 (N_40274,N_36700,N_36429);
nor U40275 (N_40275,N_38611,N_36925);
or U40276 (N_40276,N_38867,N_39085);
or U40277 (N_40277,N_38881,N_37959);
and U40278 (N_40278,N_35517,N_39275);
nor U40279 (N_40279,N_37966,N_39896);
nand U40280 (N_40280,N_36002,N_35900);
xnor U40281 (N_40281,N_38651,N_38989);
or U40282 (N_40282,N_38390,N_39000);
and U40283 (N_40283,N_39425,N_37461);
xor U40284 (N_40284,N_35093,N_37902);
nor U40285 (N_40285,N_35230,N_38345);
or U40286 (N_40286,N_38756,N_37144);
nor U40287 (N_40287,N_37390,N_36083);
nor U40288 (N_40288,N_39637,N_36987);
or U40289 (N_40289,N_35765,N_35869);
and U40290 (N_40290,N_36096,N_37146);
nor U40291 (N_40291,N_36298,N_35165);
nor U40292 (N_40292,N_38334,N_39479);
nand U40293 (N_40293,N_37822,N_39059);
and U40294 (N_40294,N_39079,N_38501);
xnor U40295 (N_40295,N_39260,N_38385);
and U40296 (N_40296,N_37258,N_38746);
nand U40297 (N_40297,N_35068,N_39367);
nand U40298 (N_40298,N_37169,N_37116);
and U40299 (N_40299,N_38483,N_35962);
nor U40300 (N_40300,N_37155,N_35226);
xor U40301 (N_40301,N_35599,N_37439);
or U40302 (N_40302,N_35663,N_38428);
nand U40303 (N_40303,N_37538,N_38369);
xnor U40304 (N_40304,N_38015,N_37435);
and U40305 (N_40305,N_37515,N_35993);
or U40306 (N_40306,N_39410,N_36849);
nor U40307 (N_40307,N_39816,N_38326);
and U40308 (N_40308,N_38195,N_36607);
nor U40309 (N_40309,N_35255,N_38780);
or U40310 (N_40310,N_37134,N_39919);
or U40311 (N_40311,N_38367,N_39321);
and U40312 (N_40312,N_35208,N_35752);
xor U40313 (N_40313,N_39250,N_37838);
nand U40314 (N_40314,N_36962,N_38591);
and U40315 (N_40315,N_35490,N_37177);
and U40316 (N_40316,N_39595,N_35698);
or U40317 (N_40317,N_35671,N_39583);
or U40318 (N_40318,N_37947,N_39156);
and U40319 (N_40319,N_38515,N_39620);
or U40320 (N_40320,N_35734,N_37464);
and U40321 (N_40321,N_38073,N_38355);
xor U40322 (N_40322,N_38272,N_38912);
or U40323 (N_40323,N_36306,N_37278);
xor U40324 (N_40324,N_39701,N_35220);
nor U40325 (N_40325,N_36238,N_36957);
or U40326 (N_40326,N_39148,N_38764);
nor U40327 (N_40327,N_36812,N_39651);
and U40328 (N_40328,N_36790,N_35604);
nor U40329 (N_40329,N_39685,N_39920);
xor U40330 (N_40330,N_35533,N_35472);
xnor U40331 (N_40331,N_37400,N_35083);
xnor U40332 (N_40332,N_36155,N_37466);
and U40333 (N_40333,N_38871,N_38713);
nor U40334 (N_40334,N_37909,N_36365);
nor U40335 (N_40335,N_37761,N_35070);
xnor U40336 (N_40336,N_37627,N_38071);
xnor U40337 (N_40337,N_35044,N_36530);
xnor U40338 (N_40338,N_35731,N_35646);
nand U40339 (N_40339,N_39633,N_38035);
nand U40340 (N_40340,N_39098,N_38788);
xor U40341 (N_40341,N_35102,N_39424);
xnor U40342 (N_40342,N_38388,N_39045);
or U40343 (N_40343,N_37492,N_35654);
or U40344 (N_40344,N_36418,N_36008);
or U40345 (N_40345,N_39471,N_38558);
and U40346 (N_40346,N_35697,N_39201);
xor U40347 (N_40347,N_37004,N_35447);
nand U40348 (N_40348,N_35219,N_38605);
xor U40349 (N_40349,N_38202,N_37920);
nor U40350 (N_40350,N_37873,N_36736);
and U40351 (N_40351,N_39688,N_37220);
nor U40352 (N_40352,N_38386,N_37593);
xor U40353 (N_40353,N_38363,N_36396);
or U40354 (N_40354,N_36878,N_37415);
xor U40355 (N_40355,N_38938,N_38358);
xnor U40356 (N_40356,N_35901,N_37019);
xor U40357 (N_40357,N_39359,N_39668);
nor U40358 (N_40358,N_39320,N_35594);
and U40359 (N_40359,N_38252,N_39699);
xnor U40360 (N_40360,N_37619,N_36035);
nor U40361 (N_40361,N_35598,N_39408);
and U40362 (N_40362,N_35353,N_38659);
or U40363 (N_40363,N_39402,N_36624);
xor U40364 (N_40364,N_35854,N_38417);
and U40365 (N_40365,N_38837,N_37103);
xnor U40366 (N_40366,N_37958,N_36786);
nor U40367 (N_40367,N_38262,N_36133);
nand U40368 (N_40368,N_36184,N_37961);
nand U40369 (N_40369,N_37605,N_39051);
or U40370 (N_40370,N_36737,N_39017);
nor U40371 (N_40371,N_39687,N_35430);
and U40372 (N_40372,N_36024,N_39318);
or U40373 (N_40373,N_35829,N_38164);
xnor U40374 (N_40374,N_36976,N_37161);
or U40375 (N_40375,N_39102,N_36794);
nor U40376 (N_40376,N_35392,N_37222);
nor U40377 (N_40377,N_36587,N_35804);
nor U40378 (N_40378,N_38962,N_38113);
nand U40379 (N_40379,N_35343,N_38711);
or U40380 (N_40380,N_39234,N_35124);
nand U40381 (N_40381,N_39554,N_39013);
or U40382 (N_40382,N_38454,N_39663);
nor U40383 (N_40383,N_36300,N_39922);
or U40384 (N_40384,N_38463,N_36704);
nor U40385 (N_40385,N_38751,N_36430);
xnor U40386 (N_40386,N_36776,N_36457);
xnor U40387 (N_40387,N_39115,N_37409);
or U40388 (N_40388,N_36491,N_35763);
and U40389 (N_40389,N_37210,N_37221);
nor U40390 (N_40390,N_38184,N_37214);
xor U40391 (N_40391,N_38768,N_36307);
or U40392 (N_40392,N_39877,N_38392);
and U40393 (N_40393,N_39934,N_37799);
and U40394 (N_40394,N_37586,N_37764);
nor U40395 (N_40395,N_38199,N_36991);
nor U40396 (N_40396,N_38444,N_39530);
and U40397 (N_40397,N_38535,N_35700);
nor U40398 (N_40398,N_39100,N_37013);
nand U40399 (N_40399,N_38342,N_39097);
xor U40400 (N_40400,N_39041,N_38959);
nand U40401 (N_40401,N_37262,N_39184);
or U40402 (N_40402,N_37908,N_36220);
or U40403 (N_40403,N_39948,N_37580);
nand U40404 (N_40404,N_37426,N_37667);
xor U40405 (N_40405,N_37049,N_39535);
nand U40406 (N_40406,N_37772,N_37706);
xnor U40407 (N_40407,N_39200,N_36846);
and U40408 (N_40408,N_39220,N_35387);
xnor U40409 (N_40409,N_36952,N_36569);
nand U40410 (N_40410,N_35791,N_38486);
nand U40411 (N_40411,N_37099,N_38280);
and U40412 (N_40412,N_38313,N_35461);
or U40413 (N_40413,N_35773,N_38323);
nand U40414 (N_40414,N_37082,N_38963);
nand U40415 (N_40415,N_35557,N_37234);
xnor U40416 (N_40416,N_37796,N_36818);
nor U40417 (N_40417,N_38141,N_35396);
xnor U40418 (N_40418,N_39729,N_35040);
nor U40419 (N_40419,N_36708,N_35309);
nand U40420 (N_40420,N_35277,N_36287);
and U40421 (N_40421,N_39468,N_37697);
nand U40422 (N_40422,N_36148,N_37292);
nor U40423 (N_40423,N_38489,N_36575);
nor U40424 (N_40424,N_37024,N_36431);
nand U40425 (N_40425,N_39894,N_39258);
nor U40426 (N_40426,N_36953,N_38759);
or U40427 (N_40427,N_37233,N_35629);
or U40428 (N_40428,N_36824,N_37713);
xor U40429 (N_40429,N_35775,N_36902);
xor U40430 (N_40430,N_37391,N_37933);
or U40431 (N_40431,N_37862,N_38378);
nor U40432 (N_40432,N_38293,N_37078);
or U40433 (N_40433,N_36562,N_38620);
xor U40434 (N_40434,N_36381,N_37917);
nand U40435 (N_40435,N_38821,N_38972);
or U40436 (N_40436,N_38411,N_35445);
and U40437 (N_40437,N_37023,N_38324);
nor U40438 (N_40438,N_38449,N_39266);
xnor U40439 (N_40439,N_35787,N_36869);
or U40440 (N_40440,N_38696,N_35875);
or U40441 (N_40441,N_38797,N_37125);
and U40442 (N_40442,N_39708,N_35754);
and U40443 (N_40443,N_36785,N_38301);
nand U40444 (N_40444,N_35579,N_38132);
nand U40445 (N_40445,N_37751,N_38924);
and U40446 (N_40446,N_35782,N_38070);
or U40447 (N_40447,N_37042,N_38236);
xnor U40448 (N_40448,N_36450,N_39809);
xnor U40449 (N_40449,N_39319,N_36397);
xnor U40450 (N_40450,N_39966,N_35679);
nand U40451 (N_40451,N_37271,N_37081);
nor U40452 (N_40452,N_37886,N_36442);
xor U40453 (N_40453,N_37630,N_37624);
nand U40454 (N_40454,N_37872,N_36473);
xor U40455 (N_40455,N_35834,N_37897);
nand U40456 (N_40456,N_38570,N_39683);
and U40457 (N_40457,N_39228,N_36523);
and U40458 (N_40458,N_36891,N_39358);
xnor U40459 (N_40459,N_37832,N_39835);
xor U40460 (N_40460,N_35336,N_37521);
xor U40461 (N_40461,N_35894,N_37759);
nor U40462 (N_40462,N_39686,N_36106);
and U40463 (N_40463,N_37463,N_39122);
and U40464 (N_40464,N_35294,N_38227);
nor U40465 (N_40465,N_36126,N_38809);
and U40466 (N_40466,N_37996,N_36980);
xor U40467 (N_40467,N_36555,N_39324);
nor U40468 (N_40468,N_37859,N_37930);
and U40469 (N_40469,N_38758,N_39020);
xor U40470 (N_40470,N_37062,N_36371);
nand U40471 (N_40471,N_39096,N_35004);
and U40472 (N_40472,N_36829,N_36197);
nand U40473 (N_40473,N_35398,N_36049);
xor U40474 (N_40474,N_37361,N_37159);
nor U40475 (N_40475,N_35980,N_38640);
nor U40476 (N_40476,N_37484,N_36482);
or U40477 (N_40477,N_39758,N_39204);
or U40478 (N_40478,N_35887,N_39393);
xor U40479 (N_40479,N_36496,N_35808);
or U40480 (N_40480,N_39052,N_36486);
and U40481 (N_40481,N_38013,N_39577);
nor U40482 (N_40482,N_37988,N_38660);
nor U40483 (N_40483,N_35069,N_38822);
nand U40484 (N_40484,N_37038,N_37393);
and U40485 (N_40485,N_36297,N_36797);
and U40486 (N_40486,N_35205,N_37806);
nand U40487 (N_40487,N_39274,N_37513);
and U40488 (N_40488,N_36440,N_35756);
xor U40489 (N_40489,N_35778,N_36820);
xnor U40490 (N_40490,N_39865,N_35870);
nor U40491 (N_40491,N_38945,N_37186);
xnor U40492 (N_40492,N_38258,N_39650);
nor U40493 (N_40493,N_35385,N_35821);
and U40494 (N_40494,N_38518,N_39837);
and U40495 (N_40495,N_35221,N_37302);
xor U40496 (N_40496,N_38650,N_39624);
or U40497 (N_40497,N_38806,N_37329);
xnor U40498 (N_40498,N_38451,N_35714);
and U40499 (N_40499,N_37392,N_35065);
nand U40500 (N_40500,N_36997,N_38169);
nand U40501 (N_40501,N_38565,N_39090);
xor U40502 (N_40502,N_37274,N_38562);
or U40503 (N_40503,N_37241,N_35361);
xor U40504 (N_40504,N_39582,N_35290);
and U40505 (N_40505,N_35969,N_37005);
nand U40506 (N_40506,N_36517,N_36567);
nand U40507 (N_40507,N_36277,N_39560);
and U40508 (N_40508,N_37404,N_39344);
nor U40509 (N_40509,N_37632,N_37972);
nand U40510 (N_40510,N_35805,N_37171);
nand U40511 (N_40511,N_37850,N_38946);
xnor U40512 (N_40512,N_36130,N_37837);
nor U40513 (N_40513,N_37721,N_38740);
nand U40514 (N_40514,N_39640,N_38863);
nor U40515 (N_40515,N_39151,N_36774);
nand U40516 (N_40516,N_36055,N_38222);
and U40517 (N_40517,N_36185,N_39507);
and U40518 (N_40518,N_37904,N_35982);
nand U40519 (N_40519,N_37411,N_37997);
or U40520 (N_40520,N_39974,N_37027);
xnor U40521 (N_40521,N_35455,N_39842);
nor U40522 (N_40522,N_37803,N_39927);
nor U40523 (N_40523,N_39520,N_36645);
or U40524 (N_40524,N_36834,N_36933);
xor U40525 (N_40525,N_35133,N_36355);
nor U40526 (N_40526,N_35750,N_37109);
nor U40527 (N_40527,N_37549,N_38541);
or U40528 (N_40528,N_35326,N_39569);
and U40529 (N_40529,N_36536,N_35368);
or U40530 (N_40530,N_35807,N_38761);
and U40531 (N_40531,N_36061,N_37863);
nor U40532 (N_40532,N_35938,N_35054);
nand U40533 (N_40533,N_35327,N_39114);
or U40534 (N_40534,N_37000,N_39243);
and U40535 (N_40535,N_38152,N_35736);
xnor U40536 (N_40536,N_38799,N_38246);
or U40537 (N_40537,N_39110,N_37265);
nor U40538 (N_40538,N_37921,N_39191);
or U40539 (N_40539,N_39951,N_38684);
or U40540 (N_40540,N_37932,N_39280);
xor U40541 (N_40541,N_37542,N_39549);
xor U40542 (N_40542,N_37623,N_37749);
nand U40543 (N_40543,N_36628,N_39747);
nand U40544 (N_40544,N_39287,N_35713);
xnor U40545 (N_40545,N_36026,N_38752);
or U40546 (N_40546,N_39263,N_36281);
nor U40547 (N_40547,N_37203,N_35259);
and U40548 (N_40548,N_38935,N_37268);
nand U40549 (N_40549,N_36999,N_37412);
nand U40550 (N_40550,N_39498,N_38892);
or U40551 (N_40551,N_35139,N_37854);
nor U40552 (N_40552,N_36285,N_35682);
or U40553 (N_40553,N_39016,N_35407);
and U40554 (N_40554,N_39245,N_39136);
and U40555 (N_40555,N_36335,N_37694);
or U40556 (N_40556,N_39627,N_38269);
nor U40557 (N_40557,N_37059,N_36696);
and U40558 (N_40558,N_39293,N_35846);
or U40559 (N_40559,N_39095,N_39439);
or U40560 (N_40560,N_39112,N_39612);
xor U40561 (N_40561,N_36843,N_39264);
xnor U40562 (N_40562,N_35439,N_36588);
or U40563 (N_40563,N_36805,N_37715);
and U40564 (N_40564,N_39962,N_39179);
xor U40565 (N_40565,N_39355,N_35064);
xor U40566 (N_40566,N_36710,N_35724);
and U40567 (N_40567,N_38057,N_38923);
nor U40568 (N_40568,N_35918,N_35371);
nor U40569 (N_40569,N_37967,N_38317);
nand U40570 (N_40570,N_37826,N_36268);
or U40571 (N_40571,N_36959,N_35333);
xor U40572 (N_40572,N_37143,N_36189);
nor U40573 (N_40573,N_37311,N_35213);
nand U40574 (N_40574,N_39940,N_35379);
or U40575 (N_40575,N_35529,N_37045);
nor U40576 (N_40576,N_35936,N_38818);
nor U40577 (N_40577,N_36791,N_39304);
nand U40578 (N_40578,N_37561,N_38904);
or U40579 (N_40579,N_38779,N_39446);
and U40580 (N_40580,N_37800,N_37244);
nand U40581 (N_40581,N_39874,N_37083);
nor U40582 (N_40582,N_37615,N_37512);
nand U40583 (N_40583,N_39124,N_35337);
nand U40584 (N_40584,N_35382,N_38894);
xor U40585 (N_40585,N_36456,N_38127);
and U40586 (N_40586,N_36894,N_37678);
or U40587 (N_40587,N_37065,N_36632);
nand U40588 (N_40588,N_36916,N_38083);
and U40589 (N_40589,N_37279,N_36616);
or U40590 (N_40590,N_38366,N_35622);
and U40591 (N_40591,N_39844,N_36935);
xor U40592 (N_40592,N_39297,N_35503);
xnor U40593 (N_40593,N_35427,N_36920);
nand U40594 (N_40594,N_37918,N_36079);
and U40595 (N_40595,N_36109,N_38617);
and U40596 (N_40596,N_39860,N_38802);
and U40597 (N_40597,N_38925,N_39754);
or U40598 (N_40598,N_38237,N_36638);
nor U40599 (N_40599,N_38049,N_37608);
nand U40600 (N_40600,N_37885,N_35028);
and U40601 (N_40601,N_39232,N_38133);
nand U40602 (N_40602,N_37883,N_36113);
xnor U40603 (N_40603,N_35725,N_38511);
or U40604 (N_40604,N_36358,N_38745);
nor U40605 (N_40605,N_37762,N_35280);
and U40606 (N_40606,N_35485,N_39031);
nor U40607 (N_40607,N_37845,N_36367);
nand U40608 (N_40608,N_35325,N_36669);
or U40609 (N_40609,N_35271,N_35012);
or U40610 (N_40610,N_37312,N_39559);
xnor U40611 (N_40611,N_36525,N_39235);
nor U40612 (N_40612,N_39982,N_35126);
or U40613 (N_40613,N_39083,N_35662);
or U40614 (N_40614,N_36242,N_39405);
nor U40615 (N_40615,N_35184,N_38075);
or U40616 (N_40616,N_35192,N_38901);
and U40617 (N_40617,N_36448,N_36543);
or U40618 (N_40618,N_36963,N_37648);
nand U40619 (N_40619,N_38023,N_35072);
nor U40620 (N_40620,N_38674,N_36292);
xnor U40621 (N_40621,N_37991,N_38581);
nand U40622 (N_40622,N_36173,N_35655);
or U40623 (N_40623,N_39253,N_37620);
or U40624 (N_40624,N_38010,N_39231);
nor U40625 (N_40625,N_36649,N_35129);
nand U40626 (N_40626,N_36261,N_37936);
and U40627 (N_40627,N_36593,N_35892);
nand U40628 (N_40628,N_35743,N_38219);
nor U40629 (N_40629,N_39238,N_37303);
nor U40630 (N_40630,N_35270,N_38920);
or U40631 (N_40631,N_39177,N_36634);
and U40632 (N_40632,N_36706,N_38008);
nor U40633 (N_40633,N_39749,N_38343);
xor U40634 (N_40634,N_35859,N_35793);
and U40635 (N_40635,N_37238,N_37669);
nand U40636 (N_40636,N_38091,N_38631);
xor U40637 (N_40637,N_36082,N_37300);
nor U40638 (N_40638,N_35998,N_36395);
and U40639 (N_40639,N_37290,N_39455);
and U40640 (N_40640,N_36380,N_39247);
or U40641 (N_40641,N_38441,N_39565);
nor U40642 (N_40642,N_36832,N_39333);
or U40643 (N_40643,N_37444,N_37821);
and U40644 (N_40644,N_39606,N_35762);
nand U40645 (N_40645,N_35674,N_38450);
or U40646 (N_40646,N_37251,N_36490);
or U40647 (N_40647,N_38485,N_36792);
nand U40648 (N_40648,N_38432,N_38194);
and U40649 (N_40649,N_35071,N_37207);
nor U40650 (N_40650,N_37626,N_39298);
or U40651 (N_40651,N_35568,N_37009);
nand U40652 (N_40652,N_38510,N_37091);
or U40653 (N_40653,N_38228,N_38738);
nor U40654 (N_40654,N_37756,N_35986);
nor U40655 (N_40655,N_37194,N_38476);
and U40656 (N_40656,N_38064,N_38043);
nor U40657 (N_40657,N_38247,N_38875);
and U40658 (N_40658,N_36563,N_35617);
or U40659 (N_40659,N_37775,N_36204);
nor U40660 (N_40660,N_39933,N_37017);
nand U40661 (N_40661,N_37742,N_38419);
nor U40662 (N_40662,N_35089,N_36120);
nand U40663 (N_40663,N_36066,N_36635);
or U40664 (N_40664,N_38079,N_35771);
nand U40665 (N_40665,N_38433,N_35051);
nand U40666 (N_40666,N_35835,N_38389);
nand U40667 (N_40667,N_37607,N_39573);
nor U40668 (N_40668,N_38214,N_35197);
or U40669 (N_40669,N_37900,N_39171);
nand U40670 (N_40670,N_39159,N_36332);
or U40671 (N_40671,N_38537,N_35975);
and U40672 (N_40672,N_39034,N_35917);
and U40673 (N_40673,N_39813,N_36847);
or U40674 (N_40674,N_36144,N_36420);
xnor U40675 (N_40675,N_36323,N_37270);
nand U40676 (N_40676,N_39669,N_37069);
or U40677 (N_40677,N_36212,N_38416);
and U40678 (N_40678,N_37992,N_36472);
nor U40679 (N_40679,N_36454,N_39423);
and U40680 (N_40680,N_39632,N_35722);
and U40681 (N_40681,N_39746,N_38259);
xnor U40682 (N_40682,N_35211,N_38950);
xor U40683 (N_40683,N_38827,N_35183);
and U40684 (N_40684,N_35074,N_39990);
nand U40685 (N_40685,N_39918,N_39536);
nor U40686 (N_40686,N_35199,N_38409);
xnor U40687 (N_40687,N_35135,N_36871);
nor U40688 (N_40688,N_35744,N_36191);
and U40689 (N_40689,N_35496,N_35943);
and U40690 (N_40690,N_39756,N_38804);
nor U40691 (N_40691,N_36734,N_35295);
and U40692 (N_40692,N_37483,N_36675);
or U40693 (N_40693,N_36922,N_36898);
or U40694 (N_40694,N_38592,N_35795);
or U40695 (N_40695,N_38406,N_37550);
nor U40696 (N_40696,N_36961,N_38287);
nor U40697 (N_40697,N_38900,N_39942);
nor U40698 (N_40698,N_37707,N_38699);
or U40699 (N_40699,N_38909,N_38186);
or U40700 (N_40700,N_37824,N_37817);
and U40701 (N_40701,N_39876,N_38890);
nor U40702 (N_40702,N_36240,N_39316);
nor U40703 (N_40703,N_37752,N_39885);
xnor U40704 (N_40704,N_35864,N_38508);
xor U40705 (N_40705,N_37324,N_36729);
nor U40706 (N_40706,N_35253,N_35890);
nand U40707 (N_40707,N_35403,N_39625);
nor U40708 (N_40708,N_38772,N_35857);
xnor U40709 (N_40709,N_36889,N_38046);
nor U40710 (N_40710,N_37090,N_38461);
xor U40711 (N_40711,N_36522,N_35061);
and U40712 (N_40712,N_37662,N_35027);
xor U40713 (N_40713,N_36755,N_38743);
nor U40714 (N_40714,N_36917,N_38503);
and U40715 (N_40715,N_39908,N_37517);
or U40716 (N_40716,N_39556,N_35491);
nor U40717 (N_40717,N_35092,N_39864);
or U40718 (N_40718,N_37685,N_36533);
or U40719 (N_40719,N_38349,N_38180);
nand U40720 (N_40720,N_35103,N_35701);
or U40721 (N_40721,N_38316,N_36165);
or U40722 (N_40722,N_39542,N_39820);
and U40723 (N_40723,N_38889,N_38142);
xnor U40724 (N_40724,N_36338,N_35688);
nand U40725 (N_40725,N_37641,N_36248);
and U40726 (N_40726,N_39593,N_38074);
or U40727 (N_40727,N_37379,N_36728);
or U40728 (N_40728,N_35690,N_38407);
xnor U40729 (N_40729,N_35893,N_39739);
or U40730 (N_40730,N_37499,N_37132);
nor U40731 (N_40731,N_35767,N_37807);
or U40732 (N_40732,N_39897,N_36186);
nand U40733 (N_40733,N_36271,N_36613);
xor U40734 (N_40734,N_35956,N_39889);
and U40735 (N_40735,N_37498,N_37217);
nor U40736 (N_40736,N_37896,N_39681);
or U40737 (N_40737,N_35712,N_36377);
nand U40738 (N_40738,N_39216,N_35648);
nor U40739 (N_40739,N_37573,N_38579);
xnor U40740 (N_40740,N_36089,N_37805);
and U40741 (N_40741,N_35037,N_38443);
and U40742 (N_40742,N_37057,N_36412);
or U40743 (N_40743,N_35876,N_36428);
or U40744 (N_40744,N_38902,N_38529);
or U40745 (N_40745,N_35038,N_39143);
nand U40746 (N_40746,N_39679,N_37809);
nand U40747 (N_40747,N_36468,N_37176);
or U40748 (N_40748,N_36756,N_37347);
nand U40749 (N_40749,N_35026,N_39846);
nor U40750 (N_40750,N_38839,N_39162);
nor U40751 (N_40751,N_38733,N_38587);
nand U40752 (N_40752,N_38442,N_39018);
nand U40753 (N_40753,N_37051,N_39489);
nor U40754 (N_40754,N_36091,N_38830);
nor U40755 (N_40755,N_38638,N_35388);
or U40756 (N_40756,N_38226,N_38190);
or U40757 (N_40757,N_36718,N_39126);
nand U40758 (N_40758,N_36828,N_36928);
and U40759 (N_40759,N_35267,N_38307);
xnor U40760 (N_40760,N_36622,N_39192);
and U40761 (N_40761,N_37131,N_38021);
xor U40762 (N_40762,N_37965,N_35531);
and U40763 (N_40763,N_37939,N_39385);
nand U40764 (N_40764,N_39538,N_35232);
xnor U40765 (N_40765,N_38990,N_35732);
nor U40766 (N_40766,N_38273,N_38786);
nor U40767 (N_40767,N_39070,N_37537);
xor U40768 (N_40768,N_35152,N_36037);
or U40769 (N_40769,N_35627,N_35895);
or U40770 (N_40770,N_36947,N_36698);
nand U40771 (N_40771,N_38408,N_37416);
nor U40772 (N_40772,N_35202,N_39642);
or U40773 (N_40773,N_38736,N_37012);
and U40774 (N_40774,N_35415,N_38848);
or U40775 (N_40775,N_35087,N_37365);
xor U40776 (N_40776,N_39241,N_38235);
xnor U40777 (N_40777,N_39599,N_36033);
and U40778 (N_40778,N_38029,N_37665);
or U40779 (N_40779,N_35042,N_35352);
and U40780 (N_40780,N_38654,N_39638);
nand U40781 (N_40781,N_38197,N_36672);
xor U40782 (N_40782,N_38767,N_38790);
and U40783 (N_40783,N_35984,N_37544);
nand U40784 (N_40784,N_37745,N_37088);
or U40785 (N_40785,N_38687,N_36312);
nor U40786 (N_40786,N_38370,N_36108);
nor U40787 (N_40787,N_39891,N_35868);
xor U40788 (N_40788,N_36614,N_35275);
xnor U40789 (N_40789,N_36435,N_36629);
nand U40790 (N_40790,N_38089,N_39925);
nand U40791 (N_40791,N_39748,N_38077);
nor U40792 (N_40792,N_39622,N_36860);
or U40793 (N_40793,N_35548,N_35134);
nand U40794 (N_40794,N_38168,N_37396);
nand U40795 (N_40795,N_35338,N_37601);
nor U40796 (N_40796,N_38668,N_36707);
xnor U40797 (N_40797,N_39527,N_37587);
or U40798 (N_40798,N_37331,N_36942);
nor U40799 (N_40799,N_35583,N_39707);
nand U40800 (N_40800,N_35342,N_37860);
xor U40801 (N_40801,N_37980,N_36589);
xnor U40802 (N_40802,N_36725,N_35412);
nor U40803 (N_40803,N_36319,N_39875);
or U40804 (N_40804,N_37766,N_35283);
nand U40805 (N_40805,N_36104,N_37198);
xor U40806 (N_40806,N_38290,N_39614);
or U40807 (N_40807,N_36138,N_39375);
and U40808 (N_40808,N_37445,N_36937);
nand U40809 (N_40809,N_39821,N_36039);
nor U40810 (N_40810,N_39511,N_37771);
and U40811 (N_40811,N_39189,N_38878);
and U40812 (N_40812,N_39438,N_36471);
or U40813 (N_40813,N_36288,N_35928);
xnor U40814 (N_40814,N_36259,N_37357);
and U40815 (N_40815,N_36566,N_38823);
xor U40816 (N_40816,N_38658,N_38059);
nor U40817 (N_40817,N_39351,N_36731);
or U40818 (N_40818,N_35784,N_37399);
nand U40819 (N_40819,N_39262,N_35729);
xnor U40820 (N_40820,N_39169,N_38336);
xor U40821 (N_40821,N_39462,N_35321);
or U40822 (N_40822,N_39296,N_38629);
xor U40823 (N_40823,N_39795,N_37205);
xor U40824 (N_40824,N_39760,N_36576);
nand U40825 (N_40825,N_36908,N_36679);
nand U40826 (N_40826,N_38480,N_36201);
nand U40827 (N_40827,N_35909,N_38491);
or U40828 (N_40828,N_37717,N_37275);
nor U40829 (N_40829,N_35845,N_35108);
nand U40830 (N_40830,N_37658,N_39597);
xnor U40831 (N_40831,N_39134,N_36016);
nand U40832 (N_40832,N_38861,N_37497);
and U40833 (N_40833,N_36840,N_36678);
nor U40834 (N_40834,N_35409,N_36912);
or U40835 (N_40835,N_37765,N_38765);
nor U40836 (N_40836,N_39117,N_38560);
nor U40837 (N_40837,N_35607,N_36789);
nand U40838 (N_40838,N_36226,N_37919);
nor U40839 (N_40839,N_37298,N_35707);
nor U40840 (N_40840,N_39444,N_36455);
or U40841 (N_40841,N_35658,N_36210);
nor U40842 (N_40842,N_38682,N_37625);
and U40843 (N_40843,N_36691,N_39400);
xnor U40844 (N_40844,N_35587,N_39714);
xor U40845 (N_40845,N_35780,N_35833);
xnor U40846 (N_40846,N_35257,N_38564);
nor U40847 (N_40847,N_35357,N_37699);
and U40848 (N_40848,N_35144,N_35676);
and U40849 (N_40849,N_39698,N_39340);
nor U40850 (N_40850,N_37340,N_36549);
xor U40851 (N_40851,N_38664,N_37579);
and U40852 (N_40852,N_38123,N_37403);
and U40853 (N_40853,N_37383,N_37342);
and U40854 (N_40854,N_37121,N_37636);
xnor U40855 (N_40855,N_35999,N_35003);
and U40856 (N_40856,N_38208,N_36667);
and U40857 (N_40857,N_35595,N_39488);
or U40858 (N_40858,N_38843,N_35196);
nand U40859 (N_40859,N_36003,N_39178);
nor U40860 (N_40860,N_36735,N_36714);
and U40861 (N_40861,N_39646,N_37695);
or U40862 (N_40862,N_36539,N_35223);
nor U40863 (N_40863,N_38308,N_36618);
nor U40864 (N_40864,N_35781,N_37767);
or U40865 (N_40865,N_35861,N_39858);
nor U40866 (N_40866,N_35643,N_36299);
xnor U40867 (N_40867,N_38858,N_39914);
or U40868 (N_40868,N_38447,N_35746);
and U40869 (N_40869,N_39140,N_37077);
or U40870 (N_40870,N_35542,N_39572);
and U40871 (N_40871,N_39890,N_36680);
or U40872 (N_40872,N_39980,N_39895);
xor U40873 (N_40873,N_35814,N_37725);
xor U40874 (N_40874,N_37583,N_38955);
nand U40875 (N_40875,N_36463,N_38807);
nand U40876 (N_40876,N_35783,N_37350);
or U40877 (N_40877,N_39492,N_38965);
and U40878 (N_40878,N_39946,N_36558);
or U40879 (N_40879,N_36551,N_36031);
xnor U40880 (N_40880,N_38048,N_39576);
nor U40881 (N_40881,N_38522,N_35950);
and U40882 (N_40882,N_39406,N_35190);
nand U40883 (N_40883,N_35452,N_37075);
nand U40884 (N_40884,N_38847,N_37204);
or U40885 (N_40885,N_35039,N_37815);
or U40886 (N_40886,N_38466,N_39943);
nor U40887 (N_40887,N_38527,N_37737);
nand U40888 (N_40888,N_36501,N_38517);
and U40889 (N_40889,N_36943,N_37158);
or U40890 (N_40890,N_37643,N_38305);
nand U40891 (N_40891,N_35289,N_37086);
and U40892 (N_40892,N_36899,N_36051);
or U40893 (N_40893,N_37705,N_36578);
and U40894 (N_40894,N_37529,N_38885);
or U40895 (N_40895,N_36595,N_36021);
nand U40896 (N_40896,N_35355,N_35122);
nor U40897 (N_40897,N_36118,N_36019);
nand U40898 (N_40898,N_38495,N_35002);
nand U40899 (N_40899,N_38887,N_37448);
xor U40900 (N_40900,N_39917,N_37346);
or U40901 (N_40901,N_37427,N_36950);
nand U40902 (N_40902,N_39752,N_36752);
and U40903 (N_40903,N_37747,N_39757);
xnor U40904 (N_40904,N_38573,N_35930);
xnor U40905 (N_40905,N_36487,N_38424);
and U40906 (N_40906,N_39312,N_37525);
or U40907 (N_40907,N_37229,N_39589);
nand U40908 (N_40908,N_39645,N_36888);
nand U40909 (N_40909,N_38453,N_35944);
nand U40910 (N_40910,N_35166,N_38730);
xor U40911 (N_40911,N_37219,N_38179);
or U40912 (N_40912,N_39145,N_36411);
or U40913 (N_40913,N_38329,N_38584);
nand U40914 (N_40914,N_37261,N_35476);
xor U40915 (N_40915,N_39089,N_39552);
and U40916 (N_40916,N_36213,N_39372);
nand U40917 (N_40917,N_38224,N_36153);
nor U40918 (N_40918,N_37887,N_36560);
and U40919 (N_40919,N_35156,N_36726);
nor U40920 (N_40920,N_38314,N_35920);
and U40921 (N_40921,N_35236,N_36655);
nor U40922 (N_40922,N_35545,N_37323);
and U40923 (N_40923,N_38886,N_35244);
nor U40924 (N_40924,N_35113,N_38174);
nor U40925 (N_40925,N_37781,N_36364);
or U40926 (N_40926,N_35478,N_35238);
or U40927 (N_40927,N_36873,N_38362);
nand U40928 (N_40928,N_37269,N_38044);
nand U40929 (N_40929,N_37946,N_36682);
xor U40930 (N_40930,N_36938,N_37474);
or U40931 (N_40931,N_37901,N_36819);
or U40932 (N_40932,N_35553,N_35080);
xor U40933 (N_40933,N_36194,N_39254);
xor U40934 (N_40934,N_37119,N_36557);
nor U40935 (N_40935,N_36492,N_39030);
xnor U40936 (N_40936,N_36351,N_38165);
xnor U40937 (N_40937,N_36224,N_39728);
nor U40938 (N_40938,N_38532,N_36926);
xor U40939 (N_40939,N_35926,N_36771);
nand U40940 (N_40940,N_37690,N_35990);
or U40941 (N_40941,N_38177,N_39215);
and U40942 (N_40942,N_35665,N_39626);
or U40943 (N_40943,N_38879,N_39722);
xnor U40944 (N_40944,N_38849,N_39533);
nor U40945 (N_40945,N_39383,N_35401);
or U40946 (N_40946,N_37559,N_39137);
and U40947 (N_40947,N_36974,N_38623);
and U40948 (N_40948,N_36310,N_35738);
and U40949 (N_40949,N_38225,N_36141);
and U40950 (N_40950,N_36673,N_35359);
or U40951 (N_40951,N_38382,N_38525);
and U40952 (N_40952,N_37877,N_38084);
or U40953 (N_40953,N_37683,N_38036);
and U40954 (N_40954,N_35254,N_38210);
or U40955 (N_40955,N_35010,N_38671);
or U40956 (N_40956,N_35747,N_38846);
nor U40957 (N_40957,N_37871,N_35057);
xnor U40958 (N_40958,N_38205,N_37784);
nor U40959 (N_40959,N_38523,N_39291);
and U40960 (N_40960,N_38803,N_38426);
nor U40961 (N_40961,N_36515,N_36264);
or U40962 (N_40962,N_37925,N_36837);
nand U40963 (N_40963,N_36156,N_36123);
xor U40964 (N_40964,N_35454,N_36012);
nor U40965 (N_40965,N_37227,N_38666);
xnor U40966 (N_40966,N_39931,N_36919);
or U40967 (N_40967,N_37033,N_35457);
nand U40968 (N_40968,N_39659,N_39164);
nor U40969 (N_40969,N_35145,N_37693);
nor U40970 (N_40970,N_37938,N_35527);
and U40971 (N_40971,N_38356,N_39753);
nor U40972 (N_40972,N_37686,N_37814);
nor U40973 (N_40973,N_35376,N_37840);
nand U40974 (N_40974,N_36739,N_38274);
or U40975 (N_40975,N_36128,N_38448);
and U40976 (N_40976,N_39249,N_35865);
nand U40977 (N_40977,N_37926,N_37644);
or U40978 (N_40978,N_35737,N_39798);
nand U40979 (N_40979,N_35558,N_35375);
xnor U40980 (N_40980,N_38114,N_39856);
or U40981 (N_40981,N_37640,N_37164);
nand U40982 (N_40982,N_37259,N_37334);
nor U40983 (N_40983,N_37700,N_39069);
xor U40984 (N_40984,N_37507,N_37056);
or U40985 (N_40985,N_38844,N_35335);
nand U40986 (N_40986,N_39567,N_37609);
nor U40987 (N_40987,N_37701,N_37410);
or U40988 (N_40988,N_36783,N_39720);
or U40989 (N_40989,N_35507,N_36074);
or U40990 (N_40990,N_38111,N_38330);
nor U40991 (N_40991,N_39154,N_36125);
nor U40992 (N_40992,N_39854,N_37792);
nor U40993 (N_40993,N_36000,N_37105);
nor U40994 (N_40994,N_39093,N_36897);
nor U40995 (N_40995,N_38090,N_39787);
xnor U40996 (N_40996,N_39193,N_37320);
nand U40997 (N_40997,N_35925,N_36467);
nand U40998 (N_40998,N_35742,N_35109);
xnor U40999 (N_40999,N_39671,N_37855);
nor U41000 (N_41000,N_39053,N_36966);
or U41001 (N_41001,N_38708,N_36556);
nand U41002 (N_41002,N_39233,N_39649);
xor U41003 (N_41003,N_36982,N_36570);
nand U41004 (N_41004,N_39021,N_36663);
nand U41005 (N_41005,N_38276,N_36716);
and U41006 (N_41006,N_39938,N_35245);
or U41007 (N_41007,N_39721,N_39901);
xnor U41008 (N_41008,N_36825,N_37848);
and U41009 (N_41009,N_35341,N_37180);
xnor U41010 (N_41010,N_35830,N_37473);
nand U41011 (N_41011,N_37007,N_35794);
xor U41012 (N_41012,N_39483,N_36896);
nor U41013 (N_41013,N_37962,N_37407);
nand U41014 (N_41014,N_39705,N_36856);
xor U41015 (N_41015,N_37642,N_39906);
nand U41016 (N_41016,N_36995,N_36662);
nor U41017 (N_41017,N_35934,N_38117);
or U41018 (N_41018,N_38268,N_39285);
xnor U41019 (N_41019,N_36750,N_38014);
or U41020 (N_41020,N_35723,N_36409);
nor U41021 (N_41021,N_37982,N_35248);
or U41022 (N_41022,N_37230,N_38796);
nor U41023 (N_41023,N_38054,N_36136);
nand U41024 (N_41024,N_37240,N_39972);
nand U41025 (N_41025,N_36841,N_39086);
and U41026 (N_41026,N_38289,N_37545);
nor U41027 (N_41027,N_38899,N_37060);
xor U41028 (N_41028,N_36437,N_38005);
or U41029 (N_41029,N_35721,N_35302);
or U41030 (N_41030,N_37459,N_39421);
xor U41031 (N_41031,N_36939,N_38159);
or U41032 (N_41032,N_36524,N_35250);
and U41033 (N_41033,N_35666,N_38655);
and U41034 (N_41034,N_37710,N_35911);
and U41035 (N_41035,N_38203,N_37612);
nand U41036 (N_41036,N_36986,N_38916);
and U41037 (N_41037,N_37030,N_38494);
nand U41038 (N_41038,N_38429,N_39113);
or U41039 (N_41039,N_36992,N_37481);
nand U41040 (N_41040,N_38766,N_35035);
and U41041 (N_41041,N_37130,N_35014);
and U41042 (N_41042,N_35132,N_37493);
and U41043 (N_41043,N_37664,N_38991);
and U41044 (N_41044,N_36370,N_36433);
nor U41045 (N_41045,N_35589,N_35366);
nor U41046 (N_41046,N_38926,N_35524);
nand U41047 (N_41047,N_35397,N_38109);
nand U41048 (N_41048,N_35997,N_38000);
nand U41049 (N_41049,N_35929,N_37754);
xnor U41050 (N_41050,N_37315,N_39101);
nand U41051 (N_41051,N_37870,N_37368);
xnor U41052 (N_41052,N_39487,N_38528);
xnor U41053 (N_41053,N_39992,N_35048);
nand U41054 (N_41054,N_39230,N_35995);
and U41055 (N_41055,N_35816,N_36764);
and U41056 (N_41056,N_39678,N_36058);
or U41057 (N_41057,N_36149,N_38988);
or U41058 (N_41058,N_36498,N_36276);
nor U41059 (N_41059,N_38748,N_38022);
or U41060 (N_41060,N_39244,N_37402);
and U41061 (N_41061,N_39010,N_38383);
and U41062 (N_41062,N_37603,N_38166);
or U41063 (N_41063,N_37592,N_39939);
or U41064 (N_41064,N_38221,N_35319);
nand U41065 (N_41065,N_36402,N_35994);
nor U41066 (N_41066,N_35475,N_39600);
xnor U41067 (N_41067,N_38204,N_36485);
xnor U41068 (N_41068,N_35904,N_39023);
xnor U41069 (N_41069,N_36948,N_35446);
and U41070 (N_41070,N_35603,N_39737);
nor U41071 (N_41071,N_39219,N_35344);
or U41072 (N_41072,N_38507,N_36179);
xnor U41073 (N_41073,N_38160,N_35084);
xor U41074 (N_41074,N_39360,N_39373);
nand U41075 (N_41075,N_37760,N_37774);
and U41076 (N_41076,N_38361,N_36559);
nand U41077 (N_41077,N_37294,N_35204);
xor U41078 (N_41078,N_37201,N_37928);
and U41079 (N_41079,N_38762,N_39568);
nand U41080 (N_41080,N_39811,N_39519);
xnor U41081 (N_41081,N_36257,N_36875);
or U41082 (N_41082,N_37798,N_35623);
and U41083 (N_41083,N_36657,N_37882);
and U41084 (N_41084,N_35467,N_37046);
nor U41085 (N_41085,N_39172,N_37267);
xnor U41086 (N_41086,N_35809,N_35941);
or U41087 (N_41087,N_35154,N_39252);
or U41088 (N_41088,N_36906,N_38634);
nor U41089 (N_41089,N_35534,N_36416);
xor U41090 (N_41090,N_36803,N_36085);
and U41091 (N_41091,N_39354,N_38295);
or U41092 (N_41092,N_35576,N_35687);
or U41093 (N_41093,N_37284,N_35931);
xnor U41094 (N_41094,N_39870,N_36744);
nor U41095 (N_41095,N_35874,N_36098);
xor U41096 (N_41096,N_35495,N_39505);
nor U41097 (N_41097,N_37950,N_37787);
nand U41098 (N_41098,N_38384,N_36617);
nand U41099 (N_41099,N_36084,N_37479);
and U41100 (N_41100,N_39562,N_38116);
nor U41101 (N_41101,N_36385,N_38201);
and U41102 (N_41102,N_38594,N_39440);
and U41103 (N_41103,N_39447,N_36260);
nand U41104 (N_41104,N_35400,N_36866);
and U41105 (N_41105,N_35656,N_36775);
nor U41106 (N_41106,N_39516,N_36289);
or U41107 (N_41107,N_35115,N_38173);
and U41108 (N_41108,N_36733,N_39779);
nor U41109 (N_41109,N_39690,N_36413);
nand U41110 (N_41110,N_37923,N_36564);
and U41111 (N_41111,N_39214,N_37843);
or U41112 (N_41112,N_38749,N_39067);
and U41113 (N_41113,N_35450,N_36526);
and U41114 (N_41114,N_37355,N_36228);
nor U41115 (N_41115,N_37114,N_35214);
xnor U41116 (N_41116,N_35130,N_38728);
nand U41117 (N_41117,N_38614,N_36510);
nand U41118 (N_41118,N_39851,N_36921);
and U41119 (N_41119,N_35354,N_38561);
nor U41120 (N_41120,N_35638,N_36330);
and U41121 (N_41121,N_36858,N_36103);
nand U41122 (N_41122,N_39074,N_36577);
xor U41123 (N_41123,N_35024,N_39345);
nor U41124 (N_41124,N_39246,N_36466);
nor U41125 (N_41125,N_39006,N_35022);
nand U41126 (N_41126,N_36504,N_39226);
nand U41127 (N_41127,N_39598,N_35404);
xor U41128 (N_41128,N_35933,N_38492);
or U41129 (N_41129,N_38354,N_37018);
xor U41130 (N_41130,N_38816,N_37139);
nand U41131 (N_41131,N_37602,N_37157);
nor U41132 (N_41132,N_39745,N_36727);
and U41133 (N_41133,N_39882,N_38656);
or U41134 (N_41134,N_35695,N_39012);
and U41135 (N_41135,N_36116,N_39957);
xor U41136 (N_41136,N_38590,N_36683);
nand U41137 (N_41137,N_36838,N_35512);
or U41138 (N_41138,N_36527,N_36460);
nand U41139 (N_41139,N_36811,N_37652);
xnor U41140 (N_41140,N_35992,N_35471);
and U41141 (N_41141,N_37940,N_37035);
or U41142 (N_41142,N_37263,N_39496);
nor U41143 (N_41143,N_38192,N_39574);
xor U41144 (N_41144,N_35339,N_38028);
nor U41145 (N_41145,N_38698,N_37235);
and U41146 (N_41146,N_36234,N_37295);
xnor U41147 (N_41147,N_37184,N_38619);
or U41148 (N_41148,N_35148,N_35642);
nand U41149 (N_41149,N_37831,N_37170);
nand U41150 (N_41150,N_36441,N_35015);
xor U41151 (N_41151,N_35983,N_35413);
or U41152 (N_41152,N_37451,N_37359);
and U41153 (N_41153,N_37440,N_39631);
xnor U41154 (N_41154,N_36474,N_35749);
nand U41155 (N_41155,N_36070,N_35350);
xnor U41156 (N_41156,N_39959,N_38018);
or U41157 (N_41157,N_36690,N_37931);
nand U41158 (N_41158,N_39508,N_36759);
nand U41159 (N_41159,N_39217,N_36529);
nand U41160 (N_41160,N_39149,N_38834);
nand U41161 (N_41161,N_39608,N_37374);
or U41162 (N_41162,N_39958,N_38050);
and U41163 (N_41163,N_37276,N_37084);
xor U41164 (N_41164,N_36137,N_36045);
nand U41165 (N_41165,N_38723,N_39848);
nand U41166 (N_41166,N_36571,N_35891);
and U41167 (N_41167,N_35862,N_36989);
nand U41168 (N_41168,N_38001,N_37942);
and U41169 (N_41169,N_36903,N_38456);
and U41170 (N_41170,N_36877,N_37063);
or U41171 (N_41171,N_35422,N_37584);
nand U41172 (N_41172,N_36376,N_35584);
or U41173 (N_41173,N_38435,N_35081);
nand U41174 (N_41174,N_38327,N_39277);
or U41175 (N_41175,N_38331,N_35235);
xnor U41176 (N_41176,N_36833,N_38047);
nand U41177 (N_41177,N_39814,N_38033);
nor U41178 (N_41178,N_35112,N_38332);
nand U41179 (N_41179,N_38625,N_36119);
or U41180 (N_41180,N_35616,N_36981);
nor U41181 (N_41181,N_39768,N_38315);
xor U41182 (N_41182,N_36626,N_38425);
or U41183 (N_41183,N_35555,N_37673);
xnor U41184 (N_41184,N_36301,N_35916);
nor U41185 (N_41185,N_38242,N_35610);
and U41186 (N_41186,N_38992,N_38178);
nand U41187 (N_41187,N_38530,N_38410);
and U41188 (N_41188,N_38138,N_35025);
or U41189 (N_41189,N_36333,N_37866);
nor U41190 (N_41190,N_38960,N_35806);
nand U41191 (N_41191,N_38239,N_38438);
nand U41192 (N_41192,N_37724,N_37851);
nor U41193 (N_41193,N_39834,N_37797);
nor U41194 (N_41194,N_38769,N_39644);
or U41195 (N_41195,N_39823,N_38041);
and U41196 (N_41196,N_38148,N_37152);
nand U41197 (N_41197,N_39610,N_36692);
nand U41198 (N_41198,N_36870,N_38175);
or U41199 (N_41199,N_35304,N_37915);
or U41200 (N_41200,N_38188,N_39969);
nand U41201 (N_41201,N_38600,N_35434);
nand U41202 (N_41202,N_37907,N_39161);
xor U41203 (N_41203,N_38430,N_35408);
xnor U41204 (N_41204,N_37684,N_35685);
xnor U41205 (N_41205,N_36022,N_35573);
nand U41206 (N_41206,N_36636,N_35813);
or U41207 (N_41207,N_35565,N_37913);
xor U41208 (N_41208,N_35098,N_39903);
and U41209 (N_41209,N_35966,N_37890);
and U41210 (N_41210,N_39365,N_36247);
xnor U41211 (N_41211,N_37734,N_35670);
nand U41212 (N_41212,N_38238,N_39138);
nor U41213 (N_41213,N_36687,N_35443);
nor U41214 (N_41214,N_35182,N_35730);
nor U41215 (N_41215,N_39328,N_36848);
and U41216 (N_41216,N_38921,N_37952);
nor U41217 (N_41217,N_36392,N_36538);
and U41218 (N_41218,N_37874,N_39601);
nor U41219 (N_41219,N_36168,N_38531);
and U41220 (N_41220,N_37129,N_36765);
or U41221 (N_41221,N_35764,N_38241);
nand U41222 (N_41222,N_35855,N_35314);
and U41223 (N_41223,N_35086,N_36347);
and U41224 (N_41224,N_36017,N_35592);
xnor U41225 (N_41225,N_39482,N_37777);
nor U41226 (N_41226,N_35785,N_37373);
nand U41227 (N_41227,N_39087,N_38421);
nor U41228 (N_41228,N_37661,N_35073);
nor U41229 (N_41229,N_36094,N_38423);
nor U41230 (N_41230,N_37536,N_38189);
nor U41231 (N_41231,N_35686,N_37716);
xnor U41232 (N_41232,N_39457,N_38554);
nor U41233 (N_41233,N_37213,N_37193);
and U41234 (N_41234,N_37172,N_36399);
xnor U41235 (N_41235,N_36823,N_39611);
nand U41236 (N_41236,N_35090,N_35819);
or U41237 (N_41237,N_35758,N_38007);
or U41238 (N_41238,N_35241,N_38229);
and U41239 (N_41239,N_35840,N_39082);
and U41240 (N_41240,N_36573,N_37367);
or U41241 (N_41241,N_35155,N_35774);
and U41242 (N_41242,N_38446,N_35575);
nand U41243 (N_41243,N_39427,N_39783);
nor U41244 (N_41244,N_35562,N_38271);
and U41245 (N_41245,N_36685,N_39038);
xor U41246 (N_41246,N_38115,N_37523);
nand U41247 (N_41247,N_38270,N_38943);
or U41248 (N_41248,N_38292,N_37344);
nand U41249 (N_41249,N_39167,N_35841);
or U41250 (N_41250,N_35494,N_37309);
nand U41251 (N_41251,N_39603,N_38283);
and U41252 (N_41252,N_35451,N_38037);
nor U41253 (N_41253,N_35552,N_38368);
nand U41254 (N_41254,N_37167,N_37505);
and U41255 (N_41255,N_36859,N_36166);
nor U41256 (N_41256,N_39309,N_37975);
or U41257 (N_41257,N_38800,N_38641);
nand U41258 (N_41258,N_38637,N_37471);
and U41259 (N_41259,N_36171,N_39947);
and U41260 (N_41260,N_37956,N_39911);
nand U41261 (N_41261,N_37924,N_39907);
nor U41262 (N_41262,N_38200,N_36713);
nor U41263 (N_41263,N_39697,N_36619);
xnor U41264 (N_41264,N_39353,N_39040);
or U41265 (N_41265,N_35540,N_39912);
nor U41266 (N_41266,N_39761,N_37613);
nand U41267 (N_41267,N_37378,N_36405);
or U41268 (N_41268,N_38306,N_35378);
and U41269 (N_41269,N_39448,N_36813);
xnor U41270 (N_41270,N_38404,N_37406);
and U41271 (N_41271,N_35021,N_38318);
or U41272 (N_41272,N_38876,N_38826);
nand U41273 (N_41273,N_36627,N_36697);
and U41274 (N_41274,N_37600,N_39667);
xor U41275 (N_41275,N_38520,N_39434);
or U41276 (N_41276,N_37712,N_38893);
nor U41277 (N_41277,N_38874,N_35620);
nand U41278 (N_41278,N_36605,N_38296);
nand U41279 (N_41279,N_37905,N_37744);
xnor U41280 (N_41280,N_36132,N_37786);
nand U41281 (N_41281,N_39613,N_35414);
nand U41282 (N_41282,N_38056,N_36424);
xnor U41283 (N_41283,N_35818,N_37053);
nor U41284 (N_41284,N_37841,N_35669);
xor U41285 (N_41285,N_36417,N_37829);
nand U41286 (N_41286,N_37590,N_38357);
and U41287 (N_41287,N_35278,N_38552);
nor U41288 (N_41288,N_39735,N_38143);
or U41289 (N_41289,N_38167,N_38707);
nand U41290 (N_41290,N_37929,N_35581);
nor U41291 (N_41291,N_37482,N_37345);
or U41292 (N_41292,N_39153,N_35316);
or U41293 (N_41293,N_37677,N_39831);
nand U41294 (N_41294,N_35606,N_35262);
and U41295 (N_41295,N_36709,N_38566);
nor U41296 (N_41296,N_36475,N_38911);
nand U41297 (N_41297,N_36427,N_37430);
nor U41298 (N_41298,N_38953,N_38932);
nand U41299 (N_41299,N_39928,N_35077);
nor U41300 (N_41300,N_36964,N_35174);
or U41301 (N_41301,N_37089,N_37118);
and U41302 (N_41302,N_35883,N_39709);
and U41303 (N_41303,N_38147,N_38864);
xnor U41304 (N_41304,N_37031,N_38526);
and U41305 (N_41305,N_36161,N_36777);
nor U41306 (N_41306,N_36198,N_39952);
or U41307 (N_41307,N_36544,N_35279);
nand U41308 (N_41308,N_38484,N_35611);
or U41309 (N_41309,N_39788,N_36258);
or U41310 (N_41310,N_38003,N_36237);
xnor U41311 (N_41311,N_36304,N_38006);
nor U41312 (N_41312,N_37178,N_37531);
nor U41313 (N_41313,N_38475,N_36164);
and U41314 (N_41314,N_35007,N_39987);
xnor U41315 (N_41315,N_35125,N_37679);
or U41316 (N_41316,N_37458,N_38154);
xnor U41317 (N_41317,N_37998,N_37232);
and U41318 (N_41318,N_35066,N_38402);
or U41319 (N_41319,N_35639,N_35194);
and U41320 (N_41320,N_37541,N_38977);
and U41321 (N_41321,N_37577,N_38076);
nor U41322 (N_41322,N_39643,N_36666);
or U41323 (N_41323,N_37245,N_38795);
nand U41324 (N_41324,N_35149,N_37124);
or U41325 (N_41325,N_35546,N_37554);
xnor U41326 (N_41326,N_35822,N_39564);
xor U41327 (N_41327,N_38754,N_39314);
nand U41328 (N_41328,N_37776,N_38207);
nor U41329 (N_41329,N_39368,N_37949);
or U41330 (N_41330,N_37691,N_35528);
nand U41331 (N_41331,N_36598,N_38244);
xnor U41332 (N_41332,N_35000,N_36907);
xnor U41333 (N_41333,N_39381,N_37633);
and U41334 (N_41334,N_37783,N_39767);
nor U41335 (N_41335,N_38521,N_37236);
and U41336 (N_41336,N_37052,N_38379);
xnor U41337 (N_41337,N_35405,N_36152);
and U41338 (N_41338,N_35683,N_39364);
nand U41339 (N_41339,N_35699,N_39796);
nand U41340 (N_41340,N_39945,N_39808);
nor U41341 (N_41341,N_39315,N_38472);
nor U41342 (N_41342,N_36689,N_39544);
or U41343 (N_41343,N_36404,N_38995);
nor U41344 (N_41344,N_36717,N_37572);
nor U41345 (N_41345,N_37450,N_35858);
xor U41346 (N_41346,N_38104,N_39076);
or U41347 (N_41347,N_35677,N_39061);
xnor U41348 (N_41348,N_38967,N_37418);
or U41349 (N_41349,N_35613,N_38172);
or U41350 (N_41350,N_39545,N_39146);
or U41351 (N_41351,N_38639,N_38724);
or U41352 (N_41352,N_39657,N_35812);
nand U41353 (N_41353,N_36421,N_39630);
nand U41354 (N_41354,N_36142,N_37788);
nand U41355 (N_41355,N_35559,N_37629);
nor U41356 (N_41356,N_38908,N_37111);
xnor U41357 (N_41357,N_38574,N_35402);
nor U41358 (N_41358,N_38794,N_36162);
xor U41359 (N_41359,N_36076,N_35323);
nand U41360 (N_41360,N_37358,N_35127);
nand U41361 (N_41361,N_35187,N_37649);
xor U41362 (N_41362,N_39514,N_37149);
xor U41363 (N_41363,N_39741,N_38182);
xor U41364 (N_41364,N_37316,N_38706);
nand U41365 (N_41365,N_39546,N_39104);
xnor U41366 (N_41366,N_36602,N_36703);
xor U41367 (N_41367,N_36408,N_35949);
nor U41368 (N_41368,N_36453,N_36770);
xnor U41369 (N_41369,N_35777,N_39997);
or U41370 (N_41370,N_38873,N_36357);
and U41371 (N_41371,N_39672,N_38100);
nand U41372 (N_41372,N_36249,N_39592);
nor U41373 (N_41373,N_36102,N_36407);
and U41374 (N_41374,N_39443,N_36369);
nand U41375 (N_41375,N_38686,N_37476);
xnor U41376 (N_41376,N_38700,N_35329);
or U41377 (N_41377,N_38813,N_37830);
and U41378 (N_41378,N_35872,N_36586);
nand U41379 (N_41379,N_35442,N_38548);
or U41380 (N_41380,N_36211,N_37516);
nor U41381 (N_41381,N_38157,N_36815);
nand U41382 (N_41382,N_35702,N_39935);
nor U41383 (N_41383,N_35058,N_36596);
and U41384 (N_41384,N_36449,N_37457);
nand U41385 (N_41385,N_38742,N_36990);
and U41386 (N_41386,N_39803,N_35888);
xor U41387 (N_41387,N_36568,N_39791);
nand U41388 (N_41388,N_37362,N_35560);
and U41389 (N_41389,N_39002,N_35564);
nor U41390 (N_41390,N_39605,N_36702);
or U41391 (N_41391,N_36390,N_37509);
and U41392 (N_41392,N_38261,N_38993);
nand U41393 (N_41393,N_36500,N_35381);
nand U41394 (N_41394,N_38613,N_38436);
and U41395 (N_41395,N_39174,N_39515);
or U41396 (N_41396,N_36112,N_39843);
xor U41397 (N_41397,N_37638,N_39330);
or U41398 (N_41398,N_37246,N_35299);
or U41399 (N_41399,N_38944,N_38585);
or U41400 (N_41400,N_36056,N_36579);
nor U41401 (N_41401,N_38098,N_36327);
or U41402 (N_41402,N_36520,N_39628);
and U41403 (N_41403,N_39983,N_39377);
nand U41404 (N_41404,N_35757,N_35566);
xor U41405 (N_41405,N_39407,N_39832);
nor U41406 (N_41406,N_36893,N_38058);
nand U41407 (N_41407,N_39893,N_35884);
nand U41408 (N_41408,N_36342,N_36398);
xor U41409 (N_41409,N_35297,N_37704);
nor U41410 (N_41410,N_36851,N_36633);
and U41411 (N_41411,N_37456,N_38897);
nor U41412 (N_41412,N_36436,N_37468);
xor U41413 (N_41413,N_36097,N_37922);
nor U41414 (N_41414,N_39165,N_36163);
or U41415 (N_41415,N_39713,N_39311);
xor U41416 (N_41416,N_39680,N_36531);
xnor U41417 (N_41417,N_38715,N_38371);
and U41418 (N_41418,N_36781,N_36205);
xor U41419 (N_41419,N_35612,N_35320);
nand U41420 (N_41420,N_35486,N_35468);
nand U41421 (N_41421,N_38970,N_38158);
xor U41422 (N_41422,N_39158,N_38547);
nor U41423 (N_41423,N_35680,N_35047);
or U41424 (N_41424,N_38234,N_37381);
and U41425 (N_41425,N_38497,N_37055);
nor U41426 (N_41426,N_37206,N_35497);
or U41427 (N_41427,N_39453,N_36230);
and U41428 (N_41428,N_39464,N_37994);
nand U41429 (N_41429,N_39883,N_36291);
xnor U41430 (N_41430,N_38859,N_36604);
and U41431 (N_41431,N_35273,N_36458);
or U41432 (N_41432,N_38927,N_38557);
and U41433 (N_41433,N_38391,N_35140);
nand U41434 (N_41434,N_39953,N_38694);
xor U41435 (N_41435,N_39586,N_37811);
or U41436 (N_41436,N_39676,N_35110);
and U41437 (N_41437,N_38599,N_38860);
and U41438 (N_41438,N_38434,N_38722);
xor U41439 (N_41439,N_39955,N_37477);
nor U41440 (N_41440,N_37387,N_37127);
nand U41441 (N_41441,N_38808,N_37394);
and U41442 (N_41442,N_37256,N_37469);
nand U41443 (N_41443,N_39118,N_39039);
xnor U41444 (N_41444,N_36223,N_39981);
or U41445 (N_41445,N_36799,N_38420);
or U41446 (N_41446,N_37472,N_39465);
nand U41447 (N_41447,N_39437,N_37003);
or U41448 (N_41448,N_36583,N_36465);
nor U41449 (N_41449,N_36046,N_37656);
xnor U41450 (N_41450,N_38612,N_36180);
and U41451 (N_41451,N_37504,N_39528);
or U41452 (N_41452,N_36592,N_36769);
nand U41453 (N_41453,N_35055,N_38066);
xor U41454 (N_41454,N_35640,N_39615);
xnor U41455 (N_41455,N_35863,N_39654);
nand U41456 (N_41456,N_39623,N_36652);
xnor U41457 (N_41457,N_35399,N_36372);
and U41458 (N_41458,N_37140,N_39744);
nor U41459 (N_41459,N_38220,N_36233);
nor U41460 (N_41460,N_36901,N_36375);
xnor U41461 (N_41461,N_38636,N_38777);
nor U41462 (N_41462,N_39786,N_37287);
or U41463 (N_41463,N_36317,N_39451);
or U41464 (N_41464,N_36386,N_37884);
and U41465 (N_41465,N_36059,N_38646);
nand U41466 (N_41466,N_36241,N_36816);
xnor U41467 (N_41467,N_38928,N_35520);
or U41468 (N_41468,N_38877,N_35101);
nand U41469 (N_41469,N_39726,N_35979);
nor U41470 (N_41470,N_35967,N_39486);
nor U41471 (N_41471,N_38067,N_39380);
nand U41472 (N_41472,N_39621,N_35973);
nand U41473 (N_41473,N_38065,N_37079);
xor U41474 (N_41474,N_36640,N_39696);
nand U41475 (N_41475,N_38870,N_35976);
and U41476 (N_41476,N_35910,N_38380);
xnor U41477 (N_41477,N_37141,N_35667);
or U41478 (N_41478,N_36488,N_38153);
xor U41479 (N_41479,N_38719,N_39971);
or U41480 (N_41480,N_39913,N_35632);
and U41481 (N_41481,N_37478,N_38954);
nand U41482 (N_41482,N_39639,N_35508);
nor U41483 (N_41483,N_37096,N_36272);
xnor U41484 (N_41484,N_36001,N_36738);
or U41485 (N_41485,N_39306,N_37337);
and U41486 (N_41486,N_36303,N_36513);
or U41487 (N_41487,N_38969,N_38412);
nor U41488 (N_41488,N_35085,N_35193);
or U41489 (N_41489,N_39075,N_38918);
nand U41490 (N_41490,N_35898,N_36107);
and U41491 (N_41491,N_36585,N_37736);
and U41492 (N_41492,N_39335,N_39839);
nor U41493 (N_41493,N_37277,N_39585);
nor U41494 (N_41494,N_39493,N_37154);
xor U41495 (N_41495,N_38359,N_35097);
and U41496 (N_41496,N_39522,N_36554);
xnor U41497 (N_41497,N_37739,N_39166);
nor U41498 (N_41498,N_35243,N_36493);
or U41499 (N_41499,N_35974,N_39736);
and U41500 (N_41500,N_37044,N_36235);
and U41501 (N_41501,N_39432,N_36207);
xor U41502 (N_41502,N_35550,N_36140);
or U41503 (N_41503,N_36814,N_39080);
or U41504 (N_41504,N_36865,N_35306);
nand U41505 (N_41505,N_36134,N_39210);
xnor U41506 (N_41506,N_36615,N_38095);
nor U41507 (N_41507,N_38347,N_35411);
nor U41508 (N_41508,N_37979,N_37506);
nor U41509 (N_41509,N_37351,N_35188);
xnor U41510 (N_41510,N_38852,N_37634);
nor U41511 (N_41511,N_36020,N_35393);
nand U41512 (N_41512,N_35317,N_35867);
xnor U41513 (N_41513,N_37987,N_38002);
xor U41514 (N_41514,N_39474,N_39655);
nand U41515 (N_41515,N_39932,N_38603);
nand U41516 (N_41516,N_39295,N_39127);
nor U41517 (N_41517,N_35820,N_37405);
or U41518 (N_41518,N_37954,N_36597);
nand U41519 (N_41519,N_37253,N_36932);
and U41520 (N_41520,N_39703,N_37533);
or U41521 (N_41521,N_35501,N_36671);
nand U41522 (N_41522,N_35169,N_36958);
nor U41523 (N_41523,N_39965,N_38661);
or U41524 (N_41524,N_37709,N_36910);
xor U41525 (N_41525,N_37558,N_35748);
nor U41526 (N_41526,N_39476,N_36129);
nand U41527 (N_41527,N_36350,N_35694);
nor U41528 (N_41528,N_36187,N_38375);
or U41529 (N_41529,N_35456,N_37564);
xor U41530 (N_41530,N_39989,N_38328);
nor U41531 (N_41531,N_36630,N_35769);
nor U41532 (N_41532,N_35631,N_36699);
or U41533 (N_41533,N_36438,N_36311);
nor U41534 (N_41534,N_36065,N_35823);
and U41535 (N_41535,N_35619,N_39763);
nor U41536 (N_41536,N_35856,N_36057);
nor U41537 (N_41537,N_38468,N_35535);
or U41538 (N_41538,N_36244,N_39190);
nand U41539 (N_41539,N_38110,N_38181);
nor U41540 (N_41540,N_36273,N_39693);
xnor U41541 (N_41541,N_38103,N_38814);
nand U41542 (N_41542,N_37064,N_35597);
xor U41543 (N_41543,N_37486,N_37491);
xnor U41544 (N_41544,N_38285,N_37876);
and U41545 (N_41545,N_37631,N_37067);
nor U41546 (N_41546,N_39641,N_37995);
or U41547 (N_41547,N_37366,N_39504);
xor U41548 (N_41548,N_37437,N_39033);
and U41549 (N_41549,N_38648,N_38635);
nand U41550 (N_41550,N_39341,N_38223);
and U41551 (N_41551,N_38679,N_37173);
xor U41552 (N_41552,N_39027,N_35921);
or U41553 (N_41553,N_35484,N_36625);
and U41554 (N_41554,N_38831,N_35885);
nand U41555 (N_41555,N_35770,N_39467);
nor U41556 (N_41556,N_36446,N_36345);
nor U41557 (N_41557,N_35421,N_38387);
xnor U41558 (N_41558,N_37034,N_38506);
or U41559 (N_41559,N_36489,N_36336);
xnor U41560 (N_41560,N_35298,N_37892);
and U41561 (N_41561,N_39399,N_36660);
nand U41562 (N_41562,N_38850,N_36892);
xnor U41563 (N_41563,N_37192,N_38102);
nor U41564 (N_41564,N_38726,N_38692);
xor U41565 (N_41565,N_38855,N_38669);
or U41566 (N_41566,N_39475,N_38572);
and U41567 (N_41567,N_36275,N_35641);
xor U41568 (N_41568,N_39861,N_35431);
xor U41569 (N_41569,N_39133,N_37868);
nor U41570 (N_41570,N_39961,N_39841);
nand U41571 (N_41571,N_38096,N_38978);
and U41572 (N_41572,N_36483,N_39207);
or U41573 (N_41573,N_39607,N_36010);
xnor U41574 (N_41574,N_35161,N_37825);
and U41575 (N_41575,N_39636,N_37218);
or U41576 (N_41576,N_38072,N_36073);
or U41577 (N_41577,N_39923,N_35111);
or U41578 (N_41578,N_39900,N_35121);
nor U41579 (N_41579,N_39976,N_38140);
nor U41580 (N_41580,N_37878,N_36007);
or U41581 (N_41581,N_38750,N_38607);
nand U41582 (N_41582,N_38556,N_36182);
and U41583 (N_41583,N_37614,N_39789);
nor U41584 (N_41584,N_35307,N_39802);
nand U41585 (N_41585,N_37790,N_39350);
xnor U41586 (N_41586,N_36052,N_39273);
or U41587 (N_41587,N_38632,N_38903);
xor U41588 (N_41588,N_38609,N_37097);
xor U41589 (N_41589,N_38533,N_35240);
xor U41590 (N_41590,N_36218,N_38559);
or U41591 (N_41591,N_39743,N_36883);
xor U41592 (N_41592,N_36684,N_36393);
nand U41593 (N_41593,N_38088,N_38107);
nor U41594 (N_41594,N_37768,N_36042);
nand U41595 (N_41595,N_36955,N_35009);
or U41596 (N_41596,N_37093,N_39094);
nor U41597 (N_41597,N_39382,N_35593);
nor U41598 (N_41598,N_36255,N_36384);
nand U41599 (N_41599,N_38755,N_37688);
and U41600 (N_41600,N_38842,N_36004);
xor U41601 (N_41601,N_38162,N_36374);
xor U41602 (N_41602,N_36280,N_39828);
or U41603 (N_41603,N_37957,N_39824);
nand U41604 (N_41604,N_37021,N_39212);
nor U41605 (N_41605,N_38277,N_39973);
and U41606 (N_41606,N_39313,N_36200);
xnor U41607 (N_41607,N_35429,N_37047);
and U41608 (N_41608,N_35234,N_37266);
nor U41609 (N_41609,N_35334,N_39003);
or U41610 (N_41610,N_37110,N_39008);
xnor U41611 (N_41611,N_37555,N_35692);
nand U41612 (N_41612,N_38016,N_35515);
nor U41613 (N_41613,N_36422,N_39937);
nor U41614 (N_41614,N_37927,N_35050);
nand U41615 (N_41615,N_35647,N_35968);
or U41616 (N_41616,N_39857,N_39270);
and U41617 (N_41617,N_37147,N_35448);
xor U41618 (N_41618,N_36884,N_38974);
or U41619 (N_41619,N_37560,N_39068);
nor U41620 (N_41620,N_38341,N_39494);
or U41621 (N_41621,N_38836,N_39307);
and U41622 (N_41622,N_36863,N_38051);
nor U41623 (N_41623,N_38126,N_36787);
xor U41624 (N_41624,N_36086,N_36373);
nand U41625 (N_41625,N_36006,N_37074);
nand U41626 (N_41626,N_39510,N_38604);
xor U41627 (N_41627,N_37168,N_37489);
nand U41628 (N_41628,N_37535,N_36887);
or U41629 (N_41629,N_35264,N_39109);
or U41630 (N_41630,N_36481,N_36767);
nand U41631 (N_41631,N_36262,N_37616);
nand U41632 (N_41632,N_37911,N_37225);
nor U41633 (N_41633,N_35274,N_38586);
xnor U41634 (N_41634,N_37953,N_35582);
or U41635 (N_41635,N_38320,N_36842);
nand U41636 (N_41636,N_37622,N_36503);
xnor U41637 (N_41637,N_39060,N_39484);
xor U41638 (N_41638,N_35498,N_37215);
nor U41639 (N_41639,N_35717,N_37527);
or U41640 (N_41640,N_35906,N_38688);
and U41641 (N_41641,N_38996,N_36027);
and U41642 (N_41642,N_36658,N_36984);
and U41643 (N_41643,N_39553,N_36537);
and U41644 (N_41644,N_35704,N_38602);
and U41645 (N_41645,N_38868,N_38608);
nor U41646 (N_41646,N_36853,N_39213);
nor U41647 (N_41647,N_36203,N_37306);
nand U41648 (N_41648,N_38121,N_37080);
and U41649 (N_41649,N_36746,N_38583);
nand U41650 (N_41650,N_39155,N_39188);
nand U41651 (N_41651,N_37508,N_37674);
nand U41652 (N_41652,N_37728,N_35239);
nand U41653 (N_41653,N_35252,N_39868);
xnor U41654 (N_41654,N_35034,N_37726);
and U41655 (N_41655,N_39121,N_36499);
and U41656 (N_41656,N_36401,N_39062);
nor U41657 (N_41657,N_36159,N_35203);
or U41658 (N_41658,N_39964,N_38119);
xnor U41659 (N_41659,N_37142,N_35544);
nand U41660 (N_41660,N_37423,N_36778);
xor U41661 (N_41661,N_39995,N_38405);
xnor U41662 (N_41662,N_39221,N_37960);
xor U41663 (N_41663,N_35739,N_37304);
or U41664 (N_41664,N_38085,N_38717);
or U41665 (N_41665,N_35258,N_37746);
xor U41666 (N_41666,N_39202,N_35614);
or U41667 (N_41667,N_35951,N_36326);
or U41668 (N_41668,N_35661,N_36459);
xnor U41669 (N_41669,N_39141,N_39322);
nand U41670 (N_41670,N_37989,N_38630);
xor U41671 (N_41671,N_38732,N_35372);
or U41672 (N_41672,N_39853,N_37072);
or U41673 (N_41673,N_39224,N_39363);
and U41674 (N_41674,N_39303,N_37528);
or U41675 (N_41675,N_37487,N_38545);
nand U41676 (N_41676,N_38120,N_36519);
and U41677 (N_41677,N_36169,N_35464);
and U41678 (N_41678,N_38782,N_37160);
nand U41679 (N_41679,N_37107,N_38683);
and U41680 (N_41680,N_36443,N_36965);
and U41681 (N_41681,N_36723,N_36183);
nor U41682 (N_41682,N_36872,N_36410);
and U41683 (N_41683,N_38374,N_35567);
xor U41684 (N_41684,N_39336,N_37778);
and U41685 (N_41685,N_35907,N_38264);
nor U41686 (N_41686,N_35924,N_38322);
or U41687 (N_41687,N_38496,N_37008);
nand U41688 (N_41688,N_39850,N_39386);
or U41689 (N_41689,N_36801,N_35023);
nor U41690 (N_41690,N_39704,N_39817);
or U41691 (N_41691,N_39617,N_36009);
or U41692 (N_41692,N_39534,N_37408);
nand U41693 (N_41693,N_39664,N_37731);
xnor U41694 (N_41694,N_35996,N_38337);
xnor U41695 (N_41695,N_39979,N_36494);
and U41696 (N_41696,N_35843,N_37364);
and U41697 (N_41697,N_38011,N_36831);
nor U41698 (N_41698,N_38129,N_37360);
nor U41699 (N_41699,N_35633,N_39986);
xnor U41700 (N_41700,N_38365,N_37061);
or U41701 (N_41701,N_36807,N_39750);
nor U41702 (N_41702,N_36971,N_39461);
nor U41703 (N_41703,N_39357,N_39547);
nor U41704 (N_41704,N_38727,N_36621);
nand U41705 (N_41705,N_35360,N_37906);
or U41706 (N_41706,N_38958,N_37981);
nor U41707 (N_41707,N_39066,N_38256);
nand U41708 (N_41708,N_39294,N_36651);
or U41709 (N_41709,N_35541,N_36099);
nand U41710 (N_41710,N_38257,N_38675);
nor U41711 (N_41711,N_36478,N_39540);
nor U41712 (N_41712,N_37595,N_35428);
xor U41713 (N_41713,N_39879,N_37755);
nor U41714 (N_41714,N_39526,N_36480);
or U41715 (N_41715,N_36954,N_37654);
xor U41716 (N_41716,N_39869,N_36826);
nor U41717 (N_41717,N_36631,N_36720);
or U41718 (N_41718,N_35029,N_35175);
xnor U41719 (N_41719,N_36325,N_37058);
and U41720 (N_41720,N_39289,N_36253);
or U41721 (N_41721,N_38034,N_39555);
nor U41722 (N_41722,N_36150,N_35438);
and U41723 (N_41723,N_35181,N_37937);
and U41724 (N_41724,N_37385,N_38396);
or U41725 (N_41725,N_37733,N_37321);
xnor U41726 (N_41726,N_38263,N_36110);
nand U41727 (N_41727,N_37151,N_38657);
xor U41728 (N_41728,N_37001,N_37611);
and U41729 (N_41729,N_38763,N_36047);
xor U41730 (N_41730,N_36852,N_36644);
nor U41731 (N_41731,N_37668,N_35082);
nor U41732 (N_41732,N_35650,N_36591);
and U41733 (N_41733,N_39120,N_37191);
and U41734 (N_41734,N_39203,N_35137);
and U41735 (N_41735,N_36378,N_39366);
or U41736 (N_41736,N_39566,N_35518);
or U41737 (N_41737,N_35033,N_39150);
and U41738 (N_41738,N_38832,N_36243);
and U41739 (N_41739,N_36366,N_38321);
and U41740 (N_41740,N_35882,N_37676);
nand U41741 (N_41741,N_37100,N_39723);
xor U41742 (N_41742,N_39926,N_37735);
xor U41743 (N_41743,N_37835,N_38477);
or U41744 (N_41744,N_36817,N_39057);
xnor U41745 (N_41745,N_38819,N_38626);
and U41746 (N_41746,N_37865,N_39196);
or U41747 (N_41747,N_37758,N_37828);
xnor U41748 (N_41748,N_38781,N_36135);
and U41749 (N_41749,N_36060,N_37763);
xnor U41750 (N_41750,N_38458,N_39805);
nor U41751 (N_41751,N_35128,N_37794);
xor U41752 (N_41752,N_38628,N_36174);
or U41753 (N_41753,N_39371,N_36915);
nor U41754 (N_41754,N_38753,N_37916);
or U41755 (N_41755,N_35347,N_36648);
and U41756 (N_41756,N_35915,N_39887);
or U41757 (N_41757,N_38582,N_37432);
xnor U41758 (N_41758,N_39880,N_39881);
nor U41759 (N_41759,N_35659,N_36751);
xnor U41760 (N_41760,N_36643,N_39106);
nor U41761 (N_41761,N_37823,N_36209);
nor U41762 (N_41762,N_35516,N_38230);
and U41763 (N_41763,N_35505,N_37104);
and U41764 (N_41764,N_39326,N_39426);
nand U41765 (N_41765,N_37382,N_35210);
xor U41766 (N_41766,N_38760,N_37228);
or U41767 (N_41767,N_36973,N_38519);
and U41768 (N_41768,N_39596,N_38690);
xnor U41769 (N_41769,N_36432,N_39765);
nand U41770 (N_41770,N_39394,N_38652);
nand U41771 (N_41771,N_38025,N_36064);
xor U41772 (N_41772,N_37462,N_36206);
nand U41773 (N_41773,N_35981,N_36368);
xor U41774 (N_41774,N_39777,N_37703);
nor U41775 (N_41775,N_37971,N_37651);
nand U41776 (N_41776,N_39135,N_39229);
nor U41777 (N_41777,N_35902,N_35514);
or U41778 (N_41778,N_36719,N_37414);
nand U41779 (N_41779,N_35180,N_39415);
or U41780 (N_41780,N_39660,N_38770);
nor U41781 (N_41781,N_39044,N_38479);
or U41782 (N_41782,N_36346,N_36772);
xnor U41783 (N_41783,N_37299,N_39418);
xnor U41784 (N_41784,N_39460,N_36387);
nor U41785 (N_41785,N_37197,N_37655);
nand U41786 (N_41786,N_37563,N_35634);
nor U41787 (N_41787,N_38144,N_38053);
and U41788 (N_41788,N_35060,N_35693);
or U41789 (N_41789,N_38414,N_36978);
nor U41790 (N_41790,N_39105,N_39261);
nand U41791 (N_41791,N_35100,N_38680);
xor U41792 (N_41792,N_38233,N_35621);
and U41793 (N_41793,N_38422,N_38097);
or U41794 (N_41794,N_39269,N_39531);
nor U41795 (N_41795,N_37540,N_35691);
and U41796 (N_41796,N_35436,N_37578);
and U41797 (N_41797,N_39517,N_38981);
and U41798 (N_41798,N_39409,N_35532);
xnor U41799 (N_41799,N_36606,N_36121);
and U41800 (N_41800,N_37702,N_36516);
or U41801 (N_41801,N_37510,N_39793);
nand U41802 (N_41802,N_35896,N_37196);
nor U41803 (N_41803,N_35011,N_36661);
xor U41804 (N_41804,N_37834,N_38785);
nor U41805 (N_41805,N_36309,N_38400);
xnor U41806 (N_41806,N_36686,N_37420);
nor U41807 (N_41807,N_38471,N_37183);
nor U41808 (N_41808,N_39692,N_39065);
or U41809 (N_41809,N_39916,N_38922);
or U41810 (N_41810,N_37738,N_36178);
xnor U41811 (N_41811,N_37136,N_35075);
nor U41812 (N_41812,N_36340,N_37199);
xnor U41813 (N_41813,N_38854,N_35094);
or U41814 (N_41814,N_36361,N_35444);
or U41815 (N_41815,N_35453,N_35726);
or U41816 (N_41816,N_37339,N_39967);
nand U41817 (N_41817,N_35136,N_39411);
xnor U41818 (N_41818,N_36356,N_39015);
nand U41819 (N_41819,N_39063,N_39255);
nand U41820 (N_41820,N_39898,N_39845);
xor U41821 (N_41821,N_35718,N_37983);
xor U41822 (N_41822,N_35117,N_37185);
nand U41823 (N_41823,N_38543,N_38712);
nand U41824 (N_41824,N_37433,N_36956);
nand U41825 (N_41825,N_39975,N_39734);
nand U41826 (N_41826,N_39968,N_37126);
xnor U41827 (N_41827,N_37522,N_39282);
and U41828 (N_41828,N_37820,N_35828);
or U41829 (N_41829,N_39417,N_38137);
or U41830 (N_41830,N_35664,N_35160);
and U41831 (N_41831,N_38824,N_39279);
nand U41832 (N_41832,N_39478,N_35189);
and U41833 (N_41833,N_36151,N_35590);
and U41834 (N_41834,N_38601,N_39048);
xnor U41835 (N_41835,N_39591,N_36623);
and U41836 (N_41836,N_38739,N_38968);
or U41837 (N_41837,N_38865,N_35510);
and U41838 (N_41838,N_37934,N_39025);
or U41839 (N_41839,N_39131,N_38340);
and U41840 (N_41840,N_35879,N_39032);
nand U41841 (N_41841,N_37551,N_36747);
and U41842 (N_41842,N_37252,N_39521);
xnor U41843 (N_41843,N_38398,N_39387);
or U41844 (N_41844,N_37015,N_36639);
nor U41845 (N_41845,N_39764,N_39209);
nand U41846 (N_41846,N_39445,N_36830);
nand U41847 (N_41847,N_39766,N_38851);
or U41848 (N_41848,N_35987,N_39160);
or U41849 (N_41849,N_39751,N_37881);
nor U41850 (N_41850,N_39205,N_39180);
and U41851 (N_41851,N_36274,N_39818);
nor U41852 (N_41852,N_35324,N_37948);
or U41853 (N_41853,N_36827,N_35300);
or U41854 (N_41854,N_38353,N_38673);
nand U41855 (N_41855,N_37354,N_35416);
and U41856 (N_41856,N_36548,N_37666);
nor U41857 (N_41857,N_36339,N_35374);
xnor U41858 (N_41858,N_36732,N_35322);
or U41859 (N_41859,N_35577,N_35365);
and U41860 (N_41860,N_35489,N_38452);
and U41861 (N_41861,N_36452,N_37332);
or U41862 (N_41862,N_39684,N_38344);
or U41863 (N_41863,N_39806,N_35465);
or U41864 (N_41864,N_37753,N_38249);
or U41865 (N_41865,N_36341,N_35563);
and U41866 (N_41866,N_37672,N_38364);
xor U41867 (N_41867,N_38232,N_39168);
xor U41868 (N_41868,N_35675,N_39042);
or U41869 (N_41869,N_35143,N_35963);
nor U41870 (N_41870,N_38251,N_39091);
xnor U41871 (N_41871,N_35331,N_39656);
nand U41872 (N_41872,N_38101,N_38703);
nor U41873 (N_41873,N_39331,N_38460);
and U41874 (N_41874,N_35237,N_39884);
nor U41875 (N_41875,N_39390,N_37793);
or U41876 (N_41876,N_35426,N_35395);
nand U41877 (N_41877,N_39420,N_39028);
and U41878 (N_41878,N_39502,N_35803);
xnor U41879 (N_41879,N_36216,N_39866);
nor U41880 (N_41880,N_39334,N_35164);
nor U41881 (N_41881,N_39904,N_36160);
xnor U41882 (N_41882,N_36270,N_35873);
nand U41883 (N_41883,N_37812,N_36111);
nand U41884 (N_41884,N_38986,N_39724);
and U41885 (N_41885,N_38771,N_37943);
nor U41886 (N_41886,N_38942,N_39208);
nor U41887 (N_41887,N_36158,N_37068);
nor U41888 (N_41888,N_37490,N_39352);
or U41889 (N_41889,N_38857,N_37029);
and U41890 (N_41890,N_35628,N_39005);
and U41891 (N_41891,N_38729,N_38798);
nor U41892 (N_41892,N_39369,N_36895);
xnor U41893 (N_41893,N_38939,N_37556);
nand U41894 (N_41894,N_36062,N_38961);
xnor U41895 (N_41895,N_36279,N_39970);
and U41896 (N_41896,N_38888,N_39054);
or U41897 (N_41897,N_37589,N_36229);
nor U41898 (N_41898,N_37681,N_35391);
nor U41899 (N_41899,N_39700,N_35207);
nand U41900 (N_41900,N_35653,N_39886);
nand U41901 (N_41901,N_35946,N_36918);
and U41902 (N_41902,N_38997,N_35195);
and U41903 (N_41903,N_36267,N_37732);
xor U41904 (N_41904,N_35367,N_38951);
and U41905 (N_41905,N_35959,N_39049);
nor U41906 (N_41906,N_39007,N_39283);
xor U41907 (N_41907,N_36349,N_39587);
nor U41908 (N_41908,N_35932,N_36069);
nor U41909 (N_41909,N_36850,N_36505);
xnor U41910 (N_41910,N_38038,N_38907);
nand U41911 (N_41911,N_39441,N_36100);
nand U41912 (N_41912,N_37289,N_39422);
and U41913 (N_41913,N_39099,N_38300);
and U41914 (N_41914,N_38118,N_35500);
xor U41915 (N_41915,N_36484,N_37163);
nand U41916 (N_41916,N_38883,N_37518);
xor U41917 (N_41917,N_39513,N_37501);
xnor U41918 (N_41918,N_39773,N_35689);
and U41919 (N_41919,N_37675,N_37039);
xnor U41920 (N_41920,N_37740,N_37682);
or U41921 (N_41921,N_35506,N_37165);
nor U41922 (N_41922,N_38470,N_38540);
nand U41923 (N_41923,N_37895,N_39523);
and U41924 (N_41924,N_38198,N_38395);
nand U41925 (N_41925,N_35905,N_38155);
and U41926 (N_41926,N_37179,N_36580);
xnor U41927 (N_41927,N_38161,N_39429);
nand U41928 (N_41928,N_35384,N_35147);
nand U41929 (N_41929,N_37488,N_39310);
xnor U41930 (N_41930,N_35652,N_35151);
xnor U41931 (N_41931,N_36743,N_39271);
nor U41932 (N_41932,N_37899,N_35881);
nor U41933 (N_41933,N_39780,N_39543);
nor U41934 (N_41934,N_37307,N_36425);
nand U41935 (N_41935,N_37002,N_37434);
and U41936 (N_41936,N_36077,N_39370);
and U41937 (N_41937,N_35798,N_37272);
nor U41938 (N_41938,N_37951,N_37604);
xor U41939 (N_41939,N_37257,N_38580);
or U41940 (N_41940,N_38266,N_39240);
xnor U41941 (N_41941,N_37857,N_36038);
or U41942 (N_41942,N_36724,N_39859);
or U41943 (N_41943,N_37708,N_36741);
or U41944 (N_41944,N_37166,N_39384);
xnor U41945 (N_41945,N_35668,N_39302);
xor U41946 (N_41946,N_38131,N_38524);
or U41947 (N_41947,N_39416,N_39491);
nand U41948 (N_41948,N_38462,N_37780);
nand U41949 (N_41949,N_39183,N_37255);
and U41950 (N_41950,N_39376,N_37016);
or U41951 (N_41951,N_35710,N_37955);
nand U41952 (N_41952,N_39525,N_39579);
or U41953 (N_41953,N_37397,N_36541);
nor U41954 (N_41954,N_39910,N_39026);
nor U41955 (N_41955,N_36305,N_35459);
nor U41956 (N_41956,N_39300,N_36582);
and U41957 (N_41957,N_39317,N_35031);
nor U41958 (N_41958,N_35466,N_38568);
or U41959 (N_41959,N_38338,N_36763);
and U41960 (N_41960,N_39361,N_38279);
nand U41961 (N_41961,N_38087,N_39251);
xor U41962 (N_41962,N_37743,N_38170);
nand U41963 (N_41963,N_39433,N_39762);
nor U41964 (N_41964,N_36175,N_36610);
xnor U41965 (N_41965,N_36294,N_38773);
nor U41966 (N_41966,N_35630,N_38243);
nor U41967 (N_41967,N_37395,N_39852);
nor U41968 (N_41968,N_36217,N_37617);
xor U41969 (N_41969,N_37216,N_38569);
or U41970 (N_41970,N_38467,N_35349);
xor U41971 (N_41971,N_35657,N_36122);
xnor U41972 (N_41972,N_39578,N_38810);
nor U41973 (N_41973,N_36914,N_36730);
nor U41974 (N_41974,N_35216,N_39157);
or U41975 (N_41975,N_38984,N_39784);
or U41976 (N_41976,N_39485,N_39092);
nand U41977 (N_41977,N_36320,N_35119);
nand U41978 (N_41978,N_39662,N_37714);
and U41979 (N_41979,N_39396,N_39227);
nand U41980 (N_41980,N_35312,N_35826);
nand U41981 (N_41981,N_37773,N_36115);
nand U41982 (N_41982,N_35185,N_38980);
xor U41983 (N_41983,N_37470,N_35848);
nand U41984 (N_41984,N_37237,N_35191);
and U41985 (N_41985,N_36874,N_35580);
xnor U41986 (N_41986,N_38286,N_36265);
nor U41987 (N_41987,N_35018,N_39186);
or U41988 (N_41988,N_39781,N_39009);
nor U41989 (N_41989,N_35247,N_35800);
and U41990 (N_41990,N_39634,N_35799);
nand U41991 (N_41991,N_38649,N_39715);
nor U41992 (N_41992,N_39223,N_38403);
and U41993 (N_41993,N_37092,N_35703);
nor U41994 (N_41994,N_35345,N_36983);
nand U41995 (N_41995,N_36447,N_37318);
and U41996 (N_41996,N_38994,N_35310);
or U41997 (N_41997,N_37050,N_38606);
nor U41998 (N_41998,N_35088,N_35096);
or U41999 (N_41999,N_39548,N_37719);
nand U42000 (N_42000,N_37442,N_37692);
nand U42001 (N_42001,N_38936,N_38709);
xor U42002 (N_42002,N_37190,N_38122);
xor U42003 (N_42003,N_37249,N_39902);
nor U42004 (N_42004,N_38275,N_37352);
nor U42005 (N_42005,N_37189,N_36705);
and U42006 (N_42006,N_35233,N_35539);
nand U42007 (N_42007,N_37650,N_39949);
nor U42008 (N_42008,N_36477,N_39772);
nand U42009 (N_42009,N_35104,N_38206);
or U42010 (N_42010,N_35903,N_39738);
nand U42011 (N_42011,N_35441,N_39978);
nand U42012 (N_42012,N_36994,N_39999);
nand U42013 (N_42013,N_36949,N_36290);
nand U42014 (N_42014,N_35474,N_38702);
and U42015 (N_42015,N_37020,N_39175);
xor U42016 (N_42016,N_35229,N_35282);
nor U42017 (N_42017,N_38791,N_36646);
or U42018 (N_42018,N_38553,N_38267);
nand U42019 (N_42019,N_38455,N_35899);
and U42020 (N_42020,N_39506,N_37223);
nand U42021 (N_42021,N_35588,N_39863);
nand U42022 (N_42022,N_37618,N_36389);
xor U42023 (N_42023,N_38294,N_36642);
nand U42024 (N_42024,N_39677,N_35866);
nor U42025 (N_42025,N_35020,N_36795);
nor U42026 (N_42026,N_37888,N_37349);
nand U42027 (N_42027,N_38662,N_39379);
xnor U42028 (N_42028,N_36225,N_39648);
nor U42029 (N_42029,N_35790,N_38957);
and U42030 (N_42030,N_39924,N_35225);
nor U42031 (N_42031,N_35681,N_37106);
and U42032 (N_42032,N_37844,N_36940);
and U42033 (N_42033,N_36470,N_38645);
and U42034 (N_42034,N_38845,N_35206);
xor U42035 (N_42035,N_38672,N_39665);
nand U42036 (N_42036,N_35176,N_39960);
and U42037 (N_42037,N_38502,N_38697);
or U42038 (N_42038,N_35272,N_35945);
or U42039 (N_42039,N_38678,N_37547);
xor U42040 (N_42040,N_38193,N_39236);
or U42041 (N_42041,N_38598,N_35853);
and U42042 (N_42042,N_39994,N_37569);
nand U42043 (N_42043,N_35423,N_36882);
or U42044 (N_42044,N_35937,N_35301);
nand U42045 (N_42045,N_37494,N_35017);
xor U42046 (N_42046,N_38278,N_38710);
xor U42047 (N_42047,N_36360,N_35163);
xor U42048 (N_42048,N_35635,N_37102);
xnor U42049 (N_42049,N_39265,N_38776);
or U42050 (N_42050,N_37120,N_38563);
nor U42051 (N_42051,N_36383,N_38106);
or U42052 (N_42052,N_36855,N_35157);
nand U42053 (N_42053,N_39050,N_35291);
and U42054 (N_42054,N_35168,N_38439);
or U42055 (N_42055,N_39905,N_35458);
and U42056 (N_42056,N_39550,N_39716);
nor U42057 (N_42057,N_38302,N_39495);
xnor U42058 (N_42058,N_35923,N_39509);
and U42059 (N_42059,N_35292,N_35432);
xnor U42060 (N_42060,N_35358,N_36078);
nand U42061 (N_42061,N_37175,N_36157);
and U42062 (N_42062,N_38288,N_36844);
xor U42063 (N_42063,N_39782,N_37327);
and U42064 (N_42064,N_39711,N_39132);
nor U42065 (N_42065,N_38372,N_36753);
xnor U42066 (N_42066,N_36975,N_36600);
nor U42067 (N_42067,N_38281,N_35624);
or U42068 (N_42068,N_39278,N_38546);
xnor U42069 (N_42069,N_36318,N_37341);
nor U42070 (N_42070,N_39774,N_37914);
or U42071 (N_42071,N_39452,N_35989);
nand U42072 (N_42072,N_35605,N_35418);
nor U42073 (N_42073,N_37174,N_38880);
xor U42074 (N_42074,N_38663,N_35424);
nand U42075 (N_42075,N_38624,N_39725);
xnor U42076 (N_42076,N_37138,N_37076);
and U42077 (N_42077,N_38381,N_35063);
or U42078 (N_42078,N_36930,N_37054);
nor U42079 (N_42079,N_38303,N_39661);
and U42080 (N_42080,N_35212,N_39616);
nand U42081 (N_42081,N_35036,N_35586);
nand U42082 (N_42082,N_35417,N_39257);
and U42083 (N_42083,N_36190,N_38906);
xnor U42084 (N_42084,N_37026,N_35935);
xor U42085 (N_42085,N_35850,N_36936);
and U42086 (N_42086,N_37343,N_37446);
nand U42087 (N_42087,N_35727,N_36913);
nand U42088 (N_42088,N_39398,N_35120);
and U42089 (N_42089,N_38335,N_39944);
nor U42090 (N_42090,N_37543,N_36029);
nor U42091 (N_42091,N_37209,N_35045);
or U42092 (N_42092,N_36011,N_36313);
or U42093 (N_42093,N_37519,N_36802);
or U42094 (N_42094,N_38377,N_36080);
and U42095 (N_42095,N_37804,N_38596);
xor U42096 (N_42096,N_36295,N_38915);
or U42097 (N_42097,N_37969,N_35942);
and U42098 (N_42098,N_38670,N_35114);
nand U42099 (N_42099,N_37849,N_36532);
xor U42100 (N_42100,N_39024,N_36609);
and U42101 (N_42101,N_35759,N_36540);
xor U42102 (N_42102,N_37594,N_36308);
and U42103 (N_42103,N_36050,N_38231);
or U42104 (N_42104,N_38789,N_35705);
xnor U42105 (N_42105,N_38964,N_36282);
nand U42106 (N_42106,N_37657,N_39064);
nor U42107 (N_42107,N_36005,N_35602);
nor U42108 (N_42108,N_39362,N_35796);
xor U42109 (N_42109,N_38309,N_37010);
nor U42110 (N_42110,N_37567,N_38032);
nor U42111 (N_42111,N_35356,N_38828);
xnor U42112 (N_42112,N_36590,N_39073);
or U42113 (N_42113,N_36214,N_36780);
nand U42114 (N_42114,N_35753,N_38956);
and U42115 (N_42115,N_38176,N_36810);
nand U42116 (N_42116,N_38298,N_35473);
nor U42117 (N_42117,N_37581,N_36758);
or U42118 (N_42118,N_35346,N_39539);
nand U42119 (N_42119,N_36924,N_37181);
or U42120 (N_42120,N_37576,N_38042);
nand U42121 (N_42121,N_35369,N_38872);
xor U42122 (N_42122,N_35827,N_39790);
nand U42123 (N_42123,N_35179,N_38024);
nand U42124 (N_42124,N_39088,N_39867);
nand U42125 (N_42125,N_35173,N_35008);
or U42126 (N_42126,N_35231,N_39292);
or U42127 (N_42127,N_37557,N_36354);
nor U42128 (N_42128,N_38431,N_35852);
nor U42129 (N_42129,N_37313,N_37066);
xor U42130 (N_42130,N_38191,N_35107);
nand U42131 (N_42131,N_35217,N_39170);
xnor U42132 (N_42132,N_36900,N_36929);
nand U42133 (N_42133,N_39532,N_38642);
or U42134 (N_42134,N_39430,N_37944);
and U42135 (N_42135,N_37606,N_37135);
or U42136 (N_42136,N_35078,N_38718);
or U42137 (N_42137,N_35460,N_36601);
nand U42138 (N_42138,N_36656,N_36518);
or U42139 (N_42139,N_36315,N_35141);
nor U42140 (N_42140,N_35585,N_39838);
and U42141 (N_42141,N_38498,N_37548);
or U42142 (N_42142,N_39199,N_38534);
xor U42143 (N_42143,N_38240,N_37539);
nand U42144 (N_42144,N_39956,N_35079);
nor U42145 (N_42145,N_38031,N_38009);
or U42146 (N_42146,N_38253,N_35118);
nand U42147 (N_42147,N_38966,N_38734);
and U42148 (N_42148,N_38914,N_39299);
xor U42149 (N_42149,N_37363,N_39431);
nand U42150 (N_42150,N_37789,N_37280);
nor U42151 (N_42151,N_39454,N_38801);
or U42152 (N_42152,N_38741,N_39058);
nand U42153 (N_42153,N_37480,N_37370);
and U42154 (N_42154,N_37570,N_36502);
nand U42155 (N_42155,N_37145,N_37314);
nand U42156 (N_42156,N_36804,N_39988);
xor U42157 (N_42157,N_36800,N_38805);
or U42158 (N_42158,N_39512,N_39801);
nand U42159 (N_42159,N_35370,N_39329);
xnor U42160 (N_42160,N_39563,N_36985);
nor U42161 (N_42161,N_35266,N_37348);
nor U42162 (N_42162,N_37945,N_36176);
xnor U42163 (N_42163,N_36599,N_36363);
nand U42164 (N_42164,N_35269,N_37935);
and U42165 (N_42165,N_38019,N_36254);
nor U42166 (N_42166,N_39288,N_36146);
nand U42167 (N_42167,N_39740,N_36546);
nand U42168 (N_42168,N_39666,N_37417);
nor U42169 (N_42169,N_35373,N_38216);
nand U42170 (N_42170,N_36677,N_38136);
and U42171 (N_42171,N_35227,N_36993);
nand U42172 (N_42172,N_36352,N_36749);
xnor U42173 (N_42173,N_38145,N_35965);
xor U42174 (N_42174,N_39043,N_39888);
nand U42175 (N_42175,N_39963,N_39873);
xor U42176 (N_42176,N_36822,N_37022);
and U42177 (N_42177,N_39847,N_39712);
nor U42178 (N_42178,N_38701,N_35348);
and U42179 (N_42179,N_37852,N_38695);
and U42180 (N_42180,N_36506,N_39197);
and U42181 (N_42181,N_38376,N_35551);
and U42182 (N_42182,N_36514,N_36434);
xor U42183 (N_42183,N_35178,N_39072);
or U42184 (N_42184,N_37208,N_38282);
or U42185 (N_42185,N_37372,N_36905);
or U42186 (N_42186,N_38094,N_38211);
and U42187 (N_42187,N_36534,N_39286);
xor U42188 (N_42188,N_35224,N_35172);
xor U42189 (N_42189,N_38108,N_35880);
xor U42190 (N_42190,N_38081,N_39480);
and U42191 (N_42191,N_39036,N_36034);
nand U42192 (N_42192,N_36344,N_38693);
or U42193 (N_42193,N_39123,N_35957);
nand U42194 (N_42194,N_38714,N_38731);
and U42195 (N_42195,N_36284,N_36809);
nor U42196 (N_42196,N_38482,N_39397);
nor U42197 (N_42197,N_35837,N_36722);
nand U42198 (N_42198,N_36988,N_37162);
nand U42199 (N_42199,N_38621,N_38401);
nand U42200 (N_42200,N_38588,N_39618);
nor U42201 (N_42201,N_36760,N_35523);
nand U42202 (N_42202,N_38397,N_38775);
nand U42203 (N_42203,N_37281,N_36124);
and U42204 (N_42204,N_37689,N_36762);
or U42205 (N_42205,N_36715,N_36969);
nand U42206 (N_42206,N_35792,N_39327);
nor U42207 (N_42207,N_36139,N_39541);
or U42208 (N_42208,N_39991,N_36779);
nor U42209 (N_42209,N_39769,N_39570);
or U42210 (N_42210,N_35519,N_36451);
or U42211 (N_42211,N_35260,N_36208);
nor U42212 (N_42212,N_39518,N_39800);
nand U42213 (N_42213,N_37748,N_39871);
nor U42214 (N_42214,N_35288,N_38882);
and U42215 (N_42215,N_35150,N_36654);
nor U42216 (N_42216,N_35052,N_35530);
nor U42217 (N_42217,N_35715,N_39242);
and U42218 (N_42218,N_35449,N_35406);
or U42219 (N_42219,N_39194,N_39694);
nor U42220 (N_42220,N_39206,N_36232);
nor U42221 (N_42221,N_36854,N_38667);
nor U42222 (N_42222,N_37985,N_35637);
nor U42223 (N_42223,N_35636,N_37231);
nand U42224 (N_42224,N_37727,N_39941);
xnor U42225 (N_42225,N_35513,N_36036);
or U42226 (N_42226,N_38593,N_35608);
nor U42227 (N_42227,N_39272,N_39794);
xnor U42228 (N_42228,N_37894,N_39954);
xor U42229 (N_42229,N_39284,N_37325);
or U42230 (N_42230,N_39019,N_37137);
nand U42231 (N_42231,N_37963,N_36177);
xnor U42232 (N_42232,N_38213,N_37133);
and U42233 (N_42233,N_39719,N_39195);
xor U42234 (N_42234,N_36227,N_35158);
nor U42235 (N_42235,N_37856,N_35615);
xor U42236 (N_42236,N_37101,N_38351);
and U42237 (N_42237,N_35186,N_37621);
and U42238 (N_42238,N_38689,N_36647);
xnor U42239 (N_42239,N_36553,N_39825);
or U42240 (N_42240,N_37475,N_36023);
nand U42241 (N_42241,N_39807,N_39584);
nor U42242 (N_42242,N_35988,N_36761);
and U42243 (N_42243,N_37273,N_35315);
nor U42244 (N_42244,N_36886,N_37025);
nand U42245 (N_42245,N_35041,N_39343);
xor U42246 (N_42246,N_36093,N_37723);
xor U42247 (N_42247,N_38784,N_37687);
xnor U42248 (N_42248,N_39301,N_38086);
and U42249 (N_42249,N_39833,N_37041);
or U42250 (N_42250,N_36542,N_35263);
nor U42251 (N_42251,N_38627,N_39826);
nand U42252 (N_42252,N_35886,N_37818);
nand U42253 (N_42253,N_36167,N_35952);
nand U42254 (N_42254,N_36462,N_39984);
or U42255 (N_42255,N_38982,N_35728);
xor U42256 (N_42256,N_38812,N_38218);
xor U42257 (N_42257,N_36324,N_39290);
nor U42258 (N_42258,N_37288,N_36620);
xnor U42259 (N_42259,N_35961,N_35249);
xnor U42260 (N_42260,N_35889,N_37496);
and U42261 (N_42261,N_35912,N_38346);
nor U42262 (N_42262,N_36145,N_35482);
and U42263 (N_42263,N_36581,N_39529);
or U42264 (N_42264,N_39497,N_38312);
xor U42265 (N_42265,N_35649,N_37973);
or U42266 (N_42266,N_36199,N_39211);
or U42267 (N_42267,N_36653,N_35256);
nand U42268 (N_42268,N_37964,N_38499);
and U42269 (N_42269,N_37453,N_39103);
or U42270 (N_42270,N_37757,N_38841);
or U42271 (N_42271,N_35462,N_39551);
and U42272 (N_42272,N_39342,N_39001);
xor U42273 (N_42273,N_38985,N_36584);
nor U42274 (N_42274,N_38644,N_38747);
and U42275 (N_42275,N_38255,N_35977);
xnor U42276 (N_42276,N_35836,N_39222);
and U42277 (N_42277,N_36075,N_36968);
nor U42278 (N_42278,N_36092,N_37565);
and U42279 (N_42279,N_37326,N_35170);
xnor U42280 (N_42280,N_35019,N_35543);
and U42281 (N_42281,N_38811,N_38474);
and U42282 (N_42282,N_38505,N_37296);
nand U42283 (N_42283,N_36032,N_37730);
and U42284 (N_42284,N_35419,N_39804);
and U42285 (N_42285,N_37182,N_38862);
nor U42286 (N_42286,N_35062,N_37526);
and U42287 (N_42287,N_36256,N_35922);
or U42288 (N_42288,N_35477,N_36353);
xnor U42289 (N_42289,N_38299,N_38536);
or U42290 (N_42290,N_38478,N_35433);
xnor U42291 (N_42291,N_35377,N_36742);
or U42292 (N_42292,N_38838,N_38622);
xnor U42293 (N_42293,N_38853,N_35095);
xor U42294 (N_42294,N_38139,N_36951);
or U42295 (N_42295,N_36748,N_38146);
and U42296 (N_42296,N_36512,N_35842);
nand U42297 (N_42297,N_39996,N_39084);
and U42298 (N_42298,N_36013,N_36067);
and U42299 (N_42299,N_39071,N_38045);
and U42300 (N_42300,N_36835,N_36509);
nor U42301 (N_42301,N_36215,N_36641);
nor U42302 (N_42302,N_37148,N_35991);
nand U42303 (N_42303,N_38248,N_38128);
or U42304 (N_42304,N_35488,N_37552);
nand U42305 (N_42305,N_37875,N_36419);
or U42306 (N_42306,N_35435,N_37802);
nor U42307 (N_42307,N_39011,N_35351);
or U42308 (N_42308,N_37861,N_36711);
and U42309 (N_42309,N_39349,N_37388);
xnor U42310 (N_42310,N_36071,N_36766);
and U42311 (N_42311,N_35960,N_38941);
nand U42312 (N_42312,N_38549,N_38112);
nand U42313 (N_42313,N_38500,N_37333);
nor U42314 (N_42314,N_37073,N_35265);
nor U42315 (N_42315,N_39561,N_39337);
or U42316 (N_42316,N_36302,N_35919);
and U42317 (N_42317,N_38676,N_36511);
xor U42318 (N_42318,N_37532,N_35251);
nand U42319 (N_42319,N_35016,N_38493);
xnor U42320 (N_42320,N_37503,N_38196);
or U42321 (N_42321,N_38610,N_38069);
or U42322 (N_42322,N_36283,N_35571);
nand U42323 (N_42323,N_39588,N_35716);
nand U42324 (N_42324,N_37438,N_36996);
or U42325 (N_42325,N_36495,N_39862);
nor U42326 (N_42326,N_38348,N_37976);
nor U42327 (N_42327,N_37660,N_39276);
xor U42328 (N_42328,N_35824,N_36095);
or U42329 (N_42329,N_39389,N_35131);
xnor U42330 (N_42330,N_39718,N_39107);
or U42331 (N_42331,N_37646,N_37500);
xor U42332 (N_42332,N_35138,N_37816);
xnor U42333 (N_42333,N_39702,N_36269);
xor U42334 (N_42334,N_38778,N_37785);
xnor U42335 (N_42335,N_36117,N_35215);
nand U42336 (N_42336,N_38437,N_39412);
nor U42337 (N_42337,N_35480,N_36479);
xnor U42338 (N_42338,N_37639,N_36188);
or U42339 (N_42339,N_35142,N_35554);
and U42340 (N_42340,N_38245,N_39187);
or U42341 (N_42341,N_35123,N_35574);
xnor U42342 (N_42342,N_39829,N_37447);
and U42343 (N_42343,N_37974,N_37310);
nor U42344 (N_42344,N_39374,N_36788);
and U42345 (N_42345,N_36193,N_36868);
or U42346 (N_42346,N_35394,N_39037);
nand U42347 (N_42347,N_39401,N_36391);
or U42348 (N_42348,N_35955,N_36101);
or U42349 (N_42349,N_37637,N_38575);
or U42350 (N_42350,N_38983,N_35953);
xor U42351 (N_42351,N_38291,N_36048);
nand U42352 (N_42352,N_36147,N_38217);
nand U42353 (N_42353,N_38615,N_36195);
and U42354 (N_42354,N_39558,N_36885);
nor U42355 (N_42355,N_35276,N_36331);
or U42356 (N_42356,N_35825,N_36637);
nor U42357 (N_42357,N_39810,N_35332);
and U42358 (N_42358,N_35760,N_35838);
or U42359 (N_42359,N_36572,N_38578);
nand U42360 (N_42360,N_38817,N_39557);
nor U42361 (N_42361,N_37239,N_39436);
nand U42362 (N_42362,N_36439,N_38487);
nand U42363 (N_42363,N_38677,N_36861);
nand U42364 (N_42364,N_37813,N_37264);
and U42365 (N_42365,N_38399,N_39524);
nand U42366 (N_42366,N_37153,N_37413);
nand U42367 (N_42367,N_35897,N_36127);
nor U42368 (N_42368,N_37467,N_36087);
or U42369 (N_42369,N_35481,N_38979);
nand U42370 (N_42370,N_39695,N_39759);
nand U42371 (N_42371,N_37441,N_36329);
and U42372 (N_42372,N_39323,N_36521);
xnor U42373 (N_42373,N_35569,N_39305);
or U42374 (N_42374,N_39776,N_37419);
or U42375 (N_42375,N_39580,N_39950);
nor U42376 (N_42376,N_38835,N_38004);
and U42377 (N_42377,N_38061,N_39469);
nor U42378 (N_42378,N_37006,N_37553);
and U42379 (N_42379,N_35914,N_35389);
or U42380 (N_42380,N_35913,N_38027);
or U42381 (N_42381,N_36880,N_35470);
or U42382 (N_42382,N_36081,N_36202);
nor U42383 (N_42383,N_37032,N_38459);
or U42384 (N_42384,N_37421,N_36170);
and U42385 (N_42385,N_35005,N_36414);
xnor U42386 (N_42386,N_37524,N_36845);
nor U42387 (N_42387,N_38026,N_35815);
and U42388 (N_42388,N_38373,N_36806);
nand U42389 (N_42389,N_38856,N_36561);
or U42390 (N_42390,N_37436,N_37779);
nor U42391 (N_42391,N_35059,N_36497);
and U42392 (N_42392,N_36608,N_39727);
or U42393 (N_42393,N_35030,N_39139);
or U42394 (N_42394,N_39732,N_38866);
xor U42395 (N_42395,N_36768,N_35483);
nor U42396 (N_42396,N_35964,N_39921);
and U42397 (N_42397,N_37711,N_36911);
nand U42398 (N_42398,N_35625,N_37653);
nor U42399 (N_42399,N_35076,N_39392);
nor U42400 (N_42400,N_37187,N_35246);
or U42401 (N_42401,N_38999,N_37123);
nand U42402 (N_42402,N_38418,N_38017);
nor U42403 (N_42403,N_36508,N_39022);
or U42404 (N_42404,N_35618,N_39116);
xor U42405 (N_42405,N_37810,N_35645);
nor U42406 (N_42406,N_39473,N_35261);
or U42407 (N_42407,N_37115,N_37449);
xnor U42408 (N_42408,N_35420,N_36403);
nor U42409 (N_42409,N_37670,N_38360);
nor U42410 (N_42410,N_39435,N_35908);
and U42411 (N_42411,N_39575,N_37680);
nand U42412 (N_42412,N_38940,N_38352);
or U42413 (N_42413,N_35561,N_35672);
nand U42414 (N_42414,N_39998,N_37301);
nand U42415 (N_42415,N_38350,N_39993);
and U42416 (N_42416,N_37647,N_35162);
xnor U42417 (N_42417,N_37847,N_36944);
or U42418 (N_42418,N_35116,N_35972);
nor U42419 (N_42419,N_36388,N_37858);
or U42420 (N_42420,N_39733,N_35810);
xnor U42421 (N_42421,N_38171,N_36784);
nor U42422 (N_42422,N_39347,N_36665);
and U42423 (N_42423,N_38078,N_36362);
or U42424 (N_42424,N_36426,N_37842);
xor U42425 (N_42425,N_37741,N_39785);
nor U42426 (N_42426,N_38616,N_38150);
xnor U42427 (N_42427,N_36594,N_35947);
nor U42428 (N_42428,N_35006,N_39836);
nand U42429 (N_42429,N_37150,N_38163);
nand U42430 (N_42430,N_35708,N_37335);
and U42431 (N_42431,N_39450,N_37108);
xor U42432 (N_42432,N_35741,N_39081);
nor U42433 (N_42433,N_37128,N_36231);
and U42434 (N_42434,N_38787,N_35706);
and U42435 (N_42435,N_38490,N_37718);
nand U42436 (N_42436,N_35046,N_37970);
and U42437 (N_42437,N_36239,N_36757);
xnor U42438 (N_42438,N_35538,N_35311);
nand U42439 (N_42439,N_35318,N_35735);
nor U42440 (N_42440,N_37465,N_39812);
nor U42441 (N_42441,N_35537,N_36798);
or U42442 (N_42442,N_36923,N_35877);
or U42443 (N_42443,N_37530,N_38665);
xnor U42444 (N_42444,N_37891,N_38720);
xnor U42445 (N_42445,N_39391,N_38393);
or U42446 (N_42446,N_37598,N_37566);
nand U42447 (N_42447,N_36469,N_37853);
and U42448 (N_42448,N_39348,N_35386);
nor U42449 (N_42449,N_38209,N_36754);
xnor U42450 (N_42450,N_37117,N_36025);
nor U42451 (N_42451,N_36014,N_35364);
and U42452 (N_42452,N_36143,N_38896);
and U42453 (N_42453,N_37514,N_38427);
xor U42454 (N_42454,N_36192,N_35549);
and U42455 (N_42455,N_38929,N_35801);
nor U42456 (N_42456,N_37729,N_37226);
or U42457 (N_42457,N_37322,N_35570);
xor U42458 (N_42458,N_37582,N_38891);
or U42459 (N_42459,N_38704,N_38998);
nor U42460 (N_42460,N_38976,N_35308);
and U42461 (N_42461,N_37317,N_36879);
nand U42462 (N_42462,N_37645,N_36444);
nor U42463 (N_42463,N_38721,N_38930);
nand U42464 (N_42464,N_38183,N_36321);
xor U42465 (N_42465,N_39691,N_38440);
nand U42466 (N_42466,N_36105,N_39706);
xnor U42467 (N_42467,N_36314,N_39899);
and U42468 (N_42468,N_39459,N_36251);
and U42469 (N_42469,N_35153,N_38931);
or U42470 (N_42470,N_37098,N_38757);
nor U42471 (N_42471,N_37369,N_39731);
and U42472 (N_42472,N_39125,N_36252);
or U42473 (N_42473,N_36836,N_36090);
nor U42474 (N_42474,N_36088,N_37869);
xnor U42475 (N_42475,N_39248,N_39590);
and U42476 (N_42476,N_39395,N_39198);
xnor U42477 (N_42477,N_38039,N_39346);
xnor U42478 (N_42478,N_37599,N_36379);
and U42479 (N_42479,N_37425,N_36334);
xnor U42480 (N_42480,N_37546,N_36114);
or U42481 (N_42481,N_35733,N_37879);
or U42482 (N_42482,N_37319,N_39682);
and U42483 (N_42483,N_37659,N_37085);
and U42484 (N_42484,N_38093,N_37028);
or U42485 (N_42485,N_36286,N_37188);
xor U42486 (N_42486,N_39144,N_37384);
and U42487 (N_42487,N_36266,N_36221);
nor U42488 (N_42488,N_36740,N_38840);
and U42489 (N_42489,N_35469,N_35673);
nand U42490 (N_42490,N_35786,N_37990);
nand U42491 (N_42491,N_35380,N_39388);
and U42492 (N_42492,N_39929,N_39413);
and U42493 (N_42493,N_36668,N_35591);
nand U42494 (N_42494,N_37424,N_39325);
nor U42495 (N_42495,N_39892,N_38149);
and U42496 (N_42496,N_35847,N_39670);
xor U42497 (N_42497,N_37596,N_39463);
or U42498 (N_42498,N_37839,N_37769);
xnor U42499 (N_42499,N_35740,N_39182);
nand U42500 (N_42500,N_37810,N_37610);
xnor U42501 (N_42501,N_37135,N_39727);
xor U42502 (N_42502,N_38791,N_37841);
or U42503 (N_42503,N_37751,N_38630);
and U42504 (N_42504,N_37044,N_35233);
nand U42505 (N_42505,N_36085,N_37555);
nor U42506 (N_42506,N_35978,N_38753);
nor U42507 (N_42507,N_36100,N_36674);
and U42508 (N_42508,N_38633,N_38659);
and U42509 (N_42509,N_37235,N_38499);
xor U42510 (N_42510,N_35725,N_35490);
nor U42511 (N_42511,N_35910,N_35038);
nand U42512 (N_42512,N_37215,N_39112);
nor U42513 (N_42513,N_35518,N_36319);
nand U42514 (N_42514,N_36143,N_38175);
nand U42515 (N_42515,N_36904,N_36794);
xnor U42516 (N_42516,N_38844,N_36420);
or U42517 (N_42517,N_39050,N_38983);
xor U42518 (N_42518,N_39592,N_39523);
nand U42519 (N_42519,N_38379,N_35881);
xnor U42520 (N_42520,N_36360,N_35908);
nand U42521 (N_42521,N_38186,N_38481);
nand U42522 (N_42522,N_38891,N_38487);
nor U42523 (N_42523,N_37102,N_35421);
nor U42524 (N_42524,N_35328,N_37932);
or U42525 (N_42525,N_36069,N_39608);
or U42526 (N_42526,N_36867,N_36519);
xor U42527 (N_42527,N_36313,N_35622);
nor U42528 (N_42528,N_35504,N_38056);
xnor U42529 (N_42529,N_39987,N_35516);
nand U42530 (N_42530,N_38707,N_39479);
or U42531 (N_42531,N_38660,N_37750);
nand U42532 (N_42532,N_39935,N_38919);
nand U42533 (N_42533,N_37063,N_39784);
xor U42534 (N_42534,N_35757,N_38549);
nand U42535 (N_42535,N_36266,N_35143);
xnor U42536 (N_42536,N_38328,N_39103);
and U42537 (N_42537,N_35811,N_35754);
nor U42538 (N_42538,N_38467,N_37872);
nor U42539 (N_42539,N_36231,N_36099);
or U42540 (N_42540,N_36651,N_38213);
nor U42541 (N_42541,N_36491,N_37201);
xnor U42542 (N_42542,N_38369,N_35108);
or U42543 (N_42543,N_36439,N_38254);
or U42544 (N_42544,N_35770,N_37420);
nand U42545 (N_42545,N_35363,N_35065);
and U42546 (N_42546,N_36364,N_37809);
nand U42547 (N_42547,N_36889,N_37137);
or U42548 (N_42548,N_39567,N_39067);
xor U42549 (N_42549,N_36424,N_37823);
nand U42550 (N_42550,N_35852,N_35112);
nand U42551 (N_42551,N_38908,N_38353);
xor U42552 (N_42552,N_36668,N_39823);
or U42553 (N_42553,N_35776,N_37285);
or U42554 (N_42554,N_35148,N_35376);
and U42555 (N_42555,N_39024,N_37638);
nor U42556 (N_42556,N_36561,N_37493);
and U42557 (N_42557,N_39860,N_37815);
nor U42558 (N_42558,N_38577,N_38513);
nand U42559 (N_42559,N_39461,N_38898);
xor U42560 (N_42560,N_36504,N_37203);
and U42561 (N_42561,N_37618,N_38010);
nand U42562 (N_42562,N_38933,N_38876);
nor U42563 (N_42563,N_36474,N_38649);
or U42564 (N_42564,N_35739,N_38151);
nand U42565 (N_42565,N_35586,N_36429);
nor U42566 (N_42566,N_37801,N_35472);
nor U42567 (N_42567,N_35762,N_37116);
or U42568 (N_42568,N_36537,N_35379);
nand U42569 (N_42569,N_37790,N_36406);
nand U42570 (N_42570,N_38083,N_37336);
or U42571 (N_42571,N_37916,N_37490);
or U42572 (N_42572,N_37114,N_39533);
or U42573 (N_42573,N_37994,N_37410);
nand U42574 (N_42574,N_38838,N_38341);
or U42575 (N_42575,N_36212,N_39779);
or U42576 (N_42576,N_35854,N_39227);
xor U42577 (N_42577,N_36149,N_38496);
nor U42578 (N_42578,N_35366,N_36155);
and U42579 (N_42579,N_38449,N_37786);
or U42580 (N_42580,N_38225,N_37402);
nor U42581 (N_42581,N_36890,N_35346);
and U42582 (N_42582,N_35752,N_36286);
xor U42583 (N_42583,N_35854,N_36380);
xnor U42584 (N_42584,N_35360,N_37996);
nor U42585 (N_42585,N_38985,N_39021);
and U42586 (N_42586,N_36721,N_36465);
nand U42587 (N_42587,N_38290,N_35064);
and U42588 (N_42588,N_37172,N_37008);
nor U42589 (N_42589,N_35488,N_36886);
nor U42590 (N_42590,N_37185,N_39549);
xor U42591 (N_42591,N_37859,N_39396);
nor U42592 (N_42592,N_38744,N_38781);
or U42593 (N_42593,N_38545,N_35443);
or U42594 (N_42594,N_38911,N_38602);
nand U42595 (N_42595,N_35582,N_38092);
nor U42596 (N_42596,N_39778,N_36715);
nand U42597 (N_42597,N_37868,N_38333);
nand U42598 (N_42598,N_38387,N_37147);
nand U42599 (N_42599,N_35726,N_37334);
xor U42600 (N_42600,N_39754,N_35142);
xor U42601 (N_42601,N_36911,N_38978);
xnor U42602 (N_42602,N_36035,N_36745);
nand U42603 (N_42603,N_39446,N_35891);
nand U42604 (N_42604,N_38475,N_36701);
xnor U42605 (N_42605,N_39507,N_39056);
nand U42606 (N_42606,N_35463,N_35894);
and U42607 (N_42607,N_37091,N_37852);
and U42608 (N_42608,N_37188,N_39443);
xor U42609 (N_42609,N_36138,N_37535);
xnor U42610 (N_42610,N_36399,N_35971);
nor U42611 (N_42611,N_38854,N_35328);
xor U42612 (N_42612,N_36619,N_37296);
xor U42613 (N_42613,N_38389,N_37575);
xor U42614 (N_42614,N_39369,N_37087);
xnor U42615 (N_42615,N_36461,N_38717);
nand U42616 (N_42616,N_38667,N_36223);
nand U42617 (N_42617,N_38424,N_37988);
nand U42618 (N_42618,N_37428,N_36425);
nand U42619 (N_42619,N_35986,N_37571);
nor U42620 (N_42620,N_39892,N_39928);
xnor U42621 (N_42621,N_38836,N_35714);
and U42622 (N_42622,N_36730,N_38760);
xor U42623 (N_42623,N_36526,N_38690);
xnor U42624 (N_42624,N_35453,N_37538);
nor U42625 (N_42625,N_37595,N_36127);
xnor U42626 (N_42626,N_36871,N_39609);
nor U42627 (N_42627,N_36358,N_35760);
or U42628 (N_42628,N_35275,N_39389);
or U42629 (N_42629,N_39181,N_35489);
nor U42630 (N_42630,N_38962,N_35172);
nand U42631 (N_42631,N_38992,N_38328);
or U42632 (N_42632,N_39713,N_38359);
nand U42633 (N_42633,N_38243,N_35561);
or U42634 (N_42634,N_37934,N_37128);
and U42635 (N_42635,N_38003,N_37495);
or U42636 (N_42636,N_38551,N_35911);
nor U42637 (N_42637,N_37666,N_37006);
or U42638 (N_42638,N_39085,N_36292);
xor U42639 (N_42639,N_36619,N_37314);
or U42640 (N_42640,N_35100,N_38550);
nor U42641 (N_42641,N_37941,N_39497);
and U42642 (N_42642,N_37961,N_39994);
nor U42643 (N_42643,N_37848,N_35396);
nand U42644 (N_42644,N_38371,N_38944);
nand U42645 (N_42645,N_36291,N_38350);
and U42646 (N_42646,N_38890,N_37604);
or U42647 (N_42647,N_37291,N_36729);
nor U42648 (N_42648,N_38979,N_37333);
or U42649 (N_42649,N_38359,N_35653);
or U42650 (N_42650,N_38622,N_37724);
or U42651 (N_42651,N_37337,N_38742);
and U42652 (N_42652,N_39969,N_35337);
or U42653 (N_42653,N_36056,N_37067);
or U42654 (N_42654,N_36286,N_39283);
xor U42655 (N_42655,N_36510,N_38113);
nor U42656 (N_42656,N_35235,N_35901);
and U42657 (N_42657,N_37263,N_35216);
and U42658 (N_42658,N_37076,N_36841);
xor U42659 (N_42659,N_37917,N_38450);
or U42660 (N_42660,N_35522,N_37172);
xnor U42661 (N_42661,N_35488,N_39607);
xnor U42662 (N_42662,N_39658,N_36438);
and U42663 (N_42663,N_36215,N_39666);
nor U42664 (N_42664,N_36288,N_35088);
xnor U42665 (N_42665,N_38923,N_37011);
and U42666 (N_42666,N_38232,N_39919);
xor U42667 (N_42667,N_37510,N_36962);
nand U42668 (N_42668,N_39886,N_36423);
or U42669 (N_42669,N_39161,N_37148);
nor U42670 (N_42670,N_39488,N_36273);
and U42671 (N_42671,N_36714,N_38324);
xnor U42672 (N_42672,N_39278,N_35788);
nor U42673 (N_42673,N_38665,N_35727);
nor U42674 (N_42674,N_35127,N_35221);
nand U42675 (N_42675,N_39704,N_37922);
xnor U42676 (N_42676,N_39257,N_35816);
nor U42677 (N_42677,N_39373,N_38927);
or U42678 (N_42678,N_36504,N_39731);
nand U42679 (N_42679,N_36397,N_36656);
and U42680 (N_42680,N_35814,N_36370);
nand U42681 (N_42681,N_38802,N_39871);
and U42682 (N_42682,N_37403,N_39993);
nand U42683 (N_42683,N_35444,N_35285);
xnor U42684 (N_42684,N_37018,N_39427);
xor U42685 (N_42685,N_36539,N_38984);
nand U42686 (N_42686,N_39336,N_36231);
nand U42687 (N_42687,N_39933,N_35638);
and U42688 (N_42688,N_35970,N_36033);
nor U42689 (N_42689,N_38389,N_37548);
nor U42690 (N_42690,N_37693,N_38772);
nand U42691 (N_42691,N_37183,N_37097);
nand U42692 (N_42692,N_35742,N_35797);
or U42693 (N_42693,N_39217,N_35487);
nand U42694 (N_42694,N_36800,N_39097);
nand U42695 (N_42695,N_35976,N_38096);
nor U42696 (N_42696,N_35009,N_38217);
xor U42697 (N_42697,N_35590,N_37134);
or U42698 (N_42698,N_37733,N_36044);
and U42699 (N_42699,N_38893,N_38188);
and U42700 (N_42700,N_39841,N_35312);
and U42701 (N_42701,N_35113,N_38254);
or U42702 (N_42702,N_36339,N_35560);
xor U42703 (N_42703,N_36675,N_36941);
and U42704 (N_42704,N_39645,N_39266);
nor U42705 (N_42705,N_38787,N_37884);
xor U42706 (N_42706,N_37053,N_39757);
nor U42707 (N_42707,N_37856,N_35529);
and U42708 (N_42708,N_38149,N_37994);
nor U42709 (N_42709,N_38237,N_39590);
nor U42710 (N_42710,N_36570,N_36278);
or U42711 (N_42711,N_37628,N_39247);
nand U42712 (N_42712,N_39228,N_38744);
nand U42713 (N_42713,N_35465,N_35039);
nand U42714 (N_42714,N_38126,N_35501);
nor U42715 (N_42715,N_36887,N_37130);
or U42716 (N_42716,N_36136,N_37337);
and U42717 (N_42717,N_39568,N_35704);
xor U42718 (N_42718,N_39270,N_37998);
nand U42719 (N_42719,N_36058,N_37963);
and U42720 (N_42720,N_35608,N_39188);
nor U42721 (N_42721,N_39639,N_35232);
nor U42722 (N_42722,N_35673,N_37546);
nor U42723 (N_42723,N_38151,N_37301);
nor U42724 (N_42724,N_39424,N_36849);
xor U42725 (N_42725,N_39023,N_38657);
nand U42726 (N_42726,N_35027,N_37538);
xor U42727 (N_42727,N_36868,N_36204);
nor U42728 (N_42728,N_37023,N_35522);
nand U42729 (N_42729,N_35323,N_39785);
nand U42730 (N_42730,N_37567,N_39607);
nand U42731 (N_42731,N_36736,N_38531);
and U42732 (N_42732,N_36029,N_38524);
and U42733 (N_42733,N_38272,N_36658);
nor U42734 (N_42734,N_36661,N_39980);
nor U42735 (N_42735,N_37430,N_38754);
or U42736 (N_42736,N_37840,N_39033);
and U42737 (N_42737,N_35486,N_36189);
nand U42738 (N_42738,N_39713,N_38710);
nand U42739 (N_42739,N_35854,N_35741);
nor U42740 (N_42740,N_39052,N_37729);
and U42741 (N_42741,N_36967,N_35007);
and U42742 (N_42742,N_37091,N_38883);
nor U42743 (N_42743,N_38127,N_35447);
and U42744 (N_42744,N_35207,N_37562);
nand U42745 (N_42745,N_35820,N_36145);
xor U42746 (N_42746,N_36342,N_36977);
xor U42747 (N_42747,N_39920,N_36996);
nor U42748 (N_42748,N_35822,N_38991);
or U42749 (N_42749,N_38415,N_36023);
nand U42750 (N_42750,N_35718,N_39133);
nand U42751 (N_42751,N_38625,N_35567);
or U42752 (N_42752,N_37742,N_38291);
nand U42753 (N_42753,N_37497,N_38916);
or U42754 (N_42754,N_37944,N_39809);
xnor U42755 (N_42755,N_38650,N_35313);
nand U42756 (N_42756,N_36464,N_35559);
or U42757 (N_42757,N_37502,N_36952);
nor U42758 (N_42758,N_37583,N_37120);
or U42759 (N_42759,N_35909,N_36494);
or U42760 (N_42760,N_38958,N_36127);
xnor U42761 (N_42761,N_35100,N_39238);
nor U42762 (N_42762,N_36601,N_38736);
nand U42763 (N_42763,N_35569,N_39561);
nand U42764 (N_42764,N_38899,N_35329);
or U42765 (N_42765,N_36762,N_38424);
and U42766 (N_42766,N_39797,N_36908);
xnor U42767 (N_42767,N_39948,N_37283);
nand U42768 (N_42768,N_36749,N_36950);
and U42769 (N_42769,N_37760,N_37691);
xor U42770 (N_42770,N_36952,N_35067);
or U42771 (N_42771,N_36045,N_36140);
xnor U42772 (N_42772,N_35572,N_37118);
nand U42773 (N_42773,N_39431,N_36678);
nand U42774 (N_42774,N_39756,N_39762);
nor U42775 (N_42775,N_37425,N_38668);
nor U42776 (N_42776,N_39828,N_37720);
or U42777 (N_42777,N_38845,N_35902);
and U42778 (N_42778,N_39942,N_37033);
nand U42779 (N_42779,N_38033,N_35186);
nand U42780 (N_42780,N_39315,N_36967);
nand U42781 (N_42781,N_35934,N_37807);
or U42782 (N_42782,N_37195,N_38624);
or U42783 (N_42783,N_35113,N_36306);
or U42784 (N_42784,N_39163,N_35389);
and U42785 (N_42785,N_35291,N_35968);
nor U42786 (N_42786,N_36323,N_35770);
nand U42787 (N_42787,N_39068,N_37306);
or U42788 (N_42788,N_35460,N_39946);
nor U42789 (N_42789,N_36823,N_37700);
xnor U42790 (N_42790,N_38420,N_36013);
or U42791 (N_42791,N_39732,N_35262);
or U42792 (N_42792,N_37119,N_37736);
xnor U42793 (N_42793,N_36453,N_36105);
and U42794 (N_42794,N_37683,N_38211);
and U42795 (N_42795,N_37964,N_38181);
and U42796 (N_42796,N_36843,N_39330);
nor U42797 (N_42797,N_39443,N_37493);
xor U42798 (N_42798,N_35113,N_38136);
nand U42799 (N_42799,N_39531,N_39088);
nor U42800 (N_42800,N_38496,N_39056);
and U42801 (N_42801,N_35197,N_37164);
and U42802 (N_42802,N_37977,N_38886);
nand U42803 (N_42803,N_38779,N_36490);
nand U42804 (N_42804,N_38450,N_37195);
and U42805 (N_42805,N_38702,N_37347);
nor U42806 (N_42806,N_37107,N_39952);
nor U42807 (N_42807,N_37825,N_35360);
nand U42808 (N_42808,N_35150,N_38355);
and U42809 (N_42809,N_39913,N_36219);
and U42810 (N_42810,N_35394,N_36770);
nor U42811 (N_42811,N_37527,N_35373);
nor U42812 (N_42812,N_38454,N_37962);
and U42813 (N_42813,N_36214,N_37218);
nand U42814 (N_42814,N_39936,N_37230);
nor U42815 (N_42815,N_37209,N_36459);
or U42816 (N_42816,N_38239,N_39442);
and U42817 (N_42817,N_36740,N_39071);
or U42818 (N_42818,N_36099,N_36477);
nand U42819 (N_42819,N_35284,N_38525);
xor U42820 (N_42820,N_35873,N_36218);
nor U42821 (N_42821,N_39796,N_35671);
xor U42822 (N_42822,N_39577,N_39748);
xnor U42823 (N_42823,N_39491,N_36251);
or U42824 (N_42824,N_35742,N_36927);
nor U42825 (N_42825,N_39512,N_38874);
nand U42826 (N_42826,N_36383,N_38277);
nand U42827 (N_42827,N_35325,N_37950);
nand U42828 (N_42828,N_39164,N_36233);
nor U42829 (N_42829,N_38425,N_38853);
nand U42830 (N_42830,N_38158,N_36626);
xnor U42831 (N_42831,N_39939,N_39597);
xnor U42832 (N_42832,N_38823,N_37698);
nand U42833 (N_42833,N_35507,N_38446);
xor U42834 (N_42834,N_38154,N_36237);
nand U42835 (N_42835,N_37473,N_36201);
nor U42836 (N_42836,N_37197,N_39460);
xor U42837 (N_42837,N_36968,N_38567);
and U42838 (N_42838,N_37555,N_36824);
or U42839 (N_42839,N_35328,N_39276);
nand U42840 (N_42840,N_36598,N_39225);
xnor U42841 (N_42841,N_38126,N_35122);
nand U42842 (N_42842,N_36054,N_37144);
nand U42843 (N_42843,N_37772,N_35435);
nand U42844 (N_42844,N_36230,N_39251);
and U42845 (N_42845,N_37009,N_38147);
and U42846 (N_42846,N_37602,N_36965);
nor U42847 (N_42847,N_36815,N_35439);
nand U42848 (N_42848,N_39242,N_37664);
nand U42849 (N_42849,N_39768,N_36828);
or U42850 (N_42850,N_37272,N_37935);
and U42851 (N_42851,N_36515,N_39723);
xnor U42852 (N_42852,N_35070,N_37944);
xnor U42853 (N_42853,N_39992,N_39905);
and U42854 (N_42854,N_36447,N_35465);
xnor U42855 (N_42855,N_38548,N_39115);
and U42856 (N_42856,N_38654,N_38514);
or U42857 (N_42857,N_36222,N_36215);
or U42858 (N_42858,N_35763,N_37911);
or U42859 (N_42859,N_36554,N_38762);
xor U42860 (N_42860,N_39229,N_37297);
or U42861 (N_42861,N_38586,N_36101);
nor U42862 (N_42862,N_39328,N_37920);
and U42863 (N_42863,N_37124,N_37157);
and U42864 (N_42864,N_35994,N_39020);
or U42865 (N_42865,N_36849,N_36806);
and U42866 (N_42866,N_37880,N_38620);
nand U42867 (N_42867,N_38778,N_37665);
xor U42868 (N_42868,N_39618,N_39274);
xor U42869 (N_42869,N_35397,N_38827);
and U42870 (N_42870,N_38034,N_35438);
and U42871 (N_42871,N_38913,N_38957);
xnor U42872 (N_42872,N_35341,N_36371);
nand U42873 (N_42873,N_35157,N_39391);
or U42874 (N_42874,N_37985,N_35325);
nand U42875 (N_42875,N_35653,N_35313);
nand U42876 (N_42876,N_38356,N_39492);
xor U42877 (N_42877,N_37378,N_35545);
xor U42878 (N_42878,N_35048,N_38515);
and U42879 (N_42879,N_36738,N_39460);
nand U42880 (N_42880,N_36772,N_35977);
or U42881 (N_42881,N_39565,N_36997);
or U42882 (N_42882,N_39088,N_36025);
or U42883 (N_42883,N_39698,N_35412);
nand U42884 (N_42884,N_35025,N_36781);
xor U42885 (N_42885,N_36239,N_39759);
xnor U42886 (N_42886,N_39895,N_36365);
and U42887 (N_42887,N_39945,N_38598);
and U42888 (N_42888,N_35643,N_38305);
xnor U42889 (N_42889,N_35960,N_37555);
and U42890 (N_42890,N_35490,N_36962);
nor U42891 (N_42891,N_36732,N_38133);
nor U42892 (N_42892,N_39515,N_39787);
or U42893 (N_42893,N_35582,N_36627);
xnor U42894 (N_42894,N_38091,N_37431);
xor U42895 (N_42895,N_35751,N_38007);
or U42896 (N_42896,N_38021,N_36351);
and U42897 (N_42897,N_39357,N_39744);
and U42898 (N_42898,N_39268,N_37669);
or U42899 (N_42899,N_36935,N_35043);
xor U42900 (N_42900,N_35013,N_39041);
or U42901 (N_42901,N_37714,N_39065);
xnor U42902 (N_42902,N_36407,N_35122);
nor U42903 (N_42903,N_39062,N_37938);
and U42904 (N_42904,N_35967,N_37103);
nor U42905 (N_42905,N_39857,N_36969);
and U42906 (N_42906,N_36049,N_38921);
nand U42907 (N_42907,N_38580,N_38683);
or U42908 (N_42908,N_36724,N_36557);
and U42909 (N_42909,N_39610,N_37347);
nand U42910 (N_42910,N_36201,N_39748);
xor U42911 (N_42911,N_39141,N_36908);
and U42912 (N_42912,N_35326,N_36260);
and U42913 (N_42913,N_38158,N_38411);
xnor U42914 (N_42914,N_38277,N_38340);
xnor U42915 (N_42915,N_39140,N_35556);
or U42916 (N_42916,N_35787,N_39238);
nor U42917 (N_42917,N_38479,N_38639);
xor U42918 (N_42918,N_37313,N_35466);
or U42919 (N_42919,N_39310,N_39510);
and U42920 (N_42920,N_35276,N_38790);
and U42921 (N_42921,N_38292,N_35145);
nor U42922 (N_42922,N_39133,N_39541);
xor U42923 (N_42923,N_35165,N_35910);
or U42924 (N_42924,N_37360,N_37708);
and U42925 (N_42925,N_39756,N_35954);
xnor U42926 (N_42926,N_38463,N_35692);
and U42927 (N_42927,N_36514,N_35603);
nor U42928 (N_42928,N_35771,N_39481);
nor U42929 (N_42929,N_37923,N_37021);
nor U42930 (N_42930,N_38930,N_37732);
and U42931 (N_42931,N_39322,N_39756);
and U42932 (N_42932,N_37753,N_37915);
xnor U42933 (N_42933,N_36477,N_36751);
and U42934 (N_42934,N_39723,N_36974);
and U42935 (N_42935,N_39055,N_35509);
xor U42936 (N_42936,N_38032,N_37845);
nor U42937 (N_42937,N_38130,N_35615);
nor U42938 (N_42938,N_35262,N_35256);
nand U42939 (N_42939,N_37486,N_37127);
nor U42940 (N_42940,N_37208,N_38147);
nor U42941 (N_42941,N_36574,N_37633);
or U42942 (N_42942,N_39868,N_36463);
or U42943 (N_42943,N_39671,N_36924);
nor U42944 (N_42944,N_36746,N_39490);
or U42945 (N_42945,N_36943,N_38779);
nand U42946 (N_42946,N_35149,N_35115);
nand U42947 (N_42947,N_36808,N_37971);
xnor U42948 (N_42948,N_35684,N_37174);
or U42949 (N_42949,N_38780,N_38279);
nand U42950 (N_42950,N_38173,N_37634);
or U42951 (N_42951,N_38663,N_37884);
xnor U42952 (N_42952,N_36493,N_39600);
or U42953 (N_42953,N_35651,N_35877);
nor U42954 (N_42954,N_36133,N_35465);
and U42955 (N_42955,N_38019,N_36394);
xnor U42956 (N_42956,N_36051,N_37123);
or U42957 (N_42957,N_37147,N_39181);
and U42958 (N_42958,N_39325,N_38736);
or U42959 (N_42959,N_36168,N_38105);
xnor U42960 (N_42960,N_36807,N_36827);
xnor U42961 (N_42961,N_38592,N_39422);
and U42962 (N_42962,N_35029,N_38163);
xor U42963 (N_42963,N_38841,N_39065);
nor U42964 (N_42964,N_35972,N_36683);
and U42965 (N_42965,N_39489,N_36987);
nor U42966 (N_42966,N_36916,N_37615);
or U42967 (N_42967,N_39186,N_35669);
nand U42968 (N_42968,N_36851,N_39677);
xnor U42969 (N_42969,N_35427,N_37557);
xor U42970 (N_42970,N_35466,N_35536);
nand U42971 (N_42971,N_37264,N_38280);
xnor U42972 (N_42972,N_37747,N_38821);
and U42973 (N_42973,N_35129,N_36180);
or U42974 (N_42974,N_37989,N_38565);
xnor U42975 (N_42975,N_37050,N_36757);
nand U42976 (N_42976,N_39589,N_35556);
nand U42977 (N_42977,N_38836,N_38412);
nor U42978 (N_42978,N_38781,N_36481);
and U42979 (N_42979,N_37040,N_39335);
xor U42980 (N_42980,N_35368,N_39767);
xor U42981 (N_42981,N_36661,N_38513);
nor U42982 (N_42982,N_38532,N_38830);
xor U42983 (N_42983,N_35730,N_38968);
nor U42984 (N_42984,N_36159,N_39421);
xnor U42985 (N_42985,N_39864,N_39210);
xor U42986 (N_42986,N_38953,N_36774);
nor U42987 (N_42987,N_36809,N_37581);
or U42988 (N_42988,N_35682,N_36313);
xnor U42989 (N_42989,N_36978,N_39552);
nand U42990 (N_42990,N_39732,N_38852);
or U42991 (N_42991,N_35987,N_38339);
nand U42992 (N_42992,N_38740,N_38693);
nor U42993 (N_42993,N_37692,N_38705);
nor U42994 (N_42994,N_36889,N_38791);
nand U42995 (N_42995,N_37525,N_36818);
nor U42996 (N_42996,N_39477,N_35455);
nor U42997 (N_42997,N_38540,N_39519);
and U42998 (N_42998,N_36876,N_39499);
nor U42999 (N_42999,N_36037,N_37244);
nor U43000 (N_43000,N_38783,N_38180);
nand U43001 (N_43001,N_39405,N_36342);
and U43002 (N_43002,N_36490,N_39949);
and U43003 (N_43003,N_37660,N_39942);
and U43004 (N_43004,N_35897,N_37125);
nand U43005 (N_43005,N_39997,N_37537);
or U43006 (N_43006,N_35882,N_37400);
or U43007 (N_43007,N_37506,N_39370);
or U43008 (N_43008,N_38223,N_38713);
xnor U43009 (N_43009,N_39521,N_38061);
or U43010 (N_43010,N_38682,N_36466);
xor U43011 (N_43011,N_37942,N_35715);
and U43012 (N_43012,N_39974,N_39634);
nand U43013 (N_43013,N_37884,N_35126);
nor U43014 (N_43014,N_36109,N_37940);
and U43015 (N_43015,N_36814,N_38945);
or U43016 (N_43016,N_35090,N_35000);
or U43017 (N_43017,N_38044,N_39217);
nand U43018 (N_43018,N_35195,N_35427);
nor U43019 (N_43019,N_36962,N_36813);
nand U43020 (N_43020,N_36320,N_39595);
nor U43021 (N_43021,N_39870,N_36882);
nand U43022 (N_43022,N_36095,N_39538);
nor U43023 (N_43023,N_36167,N_35247);
nor U43024 (N_43024,N_38998,N_36466);
nand U43025 (N_43025,N_37168,N_38922);
and U43026 (N_43026,N_35223,N_37276);
nand U43027 (N_43027,N_37564,N_37071);
nand U43028 (N_43028,N_38255,N_38594);
xor U43029 (N_43029,N_36444,N_37110);
xnor U43030 (N_43030,N_39388,N_36458);
nor U43031 (N_43031,N_36750,N_36063);
or U43032 (N_43032,N_38576,N_37798);
nor U43033 (N_43033,N_36993,N_36028);
nand U43034 (N_43034,N_38859,N_38484);
and U43035 (N_43035,N_38382,N_39043);
nand U43036 (N_43036,N_39028,N_39095);
nand U43037 (N_43037,N_35168,N_37827);
or U43038 (N_43038,N_38606,N_38557);
nand U43039 (N_43039,N_37762,N_36174);
nor U43040 (N_43040,N_38748,N_39982);
nand U43041 (N_43041,N_36827,N_35826);
and U43042 (N_43042,N_37774,N_36187);
or U43043 (N_43043,N_35683,N_36599);
xnor U43044 (N_43044,N_35372,N_36250);
nand U43045 (N_43045,N_36692,N_38654);
nand U43046 (N_43046,N_36492,N_35177);
xor U43047 (N_43047,N_38901,N_38613);
and U43048 (N_43048,N_36354,N_37702);
xnor U43049 (N_43049,N_38005,N_37542);
or U43050 (N_43050,N_37551,N_37313);
or U43051 (N_43051,N_38124,N_37038);
or U43052 (N_43052,N_37832,N_38984);
and U43053 (N_43053,N_39176,N_35524);
and U43054 (N_43054,N_37980,N_38890);
or U43055 (N_43055,N_35782,N_38902);
nor U43056 (N_43056,N_38607,N_38545);
nand U43057 (N_43057,N_39106,N_39350);
or U43058 (N_43058,N_36622,N_35612);
or U43059 (N_43059,N_39646,N_39978);
and U43060 (N_43060,N_37467,N_39595);
nor U43061 (N_43061,N_37231,N_35089);
nor U43062 (N_43062,N_37614,N_39915);
or U43063 (N_43063,N_38349,N_39112);
nand U43064 (N_43064,N_38008,N_38331);
nand U43065 (N_43065,N_37289,N_38744);
nor U43066 (N_43066,N_38641,N_39322);
xnor U43067 (N_43067,N_36771,N_35543);
or U43068 (N_43068,N_35710,N_37297);
and U43069 (N_43069,N_35687,N_39427);
nor U43070 (N_43070,N_36801,N_35372);
nor U43071 (N_43071,N_35658,N_35299);
nor U43072 (N_43072,N_37699,N_37593);
nand U43073 (N_43073,N_35708,N_37528);
nand U43074 (N_43074,N_38360,N_37681);
xnor U43075 (N_43075,N_38361,N_39403);
and U43076 (N_43076,N_37400,N_37259);
nor U43077 (N_43077,N_39819,N_35379);
xor U43078 (N_43078,N_35067,N_38499);
or U43079 (N_43079,N_38872,N_35875);
xor U43080 (N_43080,N_38202,N_36101);
xor U43081 (N_43081,N_37264,N_38783);
or U43082 (N_43082,N_35287,N_37364);
or U43083 (N_43083,N_37470,N_37021);
and U43084 (N_43084,N_38980,N_38904);
and U43085 (N_43085,N_35778,N_39433);
or U43086 (N_43086,N_35567,N_39242);
nor U43087 (N_43087,N_39786,N_36107);
and U43088 (N_43088,N_35132,N_38885);
nor U43089 (N_43089,N_38226,N_39501);
nand U43090 (N_43090,N_35841,N_35384);
nand U43091 (N_43091,N_37430,N_39494);
xnor U43092 (N_43092,N_39963,N_38955);
xnor U43093 (N_43093,N_37379,N_38461);
nand U43094 (N_43094,N_37432,N_37107);
or U43095 (N_43095,N_38626,N_36417);
nor U43096 (N_43096,N_35978,N_39635);
nor U43097 (N_43097,N_36598,N_37620);
or U43098 (N_43098,N_39506,N_39428);
and U43099 (N_43099,N_38636,N_36866);
or U43100 (N_43100,N_36679,N_37336);
nand U43101 (N_43101,N_35061,N_36993);
and U43102 (N_43102,N_39613,N_35385);
nand U43103 (N_43103,N_39041,N_35960);
xnor U43104 (N_43104,N_39771,N_36997);
nand U43105 (N_43105,N_38430,N_36284);
xnor U43106 (N_43106,N_38031,N_38976);
xnor U43107 (N_43107,N_39740,N_39496);
xor U43108 (N_43108,N_38839,N_39405);
or U43109 (N_43109,N_36167,N_38978);
xnor U43110 (N_43110,N_38282,N_37774);
or U43111 (N_43111,N_36900,N_37682);
and U43112 (N_43112,N_35212,N_39034);
nand U43113 (N_43113,N_37713,N_36485);
nand U43114 (N_43114,N_36155,N_35039);
and U43115 (N_43115,N_35003,N_37195);
nor U43116 (N_43116,N_36811,N_36540);
nand U43117 (N_43117,N_38189,N_37233);
nor U43118 (N_43118,N_37417,N_38883);
xnor U43119 (N_43119,N_35866,N_38098);
nand U43120 (N_43120,N_39707,N_38058);
nand U43121 (N_43121,N_36682,N_35794);
nand U43122 (N_43122,N_39995,N_35050);
nand U43123 (N_43123,N_39941,N_39633);
nand U43124 (N_43124,N_36425,N_35682);
nor U43125 (N_43125,N_35446,N_35171);
and U43126 (N_43126,N_39392,N_37848);
or U43127 (N_43127,N_37986,N_39148);
xor U43128 (N_43128,N_35904,N_36455);
nor U43129 (N_43129,N_36979,N_37803);
xnor U43130 (N_43130,N_36241,N_39258);
nand U43131 (N_43131,N_36980,N_37891);
or U43132 (N_43132,N_38069,N_35260);
xnor U43133 (N_43133,N_37981,N_37199);
nor U43134 (N_43134,N_35846,N_38458);
nand U43135 (N_43135,N_38818,N_37526);
xor U43136 (N_43136,N_38193,N_35061);
nor U43137 (N_43137,N_37325,N_35844);
and U43138 (N_43138,N_39900,N_37543);
or U43139 (N_43139,N_39529,N_37886);
or U43140 (N_43140,N_39356,N_35443);
nor U43141 (N_43141,N_38527,N_38265);
xnor U43142 (N_43142,N_39556,N_38616);
nand U43143 (N_43143,N_39003,N_35220);
and U43144 (N_43144,N_35334,N_36667);
xnor U43145 (N_43145,N_35703,N_39409);
nor U43146 (N_43146,N_37711,N_38374);
nor U43147 (N_43147,N_39590,N_38353);
nand U43148 (N_43148,N_36891,N_37031);
or U43149 (N_43149,N_36789,N_38258);
xor U43150 (N_43150,N_38365,N_38165);
or U43151 (N_43151,N_35160,N_39282);
nor U43152 (N_43152,N_38056,N_38852);
nor U43153 (N_43153,N_35629,N_39635);
xnor U43154 (N_43154,N_37983,N_36624);
xnor U43155 (N_43155,N_39356,N_38499);
nor U43156 (N_43156,N_37977,N_35075);
and U43157 (N_43157,N_35850,N_39264);
nand U43158 (N_43158,N_36891,N_38892);
and U43159 (N_43159,N_35350,N_36165);
xnor U43160 (N_43160,N_35509,N_36583);
or U43161 (N_43161,N_35014,N_36395);
and U43162 (N_43162,N_35302,N_38613);
and U43163 (N_43163,N_39565,N_35972);
and U43164 (N_43164,N_39971,N_39160);
nor U43165 (N_43165,N_37997,N_39431);
or U43166 (N_43166,N_39629,N_37009);
nor U43167 (N_43167,N_38647,N_38900);
nand U43168 (N_43168,N_37826,N_37894);
xor U43169 (N_43169,N_36084,N_35871);
xnor U43170 (N_43170,N_39662,N_39268);
xor U43171 (N_43171,N_36961,N_39462);
and U43172 (N_43172,N_39801,N_39620);
and U43173 (N_43173,N_39847,N_39941);
nor U43174 (N_43174,N_35102,N_36751);
or U43175 (N_43175,N_37628,N_39027);
and U43176 (N_43176,N_36785,N_35900);
and U43177 (N_43177,N_35080,N_36984);
nor U43178 (N_43178,N_36787,N_37220);
and U43179 (N_43179,N_36704,N_37572);
nand U43180 (N_43180,N_36342,N_38876);
nor U43181 (N_43181,N_36793,N_37843);
xnor U43182 (N_43182,N_37524,N_39234);
nor U43183 (N_43183,N_35150,N_37030);
and U43184 (N_43184,N_37169,N_35179);
nand U43185 (N_43185,N_38611,N_38870);
nor U43186 (N_43186,N_36690,N_35773);
nand U43187 (N_43187,N_38396,N_35898);
nand U43188 (N_43188,N_35294,N_37010);
or U43189 (N_43189,N_35033,N_37807);
or U43190 (N_43190,N_35449,N_39881);
nand U43191 (N_43191,N_37136,N_37992);
nand U43192 (N_43192,N_38309,N_36496);
and U43193 (N_43193,N_35489,N_38428);
nor U43194 (N_43194,N_37360,N_35753);
nand U43195 (N_43195,N_39633,N_38516);
or U43196 (N_43196,N_39228,N_36802);
or U43197 (N_43197,N_35608,N_36318);
nand U43198 (N_43198,N_36006,N_36038);
or U43199 (N_43199,N_36236,N_37937);
nor U43200 (N_43200,N_35918,N_37536);
nand U43201 (N_43201,N_36789,N_35388);
and U43202 (N_43202,N_35274,N_35390);
nand U43203 (N_43203,N_35898,N_39523);
nand U43204 (N_43204,N_38218,N_37721);
and U43205 (N_43205,N_37953,N_38001);
or U43206 (N_43206,N_39688,N_39934);
and U43207 (N_43207,N_39224,N_38133);
and U43208 (N_43208,N_35833,N_38342);
and U43209 (N_43209,N_35416,N_36588);
nor U43210 (N_43210,N_35122,N_39375);
nand U43211 (N_43211,N_35516,N_36232);
nand U43212 (N_43212,N_39566,N_35297);
and U43213 (N_43213,N_35582,N_35596);
nor U43214 (N_43214,N_36863,N_35955);
and U43215 (N_43215,N_39427,N_36322);
and U43216 (N_43216,N_39554,N_38103);
xnor U43217 (N_43217,N_37891,N_36122);
nand U43218 (N_43218,N_35689,N_35017);
xnor U43219 (N_43219,N_37503,N_35105);
xor U43220 (N_43220,N_39570,N_37045);
nand U43221 (N_43221,N_36725,N_36977);
and U43222 (N_43222,N_35427,N_35758);
and U43223 (N_43223,N_38616,N_37885);
or U43224 (N_43224,N_35869,N_36987);
xor U43225 (N_43225,N_35658,N_37660);
nand U43226 (N_43226,N_38580,N_35876);
nand U43227 (N_43227,N_39050,N_38767);
xnor U43228 (N_43228,N_35634,N_36670);
nand U43229 (N_43229,N_37065,N_38161);
and U43230 (N_43230,N_38073,N_39378);
xnor U43231 (N_43231,N_36368,N_38276);
or U43232 (N_43232,N_37387,N_35910);
xnor U43233 (N_43233,N_38091,N_35475);
nand U43234 (N_43234,N_37466,N_36754);
and U43235 (N_43235,N_38141,N_35349);
nand U43236 (N_43236,N_37374,N_37831);
nand U43237 (N_43237,N_37218,N_37810);
and U43238 (N_43238,N_38617,N_37262);
xor U43239 (N_43239,N_37175,N_37509);
nor U43240 (N_43240,N_35020,N_37810);
or U43241 (N_43241,N_38740,N_36482);
nor U43242 (N_43242,N_39794,N_36861);
or U43243 (N_43243,N_38087,N_39744);
or U43244 (N_43244,N_38436,N_39467);
nand U43245 (N_43245,N_39005,N_37568);
nand U43246 (N_43246,N_37497,N_38575);
xor U43247 (N_43247,N_36848,N_39269);
nor U43248 (N_43248,N_35738,N_35520);
nand U43249 (N_43249,N_37244,N_38809);
nor U43250 (N_43250,N_36580,N_37244);
nand U43251 (N_43251,N_37308,N_36580);
xnor U43252 (N_43252,N_38324,N_39425);
nand U43253 (N_43253,N_39872,N_37116);
or U43254 (N_43254,N_39307,N_36584);
or U43255 (N_43255,N_35391,N_38699);
nor U43256 (N_43256,N_36338,N_35770);
nand U43257 (N_43257,N_38827,N_35324);
nor U43258 (N_43258,N_39842,N_39555);
or U43259 (N_43259,N_36949,N_38433);
or U43260 (N_43260,N_36337,N_38594);
xor U43261 (N_43261,N_37147,N_36410);
or U43262 (N_43262,N_38857,N_35392);
or U43263 (N_43263,N_39280,N_35665);
nand U43264 (N_43264,N_38855,N_38367);
and U43265 (N_43265,N_36038,N_38692);
and U43266 (N_43266,N_37638,N_39260);
nor U43267 (N_43267,N_39714,N_39482);
nor U43268 (N_43268,N_36620,N_39949);
nand U43269 (N_43269,N_38810,N_35642);
nor U43270 (N_43270,N_35837,N_37118);
nand U43271 (N_43271,N_35140,N_38743);
and U43272 (N_43272,N_37421,N_37485);
or U43273 (N_43273,N_39473,N_35847);
or U43274 (N_43274,N_37832,N_38084);
xnor U43275 (N_43275,N_38615,N_36603);
nand U43276 (N_43276,N_38599,N_36709);
or U43277 (N_43277,N_36239,N_35088);
or U43278 (N_43278,N_35995,N_35621);
nand U43279 (N_43279,N_35220,N_39784);
nor U43280 (N_43280,N_37880,N_36229);
and U43281 (N_43281,N_35998,N_38571);
nor U43282 (N_43282,N_37984,N_36540);
nor U43283 (N_43283,N_36289,N_35010);
nand U43284 (N_43284,N_35842,N_37604);
xor U43285 (N_43285,N_37886,N_39924);
or U43286 (N_43286,N_39527,N_36115);
and U43287 (N_43287,N_38097,N_38092);
nand U43288 (N_43288,N_35065,N_37318);
or U43289 (N_43289,N_36039,N_35951);
or U43290 (N_43290,N_39522,N_38743);
nor U43291 (N_43291,N_38878,N_37995);
and U43292 (N_43292,N_35422,N_38629);
nor U43293 (N_43293,N_39106,N_39651);
or U43294 (N_43294,N_37087,N_35838);
xor U43295 (N_43295,N_35179,N_37139);
nand U43296 (N_43296,N_36767,N_39751);
or U43297 (N_43297,N_39846,N_39399);
xor U43298 (N_43298,N_35523,N_38957);
and U43299 (N_43299,N_37559,N_35232);
nand U43300 (N_43300,N_36845,N_37813);
nor U43301 (N_43301,N_35337,N_35990);
xnor U43302 (N_43302,N_39467,N_35967);
nand U43303 (N_43303,N_35391,N_35142);
xnor U43304 (N_43304,N_35425,N_38479);
and U43305 (N_43305,N_35903,N_35498);
nand U43306 (N_43306,N_38480,N_37608);
nand U43307 (N_43307,N_35450,N_36564);
or U43308 (N_43308,N_35889,N_38939);
or U43309 (N_43309,N_36264,N_35319);
xnor U43310 (N_43310,N_39112,N_36513);
nor U43311 (N_43311,N_35479,N_38631);
xnor U43312 (N_43312,N_36976,N_36934);
nor U43313 (N_43313,N_39760,N_39663);
xor U43314 (N_43314,N_37112,N_37607);
nor U43315 (N_43315,N_38580,N_35933);
and U43316 (N_43316,N_39412,N_39706);
or U43317 (N_43317,N_39140,N_39656);
or U43318 (N_43318,N_36513,N_38724);
and U43319 (N_43319,N_37546,N_35837);
and U43320 (N_43320,N_39901,N_37071);
or U43321 (N_43321,N_35005,N_36180);
or U43322 (N_43322,N_39956,N_37453);
nor U43323 (N_43323,N_37632,N_37911);
or U43324 (N_43324,N_36632,N_36774);
and U43325 (N_43325,N_35276,N_37470);
nor U43326 (N_43326,N_39294,N_38126);
nor U43327 (N_43327,N_35933,N_38244);
xor U43328 (N_43328,N_38712,N_37162);
or U43329 (N_43329,N_38740,N_38484);
and U43330 (N_43330,N_38172,N_39653);
nand U43331 (N_43331,N_37598,N_35515);
xor U43332 (N_43332,N_35283,N_35145);
nor U43333 (N_43333,N_37555,N_37075);
nand U43334 (N_43334,N_39836,N_36886);
or U43335 (N_43335,N_39112,N_35662);
nor U43336 (N_43336,N_38820,N_37919);
and U43337 (N_43337,N_37133,N_35908);
xor U43338 (N_43338,N_38083,N_36522);
nand U43339 (N_43339,N_37540,N_35730);
nor U43340 (N_43340,N_35523,N_39196);
nand U43341 (N_43341,N_35506,N_39708);
nand U43342 (N_43342,N_38935,N_39600);
nor U43343 (N_43343,N_35097,N_37337);
and U43344 (N_43344,N_36045,N_39440);
nor U43345 (N_43345,N_38925,N_37286);
and U43346 (N_43346,N_37444,N_36503);
or U43347 (N_43347,N_38036,N_36364);
and U43348 (N_43348,N_35933,N_35710);
or U43349 (N_43349,N_38516,N_39085);
nor U43350 (N_43350,N_37593,N_37508);
nand U43351 (N_43351,N_39300,N_36396);
nor U43352 (N_43352,N_39232,N_37146);
nand U43353 (N_43353,N_39584,N_36975);
and U43354 (N_43354,N_36205,N_36117);
nand U43355 (N_43355,N_37858,N_36465);
or U43356 (N_43356,N_37168,N_39572);
and U43357 (N_43357,N_35227,N_37848);
xnor U43358 (N_43358,N_37564,N_39991);
nor U43359 (N_43359,N_39043,N_39794);
nor U43360 (N_43360,N_38520,N_38801);
or U43361 (N_43361,N_36498,N_37094);
xor U43362 (N_43362,N_39770,N_36778);
and U43363 (N_43363,N_36779,N_38548);
or U43364 (N_43364,N_35253,N_35680);
xnor U43365 (N_43365,N_36491,N_36803);
nor U43366 (N_43366,N_36685,N_39322);
and U43367 (N_43367,N_39468,N_35233);
xnor U43368 (N_43368,N_37579,N_35689);
xnor U43369 (N_43369,N_38543,N_37832);
nand U43370 (N_43370,N_37453,N_38831);
nor U43371 (N_43371,N_36433,N_39477);
xnor U43372 (N_43372,N_35382,N_39651);
nor U43373 (N_43373,N_35305,N_36030);
nor U43374 (N_43374,N_36130,N_38193);
and U43375 (N_43375,N_37660,N_39823);
nor U43376 (N_43376,N_35429,N_37868);
and U43377 (N_43377,N_37843,N_38709);
and U43378 (N_43378,N_39701,N_39194);
xor U43379 (N_43379,N_37638,N_37857);
xor U43380 (N_43380,N_39024,N_36009);
or U43381 (N_43381,N_37077,N_37294);
xor U43382 (N_43382,N_36504,N_35625);
and U43383 (N_43383,N_37975,N_38241);
or U43384 (N_43384,N_36457,N_35263);
and U43385 (N_43385,N_38810,N_39566);
nor U43386 (N_43386,N_38425,N_36719);
xnor U43387 (N_43387,N_38108,N_36695);
and U43388 (N_43388,N_35583,N_36708);
xnor U43389 (N_43389,N_36511,N_39585);
nand U43390 (N_43390,N_35321,N_36826);
nand U43391 (N_43391,N_35352,N_38941);
nor U43392 (N_43392,N_35941,N_36207);
nor U43393 (N_43393,N_36618,N_39534);
or U43394 (N_43394,N_39307,N_37295);
xnor U43395 (N_43395,N_39832,N_38850);
nor U43396 (N_43396,N_38017,N_37582);
xor U43397 (N_43397,N_37383,N_35867);
xor U43398 (N_43398,N_38992,N_35138);
nand U43399 (N_43399,N_37632,N_37798);
and U43400 (N_43400,N_35331,N_35202);
or U43401 (N_43401,N_35628,N_38996);
xnor U43402 (N_43402,N_35935,N_36828);
nor U43403 (N_43403,N_39751,N_36499);
and U43404 (N_43404,N_38781,N_36869);
and U43405 (N_43405,N_36793,N_35796);
xor U43406 (N_43406,N_35990,N_39651);
nand U43407 (N_43407,N_35040,N_38460);
and U43408 (N_43408,N_36164,N_39322);
or U43409 (N_43409,N_35046,N_37400);
xor U43410 (N_43410,N_38830,N_37777);
and U43411 (N_43411,N_35516,N_39599);
xor U43412 (N_43412,N_36382,N_35279);
xnor U43413 (N_43413,N_39417,N_39731);
xor U43414 (N_43414,N_37820,N_35111);
nor U43415 (N_43415,N_37082,N_38680);
nand U43416 (N_43416,N_35648,N_35247);
xor U43417 (N_43417,N_37310,N_38187);
and U43418 (N_43418,N_36854,N_36414);
xor U43419 (N_43419,N_38857,N_36477);
nand U43420 (N_43420,N_37688,N_36847);
and U43421 (N_43421,N_38667,N_35742);
xnor U43422 (N_43422,N_38378,N_35924);
nor U43423 (N_43423,N_36204,N_39746);
xor U43424 (N_43424,N_35457,N_36599);
or U43425 (N_43425,N_35352,N_36975);
and U43426 (N_43426,N_39082,N_37293);
nand U43427 (N_43427,N_39406,N_38209);
and U43428 (N_43428,N_38920,N_37513);
nor U43429 (N_43429,N_38465,N_37146);
nor U43430 (N_43430,N_38256,N_38262);
nand U43431 (N_43431,N_36649,N_37864);
and U43432 (N_43432,N_36153,N_35576);
xor U43433 (N_43433,N_35312,N_35254);
or U43434 (N_43434,N_35561,N_39683);
xnor U43435 (N_43435,N_39022,N_36031);
nor U43436 (N_43436,N_37643,N_38519);
nor U43437 (N_43437,N_36960,N_35778);
or U43438 (N_43438,N_39200,N_39081);
or U43439 (N_43439,N_37779,N_37325);
nor U43440 (N_43440,N_36814,N_38482);
or U43441 (N_43441,N_39175,N_39070);
xor U43442 (N_43442,N_37935,N_37299);
or U43443 (N_43443,N_36181,N_39972);
and U43444 (N_43444,N_39683,N_38237);
nor U43445 (N_43445,N_36613,N_35318);
nor U43446 (N_43446,N_37963,N_38499);
and U43447 (N_43447,N_38069,N_36301);
nor U43448 (N_43448,N_36529,N_35964);
nor U43449 (N_43449,N_35992,N_37719);
nor U43450 (N_43450,N_38410,N_36712);
and U43451 (N_43451,N_35353,N_36052);
xnor U43452 (N_43452,N_38945,N_39532);
xnor U43453 (N_43453,N_39984,N_39683);
and U43454 (N_43454,N_35025,N_35703);
nor U43455 (N_43455,N_37208,N_36763);
nor U43456 (N_43456,N_37712,N_35071);
nor U43457 (N_43457,N_36583,N_38386);
nor U43458 (N_43458,N_35730,N_35384);
and U43459 (N_43459,N_39942,N_35914);
nor U43460 (N_43460,N_39246,N_39396);
or U43461 (N_43461,N_37451,N_35282);
xor U43462 (N_43462,N_35709,N_38757);
and U43463 (N_43463,N_36955,N_36024);
nand U43464 (N_43464,N_39150,N_35666);
nand U43465 (N_43465,N_36509,N_39148);
or U43466 (N_43466,N_36423,N_36072);
xor U43467 (N_43467,N_36692,N_38686);
nor U43468 (N_43468,N_35484,N_39954);
or U43469 (N_43469,N_36820,N_39937);
nand U43470 (N_43470,N_38835,N_35504);
nor U43471 (N_43471,N_37109,N_37962);
or U43472 (N_43472,N_38064,N_36544);
nand U43473 (N_43473,N_35601,N_39924);
nor U43474 (N_43474,N_38275,N_37461);
nor U43475 (N_43475,N_39789,N_39096);
or U43476 (N_43476,N_37829,N_39772);
or U43477 (N_43477,N_39272,N_35138);
nor U43478 (N_43478,N_39596,N_39557);
nor U43479 (N_43479,N_35751,N_38544);
nand U43480 (N_43480,N_36558,N_38863);
or U43481 (N_43481,N_37556,N_39303);
and U43482 (N_43482,N_36004,N_37996);
xnor U43483 (N_43483,N_38536,N_36054);
nand U43484 (N_43484,N_37176,N_37161);
nor U43485 (N_43485,N_37897,N_38928);
nor U43486 (N_43486,N_37103,N_39839);
nand U43487 (N_43487,N_38037,N_39761);
and U43488 (N_43488,N_38742,N_37335);
xnor U43489 (N_43489,N_38023,N_36446);
and U43490 (N_43490,N_39774,N_37689);
or U43491 (N_43491,N_39719,N_35906);
xor U43492 (N_43492,N_38538,N_36523);
nor U43493 (N_43493,N_37006,N_35520);
xnor U43494 (N_43494,N_38181,N_38169);
xnor U43495 (N_43495,N_36422,N_38030);
xor U43496 (N_43496,N_39263,N_37293);
xnor U43497 (N_43497,N_35614,N_36262);
xor U43498 (N_43498,N_38358,N_39437);
nor U43499 (N_43499,N_39899,N_37017);
nor U43500 (N_43500,N_37284,N_38964);
or U43501 (N_43501,N_38235,N_38228);
and U43502 (N_43502,N_37774,N_38874);
nor U43503 (N_43503,N_39575,N_35465);
nand U43504 (N_43504,N_38008,N_37728);
nor U43505 (N_43505,N_37318,N_39240);
xor U43506 (N_43506,N_37512,N_39389);
nand U43507 (N_43507,N_39594,N_38034);
nor U43508 (N_43508,N_36053,N_35204);
nor U43509 (N_43509,N_39247,N_36395);
nand U43510 (N_43510,N_36790,N_37907);
nor U43511 (N_43511,N_38798,N_39982);
xnor U43512 (N_43512,N_36884,N_38709);
nor U43513 (N_43513,N_37081,N_36326);
and U43514 (N_43514,N_38182,N_35108);
or U43515 (N_43515,N_38586,N_36267);
or U43516 (N_43516,N_38403,N_35553);
and U43517 (N_43517,N_37068,N_39122);
nand U43518 (N_43518,N_37804,N_37457);
nor U43519 (N_43519,N_37954,N_37666);
or U43520 (N_43520,N_36701,N_39609);
xnor U43521 (N_43521,N_35208,N_38003);
nand U43522 (N_43522,N_36449,N_39242);
nor U43523 (N_43523,N_36821,N_39284);
nor U43524 (N_43524,N_39913,N_38233);
or U43525 (N_43525,N_38163,N_36857);
nor U43526 (N_43526,N_39547,N_38043);
nand U43527 (N_43527,N_38383,N_38204);
nor U43528 (N_43528,N_38554,N_35733);
or U43529 (N_43529,N_35106,N_35841);
nand U43530 (N_43530,N_37997,N_39294);
and U43531 (N_43531,N_36344,N_37837);
and U43532 (N_43532,N_37784,N_37739);
or U43533 (N_43533,N_35185,N_39490);
or U43534 (N_43534,N_39773,N_39849);
and U43535 (N_43535,N_38921,N_37179);
xor U43536 (N_43536,N_35621,N_39543);
and U43537 (N_43537,N_39266,N_37802);
nand U43538 (N_43538,N_37954,N_35744);
nand U43539 (N_43539,N_36983,N_35794);
nor U43540 (N_43540,N_35471,N_35315);
nor U43541 (N_43541,N_36770,N_36487);
or U43542 (N_43542,N_38076,N_36600);
xnor U43543 (N_43543,N_37262,N_37926);
and U43544 (N_43544,N_38755,N_37944);
nor U43545 (N_43545,N_38679,N_37470);
xor U43546 (N_43546,N_37244,N_36201);
xor U43547 (N_43547,N_38628,N_36604);
or U43548 (N_43548,N_38580,N_39179);
or U43549 (N_43549,N_36917,N_36512);
nor U43550 (N_43550,N_37209,N_39373);
nand U43551 (N_43551,N_38665,N_37550);
xor U43552 (N_43552,N_36022,N_38842);
or U43553 (N_43553,N_38942,N_35021);
or U43554 (N_43554,N_36628,N_35063);
and U43555 (N_43555,N_35697,N_35182);
xor U43556 (N_43556,N_36908,N_37179);
xnor U43557 (N_43557,N_37459,N_36207);
nand U43558 (N_43558,N_39529,N_37940);
or U43559 (N_43559,N_35472,N_39283);
xor U43560 (N_43560,N_39092,N_36071);
xor U43561 (N_43561,N_36761,N_38218);
or U43562 (N_43562,N_35475,N_38714);
xor U43563 (N_43563,N_35792,N_39682);
nor U43564 (N_43564,N_38266,N_37929);
nor U43565 (N_43565,N_35246,N_35763);
nand U43566 (N_43566,N_38939,N_39173);
and U43567 (N_43567,N_36242,N_36028);
nor U43568 (N_43568,N_39549,N_38707);
nor U43569 (N_43569,N_39692,N_36070);
xnor U43570 (N_43570,N_39612,N_35735);
nor U43571 (N_43571,N_37741,N_39096);
xor U43572 (N_43572,N_38196,N_37097);
or U43573 (N_43573,N_37312,N_36941);
xor U43574 (N_43574,N_36021,N_36773);
and U43575 (N_43575,N_39171,N_36310);
and U43576 (N_43576,N_36174,N_39071);
nand U43577 (N_43577,N_37744,N_35736);
nand U43578 (N_43578,N_35661,N_38025);
xor U43579 (N_43579,N_39317,N_38008);
and U43580 (N_43580,N_35017,N_36908);
or U43581 (N_43581,N_36325,N_38519);
or U43582 (N_43582,N_37227,N_39408);
or U43583 (N_43583,N_39350,N_36579);
xor U43584 (N_43584,N_37089,N_36444);
or U43585 (N_43585,N_39052,N_37202);
or U43586 (N_43586,N_37803,N_37917);
nand U43587 (N_43587,N_39421,N_39170);
or U43588 (N_43588,N_36383,N_38574);
and U43589 (N_43589,N_39809,N_35981);
or U43590 (N_43590,N_36301,N_37571);
nor U43591 (N_43591,N_36491,N_35985);
or U43592 (N_43592,N_39377,N_38441);
nand U43593 (N_43593,N_35915,N_38989);
or U43594 (N_43594,N_39815,N_35414);
nand U43595 (N_43595,N_38625,N_39533);
nor U43596 (N_43596,N_35951,N_39997);
nand U43597 (N_43597,N_36209,N_39499);
xnor U43598 (N_43598,N_38243,N_37511);
nor U43599 (N_43599,N_35544,N_39370);
or U43600 (N_43600,N_35419,N_38784);
or U43601 (N_43601,N_37380,N_35161);
or U43602 (N_43602,N_38474,N_37230);
and U43603 (N_43603,N_36604,N_38924);
or U43604 (N_43604,N_37285,N_36152);
or U43605 (N_43605,N_38545,N_39087);
xnor U43606 (N_43606,N_37549,N_37292);
or U43607 (N_43607,N_37812,N_35114);
nor U43608 (N_43608,N_36492,N_38470);
nand U43609 (N_43609,N_37364,N_38433);
xor U43610 (N_43610,N_39724,N_37363);
nor U43611 (N_43611,N_36750,N_38802);
and U43612 (N_43612,N_39332,N_35202);
nand U43613 (N_43613,N_37200,N_38527);
xor U43614 (N_43614,N_37148,N_38167);
and U43615 (N_43615,N_37599,N_39507);
or U43616 (N_43616,N_36759,N_37522);
or U43617 (N_43617,N_37960,N_37974);
or U43618 (N_43618,N_37675,N_39366);
nor U43619 (N_43619,N_36711,N_35315);
xnor U43620 (N_43620,N_37838,N_37365);
nand U43621 (N_43621,N_37842,N_39146);
nor U43622 (N_43622,N_38689,N_38340);
nor U43623 (N_43623,N_37441,N_37606);
or U43624 (N_43624,N_36838,N_38188);
or U43625 (N_43625,N_37782,N_35790);
xor U43626 (N_43626,N_39150,N_38287);
xor U43627 (N_43627,N_37034,N_36068);
nand U43628 (N_43628,N_38814,N_37174);
and U43629 (N_43629,N_36961,N_36443);
xor U43630 (N_43630,N_38254,N_38814);
and U43631 (N_43631,N_37134,N_39825);
xor U43632 (N_43632,N_38469,N_38081);
and U43633 (N_43633,N_35936,N_38480);
nor U43634 (N_43634,N_36637,N_39377);
or U43635 (N_43635,N_39110,N_35013);
and U43636 (N_43636,N_39897,N_36875);
nor U43637 (N_43637,N_37240,N_39483);
nor U43638 (N_43638,N_36967,N_39116);
or U43639 (N_43639,N_38919,N_37454);
nor U43640 (N_43640,N_36895,N_35649);
nor U43641 (N_43641,N_37486,N_36797);
and U43642 (N_43642,N_38271,N_39081);
nor U43643 (N_43643,N_36062,N_37794);
xor U43644 (N_43644,N_38949,N_35327);
nand U43645 (N_43645,N_38570,N_36752);
nand U43646 (N_43646,N_35570,N_37183);
or U43647 (N_43647,N_37711,N_38994);
and U43648 (N_43648,N_36815,N_35845);
or U43649 (N_43649,N_38183,N_35710);
and U43650 (N_43650,N_37905,N_39434);
nor U43651 (N_43651,N_39552,N_39348);
xnor U43652 (N_43652,N_39348,N_39814);
xor U43653 (N_43653,N_39650,N_39264);
or U43654 (N_43654,N_39191,N_35361);
or U43655 (N_43655,N_35300,N_35076);
and U43656 (N_43656,N_35436,N_39478);
or U43657 (N_43657,N_39058,N_36849);
nor U43658 (N_43658,N_37253,N_36441);
nor U43659 (N_43659,N_36827,N_36272);
nor U43660 (N_43660,N_39142,N_37800);
xor U43661 (N_43661,N_39001,N_36110);
or U43662 (N_43662,N_36403,N_39314);
nor U43663 (N_43663,N_36882,N_38953);
and U43664 (N_43664,N_36531,N_39669);
and U43665 (N_43665,N_37260,N_35820);
and U43666 (N_43666,N_37743,N_39201);
and U43667 (N_43667,N_38632,N_37795);
and U43668 (N_43668,N_35874,N_35001);
xor U43669 (N_43669,N_36702,N_37209);
and U43670 (N_43670,N_36632,N_37350);
and U43671 (N_43671,N_36034,N_39889);
or U43672 (N_43672,N_38854,N_39194);
xnor U43673 (N_43673,N_35015,N_37683);
nor U43674 (N_43674,N_39293,N_35941);
or U43675 (N_43675,N_39520,N_37997);
xor U43676 (N_43676,N_35206,N_35470);
nor U43677 (N_43677,N_38065,N_38404);
xor U43678 (N_43678,N_36012,N_36069);
nand U43679 (N_43679,N_37229,N_38507);
xor U43680 (N_43680,N_38535,N_38771);
nand U43681 (N_43681,N_38944,N_36706);
or U43682 (N_43682,N_37252,N_35516);
or U43683 (N_43683,N_35517,N_37589);
and U43684 (N_43684,N_37356,N_39806);
and U43685 (N_43685,N_35580,N_37663);
xnor U43686 (N_43686,N_38971,N_37871);
and U43687 (N_43687,N_37677,N_38809);
or U43688 (N_43688,N_39580,N_36540);
nand U43689 (N_43689,N_37503,N_38796);
and U43690 (N_43690,N_37478,N_38122);
nor U43691 (N_43691,N_38125,N_38100);
and U43692 (N_43692,N_37452,N_36753);
nand U43693 (N_43693,N_39399,N_36470);
xor U43694 (N_43694,N_35100,N_39949);
nor U43695 (N_43695,N_37725,N_39544);
xor U43696 (N_43696,N_36818,N_36889);
xnor U43697 (N_43697,N_37346,N_37457);
nand U43698 (N_43698,N_36456,N_35680);
xnor U43699 (N_43699,N_38828,N_35056);
nand U43700 (N_43700,N_39452,N_39488);
or U43701 (N_43701,N_38375,N_36211);
and U43702 (N_43702,N_39669,N_36845);
nand U43703 (N_43703,N_36592,N_37583);
or U43704 (N_43704,N_36596,N_39342);
xor U43705 (N_43705,N_37179,N_37096);
nand U43706 (N_43706,N_37291,N_37175);
nor U43707 (N_43707,N_36140,N_39113);
and U43708 (N_43708,N_35317,N_38688);
nor U43709 (N_43709,N_38008,N_37447);
xor U43710 (N_43710,N_38814,N_37145);
or U43711 (N_43711,N_35686,N_39131);
and U43712 (N_43712,N_35911,N_39156);
or U43713 (N_43713,N_35293,N_37735);
xor U43714 (N_43714,N_35228,N_38500);
xor U43715 (N_43715,N_37768,N_36702);
and U43716 (N_43716,N_35621,N_38525);
xor U43717 (N_43717,N_39891,N_35980);
and U43718 (N_43718,N_38514,N_36548);
nor U43719 (N_43719,N_35311,N_35534);
xor U43720 (N_43720,N_37084,N_39913);
nor U43721 (N_43721,N_37761,N_37793);
nor U43722 (N_43722,N_39083,N_35064);
xnor U43723 (N_43723,N_38769,N_37449);
nor U43724 (N_43724,N_38047,N_35635);
and U43725 (N_43725,N_38315,N_36278);
or U43726 (N_43726,N_38935,N_36075);
nor U43727 (N_43727,N_37628,N_36619);
or U43728 (N_43728,N_35498,N_38674);
and U43729 (N_43729,N_38462,N_36919);
xnor U43730 (N_43730,N_35318,N_36162);
xnor U43731 (N_43731,N_36718,N_39964);
or U43732 (N_43732,N_39998,N_36540);
or U43733 (N_43733,N_35436,N_39684);
and U43734 (N_43734,N_38553,N_38695);
or U43735 (N_43735,N_37777,N_36743);
nand U43736 (N_43736,N_39826,N_39138);
nand U43737 (N_43737,N_39043,N_39574);
nor U43738 (N_43738,N_37643,N_35691);
or U43739 (N_43739,N_35660,N_35307);
or U43740 (N_43740,N_35490,N_37159);
xnor U43741 (N_43741,N_39052,N_37165);
nor U43742 (N_43742,N_38831,N_38128);
nand U43743 (N_43743,N_37178,N_35145);
xor U43744 (N_43744,N_38194,N_39522);
nand U43745 (N_43745,N_39302,N_36429);
nor U43746 (N_43746,N_35211,N_36033);
nand U43747 (N_43747,N_37252,N_37558);
and U43748 (N_43748,N_37715,N_35315);
xor U43749 (N_43749,N_35173,N_36957);
xor U43750 (N_43750,N_36762,N_35547);
nor U43751 (N_43751,N_36054,N_37719);
or U43752 (N_43752,N_36792,N_39145);
xnor U43753 (N_43753,N_35099,N_35676);
xor U43754 (N_43754,N_37430,N_37536);
and U43755 (N_43755,N_36075,N_37764);
nand U43756 (N_43756,N_36995,N_36100);
and U43757 (N_43757,N_36502,N_36643);
nand U43758 (N_43758,N_39130,N_38766);
and U43759 (N_43759,N_38343,N_39114);
nor U43760 (N_43760,N_36437,N_36642);
nor U43761 (N_43761,N_37316,N_36474);
nor U43762 (N_43762,N_38466,N_35285);
xor U43763 (N_43763,N_39794,N_38675);
xnor U43764 (N_43764,N_35909,N_36187);
xnor U43765 (N_43765,N_39828,N_35522);
nand U43766 (N_43766,N_39998,N_38332);
and U43767 (N_43767,N_37387,N_38487);
or U43768 (N_43768,N_38874,N_37559);
nor U43769 (N_43769,N_37183,N_36555);
and U43770 (N_43770,N_38599,N_37588);
xor U43771 (N_43771,N_38263,N_39923);
nor U43772 (N_43772,N_35992,N_39486);
xor U43773 (N_43773,N_35127,N_36473);
xor U43774 (N_43774,N_35845,N_38495);
or U43775 (N_43775,N_36415,N_36584);
nor U43776 (N_43776,N_37590,N_36935);
xnor U43777 (N_43777,N_37779,N_37907);
xnor U43778 (N_43778,N_38956,N_35088);
nor U43779 (N_43779,N_38702,N_37551);
nor U43780 (N_43780,N_37672,N_35878);
or U43781 (N_43781,N_39349,N_39896);
xnor U43782 (N_43782,N_35926,N_37487);
nand U43783 (N_43783,N_39040,N_38357);
and U43784 (N_43784,N_37815,N_39689);
and U43785 (N_43785,N_39811,N_38648);
nand U43786 (N_43786,N_36245,N_36376);
nand U43787 (N_43787,N_35391,N_36087);
xnor U43788 (N_43788,N_37743,N_39491);
nand U43789 (N_43789,N_38833,N_39086);
xor U43790 (N_43790,N_37105,N_38539);
xor U43791 (N_43791,N_37410,N_38517);
nor U43792 (N_43792,N_36368,N_36110);
and U43793 (N_43793,N_36116,N_39118);
and U43794 (N_43794,N_37776,N_39696);
nand U43795 (N_43795,N_39942,N_38177);
nand U43796 (N_43796,N_37284,N_37267);
nor U43797 (N_43797,N_35741,N_37103);
and U43798 (N_43798,N_37977,N_38193);
nor U43799 (N_43799,N_35390,N_38123);
nor U43800 (N_43800,N_36300,N_38545);
nor U43801 (N_43801,N_39061,N_39197);
nor U43802 (N_43802,N_37945,N_36685);
and U43803 (N_43803,N_39877,N_37069);
or U43804 (N_43804,N_38686,N_37315);
nor U43805 (N_43805,N_35637,N_38148);
nand U43806 (N_43806,N_36488,N_39761);
nor U43807 (N_43807,N_39491,N_36214);
xnor U43808 (N_43808,N_37707,N_38015);
xnor U43809 (N_43809,N_36546,N_38995);
or U43810 (N_43810,N_37756,N_37443);
and U43811 (N_43811,N_35642,N_39646);
or U43812 (N_43812,N_36969,N_37083);
nor U43813 (N_43813,N_37077,N_35571);
nand U43814 (N_43814,N_35016,N_36533);
nand U43815 (N_43815,N_37857,N_35039);
or U43816 (N_43816,N_37554,N_38139);
or U43817 (N_43817,N_36251,N_38241);
nand U43818 (N_43818,N_36359,N_38563);
and U43819 (N_43819,N_38678,N_35000);
xor U43820 (N_43820,N_36558,N_39963);
xor U43821 (N_43821,N_35966,N_35376);
and U43822 (N_43822,N_39018,N_35169);
nand U43823 (N_43823,N_35297,N_38423);
or U43824 (N_43824,N_35360,N_35266);
nand U43825 (N_43825,N_39672,N_35010);
nor U43826 (N_43826,N_39530,N_36897);
nor U43827 (N_43827,N_39940,N_36157);
nor U43828 (N_43828,N_39750,N_37951);
xor U43829 (N_43829,N_39436,N_35924);
nand U43830 (N_43830,N_36757,N_36767);
nor U43831 (N_43831,N_35000,N_37094);
nand U43832 (N_43832,N_38818,N_36513);
and U43833 (N_43833,N_39797,N_37402);
xnor U43834 (N_43834,N_36912,N_38101);
xor U43835 (N_43835,N_36891,N_37583);
and U43836 (N_43836,N_39015,N_37332);
or U43837 (N_43837,N_37883,N_39116);
nand U43838 (N_43838,N_35258,N_39571);
xor U43839 (N_43839,N_35814,N_36596);
or U43840 (N_43840,N_39584,N_36189);
xnor U43841 (N_43841,N_39962,N_38568);
nor U43842 (N_43842,N_37161,N_36562);
or U43843 (N_43843,N_39812,N_35694);
and U43844 (N_43844,N_38207,N_37221);
or U43845 (N_43845,N_37462,N_39660);
nor U43846 (N_43846,N_35607,N_35704);
nand U43847 (N_43847,N_36860,N_35355);
nand U43848 (N_43848,N_36533,N_36549);
and U43849 (N_43849,N_39721,N_39400);
and U43850 (N_43850,N_39283,N_36912);
xnor U43851 (N_43851,N_35203,N_38311);
xnor U43852 (N_43852,N_38238,N_38050);
nor U43853 (N_43853,N_38890,N_37951);
nand U43854 (N_43854,N_38930,N_37696);
nand U43855 (N_43855,N_37468,N_35910);
nand U43856 (N_43856,N_39432,N_35339);
or U43857 (N_43857,N_35379,N_36354);
xor U43858 (N_43858,N_35769,N_38429);
xnor U43859 (N_43859,N_37701,N_38914);
nand U43860 (N_43860,N_38155,N_37126);
and U43861 (N_43861,N_39224,N_39182);
xor U43862 (N_43862,N_37547,N_35539);
nor U43863 (N_43863,N_37412,N_36625);
and U43864 (N_43864,N_39546,N_37400);
nor U43865 (N_43865,N_38817,N_39854);
nor U43866 (N_43866,N_35024,N_39679);
or U43867 (N_43867,N_39342,N_37504);
xnor U43868 (N_43868,N_38306,N_38652);
xnor U43869 (N_43869,N_38484,N_36061);
nand U43870 (N_43870,N_38582,N_35885);
nor U43871 (N_43871,N_37947,N_39963);
and U43872 (N_43872,N_36148,N_39837);
and U43873 (N_43873,N_37289,N_38685);
and U43874 (N_43874,N_35718,N_39067);
or U43875 (N_43875,N_37630,N_39020);
nand U43876 (N_43876,N_39831,N_37238);
or U43877 (N_43877,N_36383,N_39212);
and U43878 (N_43878,N_36029,N_36185);
xor U43879 (N_43879,N_39985,N_39377);
nor U43880 (N_43880,N_36309,N_35111);
nand U43881 (N_43881,N_36884,N_36259);
nor U43882 (N_43882,N_37901,N_39525);
nor U43883 (N_43883,N_36613,N_39137);
or U43884 (N_43884,N_39575,N_37554);
or U43885 (N_43885,N_38857,N_35504);
nor U43886 (N_43886,N_36465,N_37512);
xnor U43887 (N_43887,N_36917,N_39335);
xnor U43888 (N_43888,N_38517,N_36050);
nor U43889 (N_43889,N_36941,N_37368);
nand U43890 (N_43890,N_39472,N_35705);
and U43891 (N_43891,N_36906,N_39961);
and U43892 (N_43892,N_35637,N_39483);
and U43893 (N_43893,N_38093,N_39920);
xnor U43894 (N_43894,N_37596,N_36640);
and U43895 (N_43895,N_36470,N_36407);
nor U43896 (N_43896,N_37198,N_36155);
and U43897 (N_43897,N_36213,N_37920);
xor U43898 (N_43898,N_35547,N_39281);
and U43899 (N_43899,N_39146,N_35169);
xnor U43900 (N_43900,N_38971,N_38839);
xnor U43901 (N_43901,N_36209,N_37222);
or U43902 (N_43902,N_35794,N_35979);
and U43903 (N_43903,N_35984,N_39392);
xor U43904 (N_43904,N_36146,N_39670);
nor U43905 (N_43905,N_38071,N_37646);
or U43906 (N_43906,N_35339,N_37492);
or U43907 (N_43907,N_35489,N_36897);
or U43908 (N_43908,N_36513,N_39143);
and U43909 (N_43909,N_39622,N_37182);
nor U43910 (N_43910,N_37275,N_38835);
or U43911 (N_43911,N_39261,N_39216);
nor U43912 (N_43912,N_36103,N_37487);
and U43913 (N_43913,N_39842,N_36394);
xor U43914 (N_43914,N_39786,N_36069);
or U43915 (N_43915,N_39571,N_39162);
xnor U43916 (N_43916,N_38997,N_37481);
xor U43917 (N_43917,N_38024,N_37134);
xor U43918 (N_43918,N_38032,N_35049);
xor U43919 (N_43919,N_39381,N_35730);
or U43920 (N_43920,N_37269,N_36348);
or U43921 (N_43921,N_37838,N_37240);
or U43922 (N_43922,N_35602,N_37271);
or U43923 (N_43923,N_36802,N_38262);
or U43924 (N_43924,N_35299,N_35852);
or U43925 (N_43925,N_37079,N_37362);
nor U43926 (N_43926,N_36175,N_35590);
xnor U43927 (N_43927,N_38359,N_38841);
nor U43928 (N_43928,N_38662,N_36624);
and U43929 (N_43929,N_37288,N_37205);
or U43930 (N_43930,N_37095,N_38245);
xor U43931 (N_43931,N_38903,N_38592);
xor U43932 (N_43932,N_37989,N_39804);
xnor U43933 (N_43933,N_39964,N_36424);
nand U43934 (N_43934,N_39834,N_38954);
xor U43935 (N_43935,N_36003,N_39269);
nand U43936 (N_43936,N_36847,N_35194);
nand U43937 (N_43937,N_36525,N_35941);
nand U43938 (N_43938,N_36077,N_36114);
xnor U43939 (N_43939,N_37155,N_35169);
nand U43940 (N_43940,N_35276,N_39844);
and U43941 (N_43941,N_37946,N_37385);
nand U43942 (N_43942,N_39953,N_37841);
nor U43943 (N_43943,N_36322,N_38493);
xor U43944 (N_43944,N_35706,N_38027);
xnor U43945 (N_43945,N_39565,N_36704);
nor U43946 (N_43946,N_36765,N_38528);
or U43947 (N_43947,N_37002,N_35601);
xnor U43948 (N_43948,N_35819,N_38974);
xnor U43949 (N_43949,N_38566,N_35443);
xor U43950 (N_43950,N_39366,N_35714);
xor U43951 (N_43951,N_38210,N_35734);
nand U43952 (N_43952,N_39012,N_36482);
or U43953 (N_43953,N_35858,N_37861);
nor U43954 (N_43954,N_39784,N_38641);
xor U43955 (N_43955,N_37873,N_35777);
nand U43956 (N_43956,N_39918,N_35441);
and U43957 (N_43957,N_37214,N_36606);
nor U43958 (N_43958,N_35610,N_39118);
xor U43959 (N_43959,N_36655,N_37901);
and U43960 (N_43960,N_37242,N_39411);
nor U43961 (N_43961,N_39855,N_35795);
xnor U43962 (N_43962,N_38626,N_38084);
nor U43963 (N_43963,N_39406,N_35714);
nand U43964 (N_43964,N_35705,N_36764);
or U43965 (N_43965,N_35224,N_36072);
and U43966 (N_43966,N_37906,N_38679);
and U43967 (N_43967,N_39071,N_39206);
xnor U43968 (N_43968,N_36466,N_36882);
nor U43969 (N_43969,N_37837,N_37516);
and U43970 (N_43970,N_39077,N_35396);
xor U43971 (N_43971,N_35603,N_36912);
or U43972 (N_43972,N_39328,N_39376);
or U43973 (N_43973,N_38179,N_36742);
xor U43974 (N_43974,N_35578,N_38814);
or U43975 (N_43975,N_39879,N_37731);
and U43976 (N_43976,N_35460,N_37207);
nand U43977 (N_43977,N_37536,N_36715);
xnor U43978 (N_43978,N_36194,N_35059);
nor U43979 (N_43979,N_36593,N_37070);
or U43980 (N_43980,N_37057,N_36750);
and U43981 (N_43981,N_37591,N_35254);
xor U43982 (N_43982,N_38508,N_35857);
xor U43983 (N_43983,N_37952,N_35880);
or U43984 (N_43984,N_38734,N_38255);
nand U43985 (N_43985,N_38566,N_38904);
and U43986 (N_43986,N_39317,N_36931);
xor U43987 (N_43987,N_35930,N_36471);
nand U43988 (N_43988,N_35334,N_38402);
or U43989 (N_43989,N_37822,N_36475);
xor U43990 (N_43990,N_36754,N_39350);
and U43991 (N_43991,N_35994,N_38981);
nor U43992 (N_43992,N_39764,N_39740);
nor U43993 (N_43993,N_38860,N_35404);
or U43994 (N_43994,N_38502,N_39175);
and U43995 (N_43995,N_35653,N_39848);
nor U43996 (N_43996,N_37157,N_35388);
nor U43997 (N_43997,N_38815,N_38372);
nand U43998 (N_43998,N_39581,N_35067);
and U43999 (N_43999,N_35243,N_38956);
or U44000 (N_44000,N_39382,N_36187);
and U44001 (N_44001,N_36998,N_39173);
nand U44002 (N_44002,N_37187,N_38713);
xor U44003 (N_44003,N_39294,N_37071);
and U44004 (N_44004,N_39483,N_37770);
or U44005 (N_44005,N_35114,N_36472);
nor U44006 (N_44006,N_36976,N_38866);
and U44007 (N_44007,N_37450,N_35850);
nor U44008 (N_44008,N_36147,N_35959);
nand U44009 (N_44009,N_36010,N_37169);
nand U44010 (N_44010,N_37103,N_39647);
xnor U44011 (N_44011,N_38147,N_36237);
xnor U44012 (N_44012,N_37352,N_35613);
nor U44013 (N_44013,N_39686,N_38198);
and U44014 (N_44014,N_35135,N_38841);
and U44015 (N_44015,N_35425,N_37041);
xnor U44016 (N_44016,N_36657,N_36373);
or U44017 (N_44017,N_35244,N_37400);
nand U44018 (N_44018,N_35557,N_36781);
and U44019 (N_44019,N_39055,N_39136);
nand U44020 (N_44020,N_38854,N_38371);
nor U44021 (N_44021,N_35140,N_36689);
nand U44022 (N_44022,N_37144,N_38843);
and U44023 (N_44023,N_39618,N_39306);
nor U44024 (N_44024,N_35276,N_37184);
or U44025 (N_44025,N_35098,N_36518);
and U44026 (N_44026,N_36270,N_35533);
xor U44027 (N_44027,N_35307,N_35901);
xor U44028 (N_44028,N_38042,N_36288);
nor U44029 (N_44029,N_35632,N_39451);
or U44030 (N_44030,N_35668,N_38615);
nand U44031 (N_44031,N_36625,N_39903);
and U44032 (N_44032,N_39939,N_37381);
nor U44033 (N_44033,N_35766,N_37343);
nor U44034 (N_44034,N_37293,N_35062);
nand U44035 (N_44035,N_36019,N_36989);
and U44036 (N_44036,N_39052,N_37334);
or U44037 (N_44037,N_35258,N_37508);
or U44038 (N_44038,N_38577,N_37310);
nor U44039 (N_44039,N_36089,N_38221);
and U44040 (N_44040,N_38715,N_38790);
xor U44041 (N_44041,N_36842,N_39685);
and U44042 (N_44042,N_36102,N_37258);
nand U44043 (N_44043,N_38808,N_35081);
nand U44044 (N_44044,N_35029,N_38451);
and U44045 (N_44045,N_38859,N_38377);
nor U44046 (N_44046,N_39018,N_39194);
or U44047 (N_44047,N_35752,N_38446);
or U44048 (N_44048,N_36651,N_39804);
and U44049 (N_44049,N_39735,N_39144);
and U44050 (N_44050,N_36406,N_38596);
and U44051 (N_44051,N_38893,N_37741);
or U44052 (N_44052,N_35994,N_38946);
or U44053 (N_44053,N_39845,N_39459);
nand U44054 (N_44054,N_35063,N_38646);
nand U44055 (N_44055,N_35628,N_36856);
nor U44056 (N_44056,N_37723,N_37988);
nor U44057 (N_44057,N_36531,N_39591);
nor U44058 (N_44058,N_38016,N_39898);
nor U44059 (N_44059,N_36764,N_35210);
and U44060 (N_44060,N_39432,N_35202);
and U44061 (N_44061,N_37012,N_35825);
nand U44062 (N_44062,N_38472,N_38714);
and U44063 (N_44063,N_37106,N_38569);
xor U44064 (N_44064,N_39651,N_37516);
xnor U44065 (N_44065,N_38971,N_39263);
nand U44066 (N_44066,N_35488,N_39722);
nand U44067 (N_44067,N_37793,N_38341);
and U44068 (N_44068,N_35764,N_39939);
nor U44069 (N_44069,N_36220,N_38307);
xnor U44070 (N_44070,N_38227,N_37263);
nand U44071 (N_44071,N_38430,N_37263);
xor U44072 (N_44072,N_35625,N_36120);
nand U44073 (N_44073,N_35915,N_37393);
or U44074 (N_44074,N_38886,N_36225);
nand U44075 (N_44075,N_36232,N_36540);
or U44076 (N_44076,N_37533,N_35555);
nand U44077 (N_44077,N_37365,N_36260);
nand U44078 (N_44078,N_36955,N_38757);
nand U44079 (N_44079,N_39469,N_38755);
nand U44080 (N_44080,N_38343,N_35749);
and U44081 (N_44081,N_36336,N_35140);
xnor U44082 (N_44082,N_38541,N_36904);
and U44083 (N_44083,N_38944,N_39580);
or U44084 (N_44084,N_37542,N_39036);
nand U44085 (N_44085,N_36514,N_38032);
nor U44086 (N_44086,N_37799,N_39092);
or U44087 (N_44087,N_37548,N_35062);
xor U44088 (N_44088,N_36590,N_36244);
nor U44089 (N_44089,N_39623,N_39868);
and U44090 (N_44090,N_39795,N_35490);
nand U44091 (N_44091,N_36923,N_36487);
nor U44092 (N_44092,N_37107,N_36317);
xor U44093 (N_44093,N_36565,N_37348);
xor U44094 (N_44094,N_38350,N_35938);
nand U44095 (N_44095,N_39768,N_38877);
nand U44096 (N_44096,N_39174,N_37183);
or U44097 (N_44097,N_35588,N_35600);
nand U44098 (N_44098,N_38264,N_39704);
nor U44099 (N_44099,N_36637,N_36102);
or U44100 (N_44100,N_35496,N_35924);
nor U44101 (N_44101,N_37883,N_35423);
nand U44102 (N_44102,N_39528,N_37249);
and U44103 (N_44103,N_38400,N_37209);
xor U44104 (N_44104,N_35387,N_35629);
xor U44105 (N_44105,N_37396,N_35934);
and U44106 (N_44106,N_39116,N_38987);
or U44107 (N_44107,N_35041,N_35422);
or U44108 (N_44108,N_39716,N_37104);
or U44109 (N_44109,N_38871,N_38114);
nand U44110 (N_44110,N_36167,N_39450);
nand U44111 (N_44111,N_37523,N_38777);
and U44112 (N_44112,N_38724,N_39276);
nand U44113 (N_44113,N_38663,N_37143);
and U44114 (N_44114,N_36367,N_39509);
and U44115 (N_44115,N_36423,N_39166);
or U44116 (N_44116,N_35765,N_39232);
nor U44117 (N_44117,N_39671,N_37289);
and U44118 (N_44118,N_39876,N_38518);
and U44119 (N_44119,N_38634,N_37550);
nand U44120 (N_44120,N_35378,N_37184);
nand U44121 (N_44121,N_39343,N_35132);
and U44122 (N_44122,N_38463,N_38060);
nor U44123 (N_44123,N_36945,N_36576);
nor U44124 (N_44124,N_37919,N_36344);
nand U44125 (N_44125,N_39715,N_38805);
nor U44126 (N_44126,N_36059,N_38983);
or U44127 (N_44127,N_35736,N_37619);
nand U44128 (N_44128,N_38957,N_35042);
nand U44129 (N_44129,N_38595,N_38660);
or U44130 (N_44130,N_36574,N_38377);
nor U44131 (N_44131,N_37552,N_35948);
xor U44132 (N_44132,N_36802,N_37382);
xnor U44133 (N_44133,N_36367,N_35034);
or U44134 (N_44134,N_39062,N_35358);
nand U44135 (N_44135,N_35471,N_39438);
or U44136 (N_44136,N_36320,N_35252);
nand U44137 (N_44137,N_36517,N_38882);
xor U44138 (N_44138,N_38687,N_36879);
nor U44139 (N_44139,N_39915,N_37658);
and U44140 (N_44140,N_37001,N_38914);
nor U44141 (N_44141,N_38552,N_39523);
and U44142 (N_44142,N_35695,N_39963);
or U44143 (N_44143,N_38781,N_37545);
nand U44144 (N_44144,N_36413,N_39040);
nor U44145 (N_44145,N_35678,N_39616);
and U44146 (N_44146,N_35290,N_37916);
nand U44147 (N_44147,N_35884,N_35516);
xor U44148 (N_44148,N_35152,N_37409);
xnor U44149 (N_44149,N_37367,N_35587);
nor U44150 (N_44150,N_35998,N_36998);
nand U44151 (N_44151,N_37752,N_38461);
nor U44152 (N_44152,N_35503,N_36887);
nor U44153 (N_44153,N_37530,N_37377);
xor U44154 (N_44154,N_38076,N_37031);
nor U44155 (N_44155,N_37499,N_37331);
nor U44156 (N_44156,N_38655,N_38395);
and U44157 (N_44157,N_35050,N_39444);
and U44158 (N_44158,N_37200,N_37527);
and U44159 (N_44159,N_36126,N_35090);
nand U44160 (N_44160,N_39062,N_37918);
or U44161 (N_44161,N_36011,N_35258);
xor U44162 (N_44162,N_37025,N_36462);
nor U44163 (N_44163,N_39249,N_35428);
and U44164 (N_44164,N_35205,N_38045);
or U44165 (N_44165,N_38227,N_37768);
and U44166 (N_44166,N_35278,N_35650);
xnor U44167 (N_44167,N_35154,N_39813);
or U44168 (N_44168,N_37670,N_35563);
xnor U44169 (N_44169,N_36287,N_35254);
nor U44170 (N_44170,N_37634,N_35637);
nor U44171 (N_44171,N_36320,N_37056);
or U44172 (N_44172,N_39888,N_38932);
nand U44173 (N_44173,N_37075,N_35003);
nor U44174 (N_44174,N_38774,N_38069);
and U44175 (N_44175,N_38790,N_39176);
xor U44176 (N_44176,N_38018,N_35871);
or U44177 (N_44177,N_35486,N_37688);
nor U44178 (N_44178,N_35312,N_35083);
xor U44179 (N_44179,N_35031,N_38786);
xnor U44180 (N_44180,N_35699,N_38807);
or U44181 (N_44181,N_39033,N_39607);
nor U44182 (N_44182,N_38497,N_35481);
and U44183 (N_44183,N_39454,N_37283);
and U44184 (N_44184,N_39786,N_39831);
and U44185 (N_44185,N_37688,N_37385);
xnor U44186 (N_44186,N_38288,N_38041);
and U44187 (N_44187,N_37265,N_35389);
nor U44188 (N_44188,N_35102,N_37554);
nor U44189 (N_44189,N_35007,N_39138);
nor U44190 (N_44190,N_38717,N_38281);
nand U44191 (N_44191,N_37821,N_35086);
nand U44192 (N_44192,N_39238,N_36936);
nand U44193 (N_44193,N_39272,N_39110);
nor U44194 (N_44194,N_36556,N_35152);
nor U44195 (N_44195,N_36748,N_37658);
or U44196 (N_44196,N_35611,N_39148);
and U44197 (N_44197,N_37368,N_35611);
nor U44198 (N_44198,N_37030,N_35810);
xnor U44199 (N_44199,N_39348,N_36054);
or U44200 (N_44200,N_36165,N_37657);
and U44201 (N_44201,N_36239,N_35614);
nor U44202 (N_44202,N_37435,N_39257);
or U44203 (N_44203,N_38157,N_36361);
nor U44204 (N_44204,N_38811,N_39917);
xnor U44205 (N_44205,N_39401,N_35099);
and U44206 (N_44206,N_37456,N_35735);
and U44207 (N_44207,N_35992,N_37985);
nand U44208 (N_44208,N_35016,N_37149);
or U44209 (N_44209,N_35437,N_35231);
nor U44210 (N_44210,N_39233,N_37221);
and U44211 (N_44211,N_35707,N_36011);
nor U44212 (N_44212,N_39963,N_38447);
or U44213 (N_44213,N_38119,N_35674);
and U44214 (N_44214,N_39261,N_39377);
or U44215 (N_44215,N_38804,N_38809);
nor U44216 (N_44216,N_39210,N_35792);
xnor U44217 (N_44217,N_35334,N_36492);
or U44218 (N_44218,N_36062,N_36346);
nand U44219 (N_44219,N_39885,N_38448);
nand U44220 (N_44220,N_35333,N_38127);
and U44221 (N_44221,N_36403,N_38967);
nand U44222 (N_44222,N_39758,N_36138);
nor U44223 (N_44223,N_35279,N_38045);
nand U44224 (N_44224,N_35127,N_39714);
nand U44225 (N_44225,N_36997,N_35156);
nand U44226 (N_44226,N_35823,N_35242);
or U44227 (N_44227,N_36417,N_35165);
and U44228 (N_44228,N_36977,N_39648);
nand U44229 (N_44229,N_39000,N_37295);
nand U44230 (N_44230,N_36030,N_36255);
or U44231 (N_44231,N_36033,N_38595);
or U44232 (N_44232,N_39259,N_35740);
or U44233 (N_44233,N_39478,N_37968);
or U44234 (N_44234,N_38034,N_35325);
xor U44235 (N_44235,N_36125,N_35801);
nor U44236 (N_44236,N_39993,N_35807);
nand U44237 (N_44237,N_39989,N_38555);
nor U44238 (N_44238,N_36693,N_38599);
xnor U44239 (N_44239,N_35341,N_37525);
nand U44240 (N_44240,N_36892,N_36764);
and U44241 (N_44241,N_36454,N_39442);
nor U44242 (N_44242,N_36162,N_35640);
and U44243 (N_44243,N_38885,N_36183);
xor U44244 (N_44244,N_36051,N_39911);
and U44245 (N_44245,N_37288,N_38865);
or U44246 (N_44246,N_39070,N_37192);
xor U44247 (N_44247,N_38888,N_35589);
nor U44248 (N_44248,N_39651,N_37969);
xnor U44249 (N_44249,N_36919,N_39162);
xnor U44250 (N_44250,N_36181,N_36478);
xnor U44251 (N_44251,N_35212,N_35923);
or U44252 (N_44252,N_39699,N_38064);
nand U44253 (N_44253,N_39235,N_37147);
and U44254 (N_44254,N_37572,N_36454);
xnor U44255 (N_44255,N_36892,N_36877);
or U44256 (N_44256,N_37718,N_38266);
and U44257 (N_44257,N_39974,N_35970);
or U44258 (N_44258,N_36834,N_36155);
or U44259 (N_44259,N_37735,N_36456);
or U44260 (N_44260,N_37749,N_36815);
nor U44261 (N_44261,N_36502,N_39587);
nor U44262 (N_44262,N_39666,N_35951);
nor U44263 (N_44263,N_37107,N_38728);
nor U44264 (N_44264,N_39607,N_38991);
and U44265 (N_44265,N_36392,N_37956);
and U44266 (N_44266,N_36694,N_39203);
nand U44267 (N_44267,N_38313,N_37197);
xor U44268 (N_44268,N_36170,N_36834);
nand U44269 (N_44269,N_36487,N_39232);
nand U44270 (N_44270,N_36479,N_38121);
and U44271 (N_44271,N_36893,N_39880);
nor U44272 (N_44272,N_38905,N_39434);
xor U44273 (N_44273,N_37221,N_38968);
or U44274 (N_44274,N_37956,N_35419);
or U44275 (N_44275,N_39931,N_37769);
and U44276 (N_44276,N_36283,N_36504);
xor U44277 (N_44277,N_38921,N_38379);
nor U44278 (N_44278,N_38128,N_36300);
nand U44279 (N_44279,N_37712,N_39543);
xnor U44280 (N_44280,N_35974,N_35420);
xnor U44281 (N_44281,N_36436,N_38947);
and U44282 (N_44282,N_37083,N_36699);
xor U44283 (N_44283,N_38376,N_37438);
and U44284 (N_44284,N_39227,N_39295);
or U44285 (N_44285,N_36085,N_35481);
nand U44286 (N_44286,N_35541,N_38477);
nand U44287 (N_44287,N_39899,N_36643);
xnor U44288 (N_44288,N_39487,N_38242);
xnor U44289 (N_44289,N_38965,N_36464);
nand U44290 (N_44290,N_35201,N_35949);
and U44291 (N_44291,N_36709,N_37479);
and U44292 (N_44292,N_37716,N_37655);
nand U44293 (N_44293,N_39621,N_39050);
nand U44294 (N_44294,N_35169,N_37486);
nor U44295 (N_44295,N_39989,N_37009);
or U44296 (N_44296,N_38501,N_37903);
nor U44297 (N_44297,N_37765,N_39824);
and U44298 (N_44298,N_38570,N_37827);
and U44299 (N_44299,N_35254,N_37276);
and U44300 (N_44300,N_36189,N_39289);
and U44301 (N_44301,N_38982,N_36396);
or U44302 (N_44302,N_39577,N_39954);
or U44303 (N_44303,N_35994,N_36452);
nor U44304 (N_44304,N_35972,N_36331);
xor U44305 (N_44305,N_38268,N_36516);
nand U44306 (N_44306,N_36013,N_39932);
or U44307 (N_44307,N_39109,N_38259);
nand U44308 (N_44308,N_36218,N_39625);
and U44309 (N_44309,N_37446,N_35537);
nor U44310 (N_44310,N_38925,N_36553);
and U44311 (N_44311,N_37362,N_37753);
xnor U44312 (N_44312,N_36542,N_38984);
nor U44313 (N_44313,N_36233,N_38157);
and U44314 (N_44314,N_35834,N_36847);
and U44315 (N_44315,N_38579,N_37807);
nand U44316 (N_44316,N_35583,N_37996);
nor U44317 (N_44317,N_39951,N_37119);
xnor U44318 (N_44318,N_36291,N_36703);
nand U44319 (N_44319,N_37551,N_37786);
nor U44320 (N_44320,N_39285,N_36557);
or U44321 (N_44321,N_39069,N_37270);
nand U44322 (N_44322,N_39598,N_35350);
xor U44323 (N_44323,N_39263,N_36932);
xor U44324 (N_44324,N_38585,N_37581);
or U44325 (N_44325,N_36814,N_38145);
nand U44326 (N_44326,N_38725,N_37062);
xor U44327 (N_44327,N_37965,N_35734);
xor U44328 (N_44328,N_38529,N_36562);
xnor U44329 (N_44329,N_36094,N_35741);
nor U44330 (N_44330,N_38760,N_38619);
nor U44331 (N_44331,N_39689,N_36546);
nor U44332 (N_44332,N_38123,N_38173);
nor U44333 (N_44333,N_39325,N_36137);
or U44334 (N_44334,N_36623,N_39727);
nand U44335 (N_44335,N_38842,N_39343);
or U44336 (N_44336,N_37443,N_37469);
and U44337 (N_44337,N_35362,N_38608);
nand U44338 (N_44338,N_38398,N_37307);
nor U44339 (N_44339,N_39982,N_38746);
nand U44340 (N_44340,N_35234,N_38221);
nand U44341 (N_44341,N_36519,N_37221);
nand U44342 (N_44342,N_38415,N_36217);
and U44343 (N_44343,N_35905,N_37863);
nor U44344 (N_44344,N_38311,N_38672);
nor U44345 (N_44345,N_39428,N_38919);
nand U44346 (N_44346,N_37920,N_38072);
and U44347 (N_44347,N_35222,N_35716);
and U44348 (N_44348,N_38452,N_37023);
and U44349 (N_44349,N_36572,N_38935);
or U44350 (N_44350,N_39276,N_36245);
or U44351 (N_44351,N_35620,N_37152);
nand U44352 (N_44352,N_38222,N_39024);
xnor U44353 (N_44353,N_39539,N_35818);
and U44354 (N_44354,N_39033,N_38769);
nor U44355 (N_44355,N_38590,N_35521);
nand U44356 (N_44356,N_38977,N_36792);
nor U44357 (N_44357,N_37473,N_38284);
and U44358 (N_44358,N_38772,N_37924);
xor U44359 (N_44359,N_37900,N_36434);
nand U44360 (N_44360,N_39243,N_35415);
and U44361 (N_44361,N_39584,N_36475);
nand U44362 (N_44362,N_37097,N_37108);
xnor U44363 (N_44363,N_35823,N_39030);
xnor U44364 (N_44364,N_36536,N_38073);
and U44365 (N_44365,N_37670,N_39902);
nor U44366 (N_44366,N_39024,N_39427);
and U44367 (N_44367,N_35253,N_39312);
or U44368 (N_44368,N_39432,N_36241);
nand U44369 (N_44369,N_38566,N_35863);
nand U44370 (N_44370,N_36433,N_39644);
nor U44371 (N_44371,N_37002,N_37673);
nor U44372 (N_44372,N_37988,N_37441);
nor U44373 (N_44373,N_35353,N_35718);
xor U44374 (N_44374,N_38109,N_35034);
and U44375 (N_44375,N_39610,N_38797);
nand U44376 (N_44376,N_37436,N_35348);
or U44377 (N_44377,N_36496,N_36593);
nor U44378 (N_44378,N_39970,N_37056);
or U44379 (N_44379,N_39617,N_39055);
nand U44380 (N_44380,N_36183,N_38159);
and U44381 (N_44381,N_37456,N_37121);
xor U44382 (N_44382,N_35652,N_35807);
nand U44383 (N_44383,N_37490,N_37821);
and U44384 (N_44384,N_36462,N_37946);
or U44385 (N_44385,N_36547,N_35905);
nor U44386 (N_44386,N_37642,N_36836);
nor U44387 (N_44387,N_36563,N_35603);
or U44388 (N_44388,N_39516,N_38259);
xor U44389 (N_44389,N_38321,N_39332);
or U44390 (N_44390,N_38594,N_35015);
and U44391 (N_44391,N_37624,N_38871);
nand U44392 (N_44392,N_38856,N_39179);
and U44393 (N_44393,N_36008,N_36430);
nor U44394 (N_44394,N_38886,N_35773);
nand U44395 (N_44395,N_38606,N_37583);
xor U44396 (N_44396,N_36793,N_36652);
nor U44397 (N_44397,N_39524,N_37983);
nor U44398 (N_44398,N_37163,N_38780);
xnor U44399 (N_44399,N_39558,N_37610);
and U44400 (N_44400,N_35023,N_39464);
nor U44401 (N_44401,N_37011,N_35271);
nand U44402 (N_44402,N_37217,N_36757);
and U44403 (N_44403,N_35035,N_36742);
and U44404 (N_44404,N_35313,N_39909);
and U44405 (N_44405,N_36562,N_35678);
or U44406 (N_44406,N_36205,N_38689);
nand U44407 (N_44407,N_36204,N_39678);
and U44408 (N_44408,N_39107,N_35480);
nand U44409 (N_44409,N_35690,N_37323);
xnor U44410 (N_44410,N_37404,N_37202);
nor U44411 (N_44411,N_39986,N_39731);
nor U44412 (N_44412,N_35453,N_37676);
nor U44413 (N_44413,N_37168,N_37672);
nand U44414 (N_44414,N_36141,N_38976);
or U44415 (N_44415,N_38929,N_37982);
or U44416 (N_44416,N_38555,N_38189);
and U44417 (N_44417,N_35878,N_37246);
nand U44418 (N_44418,N_38332,N_38948);
or U44419 (N_44419,N_37127,N_36455);
or U44420 (N_44420,N_35929,N_37071);
and U44421 (N_44421,N_37446,N_38308);
nor U44422 (N_44422,N_39586,N_36886);
nor U44423 (N_44423,N_39149,N_35658);
xnor U44424 (N_44424,N_39403,N_38171);
and U44425 (N_44425,N_37882,N_37179);
or U44426 (N_44426,N_35021,N_38403);
and U44427 (N_44427,N_39332,N_39306);
or U44428 (N_44428,N_38538,N_38324);
or U44429 (N_44429,N_39750,N_38140);
or U44430 (N_44430,N_38148,N_39758);
xor U44431 (N_44431,N_39905,N_36639);
and U44432 (N_44432,N_39090,N_35659);
nor U44433 (N_44433,N_36693,N_38978);
or U44434 (N_44434,N_35042,N_35009);
nor U44435 (N_44435,N_39678,N_36822);
nand U44436 (N_44436,N_35636,N_35548);
or U44437 (N_44437,N_39303,N_35711);
nand U44438 (N_44438,N_38700,N_35145);
and U44439 (N_44439,N_38077,N_36577);
xnor U44440 (N_44440,N_39519,N_38586);
xnor U44441 (N_44441,N_35325,N_39648);
and U44442 (N_44442,N_36329,N_36623);
xnor U44443 (N_44443,N_36110,N_38639);
and U44444 (N_44444,N_39088,N_35988);
xnor U44445 (N_44445,N_36471,N_39066);
or U44446 (N_44446,N_36981,N_35582);
and U44447 (N_44447,N_39782,N_39546);
xnor U44448 (N_44448,N_38937,N_36166);
nor U44449 (N_44449,N_37876,N_37914);
or U44450 (N_44450,N_38367,N_37700);
or U44451 (N_44451,N_37984,N_35263);
and U44452 (N_44452,N_37939,N_36642);
nor U44453 (N_44453,N_37765,N_39802);
and U44454 (N_44454,N_39143,N_38493);
and U44455 (N_44455,N_35577,N_38302);
or U44456 (N_44456,N_35661,N_37421);
xnor U44457 (N_44457,N_37336,N_35719);
xor U44458 (N_44458,N_37208,N_35909);
and U44459 (N_44459,N_37235,N_37074);
and U44460 (N_44460,N_38687,N_38801);
or U44461 (N_44461,N_37303,N_35717);
and U44462 (N_44462,N_36628,N_37301);
xnor U44463 (N_44463,N_36477,N_39496);
xor U44464 (N_44464,N_36812,N_36988);
or U44465 (N_44465,N_38557,N_38020);
nor U44466 (N_44466,N_39459,N_35575);
and U44467 (N_44467,N_36665,N_35306);
nor U44468 (N_44468,N_38012,N_36438);
nor U44469 (N_44469,N_38799,N_36270);
nor U44470 (N_44470,N_36516,N_37987);
and U44471 (N_44471,N_36518,N_39514);
nor U44472 (N_44472,N_38831,N_35921);
xnor U44473 (N_44473,N_38487,N_38101);
or U44474 (N_44474,N_35268,N_38664);
nand U44475 (N_44475,N_36497,N_35051);
xor U44476 (N_44476,N_35512,N_37769);
nand U44477 (N_44477,N_36818,N_35729);
and U44478 (N_44478,N_38099,N_35655);
xnor U44479 (N_44479,N_39140,N_37128);
nor U44480 (N_44480,N_35283,N_36277);
or U44481 (N_44481,N_35496,N_36852);
and U44482 (N_44482,N_38397,N_39696);
xor U44483 (N_44483,N_35294,N_35954);
nand U44484 (N_44484,N_36300,N_38030);
or U44485 (N_44485,N_36055,N_36524);
nand U44486 (N_44486,N_35263,N_38328);
and U44487 (N_44487,N_35792,N_38221);
or U44488 (N_44488,N_37187,N_35446);
xnor U44489 (N_44489,N_35042,N_35262);
and U44490 (N_44490,N_37612,N_35595);
or U44491 (N_44491,N_36821,N_36826);
and U44492 (N_44492,N_35445,N_38812);
nand U44493 (N_44493,N_38574,N_35456);
xnor U44494 (N_44494,N_35027,N_38109);
xor U44495 (N_44495,N_35987,N_39355);
xnor U44496 (N_44496,N_35116,N_39249);
and U44497 (N_44497,N_39335,N_35109);
nand U44498 (N_44498,N_38620,N_38709);
and U44499 (N_44499,N_37326,N_38047);
and U44500 (N_44500,N_38358,N_36008);
and U44501 (N_44501,N_35833,N_37230);
xnor U44502 (N_44502,N_38962,N_39461);
or U44503 (N_44503,N_35444,N_35657);
and U44504 (N_44504,N_38718,N_35776);
or U44505 (N_44505,N_35724,N_38190);
or U44506 (N_44506,N_38087,N_35767);
nor U44507 (N_44507,N_36726,N_38834);
and U44508 (N_44508,N_37862,N_36513);
nor U44509 (N_44509,N_37413,N_36416);
nand U44510 (N_44510,N_35564,N_37060);
nor U44511 (N_44511,N_38325,N_35662);
nor U44512 (N_44512,N_37036,N_35347);
nand U44513 (N_44513,N_36212,N_36035);
or U44514 (N_44514,N_39358,N_36623);
xnor U44515 (N_44515,N_35496,N_35063);
nand U44516 (N_44516,N_38270,N_35385);
or U44517 (N_44517,N_38683,N_39382);
or U44518 (N_44518,N_37402,N_38677);
or U44519 (N_44519,N_38616,N_37005);
and U44520 (N_44520,N_36069,N_37475);
nor U44521 (N_44521,N_39543,N_37353);
nand U44522 (N_44522,N_35639,N_36988);
xnor U44523 (N_44523,N_37210,N_39131);
nor U44524 (N_44524,N_35161,N_38761);
and U44525 (N_44525,N_35648,N_36640);
nor U44526 (N_44526,N_35614,N_39570);
nand U44527 (N_44527,N_39984,N_38443);
and U44528 (N_44528,N_37536,N_36010);
xnor U44529 (N_44529,N_37770,N_39181);
nor U44530 (N_44530,N_38103,N_37722);
and U44531 (N_44531,N_38098,N_37375);
nand U44532 (N_44532,N_39526,N_38003);
nand U44533 (N_44533,N_36856,N_37948);
or U44534 (N_44534,N_35267,N_38107);
or U44535 (N_44535,N_39762,N_36978);
and U44536 (N_44536,N_37635,N_37615);
nand U44537 (N_44537,N_37621,N_35844);
and U44538 (N_44538,N_38575,N_35537);
or U44539 (N_44539,N_36680,N_38188);
nand U44540 (N_44540,N_36633,N_35667);
nand U44541 (N_44541,N_38622,N_37971);
nor U44542 (N_44542,N_36008,N_36976);
xor U44543 (N_44543,N_38316,N_38870);
and U44544 (N_44544,N_36944,N_38835);
nor U44545 (N_44545,N_36414,N_36522);
or U44546 (N_44546,N_38484,N_36668);
nand U44547 (N_44547,N_39651,N_39083);
or U44548 (N_44548,N_35753,N_35313);
and U44549 (N_44549,N_36827,N_37418);
nand U44550 (N_44550,N_37338,N_36943);
nand U44551 (N_44551,N_36023,N_37562);
nor U44552 (N_44552,N_37012,N_38500);
nand U44553 (N_44553,N_39360,N_39543);
and U44554 (N_44554,N_37739,N_39813);
and U44555 (N_44555,N_38755,N_37420);
nor U44556 (N_44556,N_35041,N_39181);
nor U44557 (N_44557,N_38070,N_39014);
xor U44558 (N_44558,N_35924,N_38055);
nor U44559 (N_44559,N_39396,N_38647);
xor U44560 (N_44560,N_35708,N_38737);
and U44561 (N_44561,N_36152,N_38103);
and U44562 (N_44562,N_39700,N_35652);
xnor U44563 (N_44563,N_35814,N_38894);
xor U44564 (N_44564,N_37511,N_37072);
xor U44565 (N_44565,N_37121,N_39763);
or U44566 (N_44566,N_35308,N_35695);
or U44567 (N_44567,N_38224,N_36331);
and U44568 (N_44568,N_35952,N_36978);
or U44569 (N_44569,N_35901,N_38705);
and U44570 (N_44570,N_37575,N_35570);
and U44571 (N_44571,N_36851,N_39219);
and U44572 (N_44572,N_35217,N_35968);
nor U44573 (N_44573,N_35710,N_39376);
nand U44574 (N_44574,N_38610,N_39495);
and U44575 (N_44575,N_36171,N_35060);
and U44576 (N_44576,N_35813,N_38626);
or U44577 (N_44577,N_39542,N_36464);
xor U44578 (N_44578,N_39135,N_39128);
or U44579 (N_44579,N_35979,N_38967);
xnor U44580 (N_44580,N_39555,N_38049);
nand U44581 (N_44581,N_37345,N_35228);
nor U44582 (N_44582,N_38551,N_39051);
nor U44583 (N_44583,N_35991,N_38115);
or U44584 (N_44584,N_38166,N_36340);
and U44585 (N_44585,N_37530,N_39274);
or U44586 (N_44586,N_35342,N_37928);
nor U44587 (N_44587,N_36438,N_35912);
or U44588 (N_44588,N_35712,N_38153);
or U44589 (N_44589,N_36354,N_38241);
nor U44590 (N_44590,N_38947,N_36728);
or U44591 (N_44591,N_39106,N_36295);
and U44592 (N_44592,N_35425,N_35377);
nand U44593 (N_44593,N_36100,N_37986);
nor U44594 (N_44594,N_36493,N_35829);
or U44595 (N_44595,N_36334,N_37659);
and U44596 (N_44596,N_39445,N_38584);
or U44597 (N_44597,N_36789,N_35763);
nor U44598 (N_44598,N_35502,N_36595);
nand U44599 (N_44599,N_37769,N_39100);
xor U44600 (N_44600,N_39480,N_36239);
and U44601 (N_44601,N_36981,N_37597);
xnor U44602 (N_44602,N_38491,N_35811);
and U44603 (N_44603,N_35247,N_35572);
or U44604 (N_44604,N_38454,N_35698);
nor U44605 (N_44605,N_38948,N_37529);
or U44606 (N_44606,N_39264,N_36408);
nor U44607 (N_44607,N_35472,N_37656);
and U44608 (N_44608,N_37379,N_37511);
nand U44609 (N_44609,N_36902,N_37052);
and U44610 (N_44610,N_36247,N_39554);
xor U44611 (N_44611,N_36493,N_39245);
or U44612 (N_44612,N_37962,N_37816);
nor U44613 (N_44613,N_36398,N_39910);
nand U44614 (N_44614,N_39371,N_36374);
nand U44615 (N_44615,N_37740,N_38416);
or U44616 (N_44616,N_37212,N_37078);
nor U44617 (N_44617,N_39028,N_38612);
xnor U44618 (N_44618,N_35260,N_38477);
nor U44619 (N_44619,N_37600,N_39728);
and U44620 (N_44620,N_35624,N_37202);
xor U44621 (N_44621,N_35603,N_35038);
nand U44622 (N_44622,N_38654,N_36652);
nand U44623 (N_44623,N_37740,N_38768);
nor U44624 (N_44624,N_38935,N_36997);
xor U44625 (N_44625,N_39555,N_36231);
nor U44626 (N_44626,N_36517,N_38163);
nand U44627 (N_44627,N_36284,N_35062);
and U44628 (N_44628,N_37606,N_36559);
xor U44629 (N_44629,N_37447,N_36388);
and U44630 (N_44630,N_36066,N_37564);
and U44631 (N_44631,N_38402,N_36814);
and U44632 (N_44632,N_36167,N_39002);
xnor U44633 (N_44633,N_39807,N_39849);
nand U44634 (N_44634,N_36037,N_38498);
nor U44635 (N_44635,N_36952,N_35819);
and U44636 (N_44636,N_36420,N_36852);
nor U44637 (N_44637,N_37944,N_35534);
or U44638 (N_44638,N_39453,N_39029);
nand U44639 (N_44639,N_37326,N_38032);
xnor U44640 (N_44640,N_38062,N_38219);
or U44641 (N_44641,N_35338,N_36758);
xor U44642 (N_44642,N_35449,N_35288);
and U44643 (N_44643,N_37204,N_39660);
and U44644 (N_44644,N_39667,N_38502);
xnor U44645 (N_44645,N_39429,N_35938);
nand U44646 (N_44646,N_39409,N_37795);
nand U44647 (N_44647,N_37666,N_38243);
nand U44648 (N_44648,N_38027,N_39381);
xnor U44649 (N_44649,N_39467,N_36211);
nor U44650 (N_44650,N_35020,N_38009);
nor U44651 (N_44651,N_39069,N_36638);
nor U44652 (N_44652,N_35594,N_37019);
xor U44653 (N_44653,N_38539,N_38989);
and U44654 (N_44654,N_37102,N_35104);
or U44655 (N_44655,N_38878,N_36354);
xnor U44656 (N_44656,N_35849,N_37844);
nor U44657 (N_44657,N_38586,N_37119);
xor U44658 (N_44658,N_35590,N_37659);
and U44659 (N_44659,N_38172,N_35171);
and U44660 (N_44660,N_35434,N_38995);
xor U44661 (N_44661,N_36475,N_36694);
nand U44662 (N_44662,N_36754,N_38542);
nand U44663 (N_44663,N_38519,N_39793);
or U44664 (N_44664,N_35666,N_35140);
or U44665 (N_44665,N_35046,N_39913);
nor U44666 (N_44666,N_37359,N_35948);
xor U44667 (N_44667,N_38303,N_39973);
nor U44668 (N_44668,N_37987,N_38120);
nor U44669 (N_44669,N_39659,N_35430);
and U44670 (N_44670,N_37965,N_37743);
or U44671 (N_44671,N_36082,N_38457);
and U44672 (N_44672,N_39559,N_38283);
and U44673 (N_44673,N_35492,N_39195);
and U44674 (N_44674,N_37983,N_38796);
xor U44675 (N_44675,N_37623,N_38159);
xor U44676 (N_44676,N_37463,N_35029);
or U44677 (N_44677,N_37840,N_38544);
nor U44678 (N_44678,N_38089,N_38225);
or U44679 (N_44679,N_38264,N_39247);
xor U44680 (N_44680,N_35051,N_36324);
xor U44681 (N_44681,N_37434,N_38422);
xor U44682 (N_44682,N_37146,N_37554);
nor U44683 (N_44683,N_35061,N_39998);
nor U44684 (N_44684,N_36128,N_38987);
nor U44685 (N_44685,N_39131,N_39488);
nor U44686 (N_44686,N_36775,N_37782);
and U44687 (N_44687,N_35572,N_39942);
xnor U44688 (N_44688,N_36016,N_35161);
xnor U44689 (N_44689,N_36586,N_37623);
xnor U44690 (N_44690,N_39553,N_36478);
nor U44691 (N_44691,N_39533,N_37595);
nand U44692 (N_44692,N_37271,N_38454);
nor U44693 (N_44693,N_35107,N_39080);
nand U44694 (N_44694,N_38323,N_38477);
xor U44695 (N_44695,N_36386,N_35344);
nor U44696 (N_44696,N_36601,N_37564);
nand U44697 (N_44697,N_38276,N_37698);
xor U44698 (N_44698,N_35934,N_38322);
xnor U44699 (N_44699,N_36478,N_36283);
or U44700 (N_44700,N_38833,N_36001);
nor U44701 (N_44701,N_38014,N_39408);
or U44702 (N_44702,N_36472,N_38514);
xor U44703 (N_44703,N_36768,N_35979);
xnor U44704 (N_44704,N_38194,N_35197);
nor U44705 (N_44705,N_36721,N_35913);
xnor U44706 (N_44706,N_37384,N_36996);
xor U44707 (N_44707,N_39801,N_39809);
nor U44708 (N_44708,N_39647,N_36612);
nor U44709 (N_44709,N_38754,N_36395);
or U44710 (N_44710,N_39826,N_38731);
or U44711 (N_44711,N_35097,N_35585);
and U44712 (N_44712,N_36644,N_38002);
nor U44713 (N_44713,N_37037,N_36258);
nor U44714 (N_44714,N_39267,N_37698);
and U44715 (N_44715,N_38547,N_37171);
nor U44716 (N_44716,N_39673,N_39054);
nor U44717 (N_44717,N_37935,N_38334);
xor U44718 (N_44718,N_38502,N_38024);
and U44719 (N_44719,N_39390,N_37115);
nand U44720 (N_44720,N_36862,N_36596);
nand U44721 (N_44721,N_38668,N_39826);
and U44722 (N_44722,N_38410,N_35126);
xnor U44723 (N_44723,N_35363,N_35594);
nand U44724 (N_44724,N_37883,N_38088);
and U44725 (N_44725,N_37501,N_38459);
and U44726 (N_44726,N_38626,N_39316);
nand U44727 (N_44727,N_36468,N_39593);
nor U44728 (N_44728,N_36724,N_35947);
xor U44729 (N_44729,N_35023,N_38635);
nand U44730 (N_44730,N_35399,N_35506);
and U44731 (N_44731,N_39475,N_38647);
or U44732 (N_44732,N_36557,N_39536);
nor U44733 (N_44733,N_35149,N_37966);
and U44734 (N_44734,N_35372,N_35520);
xnor U44735 (N_44735,N_35493,N_36022);
or U44736 (N_44736,N_37554,N_39721);
nand U44737 (N_44737,N_35216,N_36532);
nand U44738 (N_44738,N_39668,N_37562);
nor U44739 (N_44739,N_35464,N_39665);
xor U44740 (N_44740,N_37617,N_36693);
nor U44741 (N_44741,N_39948,N_38864);
nor U44742 (N_44742,N_36482,N_35165);
xnor U44743 (N_44743,N_38859,N_37371);
and U44744 (N_44744,N_37343,N_39524);
xor U44745 (N_44745,N_36866,N_36983);
nor U44746 (N_44746,N_37158,N_39547);
nand U44747 (N_44747,N_35548,N_37338);
or U44748 (N_44748,N_37308,N_38406);
and U44749 (N_44749,N_35036,N_35166);
or U44750 (N_44750,N_35507,N_39912);
xor U44751 (N_44751,N_36830,N_37173);
xnor U44752 (N_44752,N_39016,N_35553);
nor U44753 (N_44753,N_38368,N_38994);
and U44754 (N_44754,N_36548,N_36275);
nor U44755 (N_44755,N_37576,N_38840);
or U44756 (N_44756,N_39214,N_36906);
nand U44757 (N_44757,N_39354,N_39917);
or U44758 (N_44758,N_39241,N_37577);
nand U44759 (N_44759,N_37855,N_38993);
nand U44760 (N_44760,N_36837,N_38374);
or U44761 (N_44761,N_35999,N_38179);
nand U44762 (N_44762,N_39263,N_36143);
nand U44763 (N_44763,N_35796,N_37932);
nor U44764 (N_44764,N_35597,N_36741);
and U44765 (N_44765,N_36317,N_37216);
xor U44766 (N_44766,N_39929,N_35607);
nand U44767 (N_44767,N_39845,N_38798);
and U44768 (N_44768,N_38459,N_39446);
xnor U44769 (N_44769,N_37219,N_37215);
or U44770 (N_44770,N_39648,N_36750);
nor U44771 (N_44771,N_35900,N_38588);
nor U44772 (N_44772,N_36012,N_38995);
xnor U44773 (N_44773,N_38149,N_38009);
and U44774 (N_44774,N_39662,N_35572);
nor U44775 (N_44775,N_36527,N_36895);
xnor U44776 (N_44776,N_38005,N_39423);
or U44777 (N_44777,N_36346,N_35271);
nor U44778 (N_44778,N_37693,N_39085);
and U44779 (N_44779,N_38070,N_38096);
nand U44780 (N_44780,N_36304,N_36772);
nor U44781 (N_44781,N_36531,N_39570);
nand U44782 (N_44782,N_38301,N_37185);
nand U44783 (N_44783,N_39809,N_37332);
nor U44784 (N_44784,N_37362,N_35689);
xor U44785 (N_44785,N_39857,N_38048);
nand U44786 (N_44786,N_35286,N_36173);
or U44787 (N_44787,N_37291,N_37439);
and U44788 (N_44788,N_35880,N_39353);
nand U44789 (N_44789,N_36051,N_35098);
xnor U44790 (N_44790,N_35396,N_35775);
nor U44791 (N_44791,N_38521,N_35094);
nand U44792 (N_44792,N_36764,N_36217);
and U44793 (N_44793,N_35967,N_35266);
nor U44794 (N_44794,N_39442,N_36209);
and U44795 (N_44795,N_37296,N_39348);
or U44796 (N_44796,N_38817,N_37354);
nand U44797 (N_44797,N_36514,N_39668);
nand U44798 (N_44798,N_38968,N_37380);
nand U44799 (N_44799,N_39597,N_36762);
nor U44800 (N_44800,N_38786,N_38096);
nand U44801 (N_44801,N_37909,N_36990);
nand U44802 (N_44802,N_38484,N_39892);
or U44803 (N_44803,N_35887,N_39841);
or U44804 (N_44804,N_37391,N_39029);
xnor U44805 (N_44805,N_37247,N_35151);
nand U44806 (N_44806,N_37085,N_36283);
and U44807 (N_44807,N_35852,N_38766);
xor U44808 (N_44808,N_38874,N_35925);
or U44809 (N_44809,N_36756,N_35703);
nand U44810 (N_44810,N_39440,N_35719);
and U44811 (N_44811,N_39560,N_35759);
and U44812 (N_44812,N_39868,N_38123);
and U44813 (N_44813,N_35611,N_39633);
nand U44814 (N_44814,N_35106,N_38910);
or U44815 (N_44815,N_37822,N_38848);
and U44816 (N_44816,N_38779,N_39456);
nor U44817 (N_44817,N_35806,N_38710);
and U44818 (N_44818,N_38890,N_37647);
and U44819 (N_44819,N_38040,N_39463);
xor U44820 (N_44820,N_36104,N_37197);
nor U44821 (N_44821,N_38370,N_38690);
xnor U44822 (N_44822,N_39905,N_35424);
nand U44823 (N_44823,N_38945,N_35731);
and U44824 (N_44824,N_39959,N_38799);
nand U44825 (N_44825,N_38200,N_35282);
or U44826 (N_44826,N_35858,N_38674);
nor U44827 (N_44827,N_36230,N_35993);
nor U44828 (N_44828,N_39145,N_36310);
or U44829 (N_44829,N_35203,N_36100);
or U44830 (N_44830,N_37906,N_37242);
or U44831 (N_44831,N_39456,N_36193);
nand U44832 (N_44832,N_36856,N_38919);
nand U44833 (N_44833,N_38558,N_37944);
xor U44834 (N_44834,N_36594,N_39715);
nor U44835 (N_44835,N_37240,N_37770);
nand U44836 (N_44836,N_39570,N_38022);
and U44837 (N_44837,N_39232,N_38019);
and U44838 (N_44838,N_39182,N_35918);
nor U44839 (N_44839,N_37736,N_36707);
xnor U44840 (N_44840,N_35556,N_39131);
nand U44841 (N_44841,N_37095,N_35466);
and U44842 (N_44842,N_37182,N_37634);
nor U44843 (N_44843,N_36087,N_35996);
or U44844 (N_44844,N_36817,N_36425);
or U44845 (N_44845,N_35099,N_35334);
xor U44846 (N_44846,N_39083,N_37501);
xnor U44847 (N_44847,N_36120,N_35401);
nor U44848 (N_44848,N_36052,N_37265);
nand U44849 (N_44849,N_35538,N_39831);
nand U44850 (N_44850,N_39715,N_37308);
nand U44851 (N_44851,N_39200,N_38403);
nand U44852 (N_44852,N_38524,N_37250);
xor U44853 (N_44853,N_39740,N_36135);
nor U44854 (N_44854,N_37128,N_36489);
and U44855 (N_44855,N_39604,N_37900);
nor U44856 (N_44856,N_39731,N_36298);
nor U44857 (N_44857,N_38975,N_36762);
nor U44858 (N_44858,N_36330,N_39044);
and U44859 (N_44859,N_36970,N_37326);
or U44860 (N_44860,N_37465,N_37789);
xnor U44861 (N_44861,N_36675,N_38046);
and U44862 (N_44862,N_38712,N_35330);
or U44863 (N_44863,N_35874,N_38139);
nand U44864 (N_44864,N_37684,N_38597);
xor U44865 (N_44865,N_38779,N_38081);
nor U44866 (N_44866,N_35252,N_38191);
and U44867 (N_44867,N_36328,N_38217);
or U44868 (N_44868,N_37106,N_38489);
or U44869 (N_44869,N_36737,N_37880);
or U44870 (N_44870,N_39496,N_38262);
and U44871 (N_44871,N_37598,N_36459);
or U44872 (N_44872,N_39717,N_38474);
xnor U44873 (N_44873,N_37261,N_37048);
xor U44874 (N_44874,N_39364,N_39179);
xor U44875 (N_44875,N_37126,N_38708);
nand U44876 (N_44876,N_35440,N_38570);
xnor U44877 (N_44877,N_39283,N_35937);
and U44878 (N_44878,N_35367,N_36183);
and U44879 (N_44879,N_39615,N_35000);
xnor U44880 (N_44880,N_39320,N_36879);
and U44881 (N_44881,N_39990,N_37748);
nor U44882 (N_44882,N_39211,N_36919);
or U44883 (N_44883,N_37487,N_36467);
nand U44884 (N_44884,N_38775,N_35028);
xor U44885 (N_44885,N_36188,N_36607);
nor U44886 (N_44886,N_35726,N_38342);
nand U44887 (N_44887,N_37711,N_37444);
xor U44888 (N_44888,N_38897,N_35685);
nor U44889 (N_44889,N_36955,N_39465);
nand U44890 (N_44890,N_39461,N_39004);
nand U44891 (N_44891,N_37870,N_35439);
nor U44892 (N_44892,N_39148,N_39386);
or U44893 (N_44893,N_39738,N_36743);
nor U44894 (N_44894,N_36635,N_37915);
xnor U44895 (N_44895,N_39837,N_35966);
xnor U44896 (N_44896,N_38929,N_38145);
nand U44897 (N_44897,N_36434,N_38239);
or U44898 (N_44898,N_36690,N_39748);
nor U44899 (N_44899,N_37284,N_39943);
or U44900 (N_44900,N_38965,N_35274);
or U44901 (N_44901,N_38750,N_35311);
nand U44902 (N_44902,N_39654,N_36034);
xnor U44903 (N_44903,N_35439,N_39176);
and U44904 (N_44904,N_36271,N_39983);
nand U44905 (N_44905,N_37963,N_37596);
xor U44906 (N_44906,N_39292,N_37956);
or U44907 (N_44907,N_38421,N_37854);
and U44908 (N_44908,N_36244,N_37703);
or U44909 (N_44909,N_38782,N_38477);
or U44910 (N_44910,N_39811,N_35886);
nand U44911 (N_44911,N_37666,N_36012);
and U44912 (N_44912,N_38368,N_35393);
nor U44913 (N_44913,N_37864,N_39433);
and U44914 (N_44914,N_37489,N_38299);
nand U44915 (N_44915,N_37866,N_36375);
nand U44916 (N_44916,N_39392,N_37372);
xnor U44917 (N_44917,N_38404,N_38557);
nand U44918 (N_44918,N_35001,N_39046);
nand U44919 (N_44919,N_39675,N_38707);
and U44920 (N_44920,N_37923,N_35914);
and U44921 (N_44921,N_38007,N_36810);
and U44922 (N_44922,N_38585,N_38281);
or U44923 (N_44923,N_37145,N_37596);
nand U44924 (N_44924,N_38020,N_37698);
or U44925 (N_44925,N_39030,N_39191);
nor U44926 (N_44926,N_39741,N_36791);
nand U44927 (N_44927,N_37904,N_39046);
nand U44928 (N_44928,N_39248,N_39952);
nand U44929 (N_44929,N_36628,N_35880);
and U44930 (N_44930,N_39486,N_38066);
nand U44931 (N_44931,N_38191,N_36852);
nor U44932 (N_44932,N_35573,N_38520);
nand U44933 (N_44933,N_37644,N_36486);
xnor U44934 (N_44934,N_37787,N_37160);
nor U44935 (N_44935,N_37747,N_38521);
or U44936 (N_44936,N_37365,N_38110);
and U44937 (N_44937,N_38395,N_38748);
or U44938 (N_44938,N_38050,N_36411);
or U44939 (N_44939,N_38527,N_37588);
and U44940 (N_44940,N_35703,N_38149);
xor U44941 (N_44941,N_38025,N_38124);
nand U44942 (N_44942,N_35203,N_37330);
or U44943 (N_44943,N_38105,N_39249);
nor U44944 (N_44944,N_38740,N_38346);
nand U44945 (N_44945,N_38237,N_39170);
and U44946 (N_44946,N_36031,N_37202);
xnor U44947 (N_44947,N_35788,N_39163);
or U44948 (N_44948,N_36145,N_37408);
and U44949 (N_44949,N_38757,N_39478);
nand U44950 (N_44950,N_36091,N_37296);
xnor U44951 (N_44951,N_38080,N_35744);
xnor U44952 (N_44952,N_35943,N_37151);
xnor U44953 (N_44953,N_39307,N_39502);
nand U44954 (N_44954,N_39250,N_36861);
nand U44955 (N_44955,N_36077,N_39185);
and U44956 (N_44956,N_36937,N_37277);
xor U44957 (N_44957,N_38123,N_37856);
nor U44958 (N_44958,N_39711,N_38275);
and U44959 (N_44959,N_36749,N_39573);
nand U44960 (N_44960,N_39092,N_35864);
or U44961 (N_44961,N_39682,N_35935);
nor U44962 (N_44962,N_38189,N_39510);
nand U44963 (N_44963,N_36879,N_36039);
or U44964 (N_44964,N_39470,N_39610);
xnor U44965 (N_44965,N_37485,N_36441);
xor U44966 (N_44966,N_37513,N_39813);
nor U44967 (N_44967,N_36450,N_39294);
xor U44968 (N_44968,N_36211,N_37047);
nand U44969 (N_44969,N_39520,N_37876);
and U44970 (N_44970,N_39564,N_39134);
or U44971 (N_44971,N_35792,N_35689);
and U44972 (N_44972,N_37597,N_35501);
nor U44973 (N_44973,N_38171,N_35914);
or U44974 (N_44974,N_38417,N_38795);
xnor U44975 (N_44975,N_38150,N_35540);
nor U44976 (N_44976,N_37224,N_39730);
or U44977 (N_44977,N_37386,N_35229);
and U44978 (N_44978,N_39528,N_38003);
and U44979 (N_44979,N_38252,N_39321);
nor U44980 (N_44980,N_38572,N_38691);
xnor U44981 (N_44981,N_35756,N_35248);
nor U44982 (N_44982,N_35783,N_38447);
and U44983 (N_44983,N_37100,N_39298);
and U44984 (N_44984,N_37429,N_39380);
and U44985 (N_44985,N_35008,N_39283);
xnor U44986 (N_44986,N_37615,N_38139);
nand U44987 (N_44987,N_37145,N_36435);
nand U44988 (N_44988,N_38241,N_36958);
xnor U44989 (N_44989,N_37433,N_38370);
or U44990 (N_44990,N_37294,N_35814);
and U44991 (N_44991,N_38240,N_39672);
nor U44992 (N_44992,N_35614,N_38234);
or U44993 (N_44993,N_39602,N_36182);
nand U44994 (N_44994,N_35800,N_39942);
or U44995 (N_44995,N_38574,N_38491);
nor U44996 (N_44996,N_37654,N_36850);
xor U44997 (N_44997,N_35647,N_39389);
and U44998 (N_44998,N_36443,N_36783);
nor U44999 (N_44999,N_37293,N_38518);
nor U45000 (N_45000,N_42941,N_41762);
or U45001 (N_45001,N_41385,N_40431);
nor U45002 (N_45002,N_40896,N_41590);
nand U45003 (N_45003,N_43780,N_40312);
nor U45004 (N_45004,N_41063,N_42136);
nand U45005 (N_45005,N_41391,N_42653);
nor U45006 (N_45006,N_44280,N_42746);
or U45007 (N_45007,N_44665,N_40861);
nand U45008 (N_45008,N_43283,N_41470);
or U45009 (N_45009,N_40919,N_43866);
and U45010 (N_45010,N_40239,N_44300);
nor U45011 (N_45011,N_42438,N_44456);
and U45012 (N_45012,N_42801,N_41288);
xnor U45013 (N_45013,N_43830,N_40955);
nor U45014 (N_45014,N_43470,N_44038);
nand U45015 (N_45015,N_41071,N_42970);
xnor U45016 (N_45016,N_40951,N_40093);
xor U45017 (N_45017,N_42270,N_41813);
nand U45018 (N_45018,N_42637,N_40615);
nand U45019 (N_45019,N_43654,N_40260);
and U45020 (N_45020,N_43720,N_41963);
and U45021 (N_45021,N_44970,N_43106);
and U45022 (N_45022,N_42243,N_41557);
nand U45023 (N_45023,N_41347,N_40676);
xor U45024 (N_45024,N_43137,N_40787);
xnor U45025 (N_45025,N_40458,N_43526);
nand U45026 (N_45026,N_42093,N_40317);
nand U45027 (N_45027,N_43399,N_44897);
and U45028 (N_45028,N_40358,N_41792);
and U45029 (N_45029,N_43394,N_40927);
xor U45030 (N_45030,N_43496,N_43999);
and U45031 (N_45031,N_44940,N_42635);
xnor U45032 (N_45032,N_41240,N_42834);
or U45033 (N_45033,N_43902,N_41205);
or U45034 (N_45034,N_40820,N_44728);
or U45035 (N_45035,N_43338,N_41969);
nor U45036 (N_45036,N_42052,N_43737);
or U45037 (N_45037,N_41147,N_42462);
nor U45038 (N_45038,N_43497,N_40945);
or U45039 (N_45039,N_43628,N_41647);
nand U45040 (N_45040,N_42456,N_42795);
nand U45041 (N_45041,N_42115,N_42512);
nor U45042 (N_45042,N_42631,N_42691);
or U45043 (N_45043,N_44944,N_40717);
xnor U45044 (N_45044,N_42302,N_41660);
xor U45045 (N_45045,N_42851,N_40072);
nor U45046 (N_45046,N_42586,N_42413);
or U45047 (N_45047,N_44269,N_43082);
and U45048 (N_45048,N_44289,N_44333);
xnor U45049 (N_45049,N_41268,N_44595);
xor U45050 (N_45050,N_42471,N_40636);
nor U45051 (N_45051,N_40759,N_41734);
nand U45052 (N_45052,N_41508,N_44208);
or U45053 (N_45053,N_41368,N_43589);
nand U45054 (N_45054,N_42830,N_42117);
xnor U45055 (N_45055,N_40572,N_41922);
nor U45056 (N_45056,N_42472,N_44635);
nand U45057 (N_45057,N_42569,N_44015);
xnor U45058 (N_45058,N_41487,N_41767);
nor U45059 (N_45059,N_42762,N_41970);
or U45060 (N_45060,N_44697,N_40825);
xor U45061 (N_45061,N_42086,N_40757);
or U45062 (N_45062,N_44872,N_42181);
or U45063 (N_45063,N_40700,N_44692);
nor U45064 (N_45064,N_41124,N_44762);
or U45065 (N_45065,N_43693,N_42233);
nor U45066 (N_45066,N_43197,N_41296);
xnor U45067 (N_45067,N_42773,N_41967);
or U45068 (N_45068,N_42336,N_43371);
and U45069 (N_45069,N_44524,N_40149);
and U45070 (N_45070,N_40224,N_42999);
xnor U45071 (N_45071,N_44436,N_44474);
and U45072 (N_45072,N_40283,N_42210);
nor U45073 (N_45073,N_43125,N_43224);
nand U45074 (N_45074,N_44854,N_42615);
or U45075 (N_45075,N_41444,N_41014);
or U45076 (N_45076,N_41087,N_44032);
xnor U45077 (N_45077,N_41153,N_41715);
nor U45078 (N_45078,N_42397,N_40301);
xnor U45079 (N_45079,N_41214,N_40668);
and U45080 (N_45080,N_44306,N_43630);
or U45081 (N_45081,N_41742,N_43129);
nor U45082 (N_45082,N_40745,N_42562);
nor U45083 (N_45083,N_44618,N_44473);
nand U45084 (N_45084,N_44251,N_44139);
or U45085 (N_45085,N_42262,N_42351);
and U45086 (N_45086,N_44347,N_42113);
or U45087 (N_45087,N_44416,N_40021);
nand U45088 (N_45088,N_44562,N_41149);
nand U45089 (N_45089,N_40444,N_42257);
and U45090 (N_45090,N_42112,N_40735);
nand U45091 (N_45091,N_41882,N_43366);
or U45092 (N_45092,N_42700,N_43325);
nor U45093 (N_45093,N_43282,N_44846);
nor U45094 (N_45094,N_42187,N_40201);
xnor U45095 (N_45095,N_42904,N_40263);
nand U45096 (N_45096,N_40567,N_42287);
or U45097 (N_45097,N_43947,N_43181);
xor U45098 (N_45098,N_44177,N_40988);
nand U45099 (N_45099,N_42687,N_41401);
or U45100 (N_45100,N_43350,N_44200);
or U45101 (N_45101,N_43518,N_43736);
or U45102 (N_45102,N_44369,N_42249);
and U45103 (N_45103,N_44112,N_42053);
and U45104 (N_45104,N_41408,N_40216);
nand U45105 (N_45105,N_43632,N_42502);
xor U45106 (N_45106,N_43735,N_44540);
xnor U45107 (N_45107,N_41726,N_42190);
or U45108 (N_45108,N_41949,N_41561);
nor U45109 (N_45109,N_40142,N_43059);
xnor U45110 (N_45110,N_43126,N_44935);
xor U45111 (N_45111,N_40899,N_40023);
or U45112 (N_45112,N_40950,N_43533);
nand U45113 (N_45113,N_42792,N_40967);
or U45114 (N_45114,N_42808,N_43367);
xor U45115 (N_45115,N_42650,N_44435);
or U45116 (N_45116,N_41155,N_43025);
xor U45117 (N_45117,N_41649,N_40491);
xor U45118 (N_45118,N_44817,N_42704);
nand U45119 (N_45119,N_40114,N_40248);
or U45120 (N_45120,N_42370,N_40859);
or U45121 (N_45121,N_40590,N_44071);
and U45122 (N_45122,N_42170,N_42162);
xnor U45123 (N_45123,N_43670,N_41950);
or U45124 (N_45124,N_42060,N_41816);
nand U45125 (N_45125,N_42359,N_40771);
nor U45126 (N_45126,N_40936,N_43638);
nand U45127 (N_45127,N_42987,N_41801);
nand U45128 (N_45128,N_42638,N_43853);
nor U45129 (N_45129,N_43984,N_40760);
xnor U45130 (N_45130,N_40067,N_41624);
xnor U45131 (N_45131,N_40664,N_42936);
and U45132 (N_45132,N_44245,N_41775);
nor U45133 (N_45133,N_41379,N_40185);
and U45134 (N_45134,N_40229,N_44033);
and U45135 (N_45135,N_41419,N_43202);
nor U45136 (N_45136,N_42744,N_42309);
or U45137 (N_45137,N_40698,N_43817);
nand U45138 (N_45138,N_40543,N_42361);
nand U45139 (N_45139,N_42515,N_44201);
and U45140 (N_45140,N_41946,N_43214);
xor U45141 (N_45141,N_44716,N_41743);
and U45142 (N_45142,N_42558,N_40715);
nand U45143 (N_45143,N_44604,N_42924);
nand U45144 (N_45144,N_44822,N_40837);
xnor U45145 (N_45145,N_43225,N_41681);
nor U45146 (N_45146,N_43344,N_40970);
xor U45147 (N_45147,N_41522,N_43631);
and U45148 (N_45148,N_40827,N_41261);
xor U45149 (N_45149,N_40932,N_40391);
and U45150 (N_45150,N_42372,N_42278);
nor U45151 (N_45151,N_43748,N_42894);
nor U45152 (N_45152,N_44580,N_41892);
and U45153 (N_45153,N_44429,N_44180);
nor U45154 (N_45154,N_41777,N_41981);
nand U45155 (N_45155,N_42717,N_44099);
and U45156 (N_45156,N_43802,N_42193);
nor U45157 (N_45157,N_43969,N_44359);
nor U45158 (N_45158,N_43369,N_44262);
nor U45159 (N_45159,N_41115,N_42793);
nand U45160 (N_45160,N_40345,N_43647);
and U45161 (N_45161,N_42791,N_40066);
nand U45162 (N_45162,N_40087,N_40480);
or U45163 (N_45163,N_44956,N_43359);
or U45164 (N_45164,N_43188,N_43039);
nand U45165 (N_45165,N_43103,N_41366);
nor U45166 (N_45166,N_44044,N_40349);
and U45167 (N_45167,N_40853,N_43566);
xor U45168 (N_45168,N_40915,N_44478);
or U45169 (N_45169,N_44643,N_44081);
nand U45170 (N_45170,N_40037,N_41984);
xnor U45171 (N_45171,N_44975,N_40638);
and U45172 (N_45172,N_44971,N_44838);
and U45173 (N_45173,N_42268,N_40714);
xor U45174 (N_45174,N_42495,N_41934);
nand U45175 (N_45175,N_41693,N_41815);
nor U45176 (N_45176,N_42223,N_44093);
nand U45177 (N_45177,N_42751,N_43576);
nand U45178 (N_45178,N_40725,N_41502);
nand U45179 (N_45179,N_41553,N_43121);
or U45180 (N_45180,N_44060,N_42568);
nor U45181 (N_45181,N_44632,N_40669);
nand U45182 (N_45182,N_40310,N_41409);
or U45183 (N_45183,N_40790,N_41318);
nor U45184 (N_45184,N_41266,N_43538);
nor U45185 (N_45185,N_44482,N_41988);
and U45186 (N_45186,N_40098,N_40257);
xnor U45187 (N_45187,N_41944,N_43959);
xnor U45188 (N_45188,N_41940,N_43781);
xor U45189 (N_45189,N_40267,N_40702);
or U45190 (N_45190,N_42705,N_42885);
nand U45191 (N_45191,N_40075,N_42730);
nor U45192 (N_45192,N_42364,N_44963);
xor U45193 (N_45193,N_41571,N_40435);
nand U45194 (N_45194,N_41051,N_40404);
nand U45195 (N_45195,N_40238,N_44118);
nor U45196 (N_45196,N_40370,N_44009);
xor U45197 (N_45197,N_43926,N_41622);
nand U45198 (N_45198,N_43938,N_43045);
xor U45199 (N_45199,N_44465,N_41180);
xor U45200 (N_45200,N_42982,N_41628);
and U45201 (N_45201,N_44171,N_41304);
nand U45202 (N_45202,N_43248,N_43149);
and U45203 (N_45203,N_41723,N_41298);
or U45204 (N_45204,N_41231,N_43998);
nor U45205 (N_45205,N_41370,N_42642);
xor U45206 (N_45206,N_40335,N_41835);
nor U45207 (N_45207,N_41161,N_43711);
nand U45208 (N_45208,N_40971,N_40848);
nand U45209 (N_45209,N_43501,N_42483);
and U45210 (N_45210,N_41454,N_42748);
xnor U45211 (N_45211,N_40459,N_43118);
xnor U45212 (N_45212,N_44389,N_44973);
nand U45213 (N_45213,N_44159,N_44902);
or U45214 (N_45214,N_41962,N_43411);
and U45215 (N_45215,N_42977,N_43457);
and U45216 (N_45216,N_40105,N_43491);
nand U45217 (N_45217,N_44727,N_44192);
nor U45218 (N_45218,N_41461,N_41684);
nand U45219 (N_45219,N_41621,N_42334);
nor U45220 (N_45220,N_44880,N_44431);
or U45221 (N_45221,N_42485,N_44411);
and U45222 (N_45222,N_41250,N_41668);
and U45223 (N_45223,N_43459,N_43981);
and U45224 (N_45224,N_43458,N_40772);
nor U45225 (N_45225,N_43275,N_42360);
or U45226 (N_45226,N_44253,N_43398);
or U45227 (N_45227,N_44212,N_41282);
xor U45228 (N_45228,N_40095,N_44368);
xor U45229 (N_45229,N_41467,N_44041);
nor U45230 (N_45230,N_44862,N_41905);
nor U45231 (N_45231,N_43029,N_43562);
nand U45232 (N_45232,N_42685,N_40078);
or U45233 (N_45233,N_41039,N_43657);
nor U45234 (N_45234,N_40341,N_44030);
xnor U45235 (N_45235,N_43838,N_43454);
or U45236 (N_45236,N_44448,N_44188);
and U45237 (N_45237,N_40050,N_40205);
nor U45238 (N_45238,N_44185,N_40278);
or U45239 (N_45239,N_41334,N_42988);
or U45240 (N_45240,N_40150,N_40054);
nand U45241 (N_45241,N_42037,N_42484);
nand U45242 (N_45242,N_41840,N_41993);
and U45243 (N_45243,N_42218,N_44608);
nand U45244 (N_45244,N_43370,N_40268);
xnor U45245 (N_45245,N_43060,N_43922);
and U45246 (N_45246,N_40764,N_42134);
xor U45247 (N_45247,N_40166,N_40693);
nand U45248 (N_45248,N_44860,N_40364);
xnor U45249 (N_45249,N_40195,N_42716);
nand U45250 (N_45250,N_40289,N_43081);
and U45251 (N_45251,N_43074,N_43556);
and U45252 (N_45252,N_41773,N_43320);
xor U45253 (N_45253,N_40610,N_41400);
xnor U45254 (N_45254,N_42902,N_44736);
or U45255 (N_45255,N_42958,N_42414);
xnor U45256 (N_45256,N_40875,N_42008);
nand U45257 (N_45257,N_40934,N_41437);
nor U45258 (N_45258,N_41802,N_44348);
xor U45259 (N_45259,N_43688,N_43784);
nor U45260 (N_45260,N_43757,N_43294);
xnor U45261 (N_45261,N_40536,N_40938);
xnor U45262 (N_45262,N_42064,N_42989);
xor U45263 (N_45263,N_40448,N_44903);
xnor U45264 (N_45264,N_42587,N_42421);
nand U45265 (N_45265,N_44248,N_43226);
nand U45266 (N_45266,N_43531,N_44377);
nand U45267 (N_45267,N_41024,N_43582);
nor U45268 (N_45268,N_42927,N_41337);
and U45269 (N_45269,N_44585,N_42247);
nand U45270 (N_45270,N_43343,N_40100);
nand U45271 (N_45271,N_40152,N_44126);
and U45272 (N_45272,N_43260,N_41291);
and U45273 (N_45273,N_40477,N_43009);
nand U45274 (N_45274,N_41355,N_43528);
xor U45275 (N_45275,N_40911,N_43416);
nor U45276 (N_45276,N_40261,N_44357);
and U45277 (N_45277,N_41852,N_41771);
nor U45278 (N_45278,N_41617,N_41045);
or U45279 (N_45279,N_42627,N_41806);
nand U45280 (N_45280,N_43641,N_40868);
and U45281 (N_45281,N_40390,N_42046);
nor U45282 (N_45282,N_40846,N_44390);
and U45283 (N_45283,N_40338,N_42632);
nor U45284 (N_45284,N_44628,N_41193);
nand U45285 (N_45285,N_40116,N_44645);
and U45286 (N_45286,N_44680,N_44847);
or U45287 (N_45287,N_43982,N_41332);
or U45288 (N_45288,N_44741,N_40344);
xor U45289 (N_45289,N_40797,N_44802);
nand U45290 (N_45290,N_40786,N_43919);
or U45291 (N_45291,N_43179,N_40946);
or U45292 (N_45292,N_40887,N_41455);
nand U45293 (N_45293,N_43231,N_42141);
and U45294 (N_45294,N_40056,N_43148);
nand U45295 (N_45295,N_44052,N_44361);
nor U45296 (N_45296,N_44577,N_40769);
and U45297 (N_45297,N_40704,N_44063);
nor U45298 (N_45298,N_40677,N_42812);
nand U45299 (N_45299,N_44279,N_43951);
nor U45300 (N_45300,N_43418,N_40972);
xor U45301 (N_45301,N_43395,N_40481);
and U45302 (N_45302,N_41381,N_42435);
xor U45303 (N_45303,N_43574,N_41744);
nand U45304 (N_45304,N_40619,N_42279);
nand U45305 (N_45305,N_41386,N_40627);
and U45306 (N_45306,N_41070,N_44710);
or U45307 (N_45307,N_44203,N_41239);
and U45308 (N_45308,N_40751,N_40778);
nor U45309 (N_45309,N_42550,N_43808);
nor U45310 (N_45310,N_43384,N_44241);
nand U45311 (N_45311,N_41781,N_40197);
and U45312 (N_45312,N_42025,N_42585);
and U45313 (N_45313,N_42544,N_42583);
and U45314 (N_45314,N_41348,N_42592);
or U45315 (N_45315,N_40531,N_44107);
or U45316 (N_45316,N_43506,N_44437);
xor U45317 (N_45317,N_42817,N_43168);
and U45318 (N_45318,N_40383,N_43228);
and U45319 (N_45319,N_44529,N_40975);
nor U45320 (N_45320,N_43358,N_44045);
xnor U45321 (N_45321,N_44109,N_43667);
or U45322 (N_45322,N_43712,N_40532);
or U45323 (N_45323,N_43655,N_43656);
xor U45324 (N_45324,N_40112,N_41344);
and U45325 (N_45325,N_40001,N_43405);
and U45326 (N_45326,N_44138,N_42572);
or U45327 (N_45327,N_44864,N_42844);
xor U45328 (N_45328,N_41476,N_41639);
nor U45329 (N_45329,N_43776,N_41229);
xor U45330 (N_45330,N_42580,N_43747);
and U45331 (N_45331,N_42680,N_41544);
nor U45332 (N_45332,N_43024,N_42840);
or U45333 (N_45333,N_44210,N_42165);
nand U45334 (N_45334,N_41083,N_40443);
xor U45335 (N_45335,N_42330,N_40523);
nor U45336 (N_45336,N_42657,N_41152);
or U45337 (N_45337,N_43990,N_40012);
nor U45338 (N_45338,N_41791,N_41827);
nor U45339 (N_45339,N_43852,N_42600);
xor U45340 (N_45340,N_40298,N_43334);
xor U45341 (N_45341,N_44219,N_43683);
nor U45342 (N_45342,N_43699,N_44085);
or U45343 (N_45343,N_40277,N_40159);
nand U45344 (N_45344,N_40940,N_41423);
or U45345 (N_45345,N_42822,N_40094);
or U45346 (N_45346,N_44647,N_42384);
nor U45347 (N_45347,N_40371,N_40897);
nor U45348 (N_45348,N_44922,N_42248);
and U45349 (N_45349,N_43005,N_41997);
and U45350 (N_45350,N_41146,N_43704);
or U45351 (N_45351,N_41914,N_42103);
xor U45352 (N_45352,N_42080,N_41085);
and U45353 (N_45353,N_41938,N_41587);
and U45354 (N_45354,N_43162,N_44329);
nand U45355 (N_45355,N_42481,N_44891);
nand U45356 (N_45356,N_42332,N_42229);
nor U45357 (N_45357,N_44867,N_40929);
nand U45358 (N_45358,N_41450,N_40992);
and U45359 (N_45359,N_43002,N_42007);
xnor U45360 (N_45360,N_40752,N_44278);
nand U45361 (N_45361,N_43831,N_42777);
nor U45362 (N_45362,N_44589,N_44384);
and U45363 (N_45363,N_44855,N_43382);
and U45364 (N_45364,N_43105,N_42898);
nor U45365 (N_45365,N_40308,N_42644);
and U45366 (N_45366,N_40128,N_41463);
xnor U45367 (N_45367,N_40770,N_41828);
or U45368 (N_45368,N_44826,N_41549);
and U45369 (N_45369,N_41688,N_43408);
and U45370 (N_45370,N_40419,N_43027);
or U45371 (N_45371,N_40518,N_43452);
or U45372 (N_45372,N_43575,N_41412);
nor U45373 (N_45373,N_41689,N_41739);
xnor U45374 (N_45374,N_42900,N_44412);
or U45375 (N_45375,N_44931,N_41211);
nand U45376 (N_45376,N_41812,N_44001);
and U45377 (N_45377,N_43883,N_43098);
nand U45378 (N_45378,N_44307,N_44655);
or U45379 (N_45379,N_42827,N_42617);
nor U45380 (N_45380,N_43598,N_40234);
or U45381 (N_45381,N_41328,N_44950);
nand U45382 (N_45382,N_44504,N_41089);
or U45383 (N_45383,N_41746,N_42918);
nand U45384 (N_45384,N_43288,N_43966);
and U45385 (N_45385,N_42608,N_40305);
or U45386 (N_45386,N_41595,N_43347);
or U45387 (N_45387,N_44488,N_42677);
nand U45388 (N_45388,N_40004,N_44754);
and U45389 (N_45389,N_44191,N_40608);
xor U45390 (N_45390,N_43665,N_40549);
xor U45391 (N_45391,N_44545,N_42298);
nor U45392 (N_45392,N_40139,N_44483);
or U45393 (N_45393,N_42156,N_40879);
or U45394 (N_45394,N_40813,N_42802);
and U45395 (N_45395,N_43270,N_41800);
nor U45396 (N_45396,N_43013,N_44806);
xor U45397 (N_45397,N_42625,N_43007);
xor U45398 (N_45398,N_44681,N_41360);
nand U45399 (N_45399,N_43186,N_44338);
and U45400 (N_45400,N_43507,N_43573);
nand U45401 (N_45401,N_43061,N_41990);
xnor U45402 (N_45402,N_40791,N_40161);
nor U45403 (N_45403,N_41046,N_43836);
xor U45404 (N_45404,N_42574,N_40379);
nand U45405 (N_45405,N_44297,N_43389);
or U45406 (N_45406,N_41507,N_40131);
and U45407 (N_45407,N_43298,N_44987);
nor U45408 (N_45408,N_41367,N_40104);
or U45409 (N_45409,N_42910,N_44160);
xor U45410 (N_45410,N_42534,N_44325);
nand U45411 (N_45411,N_40452,N_40653);
xor U45412 (N_45412,N_40434,N_41503);
nor U45413 (N_45413,N_40099,N_44719);
xnor U45414 (N_45414,N_40713,N_40027);
xor U45415 (N_45415,N_42752,N_43925);
xnor U45416 (N_45416,N_42595,N_43714);
nor U45417 (N_45417,N_42137,N_40961);
xnor U45418 (N_45418,N_43602,N_43687);
and U45419 (N_45419,N_44974,N_44827);
and U45420 (N_45420,N_43851,N_41896);
nor U45421 (N_45421,N_41469,N_40577);
and U45422 (N_45422,N_44277,N_40160);
nand U45423 (N_45423,N_40175,N_40976);
nand U45424 (N_45424,N_42794,N_43662);
or U45425 (N_45425,N_44108,N_42643);
nor U45426 (N_45426,N_44290,N_44737);
xor U45427 (N_45427,N_43522,N_42565);
or U45428 (N_45428,N_43284,N_44764);
or U45429 (N_45429,N_40336,N_40040);
xnor U45430 (N_45430,N_43601,N_42199);
nand U45431 (N_45431,N_44875,N_40429);
nor U45432 (N_45432,N_44965,N_44335);
nand U45433 (N_45433,N_43119,N_42452);
nor U45434 (N_45434,N_40965,N_43274);
xor U45435 (N_45435,N_40123,N_42538);
nand U45436 (N_45436,N_43678,N_40252);
nor U45437 (N_45437,N_40593,N_43837);
nor U45438 (N_45438,N_41558,N_41378);
xor U45439 (N_45439,N_44567,N_44639);
nand U45440 (N_45440,N_40952,N_40513);
xor U45441 (N_45441,N_42449,N_41172);
xnor U45442 (N_45442,N_43327,N_43595);
and U45443 (N_45443,N_42504,N_41208);
or U45444 (N_45444,N_40993,N_43096);
nand U45445 (N_45445,N_40376,N_41420);
and U45446 (N_45446,N_41310,N_42208);
and U45447 (N_45447,N_44767,N_42041);
xor U45448 (N_45448,N_44927,N_43640);
and U45449 (N_45449,N_43484,N_44910);
nand U45450 (N_45450,N_40734,N_44418);
nor U45451 (N_45451,N_41652,N_40284);
or U45452 (N_45452,N_44076,N_42873);
nand U45453 (N_45453,N_41279,N_41442);
xnor U45454 (N_45454,N_40401,N_40985);
nor U45455 (N_45455,N_44649,N_41207);
nor U45456 (N_45456,N_43431,N_40101);
and U45457 (N_45457,N_40247,N_42559);
nor U45458 (N_45458,N_42076,N_44501);
nand U45459 (N_45459,N_40605,N_42191);
nor U45460 (N_45460,N_42919,N_44292);
xnor U45461 (N_45461,N_43471,N_41618);
or U45462 (N_45462,N_44536,N_41714);
nor U45463 (N_45463,N_42766,N_42633);
and U45464 (N_45464,N_42509,N_41518);
nand U45465 (N_45465,N_43768,N_42567);
xnor U45466 (N_45466,N_40374,N_41478);
nand U45467 (N_45467,N_44257,N_43798);
xnor U45468 (N_45468,N_42679,N_42189);
or U45469 (N_45469,N_40890,N_42916);
xnor U45470 (N_45470,N_44147,N_43324);
nand U45471 (N_45471,N_40189,N_40509);
nand U45472 (N_45472,N_40243,N_41661);
or U45473 (N_45473,N_41226,N_40894);
nor U45474 (N_45474,N_42124,N_43856);
xor U45475 (N_45475,N_42096,N_40685);
nor U45476 (N_45476,N_41778,N_41662);
nand U45477 (N_45477,N_42930,N_43286);
nor U45478 (N_45478,N_41104,N_42549);
and U45479 (N_45479,N_42804,N_40712);
nand U45480 (N_45480,N_40096,N_42526);
nor U45481 (N_45481,N_44682,N_42668);
or U45482 (N_45482,N_42415,N_40461);
xnor U45483 (N_45483,N_42159,N_43049);
nor U45484 (N_45484,N_41000,N_40217);
and U45485 (N_45485,N_43668,N_41019);
or U45486 (N_45486,N_40529,N_41441);
xnor U45487 (N_45487,N_44928,N_44223);
nor U45488 (N_45488,N_43510,N_44214);
or U45489 (N_45489,N_41608,N_44600);
or U45490 (N_45490,N_41269,N_44759);
and U45491 (N_45491,N_43462,N_44010);
xnor U45492 (N_45492,N_44709,N_43065);
xnor U45493 (N_45493,N_42255,N_41127);
nand U45494 (N_45494,N_44858,N_40015);
nand U45495 (N_45495,N_41982,N_41148);
or U45496 (N_45496,N_41731,N_41186);
nor U45497 (N_45497,N_40031,N_40865);
nor U45498 (N_45498,N_40287,N_44264);
xnor U45499 (N_45499,N_44857,N_44851);
nor U45500 (N_45500,N_41586,N_43733);
nand U45501 (N_45501,N_41234,N_41883);
xnor U45502 (N_45502,N_42290,N_43814);
and U45503 (N_45503,N_40880,N_44319);
xor U45504 (N_45504,N_42036,N_42967);
nor U45505 (N_45505,N_43960,N_44392);
and U45506 (N_45506,N_42828,N_42441);
or U45507 (N_45507,N_44984,N_40228);
nor U45508 (N_45508,N_43043,N_43287);
nor U45509 (N_45509,N_42678,N_40068);
or U45510 (N_45510,N_42349,N_41879);
xnor U45511 (N_45511,N_40339,N_44703);
xnor U45512 (N_45512,N_43758,N_41833);
and U45513 (N_45513,N_42138,N_40184);
xor U45514 (N_45514,N_42698,N_44345);
or U45515 (N_45515,N_42017,N_41033);
nor U45516 (N_45516,N_44605,N_42394);
nand U45517 (N_45517,N_43376,N_44301);
and U45518 (N_45518,N_41999,N_44516);
and U45519 (N_45519,N_40446,N_41110);
nand U45520 (N_45520,N_41169,N_41659);
and U45521 (N_45521,N_40039,N_40439);
nor U45522 (N_45522,N_42390,N_40746);
or U45523 (N_45523,N_44029,N_40486);
nand U45524 (N_45524,N_42133,N_43372);
or U45525 (N_45525,N_44000,N_41403);
and U45526 (N_45526,N_40183,N_44820);
xnor U45527 (N_45527,N_43604,N_41525);
or U45528 (N_45528,N_40025,N_42892);
xor U45529 (N_45529,N_43700,N_41768);
nor U45530 (N_45530,N_43142,N_44444);
and U45531 (N_45531,N_43872,N_42021);
nor U45532 (N_45532,N_42288,N_41144);
nor U45533 (N_45533,N_43983,N_44624);
and U45534 (N_45534,N_44355,N_42754);
nor U45535 (N_45535,N_42701,N_42624);
and U45536 (N_45536,N_42163,N_44906);
nor U45537 (N_45537,N_40688,N_44244);
xnor U45538 (N_45538,N_43708,N_43322);
nor U45539 (N_45539,N_43440,N_41238);
and U45540 (N_45540,N_40290,N_40330);
nand U45541 (N_45541,N_42373,N_42546);
or U45542 (N_45542,N_42564,N_40070);
nor U45543 (N_45543,N_44371,N_44695);
and U45544 (N_45544,N_43611,N_40500);
nand U45545 (N_45545,N_40118,N_41646);
or U45546 (N_45546,N_44053,N_44422);
or U45547 (N_45547,N_42157,N_43341);
nor U45548 (N_45548,N_44263,N_41430);
and U45549 (N_45549,N_42183,N_44901);
nor U45550 (N_45550,N_44314,N_44117);
or U45551 (N_45551,N_42114,N_40920);
nor U45552 (N_45552,N_41290,N_42294);
nand U45553 (N_45553,N_42536,N_42448);
and U45554 (N_45554,N_41458,N_44449);
and U45555 (N_45555,N_43740,N_41050);
nor U45556 (N_45556,N_41218,N_41655);
nor U45557 (N_45557,N_41656,N_41697);
and U45558 (N_45558,N_42012,N_44837);
nand U45559 (N_45559,N_42805,N_42186);
nand U45560 (N_45560,N_40755,N_43880);
or U45561 (N_45561,N_40737,N_40466);
or U45562 (N_45562,N_40506,N_43349);
xor U45563 (N_45563,N_44120,N_41850);
xnor U45564 (N_45564,N_43702,N_41594);
xor U45565 (N_45565,N_43777,N_40575);
or U45566 (N_45566,N_40013,N_44268);
or U45567 (N_45567,N_40503,N_40042);
nand U45568 (N_45568,N_43815,N_42139);
nor U45569 (N_45569,N_40222,N_44288);
nor U45570 (N_45570,N_40561,N_42200);
nand U45571 (N_45571,N_42613,N_41588);
xor U45572 (N_45572,N_44656,N_43041);
nor U45573 (N_45573,N_44097,N_44266);
or U45574 (N_45574,N_40538,N_43330);
nor U45575 (N_45575,N_42128,N_44731);
nor U45576 (N_45576,N_44243,N_41041);
nand U45577 (N_45577,N_43243,N_44207);
nand U45578 (N_45578,N_41300,N_40912);
nor U45579 (N_45579,N_44240,N_44561);
or U45580 (N_45580,N_40885,N_44360);
and U45581 (N_45581,N_44293,N_41956);
and U45582 (N_45582,N_40570,N_41579);
nor U45583 (N_45583,N_42105,N_40192);
nor U45584 (N_45584,N_42932,N_41388);
nor U45585 (N_45585,N_43812,N_41889);
nor U45586 (N_45586,N_40959,N_43268);
nor U45587 (N_45587,N_40510,N_43077);
nor U45588 (N_45588,N_40384,N_44458);
xnor U45589 (N_45589,N_41129,N_42855);
or U45590 (N_45590,N_41177,N_41601);
nor U45591 (N_45591,N_43238,N_41585);
xor U45592 (N_45592,N_41163,N_41053);
and U45593 (N_45593,N_40821,N_41884);
nor U45594 (N_45594,N_44471,N_43003);
nand U45595 (N_45595,N_40155,N_43042);
nor U45596 (N_45596,N_40280,N_42310);
nor U45597 (N_45597,N_44492,N_44166);
xor U45598 (N_45598,N_43239,N_40483);
nand U45599 (N_45599,N_40732,N_41320);
nand U45600 (N_45600,N_40162,N_42837);
or U45601 (N_45601,N_44946,N_41765);
and U45602 (N_45602,N_40493,N_44662);
or U45603 (N_45603,N_43646,N_42272);
xnor U45604 (N_45604,N_40332,N_44869);
nor U45605 (N_45605,N_44904,N_42355);
or U45606 (N_45606,N_40022,N_42980);
xnor U45607 (N_45607,N_42724,N_44842);
xnor U45608 (N_45608,N_42590,N_41707);
xnor U45609 (N_45609,N_44381,N_44844);
nand U45610 (N_45610,N_43558,N_40630);
nand U45611 (N_45611,N_44494,N_44530);
nand U45612 (N_45612,N_41825,N_43557);
nor U45613 (N_45613,N_43807,N_40451);
and U45614 (N_45614,N_44047,N_40881);
xnor U45615 (N_45615,N_44190,N_44989);
nor U45616 (N_45616,N_40181,N_41432);
nor U45617 (N_45617,N_40190,N_40966);
and U45618 (N_45618,N_43594,N_43548);
nand U45619 (N_45619,N_43300,N_41182);
or U45620 (N_45620,N_41359,N_43517);
and U45621 (N_45621,N_42070,N_43267);
nand U45622 (N_45622,N_43277,N_40811);
and U45623 (N_45623,N_41735,N_42815);
or U45624 (N_45624,N_42630,N_43846);
nand U45625 (N_45625,N_40014,N_42772);
or U45626 (N_45626,N_43824,N_41843);
xnor U45627 (N_45627,N_41477,N_42029);
or U45628 (N_45628,N_43881,N_40030);
and U45629 (N_45629,N_42753,N_44918);
nand U45630 (N_45630,N_44783,N_42706);
xor U45631 (N_45631,N_44821,N_40504);
xor U45632 (N_45632,N_41043,N_44852);
or U45633 (N_45633,N_40053,N_41361);
and U45634 (N_45634,N_44405,N_40347);
nor U45635 (N_45635,N_42154,N_42220);
and U45636 (N_45636,N_44337,N_40847);
xnor U45637 (N_45637,N_44853,N_43161);
xnor U45638 (N_45638,N_40580,N_42432);
nor U45639 (N_45639,N_43052,N_41237);
xor U45640 (N_45640,N_43884,N_41837);
or U45641 (N_45641,N_41682,N_42450);
xnor U45642 (N_45642,N_40227,N_40350);
nor U45643 (N_45643,N_43805,N_44539);
xnor U45644 (N_45644,N_42106,N_43848);
xnor U45645 (N_45645,N_42878,N_40065);
nor U45646 (N_45646,N_42923,N_40501);
and U45647 (N_45647,N_40695,N_43482);
nor U45648 (N_45648,N_40315,N_43075);
xor U45649 (N_45649,N_40253,N_42392);
xnor U45650 (N_45650,N_43621,N_43835);
and U45651 (N_45651,N_44457,N_40692);
or U45652 (N_45652,N_42674,N_40711);
or U45653 (N_45653,N_41831,N_41836);
nand U45654 (N_45654,N_44362,N_40839);
nor U45655 (N_45655,N_40595,N_41976);
xor U45656 (N_45656,N_43144,N_42770);
nand U45657 (N_45657,N_43140,N_41106);
or U45658 (N_45658,N_42482,N_44550);
and U45659 (N_45659,N_44890,N_43992);
nor U45660 (N_45660,N_41559,N_41729);
or U45661 (N_45661,N_40264,N_42602);
nor U45662 (N_45662,N_41456,N_42479);
and U45663 (N_45663,N_44939,N_43906);
xor U45664 (N_45664,N_43738,N_42296);
or U45665 (N_45665,N_43825,N_43729);
and U45666 (N_45666,N_43054,N_43578);
or U45667 (N_45667,N_40878,N_43965);
xor U45668 (N_45668,N_44913,N_40514);
or U45669 (N_45669,N_40485,N_43653);
nand U45670 (N_45670,N_44028,N_42049);
nand U45671 (N_45671,N_44886,N_44417);
nor U45672 (N_45672,N_44815,N_41059);
or U45673 (N_45673,N_44014,N_43177);
xnor U45674 (N_45674,N_42789,N_42655);
nand U45675 (N_45675,N_40479,N_41040);
or U45676 (N_45676,N_42524,N_44522);
or U45677 (N_45677,N_42347,N_41541);
nand U45678 (N_45678,N_43314,N_42460);
xor U45679 (N_45679,N_42629,N_42196);
nor U45680 (N_45680,N_44581,N_43069);
or U45681 (N_45681,N_40609,N_43469);
or U45682 (N_45682,N_41297,N_40623);
xor U45683 (N_45683,N_43219,N_42850);
or U45684 (N_45684,N_40049,N_42365);
or U45685 (N_45685,N_41597,N_42785);
and U45686 (N_45686,N_42758,N_44083);
or U45687 (N_45687,N_40795,N_41506);
or U45688 (N_45688,N_42035,N_41686);
and U45689 (N_45689,N_41338,N_40213);
and U45690 (N_45690,N_41716,N_40469);
nor U45691 (N_45691,N_44309,N_43873);
nand U45692 (N_45692,N_40979,N_42260);
xor U45693 (N_45693,N_43053,N_42889);
nand U45694 (N_45694,N_42516,N_40884);
and U45695 (N_45695,N_43596,N_43414);
or U45696 (N_45696,N_41788,N_44340);
and U45697 (N_45697,N_40858,N_43794);
or U45698 (N_45698,N_41351,N_43915);
nand U45699 (N_45699,N_43783,N_41174);
nor U45700 (N_45700,N_42267,N_44049);
xor U45701 (N_45701,N_44531,N_44775);
and U45702 (N_45702,N_41440,N_44977);
nand U45703 (N_45703,N_40789,N_42712);
or U45704 (N_45704,N_40522,N_44031);
nor U45705 (N_45705,N_41308,N_42503);
nand U45706 (N_45706,N_44740,N_40804);
xor U45707 (N_45707,N_41044,N_40862);
nand U45708 (N_45708,N_43281,N_40389);
xor U45709 (N_45709,N_41978,N_41994);
nand U45710 (N_45710,N_40079,N_43272);
xnor U45711 (N_45711,N_40288,N_40029);
nor U45712 (N_45712,N_42960,N_44102);
or U45713 (N_45713,N_42589,N_41598);
nor U45714 (N_45714,N_42733,N_41880);
or U45715 (N_45715,N_40662,N_44176);
and U45716 (N_45716,N_43860,N_40723);
or U45717 (N_45717,N_42321,N_44660);
and U45718 (N_45718,N_44919,N_43401);
nor U45719 (N_45719,N_43636,N_44850);
nor U45720 (N_45720,N_44959,N_43232);
xor U45721 (N_45721,N_43692,N_41079);
nor U45722 (N_45722,N_43310,N_41568);
and U45723 (N_45723,N_41841,N_40084);
xor U45724 (N_45724,N_41317,N_44463);
nor U45725 (N_45725,N_42771,N_40511);
nor U45726 (N_45726,N_44489,N_41803);
or U45727 (N_45727,N_41210,N_40622);
or U45728 (N_45728,N_42514,N_40552);
nand U45729 (N_45729,N_43732,N_44146);
xor U45730 (N_45730,N_42033,N_42002);
or U45731 (N_45731,N_43745,N_42250);
nor U45732 (N_45732,N_41462,N_44321);
xnor U45733 (N_45733,N_43034,N_40090);
nand U45734 (N_45734,N_40119,N_40691);
nand U45735 (N_45735,N_44803,N_40916);
and U45736 (N_45736,N_43936,N_43165);
or U45737 (N_45737,N_40729,N_43336);
nand U45738 (N_45738,N_44296,N_43789);
nor U45739 (N_45739,N_44218,N_40334);
or U45740 (N_45740,N_41986,N_44768);
xnor U45741 (N_45741,N_41284,N_42055);
and U45742 (N_45742,N_40618,N_40957);
nand U45743 (N_45743,N_43451,N_42155);
xor U45744 (N_45744,N_44391,N_44629);
and U45745 (N_45745,N_40867,N_42824);
nand U45746 (N_45746,N_44238,N_40415);
xnor U45747 (N_45747,N_40058,N_43910);
and U45748 (N_45748,N_43585,N_41060);
nor U45749 (N_45749,N_44808,N_44760);
nor U45750 (N_45750,N_41785,N_43658);
nand U45751 (N_45751,N_43271,N_41856);
and U45752 (N_45752,N_41315,N_42284);
and U45753 (N_45753,N_43173,N_44415);
xor U45754 (N_45754,N_40624,N_43524);
nand U45755 (N_45755,N_41064,N_42291);
or U45756 (N_45756,N_41719,N_40968);
or U45757 (N_45757,N_40061,N_41865);
nand U45758 (N_45758,N_41728,N_44487);
nor U45759 (N_45759,N_40036,N_42554);
nor U45760 (N_45760,N_44769,N_44315);
nand U45761 (N_45761,N_42901,N_41718);
or U45762 (N_45762,N_44370,N_42577);
or U45763 (N_45763,N_41005,N_43167);
and U45764 (N_45764,N_40731,N_43549);
xor U45765 (N_45765,N_42956,N_44452);
nor U45766 (N_45766,N_40046,N_40864);
xor U45767 (N_45767,N_42273,N_44763);
xor U45768 (N_45768,N_44098,N_42945);
nand U45769 (N_45769,N_43266,N_43756);
and U45770 (N_45770,N_41654,N_42561);
and U45771 (N_45771,N_42358,N_42654);
or U45772 (N_45772,N_40579,N_43461);
and U45773 (N_45773,N_41627,N_41709);
xnor U45774 (N_45774,N_44385,N_41221);
and U45775 (N_45775,N_40194,N_44270);
or U45776 (N_45776,N_43057,N_43381);
nand U45777 (N_45777,N_42870,N_42201);
nand U45778 (N_45778,N_40476,N_43079);
nor U45779 (N_45779,N_41796,N_40944);
and U45780 (N_45780,N_43363,N_42348);
or U45781 (N_45781,N_41394,N_42614);
nand U45782 (N_45782,N_44477,N_44088);
xor U45783 (N_45783,N_40733,N_41853);
nor U45784 (N_45784,N_44442,N_44254);
nand U45785 (N_45785,N_42715,N_40032);
nor U45786 (N_45786,N_42313,N_44090);
nor U45787 (N_45787,N_42027,N_43890);
nor U45788 (N_45788,N_41973,N_41648);
nand U45789 (N_45789,N_42821,N_41075);
nor U45790 (N_45790,N_44597,N_42090);
nor U45791 (N_45791,N_42739,N_40611);
nand U45792 (N_45792,N_40487,N_43945);
and U45793 (N_45793,N_41415,N_40470);
and U45794 (N_45794,N_43993,N_40974);
nand U45795 (N_45795,N_40127,N_40620);
or U45796 (N_45796,N_44182,N_43801);
nand U45797 (N_45797,N_40694,N_43511);
nand U45798 (N_45798,N_44999,N_44572);
xnor U45799 (N_45799,N_43100,N_40600);
xor U45800 (N_45800,N_44598,N_43785);
nor U45801 (N_45801,N_40766,N_43725);
nand U45802 (N_45802,N_43988,N_43033);
and U45803 (N_45803,N_42380,N_40482);
xor U45804 (N_45804,N_44893,N_44997);
and U45805 (N_45805,N_40062,N_42297);
nand U45806 (N_45806,N_42972,N_42326);
nand U45807 (N_45807,N_40199,N_44054);
nand U45808 (N_45808,N_42068,N_44861);
or U45809 (N_45809,N_41327,N_40241);
nor U45810 (N_45810,N_44801,N_44823);
or U45811 (N_45811,N_44236,N_43478);
nand U45812 (N_45812,N_44222,N_43070);
nand U45813 (N_45813,N_43942,N_43709);
nand U45814 (N_45814,N_43674,N_41509);
and U45815 (N_45815,N_43127,N_40560);
or U45816 (N_45816,N_42845,N_42465);
or U45817 (N_45817,N_42710,N_44654);
nor U45818 (N_45818,N_41082,N_41451);
xnor U45819 (N_45819,N_44103,N_40377);
or U45820 (N_45820,N_41393,N_42636);
and U45821 (N_45821,N_40134,N_43914);
nor U45822 (N_45822,N_40687,N_43778);
or U45823 (N_45823,N_42610,N_41013);
xor U45824 (N_45824,N_41145,N_41694);
and U45825 (N_45825,N_40019,N_42798);
nor U45826 (N_45826,N_44617,N_41278);
and U45827 (N_45827,N_42891,N_43251);
or U45828 (N_45828,N_40490,N_40064);
and U45829 (N_45829,N_41974,N_42520);
nand U45830 (N_45830,N_44326,N_40925);
or U45831 (N_45831,N_42399,N_40763);
xnor U45832 (N_45832,N_44127,N_41339);
xor U45833 (N_45833,N_42968,N_43245);
and U45834 (N_45834,N_41322,N_41436);
xnor U45835 (N_45835,N_43176,N_44547);
xnor U45836 (N_45836,N_44413,N_41468);
nand U45837 (N_45837,N_44610,N_40203);
and U45838 (N_45838,N_41142,N_40307);
nand U45839 (N_45839,N_44170,N_42030);
nor U45840 (N_45840,N_44072,N_41512);
xor U45841 (N_45841,N_42171,N_40933);
nor U45842 (N_45842,N_40211,N_40697);
xor U45843 (N_45843,N_40320,N_43155);
and U45844 (N_45844,N_42859,N_40775);
nand U45845 (N_45845,N_42261,N_44729);
nand U45846 (N_45846,N_41314,N_44178);
nor U45847 (N_45847,N_43015,N_43726);
nand U45848 (N_45848,N_40877,N_40086);
xor U45849 (N_45849,N_42899,N_41492);
and U45850 (N_45850,N_41885,N_42315);
xor U45851 (N_45851,N_44220,N_42341);
and U45852 (N_45852,N_41797,N_42406);
xnor U45853 (N_45853,N_41630,N_43445);
or U45854 (N_45854,N_44451,N_44670);
nor U45855 (N_45855,N_41103,N_41642);
xor U45856 (N_45856,N_41555,N_41349);
nand U45857 (N_45857,N_42907,N_41185);
nand U45858 (N_45858,N_40011,N_40863);
xnor U45859 (N_45859,N_43542,N_42807);
nand U45860 (N_45860,N_40423,N_43422);
nor U45861 (N_45861,N_42681,N_43437);
nand U45862 (N_45862,N_42799,N_44866);
xor U45863 (N_45863,N_40109,N_41674);
or U45864 (N_45864,N_43894,N_40220);
nor U45865 (N_45865,N_44265,N_42467);
xor U45866 (N_45866,N_44507,N_43722);
xnor U45867 (N_45867,N_40991,N_43293);
or U45868 (N_45868,N_42944,N_44189);
nor U45869 (N_45869,N_42345,N_44007);
nor U45870 (N_45870,N_42506,N_42120);
nand U45871 (N_45871,N_43374,N_42492);
nand U45872 (N_45872,N_41871,N_41294);
nand U45873 (N_45873,N_42072,N_41286);
nand U45874 (N_45874,N_42011,N_42266);
and U45875 (N_45875,N_43302,N_43185);
xor U45876 (N_45876,N_43295,N_44859);
or U45877 (N_45877,N_40057,N_40291);
and U45878 (N_45878,N_44105,N_40834);
nor U45879 (N_45879,N_40133,N_44593);
nor U45880 (N_45880,N_44017,N_41323);
nand U45881 (N_45881,N_41533,N_41918);
or U45882 (N_45882,N_40709,N_42340);
xor U45883 (N_45883,N_40785,N_42742);
nor U45884 (N_45884,N_41727,N_41126);
and U45885 (N_45885,N_43673,N_40588);
or U45886 (N_45886,N_40851,N_43236);
nor U45887 (N_45887,N_41287,N_44702);
nand U45888 (N_45888,N_42939,N_42023);
and U45889 (N_45889,N_44137,N_44568);
nor U45890 (N_45890,N_41398,N_42256);
nor U45891 (N_45891,N_40521,N_42557);
and U45892 (N_45892,N_41354,N_44732);
nor U45893 (N_45893,N_40960,N_40296);
nand U45894 (N_45894,N_43690,N_42042);
nor U45895 (N_45895,N_44046,N_40829);
nor U45896 (N_45896,N_41263,N_40554);
xor U45897 (N_45897,N_41445,N_42311);
nor U45898 (N_45898,N_43697,N_43624);
nand U45899 (N_45899,N_43811,N_44983);
nor U45900 (N_45900,N_43719,N_43138);
xor U45901 (N_45901,N_43623,N_41807);
or U45902 (N_45902,N_44205,N_40375);
and U45903 (N_45903,N_44816,N_41948);
or U45904 (N_45904,N_43967,N_43351);
and U45905 (N_45905,N_42490,N_41977);
and U45906 (N_45906,N_41413,N_44446);
nor U45907 (N_45907,N_43760,N_41216);
nor U45908 (N_45908,N_42869,N_41167);
xor U45909 (N_45909,N_42829,N_44650);
xor U45910 (N_45910,N_40449,N_42607);
and U45911 (N_45911,N_44394,N_42926);
nor U45912 (N_45912,N_40905,N_41204);
xor U45913 (N_45913,N_43908,N_44419);
nor U45914 (N_45914,N_43752,N_41066);
or U45915 (N_45915,N_40969,N_42044);
xnor U45916 (N_45916,N_41253,N_40652);
nor U45917 (N_45917,N_41134,N_40005);
xnor U45918 (N_45918,N_43474,N_42283);
or U45919 (N_45919,N_40995,N_40643);
nor U45920 (N_45920,N_40686,N_42883);
nand U45921 (N_45921,N_41181,N_41680);
xor U45922 (N_45922,N_43682,N_40672);
or U45923 (N_45923,N_40055,N_44231);
and U45924 (N_45924,N_40831,N_43717);
nor U45925 (N_45925,N_41158,N_41399);
nor U45926 (N_45926,N_41581,N_42849);
or U45927 (N_45927,N_42318,N_40900);
xnor U45928 (N_45928,N_41418,N_41254);
or U45929 (N_45929,N_43456,N_44064);
and U45930 (N_45930,N_42205,N_42496);
and U45931 (N_45931,N_44996,N_41876);
xor U45932 (N_45932,N_40781,N_44549);
and U45933 (N_45933,N_41898,N_42925);
and U45934 (N_45934,N_43597,N_40266);
nand U45935 (N_45935,N_40659,N_42116);
xnor U45936 (N_45936,N_41201,N_44425);
nor U45937 (N_45937,N_40654,N_42148);
and U45938 (N_45938,N_42217,N_41954);
and U45939 (N_45939,N_42560,N_44514);
nor U45940 (N_45940,N_44998,N_43953);
or U45941 (N_45941,N_44078,N_41805);
and U45942 (N_45942,N_40841,N_41721);
xor U45943 (N_45943,N_43379,N_42646);
nand U45944 (N_45944,N_43104,N_43095);
xor U45945 (N_45945,N_44154,N_40165);
or U45946 (N_45946,N_43430,N_42305);
xor U45947 (N_45947,N_42511,N_43220);
xnor U45948 (N_45948,N_44599,N_42709);
nor U45949 (N_45949,N_40767,N_40474);
and U45950 (N_45950,N_44106,N_40180);
and U45951 (N_45951,N_42439,N_40660);
nand U45952 (N_45952,N_43279,N_41443);
or U45953 (N_45953,N_41472,N_44184);
nor U45954 (N_45954,N_41081,N_44155);
nor U45955 (N_45955,N_42984,N_40388);
nor U45956 (N_45956,N_41893,N_41277);
or U45957 (N_45957,N_42173,N_42182);
and U45958 (N_45958,N_42239,N_42172);
nand U45959 (N_45959,N_44476,N_40512);
and U45960 (N_45960,N_42996,N_42623);
nand U45961 (N_45961,N_42696,N_40403);
xnor U45962 (N_45962,N_43570,N_42510);
nor U45963 (N_45963,N_41848,N_44881);
nand U45964 (N_45964,N_41582,N_44537);
nand U45965 (N_45965,N_43930,N_43290);
xor U45966 (N_45966,N_41078,N_40958);
nor U45967 (N_45967,N_43553,N_41529);
nor U45968 (N_45968,N_44590,N_41480);
nor U45969 (N_45969,N_41578,N_43479);
nor U45970 (N_45970,N_41623,N_41072);
xor U45971 (N_45971,N_43262,N_40909);
xnor U45972 (N_45972,N_41845,N_44036);
nand U45973 (N_45973,N_40255,N_42398);
nand U45974 (N_45974,N_43540,N_41971);
or U45975 (N_45975,N_44784,N_41776);
or U45976 (N_45976,N_40824,N_43345);
or U45977 (N_45977,N_41246,N_44573);
or U45978 (N_45978,N_43975,N_44896);
xor U45979 (N_45979,N_40530,N_42662);
xnor U45980 (N_45980,N_43285,N_43301);
xnor U45981 (N_45981,N_40661,N_42185);
nand U45982 (N_45982,N_40599,N_44651);
or U45983 (N_45983,N_43160,N_41653);
xnor U45984 (N_45984,N_43571,N_40589);
or U45985 (N_45985,N_41154,N_44490);
and U45986 (N_45986,N_42251,N_43154);
or U45987 (N_45987,N_40016,N_44726);
xnor U45988 (N_45988,N_41460,N_40621);
xor U45989 (N_45989,N_44070,N_44938);
xor U45990 (N_45990,N_41808,N_43854);
nor U45991 (N_45991,N_43020,N_42521);
and U45992 (N_45992,N_42693,N_44302);
or U45993 (N_45993,N_42985,N_43944);
and U45994 (N_45994,N_43150,N_40245);
nor U45995 (N_45995,N_42431,N_42880);
nand U45996 (N_45996,N_42469,N_40045);
nor U45997 (N_45997,N_40726,N_42178);
nand U45998 (N_45998,N_42816,N_40574);
nor U45999 (N_45999,N_43521,N_43561);
and U46000 (N_46000,N_44006,N_42014);
or U46001 (N_46001,N_42274,N_42876);
nor U46002 (N_46002,N_40604,N_41055);
and U46003 (N_46003,N_42048,N_42527);
xnor U46004 (N_46004,N_41090,N_44094);
nor U46005 (N_46005,N_42031,N_42952);
xnor U46006 (N_46006,N_43928,N_40323);
xor U46007 (N_46007,N_43937,N_43048);
nor U46008 (N_46008,N_43978,N_43940);
nand U46009 (N_46009,N_40442,N_44346);
nor U46010 (N_46010,N_42675,N_44962);
nand U46011 (N_46011,N_40810,N_40924);
and U46012 (N_46012,N_42418,N_43899);
nand U46013 (N_46013,N_41321,N_41717);
nand U46014 (N_46014,N_41704,N_43833);
xnor U46015 (N_46015,N_44899,N_44475);
and U46016 (N_46016,N_44791,N_41384);
and U46017 (N_46017,N_43348,N_41710);
nor U46018 (N_46018,N_41108,N_44735);
or U46019 (N_46019,N_40313,N_41583);
xnor U46020 (N_46020,N_41706,N_40870);
or U46021 (N_46021,N_40923,N_42241);
nand U46022 (N_46022,N_44164,N_42097);
nor U46023 (N_46023,N_42872,N_44461);
or U46024 (N_46024,N_44388,N_41685);
xnor U46025 (N_46025,N_44787,N_44535);
xnor U46026 (N_46026,N_41222,N_44310);
nand U46027 (N_46027,N_40328,N_44879);
nor U46028 (N_46028,N_40314,N_44711);
or U46029 (N_46029,N_43976,N_42056);
nor U46030 (N_46030,N_44895,N_42865);
nor U46031 (N_46031,N_40354,N_42019);
nor U46032 (N_46032,N_41135,N_41910);
and U46033 (N_46033,N_43948,N_44747);
nor U46034 (N_46034,N_44299,N_41924);
nor U46035 (N_46035,N_43568,N_40405);
and U46036 (N_46036,N_43269,N_41666);
nor U46037 (N_46037,N_41389,N_42728);
and U46038 (N_46038,N_43396,N_41753);
xor U46039 (N_46039,N_42152,N_41259);
xnor U46040 (N_46040,N_43109,N_40108);
and U46041 (N_46041,N_42263,N_43774);
nor U46042 (N_46042,N_42747,N_44150);
and U46043 (N_46043,N_42429,N_43891);
and U46044 (N_46044,N_44438,N_42057);
xor U46045 (N_46045,N_43855,N_44055);
xor U46046 (N_46046,N_44156,N_42998);
nor U46047 (N_46047,N_41048,N_41109);
nand U46048 (N_46048,N_42593,N_40088);
nand U46049 (N_46049,N_42866,N_40106);
or U46050 (N_46050,N_42216,N_40922);
and U46051 (N_46051,N_40225,N_41012);
nor U46052 (N_46052,N_40074,N_41427);
nand U46053 (N_46053,N_44584,N_41183);
and U46054 (N_46054,N_44870,N_41027);
and U46055 (N_46055,N_41820,N_41572);
and U46056 (N_46056,N_44756,N_44016);
and U46057 (N_46057,N_42325,N_44024);
xnor U46058 (N_46058,N_43090,N_43443);
nand U46059 (N_46059,N_43297,N_42246);
nand U46060 (N_46060,N_40343,N_41878);
or U46061 (N_46061,N_41113,N_44830);
and U46062 (N_46062,N_43742,N_43012);
nand U46063 (N_46063,N_42476,N_42721);
or U46064 (N_46064,N_44627,N_40472);
or U46065 (N_46065,N_40634,N_40902);
or U46066 (N_46066,N_43215,N_44505);
nand U46067 (N_46067,N_42018,N_44924);
xor U46068 (N_46068,N_42265,N_44707);
nand U46069 (N_46069,N_41136,N_42195);
and U46070 (N_46070,N_40450,N_42897);
nand U46071 (N_46071,N_43956,N_40010);
or U46072 (N_46072,N_41292,N_44911);
and U46073 (N_46073,N_44952,N_43900);
xor U46074 (N_46074,N_42995,N_42402);
nor U46075 (N_46075,N_42463,N_41929);
and U46076 (N_46076,N_43441,N_44144);
or U46077 (N_46077,N_40935,N_42639);
nand U46078 (N_46078,N_40835,N_44742);
and U46079 (N_46079,N_42238,N_43483);
nand U46080 (N_46080,N_43240,N_42391);
xor U46081 (N_46081,N_43409,N_44322);
nor U46082 (N_46082,N_40186,N_42622);
xor U46083 (N_46083,N_40113,N_41224);
or U46084 (N_46084,N_43565,N_43423);
nand U46085 (N_46085,N_42842,N_41074);
nand U46086 (N_46086,N_41225,N_44305);
xnor U46087 (N_46087,N_41313,N_43546);
and U46088 (N_46088,N_41330,N_42079);
nor U46089 (N_46089,N_41937,N_40235);
or U46090 (N_46090,N_44519,N_41464);
or U46091 (N_46091,N_43194,N_40673);
and U46092 (N_46092,N_40553,N_42396);
nor U46093 (N_46093,N_42280,N_42051);
xor U46094 (N_46094,N_43968,N_43917);
and U46095 (N_46095,N_42304,N_42722);
or U46096 (N_46096,N_40684,N_43605);
or U46097 (N_46097,N_42723,N_41592);
xor U46098 (N_46098,N_40901,N_44276);
xor U46099 (N_46099,N_41531,N_42991);
xnor U46100 (N_46100,N_43253,N_40699);
or U46101 (N_46101,N_42130,N_43676);
xor U46102 (N_46102,N_44386,N_41606);
xnor U46103 (N_46103,N_42584,N_41631);
nand U46104 (N_46104,N_43051,N_44679);
xnor U46105 (N_46105,N_43026,N_43368);
nand U46106 (N_46106,N_44133,N_42235);
nand U46107 (N_46107,N_43759,N_42906);
nand U46108 (N_46108,N_41758,N_44982);
xor U46109 (N_46109,N_42150,N_42194);
and U46110 (N_46110,N_40989,N_44750);
and U46111 (N_46111,N_43046,N_40550);
xnor U46112 (N_46112,N_43428,N_42209);
nand U46113 (N_46113,N_44272,N_41917);
nor U46114 (N_46114,N_42028,N_44863);
and U46115 (N_46115,N_44833,N_44559);
xor U46116 (N_46116,N_41471,N_42566);
or U46117 (N_46117,N_43645,N_42437);
xor U46118 (N_46118,N_44342,N_40597);
or U46119 (N_46119,N_41679,N_43679);
nor U46120 (N_46120,N_40891,N_43464);
or U46121 (N_46121,N_42981,N_41038);
nand U46122 (N_46122,N_42317,N_42671);
xor U46123 (N_46123,N_42203,N_44111);
or U46124 (N_46124,N_42295,N_43352);
xor U46125 (N_46125,N_44641,N_41084);
and U46126 (N_46126,N_41374,N_43870);
nor U46127 (N_46127,N_42505,N_41560);
nor U46128 (N_46128,N_40176,N_44874);
xnor U46129 (N_46129,N_40418,N_41966);
and U46130 (N_46130,N_42743,N_40392);
xnor U46131 (N_46131,N_40324,N_40986);
and U46132 (N_46132,N_44404,N_44588);
or U46133 (N_46133,N_42075,N_43073);
and U46134 (N_46134,N_44565,N_43991);
nor U46135 (N_46135,N_44712,N_41580);
xnor U46136 (N_46136,N_40537,N_43449);
nand U46137 (N_46137,N_43943,N_43211);
and U46138 (N_46138,N_44986,N_41267);
nor U46139 (N_46139,N_42101,N_40601);
or U46140 (N_46140,N_44758,N_44432);
nor U46141 (N_46141,N_40048,N_40738);
xor U46142 (N_46142,N_41485,N_42819);
nor U46143 (N_46143,N_44067,N_41897);
nor U46144 (N_46144,N_43713,N_44630);
and U46145 (N_46145,N_44470,N_40883);
and U46146 (N_46146,N_41137,N_44503);
and U46147 (N_46147,N_43084,N_42322);
or U46148 (N_46148,N_41741,N_42942);
nand U46149 (N_46149,N_44023,N_41490);
and U46150 (N_46150,N_43820,N_41764);
or U46151 (N_46151,N_42168,N_42811);
xnor U46152 (N_46152,N_42523,N_40703);
nor U46153 (N_46153,N_40581,N_43850);
nor U46154 (N_46154,N_41919,N_43828);
or U46155 (N_46155,N_44972,N_41140);
or U46156 (N_46156,N_40964,N_40428);
or U46157 (N_46157,N_40463,N_41699);
xnor U46158 (N_46158,N_42518,N_40816);
or U46159 (N_46159,N_44037,N_42388);
and U46160 (N_46160,N_43066,N_44400);
or U46161 (N_46161,N_41364,N_42335);
and U46162 (N_46162,N_41105,N_42222);
nand U46163 (N_46163,N_42069,N_41255);
or U46164 (N_46164,N_44981,N_43888);
nor U46165 (N_46165,N_40889,N_43191);
or U46166 (N_46166,N_43204,N_44797);
or U46167 (N_46167,N_44699,N_44878);
nand U46168 (N_46168,N_40259,N_41176);
nand U46169 (N_46169,N_41784,N_44382);
nand U46170 (N_46170,N_44230,N_43703);
and U46171 (N_46171,N_40730,N_40453);
nand U46172 (N_46172,N_41036,N_40223);
nand U46173 (N_46173,N_40613,N_44925);
xor U46174 (N_46174,N_41362,N_43183);
or U46175 (N_46175,N_44905,N_44733);
nand U46176 (N_46176,N_40135,N_43728);
nor U46177 (N_46177,N_42666,N_41065);
or U46178 (N_46178,N_40191,N_42665);
or U46179 (N_46179,N_40083,N_41769);
nor U46180 (N_46180,N_44722,N_41011);
or U46181 (N_46181,N_42606,N_40545);
xor U46182 (N_46182,N_41869,N_44119);
xnor U46183 (N_46183,N_44558,N_41713);
nor U46184 (N_46184,N_44145,N_40583);
xor U46185 (N_46185,N_43727,N_41067);
or U46186 (N_46186,N_44174,N_40519);
and U46187 (N_46187,N_40679,N_43652);
nand U46188 (N_46188,N_42010,N_44454);
or U46189 (N_46189,N_44502,N_43056);
nor U46190 (N_46190,N_40898,N_42594);
nor U46191 (N_46191,N_43791,N_40943);
xor U46192 (N_46192,N_43772,N_44757);
nand U46193 (N_46193,N_42428,N_42259);
or U46194 (N_46194,N_40882,N_44043);
nor U46195 (N_46195,N_43361,N_44557);
nand U46196 (N_46196,N_43196,N_43859);
and U46197 (N_46197,N_42161,N_42692);
and U46198 (N_46198,N_42861,N_42306);
nor U46199 (N_46199,N_43979,N_41431);
nand U46200 (N_46200,N_44751,N_41991);
nor U46201 (N_46201,N_41829,N_44187);
or U46202 (N_46202,N_42501,N_40207);
xnor U46203 (N_46203,N_41591,N_43724);
and U46204 (N_46204,N_41459,N_40793);
nand U46205 (N_46205,N_43331,N_40494);
nand U46206 (N_46206,N_44781,N_40866);
nand U46207 (N_46207,N_40215,N_44075);
xor U46208 (N_46208,N_43170,N_42645);
and U46209 (N_46209,N_41299,N_44794);
and U46210 (N_46210,N_43739,N_43050);
xnor U46211 (N_46211,N_40667,N_43083);
xor U46212 (N_46212,N_40639,N_43101);
nand U46213 (N_46213,N_42555,N_44985);
xnor U46214 (N_46214,N_44168,N_43877);
nand U46215 (N_46215,N_40520,N_43257);
xor U46216 (N_46216,N_43273,N_41120);
and U46217 (N_46217,N_40407,N_43447);
nor U46218 (N_46218,N_43001,N_44715);
nor U46219 (N_46219,N_41439,N_44954);
nand U46220 (N_46220,N_40353,N_44527);
xnor U46221 (N_46221,N_42519,N_43058);
and U46222 (N_46222,N_41605,N_41264);
xnor U46223 (N_46223,N_43971,N_40168);
xnor U46224 (N_46224,N_42750,N_41987);
nand U46225 (N_46225,N_44114,N_42131);
nand U46226 (N_46226,N_40233,N_41770);
nor U46227 (N_46227,N_40402,N_43581);
and U46228 (N_46228,N_41405,N_44614);
xor U46229 (N_46229,N_41175,N_41170);
and U46230 (N_46230,N_41190,N_43834);
and U46231 (N_46231,N_43353,N_43152);
nor U46232 (N_46232,N_41838,N_43878);
nor U46233 (N_46233,N_43514,N_43731);
nand U46234 (N_46234,N_43187,N_43435);
nand U46235 (N_46235,N_40269,N_44396);
xor U46236 (N_46236,N_41755,N_42440);
and U46237 (N_46237,N_43547,N_43309);
xor U46238 (N_46238,N_44149,N_43438);
and U46239 (N_46239,N_41007,N_44217);
xor U46240 (N_46240,N_42810,N_40856);
xor U46241 (N_46241,N_40204,N_40949);
or U46242 (N_46242,N_44433,N_40351);
xnor U46243 (N_46243,N_42601,N_40603);
nand U46244 (N_46244,N_43620,N_44420);
nand U46245 (N_46245,N_41213,N_43397);
and U46246 (N_46246,N_43896,N_43694);
nor U46247 (N_46247,N_40626,N_40727);
nor U46248 (N_46248,N_42731,N_41677);
or U46249 (N_46249,N_44317,N_42368);
or U46250 (N_46250,N_42497,N_43946);
and U46251 (N_46251,N_41798,N_40265);
nor U46252 (N_46252,N_42634,N_41887);
nand U46253 (N_46253,N_40533,N_42992);
nor U46254 (N_46254,N_43467,N_43446);
nor U46255 (N_46255,N_40998,N_41868);
nor U46256 (N_46256,N_44687,N_41111);
and U46257 (N_46257,N_44796,N_40765);
nor U46258 (N_46258,N_43898,N_43115);
and U46259 (N_46259,N_43529,N_43465);
or U46260 (N_46260,N_43642,N_43841);
nor U46261 (N_46261,N_41832,N_40292);
or U46262 (N_46262,N_42954,N_41786);
nor U46263 (N_46263,N_40172,N_40357);
nor U46264 (N_46264,N_40295,N_43139);
or U46265 (N_46265,N_41482,N_41209);
or U46266 (N_46266,N_43190,N_40417);
nand U46267 (N_46267,N_41307,N_42470);
and U46268 (N_46268,N_42381,N_44211);
nand U46269 (N_46269,N_44087,N_44173);
nor U46270 (N_46270,N_44948,N_40559);
or U46271 (N_46271,N_41383,N_42362);
or U46272 (N_46272,N_44073,N_40311);
or U46273 (N_46273,N_40774,N_40526);
xor U46274 (N_46274,N_43486,N_43537);
and U46275 (N_46275,N_42854,N_40741);
xnor U46276 (N_46276,N_40044,N_41881);
nor U46277 (N_46277,N_44466,N_40815);
and U46278 (N_46278,N_44621,N_42005);
xnor U46279 (N_46279,N_40082,N_41759);
and U46280 (N_46280,N_42966,N_44631);
nand U46281 (N_46281,N_40398,N_42207);
xor U46282 (N_46282,N_42735,N_44313);
or U46283 (N_46283,N_42911,N_40701);
nor U46284 (N_46284,N_43710,N_43572);
or U46285 (N_46285,N_40306,N_43498);
and U46286 (N_46286,N_42697,N_43315);
and U46287 (N_46287,N_41410,N_42094);
nand U46288 (N_46288,N_41687,N_41179);
nor U46289 (N_46289,N_44805,N_44022);
nor U46290 (N_46290,N_42813,N_43303);
or U46291 (N_46291,N_42860,N_41260);
and U46292 (N_46292,N_42779,N_44424);
nand U46293 (N_46293,N_44877,N_44818);
and U46294 (N_46294,N_42242,N_42672);
and U46295 (N_46295,N_41643,N_42543);
and U46296 (N_46296,N_41782,N_43477);
xor U46297 (N_46297,N_42598,N_42711);
nor U46298 (N_46298,N_41855,N_44101);
nor U46299 (N_46299,N_41184,N_43509);
and U46300 (N_46300,N_42065,N_42670);
or U46301 (N_46301,N_40047,N_41589);
xor U46302 (N_46302,N_42174,N_41031);
xor U46303 (N_46303,N_44026,N_40681);
nor U46304 (N_46304,N_44587,N_41289);
nand U46305 (N_46305,N_43664,N_42333);
nor U46306 (N_46306,N_40544,N_42699);
nand U46307 (N_46307,N_42374,N_43010);
and U46308 (N_46308,N_43011,N_43519);
and U46309 (N_46309,N_42331,N_40602);
nor U46310 (N_46310,N_44318,N_42713);
or U46311 (N_46311,N_40573,N_44718);
or U46312 (N_46312,N_42100,N_43686);
nor U46313 (N_46313,N_41196,N_40299);
xor U46314 (N_46314,N_41057,N_42480);
nor U46315 (N_46315,N_41610,N_43171);
nand U46316 (N_46316,N_42852,N_41899);
xnor U46317 (N_46317,N_44892,N_43885);
xor U46318 (N_46318,N_41567,N_44271);
xnor U46319 (N_46319,N_40249,N_44216);
nor U46320 (N_46320,N_42971,N_44261);
or U46321 (N_46321,N_41902,N_43258);
and U46322 (N_46322,N_42796,N_42382);
or U46323 (N_46323,N_42459,N_44316);
and U46324 (N_46324,N_41760,N_41626);
nand U46325 (N_46325,N_40275,N_40705);
or U46326 (N_46326,N_41273,N_40200);
and U46327 (N_46327,N_44967,N_44408);
xor U46328 (N_46328,N_43329,N_41021);
nor U46329 (N_46329,N_42354,N_44169);
or U46330 (N_46330,N_40739,N_44865);
or U46331 (N_46331,N_44934,N_43903);
xor U46332 (N_46332,N_43905,N_40076);
nand U46333 (N_46333,N_40495,N_44644);
or U46334 (N_46334,N_42993,N_43716);
xor U46335 (N_46335,N_41596,N_40516);
nand U46336 (N_46336,N_40489,N_43216);
xor U46337 (N_46337,N_42466,N_42659);
and U46338 (N_46338,N_42303,N_40366);
nor U46339 (N_46339,N_40107,N_42225);
nand U46340 (N_46340,N_44221,N_40231);
or U46341 (N_46341,N_43613,N_42292);
or U46342 (N_46342,N_42343,N_42077);
or U46343 (N_46343,N_41671,N_42301);
xor U46344 (N_46344,N_42663,N_43843);
nand U46345 (N_46345,N_41678,N_42660);
nand U46346 (N_46346,N_42219,N_41779);
nor U46347 (N_46347,N_42955,N_42425);
xor U46348 (N_46348,N_43755,N_44612);
and U46349 (N_46349,N_42389,N_44048);
or U46350 (N_46350,N_43563,N_41722);
nand U46351 (N_46351,N_43180,N_40360);
nand U46352 (N_46352,N_44942,N_44287);
or U46353 (N_46353,N_41625,N_42947);
nand U46354 (N_46354,N_42950,N_41703);
xnor U46355 (N_46355,N_40983,N_40708);
nor U46356 (N_46356,N_41452,N_40724);
or U46357 (N_46357,N_40505,N_41448);
and U46358 (N_46358,N_43858,N_43995);
or U46359 (N_46359,N_44209,N_44378);
and U46360 (N_46360,N_43543,N_42024);
nor U46361 (N_46361,N_41447,N_40582);
nand U46362 (N_46362,N_44620,N_41396);
xor U46363 (N_46363,N_41496,N_41957);
nor U46364 (N_46364,N_41593,N_42198);
nand U46365 (N_46365,N_41453,N_43707);
or U46366 (N_46366,N_40156,N_44701);
or U46367 (N_46367,N_42353,N_41203);
nor U46368 (N_46368,N_42573,N_42034);
nand U46369 (N_46369,N_41369,N_40773);
or U46370 (N_46370,N_44066,N_44074);
or U46371 (N_46371,N_44945,N_43924);
nor U46372 (N_46372,N_41150,N_41545);
and U46373 (N_46373,N_40499,N_42597);
xnor U46374 (N_46374,N_41188,N_44674);
and U46375 (N_46375,N_42300,N_43813);
xor U46376 (N_46376,N_40670,N_43318);
and U46377 (N_46377,N_41435,N_41131);
nand U46378 (N_46378,N_43845,N_41035);
nand U46379 (N_46379,N_44898,N_41009);
and U46380 (N_46380,N_44966,N_42797);
xor U46381 (N_46381,N_41965,N_44095);
nand U46382 (N_46382,N_44799,N_43291);
xor U46383 (N_46383,N_40614,N_40555);
or U46384 (N_46384,N_42451,N_41599);
xnor U46385 (N_46385,N_43385,N_41740);
nor U46386 (N_46386,N_41426,N_42786);
nand U46387 (N_46387,N_43022,N_44690);
nor U46388 (N_46388,N_40085,N_43489);
and U46389 (N_46389,N_40219,N_41097);
nor U46390 (N_46390,N_41356,N_44089);
and U46391 (N_46391,N_40696,N_41691);
or U46392 (N_46392,N_40822,N_40478);
and U46393 (N_46393,N_43627,N_42123);
nand U46394 (N_46394,N_44569,N_44172);
xor U46395 (N_46395,N_43701,N_41692);
or U46396 (N_46396,N_43819,N_44079);
nand U46397 (N_46397,N_41206,N_40818);
nor U46398 (N_46398,N_42895,N_43192);
and U46399 (N_46399,N_43912,N_41165);
and U46400 (N_46400,N_42908,N_42893);
nor U46401 (N_46401,N_42831,N_41830);
nor U46402 (N_46402,N_43453,N_43765);
nand U46403 (N_46403,N_41537,N_42063);
or U46404 (N_46404,N_43544,N_40843);
nand U46405 (N_46405,N_43332,N_40043);
nand U46406 (N_46406,N_40517,N_40467);
and U46407 (N_46407,N_43608,N_44845);
nand U46408 (N_46408,N_44658,N_44273);
xnor U46409 (N_46409,N_43328,N_44921);
and U46410 (N_46410,N_41874,N_42856);
and U46411 (N_46411,N_40171,N_43305);
xnor U46412 (N_46412,N_43312,N_44213);
xor U46413 (N_46413,N_43364,N_42784);
nor U46414 (N_46414,N_40363,N_40982);
and U46415 (N_46415,N_43954,N_41202);
xor U46416 (N_46416,N_44480,N_43651);
xor U46417 (N_46417,N_40651,N_43897);
xnor U46418 (N_46418,N_40987,N_40368);
xor U46419 (N_46419,N_41281,N_41017);
nand U46420 (N_46420,N_41073,N_44414);
and U46421 (N_46421,N_42489,N_40984);
or U46422 (N_46422,N_43319,N_42180);
and U46423 (N_46423,N_42167,N_43617);
nand U46424 (N_46424,N_44738,N_44810);
xor U46425 (N_46425,N_41676,N_40546);
nor U46426 (N_46426,N_43530,N_43600);
nand U46427 (N_46427,N_41619,N_40612);
or U46428 (N_46428,N_43767,N_44469);
nand U46429 (N_46429,N_40740,N_41343);
nand U46430 (N_46430,N_43695,N_40262);
xor U46431 (N_46431,N_41004,N_42531);
xor U46432 (N_46432,N_40799,N_40445);
nor U46433 (N_46433,N_43040,N_43508);
or U46434 (N_46434,N_40838,N_43468);
or U46435 (N_46435,N_40000,N_42965);
nand U46436 (N_46436,N_41600,N_43746);
and U46437 (N_46437,N_41495,N_40413);
or U46438 (N_46438,N_40430,N_41098);
xor U46439 (N_46439,N_41335,N_44364);
xnor U46440 (N_46440,N_40563,N_43822);
xor U46441 (N_46441,N_43134,N_41096);
xor U46442 (N_46442,N_42367,N_40426);
xnor U46443 (N_46443,N_43055,N_44746);
nor U46444 (N_46444,N_44376,N_42618);
and U46445 (N_46445,N_44499,N_43108);
xor U46446 (N_46446,N_44151,N_40980);
xor U46447 (N_46447,N_42160,N_42083);
nor U46448 (N_46448,N_43413,N_41861);
nand U46449 (N_46449,N_41139,N_43986);
xnor U46450 (N_46450,N_44917,N_40214);
nor U46451 (N_46451,N_41258,N_43750);
nand U46452 (N_46452,N_43832,N_40857);
xor U46453 (N_46453,N_41125,N_44575);
nand U46454 (N_46454,N_41528,N_40586);
or U46455 (N_46455,N_40256,N_41733);
or U46456 (N_46456,N_43844,N_43952);
xor U46457 (N_46457,N_43901,N_44467);
or U46458 (N_46458,N_40819,N_41904);
nand U46459 (N_46459,N_43094,N_44232);
or U46460 (N_46460,N_42153,N_44403);
nand U46461 (N_46461,N_43193,N_44464);
or U46462 (N_46462,N_43955,N_43661);
and U46463 (N_46463,N_44399,N_40026);
xnor U46464 (N_46464,N_42886,N_44991);
nand U46465 (N_46465,N_41342,N_44615);
nor U46466 (N_46466,N_43313,N_41675);
and U46467 (N_46467,N_44005,N_41658);
xnor U46468 (N_46468,N_41730,N_41566);
and U46469 (N_46469,N_40158,N_42102);
xnor U46470 (N_46470,N_41433,N_43504);
nand U46471 (N_46471,N_40441,N_43158);
nand U46472 (N_46472,N_44583,N_41244);
nand U46473 (N_46473,N_41516,N_41737);
nand U46474 (N_46474,N_42738,N_44606);
or U46475 (N_46475,N_40876,N_42725);
or U46476 (N_46476,N_41603,N_44260);
nor U46477 (N_46477,N_43023,N_44993);
and U46478 (N_46478,N_40872,N_42714);
nor U46479 (N_46479,N_40742,N_44980);
xor U46480 (N_46480,N_44486,N_44235);
nand U46481 (N_46481,N_42765,N_42099);
nand U46482 (N_46482,N_43842,N_43927);
xnor U46483 (N_46483,N_43321,N_43354);
xor U46484 (N_46484,N_44116,N_40632);
or U46485 (N_46485,N_40122,N_44284);
nor U46486 (N_46486,N_44592,N_44397);
and U46487 (N_46487,N_41293,N_40576);
or U46488 (N_46488,N_43250,N_44790);
xnor U46489 (N_46489,N_41953,N_42729);
or U46490 (N_46490,N_41964,N_42740);
and U46491 (N_46491,N_40749,N_40322);
nand U46492 (N_46492,N_43147,N_44909);
nor U46493 (N_46493,N_41301,N_43230);
nor U46494 (N_46494,N_43974,N_42227);
nand U46495 (N_46495,N_42458,N_44323);
xor U46496 (N_46496,N_44976,N_40647);
nand U46497 (N_46497,N_40527,N_40052);
xnor U46498 (N_46498,N_43523,N_41390);
or U46499 (N_46499,N_42581,N_42430);
or U46500 (N_46500,N_42045,N_42778);
xnor U46501 (N_46501,N_42839,N_40333);
and U46502 (N_46502,N_41872,N_41414);
nand U46503 (N_46503,N_42500,N_40024);
xor U46504 (N_46504,N_42085,N_42363);
xor U46505 (N_46505,N_44324,N_43629);
nand U46506 (N_46506,N_42825,N_41907);
nand U46507 (N_46507,N_43909,N_43865);
xnor U46508 (N_46508,N_43175,N_43887);
xnor U46509 (N_46509,N_42454,N_41166);
xor U46510 (N_46510,N_43072,N_42177);
or U46511 (N_46511,N_44636,N_40325);
or U46512 (N_46512,N_40381,N_41316);
or U46513 (N_46513,N_42727,N_40977);
or U46514 (N_46514,N_44491,N_41701);
xnor U46515 (N_46515,N_43769,N_42513);
nor U46516 (N_46516,N_41086,N_40258);
and U46517 (N_46517,N_43388,N_40908);
and U46518 (N_46518,N_41037,N_41251);
nand U46519 (N_46519,N_42419,N_40425);
or U46520 (N_46520,N_44258,N_43019);
or U46521 (N_46521,N_44714,N_41542);
or U46522 (N_46522,N_44493,N_41187);
or U46523 (N_46523,N_44136,N_40492);
and U46524 (N_46524,N_44576,N_40753);
and U46525 (N_46525,N_44002,N_41303);
and U46526 (N_46526,N_41232,N_43875);
or U46527 (N_46527,N_40091,N_40273);
nor U46528 (N_46528,N_40080,N_40592);
and U46529 (N_46529,N_44555,N_40852);
or U46530 (N_46530,N_44124,N_42461);
or U46531 (N_46531,N_42551,N_41866);
or U46532 (N_46532,N_41404,N_41510);
nand U46533 (N_46533,N_40281,N_40382);
nand U46534 (N_46534,N_43063,N_43972);
xor U46535 (N_46535,N_40077,N_43635);
nor U46536 (N_46536,N_43644,N_44669);
or U46537 (N_46537,N_44657,N_41551);
nor U46538 (N_46538,N_40994,N_42078);
and U46539 (N_46539,N_40678,N_44027);
xor U46540 (N_46540,N_43463,N_42299);
or U46541 (N_46541,N_40840,N_43089);
xnor U46542 (N_46542,N_40348,N_42346);
xnor U46543 (N_46543,N_43799,N_41305);
nor U46544 (N_46544,N_43017,N_41916);
nand U46545 (N_46545,N_44882,N_42486);
nand U46546 (N_46546,N_40498,N_44785);
xor U46547 (N_46547,N_44498,N_40416);
nand U46548 (N_46548,N_44889,N_42734);
and U46549 (N_46549,N_40319,N_41521);
nor U46550 (N_46550,N_43913,N_43797);
and U46551 (N_46551,N_44013,N_43616);
and U46552 (N_46552,N_40792,N_44226);
nand U46553 (N_46553,N_44304,N_42179);
nand U46554 (N_46554,N_40157,N_43660);
or U46555 (N_46555,N_42000,N_44688);
nor U46556 (N_46556,N_44247,N_40081);
and U46557 (N_46557,N_43375,N_43958);
nand U46558 (N_46558,N_43178,N_41862);
xor U46559 (N_46559,N_41192,N_42328);
nor U46560 (N_46560,N_41357,N_40020);
xor U46561 (N_46561,N_44229,N_40182);
and U46562 (N_46562,N_44672,N_43199);
xnor U46563 (N_46563,N_44407,N_41844);
nand U46564 (N_46564,N_40018,N_41377);
nand U46565 (N_46565,N_44050,N_44786);
nand U46566 (N_46566,N_44227,N_43254);
and U46567 (N_46567,N_42477,N_40800);
and U46568 (N_46568,N_40196,N_43403);
nand U46569 (N_46569,N_42934,N_40812);
nor U46570 (N_46570,N_42937,N_42694);
and U46571 (N_46571,N_44455,N_43718);
and U46572 (N_46572,N_42763,N_43217);
xor U46573 (N_46573,N_43876,N_43085);
or U46574 (N_46574,N_41607,N_42234);
and U46575 (N_46575,N_40254,N_43551);
or U46576 (N_46576,N_41891,N_44193);
xor U46577 (N_46577,N_41667,N_44363);
and U46578 (N_46578,N_41672,N_44995);
xnor U46579 (N_46579,N_40164,N_41754);
xnor U46580 (N_46580,N_43174,N_41198);
nor U46581 (N_46581,N_41346,N_42764);
nor U46582 (N_46582,N_42487,N_43151);
nand U46583 (N_46583,N_42539,N_40502);
or U46584 (N_46584,N_40683,N_44586);
nor U46585 (N_46585,N_43086,N_41030);
nor U46586 (N_46586,N_40515,N_41025);
nand U46587 (N_46587,N_42188,N_44607);
or U46588 (N_46588,N_41847,N_44186);
and U46589 (N_46589,N_40237,N_41245);
or U46590 (N_46590,N_44675,N_42071);
xor U46591 (N_46591,N_42621,N_43421);
xor U46592 (N_46592,N_42768,N_44525);
xor U46593 (N_46593,N_40153,N_43810);
or U46594 (N_46594,N_44884,N_42652);
xnor U46595 (N_46595,N_42039,N_44113);
nor U46596 (N_46596,N_44684,N_44336);
nor U46597 (N_46597,N_43829,N_44128);
nand U46598 (N_46598,N_40886,N_44574);
nor U46599 (N_46599,N_42868,N_44246);
and U46600 (N_46600,N_42129,N_44406);
or U46601 (N_46601,N_44800,N_41270);
nor U46602 (N_46602,N_42884,N_42224);
nor U46603 (N_46603,N_42316,N_44430);
or U46604 (N_46604,N_41941,N_44250);
and U46605 (N_46605,N_40309,N_43080);
nand U46606 (N_46606,N_44204,N_40706);
xor U46607 (N_46607,N_41429,N_43961);
and U46608 (N_46608,N_42164,N_44663);
nand U46609 (N_46609,N_43534,N_43663);
and U46610 (N_46610,N_44766,N_41194);
nor U46611 (N_46611,N_43383,N_40126);
nor U46612 (N_46612,N_41851,N_42062);
and U46613 (N_46613,N_44135,N_40455);
nand U46614 (N_46614,N_42197,N_42122);
or U46615 (N_46615,N_44744,N_41223);
or U46616 (N_46616,N_40903,N_43335);
nor U46617 (N_46617,N_42963,N_44447);
or U46618 (N_46618,N_40644,N_41751);
or U46619 (N_46619,N_41524,N_43786);
and U46620 (N_46620,N_41858,N_43771);
or U46621 (N_46621,N_42957,N_44035);
xnor U46622 (N_46622,N_41602,N_40286);
xor U46623 (N_46623,N_41763,N_43111);
nor U46624 (N_46624,N_44873,N_41673);
or U46625 (N_46625,N_43064,N_43795);
xor U46626 (N_46626,N_42104,N_40762);
xor U46627 (N_46627,N_42091,N_42499);
nand U46628 (N_46628,N_43977,N_42943);
nor U46629 (N_46629,N_44202,N_40587);
nor U46630 (N_46630,N_44395,N_42110);
nor U46631 (N_46631,N_42424,N_43356);
and U46632 (N_46632,N_40823,N_44839);
and U46633 (N_46633,N_43246,N_41552);
or U46634 (N_46634,N_41752,N_43763);
nor U46635 (N_46635,N_41392,N_42426);
or U46636 (N_46636,N_42690,N_40028);
xor U46637 (N_46637,N_41747,N_41886);
nand U46638 (N_46638,N_43340,N_40051);
nand U46639 (N_46639,N_40110,N_42232);
and U46640 (N_46640,N_44795,N_42537);
nand U46641 (N_46641,N_43037,N_40132);
nor U46642 (N_46642,N_44914,N_41890);
xnor U46643 (N_46643,N_41068,N_41498);
xor U46644 (N_46644,N_44678,N_40997);
and U46645 (N_46645,N_40471,N_44131);
nor U46646 (N_46646,N_41499,N_44704);
and U46647 (N_46647,N_40780,N_40782);
and U46648 (N_46648,N_40369,N_41535);
nand U46649 (N_46649,N_44979,N_44625);
or U46650 (N_46650,N_41272,N_44134);
nand U46651 (N_46651,N_40117,N_44479);
nand U46652 (N_46652,N_41748,N_40226);
xor U46653 (N_46653,N_44521,N_43227);
nor U46654 (N_46654,N_43130,N_40754);
or U46655 (N_46655,N_40400,N_40633);
nor U46656 (N_46656,N_40209,N_43404);
nand U46657 (N_46657,N_42050,N_43689);
and U46658 (N_46658,N_40069,N_40063);
nand U46659 (N_46659,N_41810,N_40568);
or U46660 (N_46660,N_42132,N_42669);
and U46661 (N_46661,N_40202,N_41641);
nor U46662 (N_46662,N_41888,N_41979);
and U46663 (N_46663,N_43586,N_40414);
xnor U46664 (N_46664,N_40097,N_40756);
nand U46665 (N_46665,N_43639,N_44421);
or U46666 (N_46666,N_44428,N_41636);
or U46667 (N_46667,N_44328,N_43864);
xor U46668 (N_46668,N_42783,N_44951);
nand U46669 (N_46669,N_41028,N_43241);
or U46670 (N_46670,N_43584,N_43867);
or U46671 (N_46671,N_43355,N_40635);
xnor U46672 (N_46672,N_41094,N_41422);
nor U46673 (N_46673,N_42020,N_41138);
or U46674 (N_46674,N_43889,N_40596);
or U46675 (N_46675,N_40386,N_42640);
nand U46676 (N_46676,N_44125,N_44379);
nand U46677 (N_46677,N_42535,N_41995);
or U46678 (N_46678,N_44957,N_44804);
and U46679 (N_46679,N_43599,N_44443);
or U46680 (N_46680,N_41712,N_44673);
nor U46681 (N_46681,N_40874,N_41493);
nand U46682 (N_46682,N_44613,N_40569);
or U46683 (N_46683,N_43895,N_43744);
nand U46684 (N_46684,N_41554,N_42790);
and U46685 (N_46685,N_40721,N_40297);
nor U46686 (N_46686,N_43494,N_41921);
xnor U46687 (N_46687,N_41319,N_40625);
and U46688 (N_46688,N_40606,N_43417);
nor U46689 (N_46689,N_44012,N_40720);
or U46690 (N_46690,N_44748,N_41927);
or U46691 (N_46691,N_42596,N_43839);
xor U46692 (N_46692,N_44059,N_43816);
xnor U46693 (N_46693,N_40465,N_42206);
and U46694 (N_46694,N_44167,N_40947);
nor U46695 (N_46695,N_44626,N_44025);
nor U46696 (N_46696,N_44633,N_43626);
or U46697 (N_46697,N_44496,N_43793);
or U46698 (N_46698,N_43030,N_44883);
or U46699 (N_46699,N_43392,N_42767);
and U46700 (N_46700,N_41230,N_43933);
nand U46701 (N_46701,N_40807,N_42761);
xor U46702 (N_46702,N_42084,N_43893);
and U46703 (N_46703,N_42386,N_41514);
or U46704 (N_46704,N_41233,N_41945);
nand U46705 (N_46705,N_44374,N_41197);
xnor U46706 (N_46706,N_42832,N_44096);
xor U46707 (N_46707,N_41080,N_44061);
xor U46708 (N_46708,N_44383,N_41479);
nor U46709 (N_46709,N_44868,N_40779);
and U46710 (N_46710,N_41421,N_42835);
nor U46711 (N_46711,N_40524,N_40170);
or U46712 (N_46712,N_44312,N_41018);
nor U46713 (N_46713,N_44664,N_44161);
or U46714 (N_46714,N_41947,N_43044);
nand U46715 (N_46715,N_40921,N_44398);
or U46716 (N_46716,N_44283,N_41611);
nand U46717 (N_46717,N_43460,N_40270);
and U46718 (N_46718,N_41123,N_41280);
nand U46719 (N_46719,N_40408,N_40361);
xnor U46720 (N_46720,N_44445,N_40564);
nand U46721 (N_46721,N_43146,N_44648);
nand U46722 (N_46722,N_40617,N_44774);
nand U46723 (N_46723,N_44267,N_43485);
nand U46724 (N_46724,N_42620,N_44373);
or U46725 (N_46725,N_44042,N_43110);
xnor U46726 (N_46726,N_40385,N_40710);
or U46727 (N_46727,N_43032,N_42377);
or U46728 (N_46728,N_42556,N_42879);
nand U46729 (N_46729,N_44907,N_43067);
nand U46730 (N_46730,N_43770,N_40594);
xor U46731 (N_46731,N_43741,N_44779);
nor U46732 (N_46732,N_41100,N_41877);
or U46733 (N_46733,N_40342,N_41895);
or U46734 (N_46734,N_44341,N_44020);
nand U46735 (N_46735,N_41959,N_40768);
nor U46736 (N_46736,N_42563,N_44563);
nand U46737 (N_46737,N_41483,N_44691);
nor U46738 (N_46738,N_40038,N_42254);
nor U46739 (N_46739,N_42611,N_41943);
and U46740 (N_46740,N_44380,N_41536);
xor U46741 (N_46741,N_44777,N_44367);
nand U46742 (N_46742,N_44065,N_43304);
nor U46743 (N_46743,N_44291,N_43200);
xnor U46744 (N_46744,N_41955,N_42619);
xor U46745 (N_46745,N_43087,N_41857);
and U46746 (N_46746,N_43436,N_40826);
and U46747 (N_46747,N_44091,N_40393);
xor U46748 (N_46748,N_44409,N_42446);
xnor U46749 (N_46749,N_42922,N_43882);
and U46750 (N_46750,N_44402,N_41664);
nand U46751 (N_46751,N_42411,N_44534);
xnor U46752 (N_46752,N_43280,N_44215);
or U46753 (N_46753,N_42289,N_43380);
xor U46754 (N_46754,N_42881,N_44541);
and U46755 (N_46755,N_42776,N_40387);
nor U46756 (N_46756,N_41570,N_40716);
xor U46757 (N_46757,N_43091,N_40271);
or U46758 (N_46758,N_44423,N_41708);
and U46759 (N_46759,N_40578,N_40682);
nor U46760 (N_46760,N_42410,N_41262);
or U46761 (N_46761,N_42994,N_40151);
and U46762 (N_46762,N_43696,N_40367);
or U46763 (N_46763,N_41749,N_43068);
or U46764 (N_46764,N_43323,N_40457);
and U46765 (N_46765,N_42240,N_43205);
nor U46766 (N_46766,N_44344,N_41515);
xor U46767 (N_46767,N_40996,N_44856);
or U46768 (N_46768,N_42151,N_43133);
nand U46769 (N_46769,N_44092,N_44947);
xnor U46770 (N_46770,N_44311,N_42871);
nand U46771 (N_46771,N_44778,N_41283);
and U46772 (N_46772,N_43939,N_42649);
nor U46773 (N_46773,N_42404,N_42915);
nor U46774 (N_46774,N_43754,N_43047);
and U46775 (N_46775,N_42329,N_42434);
nor U46776 (N_46776,N_41783,N_43221);
xnor U46777 (N_46777,N_40744,N_40776);
and U46778 (N_46778,N_40674,N_41352);
xnor U46779 (N_46779,N_44110,N_41215);
nor U46780 (N_46780,N_40842,N_43590);
and U46781 (N_46781,N_44677,N_40525);
xor U46782 (N_46782,N_41826,N_40198);
or U46783 (N_46783,N_41276,N_43796);
xnor U46784 (N_46784,N_42204,N_42759);
or U46785 (N_46785,N_40999,N_42286);
xnor U46786 (N_46786,N_44365,N_41756);
nor U46787 (N_46787,N_44871,N_41576);
or U46788 (N_46788,N_44929,N_42111);
or U46789 (N_46789,N_44249,N_42047);
and U46790 (N_46790,N_42591,N_41634);
nor U46791 (N_46791,N_43775,N_43823);
or U46792 (N_46792,N_44776,N_43809);
nor U46793 (N_46793,N_43527,N_40904);
nor U46794 (N_46794,N_43920,N_44434);
nor U46795 (N_46795,N_43102,N_41457);
and U46796 (N_46796,N_43255,N_41669);
nor U46797 (N_46797,N_40748,N_40137);
and U46798 (N_46798,N_44148,N_43941);
or U46799 (N_46799,N_40454,N_43386);
nor U46800 (N_46800,N_40836,N_42628);
nand U46801 (N_46801,N_43669,N_40671);
xor U46802 (N_46802,N_41333,N_42522);
or U46803 (N_46803,N_42940,N_42732);
or U46804 (N_46804,N_44831,N_44281);
nand U46805 (N_46805,N_41644,N_43536);
nor U46806 (N_46806,N_40365,N_41114);
nand U46807 (N_46807,N_40475,N_43208);
and U46808 (N_46808,N_42857,N_41839);
nand U46809 (N_46809,N_42395,N_43950);
or U46810 (N_46810,N_42202,N_41989);
nor U46811 (N_46811,N_44372,N_40649);
or U46812 (N_46812,N_41911,N_42338);
and U46813 (N_46813,N_42145,N_41010);
nor U46814 (N_46814,N_42826,N_42975);
nor U46815 (N_46815,N_41220,N_41616);
nor U46816 (N_46816,N_43210,N_41620);
or U46817 (N_46817,N_41928,N_44659);
and U46818 (N_46818,N_43346,N_44668);
or U46819 (N_46819,N_40540,N_43490);
nor U46820 (N_46820,N_41794,N_40395);
nand U46821 (N_46821,N_40373,N_41780);
and U46822 (N_46822,N_41615,N_40528);
and U46823 (N_46823,N_44835,N_41909);
nand U46824 (N_46824,N_44642,N_43874);
or U46825 (N_46825,N_41992,N_43427);
and U46826 (N_46826,N_42874,N_44646);
or U46827 (N_46827,N_44843,N_41023);
nand U46828 (N_46828,N_40246,N_42782);
xnor U46829 (N_46829,N_40962,N_43806);
nor U46830 (N_46830,N_43871,N_42427);
nor U46831 (N_46831,N_43264,N_44275);
nor U46832 (N_46832,N_43448,N_44933);
nor U46833 (N_46833,N_43276,N_41700);
and U46834 (N_46834,N_43393,N_43520);
and U46835 (N_46835,N_43560,N_42371);
and U46836 (N_46836,N_41736,N_40507);
or U46837 (N_46837,N_43420,N_43800);
xnor U46838 (N_46838,N_44352,N_44294);
and U46839 (N_46839,N_43792,N_42689);
nor U46840 (N_46840,N_41501,N_41523);
nor U46841 (N_46841,N_40293,N_41119);
nor U46842 (N_46842,N_42147,N_41302);
or U46843 (N_46843,N_41199,N_40460);
nor U46844 (N_46844,N_41311,N_42230);
or U46845 (N_46845,N_43195,N_40640);
nor U46846 (N_46846,N_40432,N_42896);
xor U46847 (N_46847,N_44676,N_40556);
xor U46848 (N_46848,N_44393,N_42127);
or U46849 (N_46849,N_40188,N_44792);
nand U46850 (N_46850,N_42264,N_41951);
nor U46851 (N_46851,N_43292,N_41143);
and U46852 (N_46852,N_41132,N_42920);
and U46853 (N_46853,N_40978,N_41032);
nand U46854 (N_46854,N_41497,N_43132);
or U46855 (N_46855,N_43145,N_40397);
xnor U46856 (N_46856,N_43931,N_44132);
nor U46857 (N_46857,N_40917,N_43099);
or U46858 (N_46858,N_41228,N_44591);
and U46859 (N_46859,N_42271,N_42387);
and U46860 (N_46860,N_42774,N_43879);
and U46861 (N_46861,N_43861,N_40436);
nor U46862 (N_46862,N_43721,N_40169);
nand U46863 (N_46863,N_41162,N_42757);
nor U46864 (N_46864,N_43723,N_43378);
nor U46865 (N_46865,N_41975,N_42726);
nand U46866 (N_46866,N_40844,N_44689);
xor U46867 (N_46867,N_43907,N_44462);
nand U46868 (N_46868,N_43734,N_40973);
nand U46869 (N_46869,N_43705,N_42656);
xor U46870 (N_46870,N_44003,N_44034);
xnor U46871 (N_46871,N_40658,N_44915);
nor U46872 (N_46872,N_43189,N_40798);
nand U46873 (N_46873,N_43862,N_43031);
and U46874 (N_46874,N_44930,N_44828);
and U46875 (N_46875,N_41936,N_44375);
xor U46876 (N_46876,N_43559,N_43360);
or U46877 (N_46877,N_43076,N_43788);
nor U46878 (N_46878,N_40571,N_43244);
and U46879 (N_46879,N_43934,N_41274);
and U46880 (N_46880,N_40242,N_44518);
nand U46881 (N_46881,N_40893,N_43455);
or U46882 (N_46882,N_40805,N_43289);
xor U46883 (N_46883,N_40300,N_40910);
xor U46884 (N_46884,N_42095,N_43625);
and U46885 (N_46885,N_44062,N_43357);
nand U46886 (N_46886,N_43592,N_40089);
nand U46887 (N_46887,N_42417,N_42755);
nor U46888 (N_46888,N_40914,N_44068);
nor U46889 (N_46889,N_43764,N_43579);
or U46890 (N_46890,N_43619,N_42688);
or U46891 (N_46891,N_42054,N_44495);
or U46892 (N_46892,N_42058,N_40926);
and U46893 (N_46893,N_43516,N_40642);
xnor U46894 (N_46894,N_41363,N_42978);
xor U46895 (N_46895,N_40832,N_41049);
and U46896 (N_46896,N_42882,N_42846);
or U46897 (N_46897,N_42990,N_41365);
nor U46898 (N_46898,N_44497,N_41475);
and U46899 (N_46899,N_44885,N_43373);
nand U46900 (N_46900,N_40873,N_40913);
or U46901 (N_46901,N_44252,N_44960);
or U46902 (N_46902,N_40409,N_44153);
and U46903 (N_46903,N_43265,N_43962);
nand U46904 (N_46904,N_42040,N_41200);
and U46905 (N_46905,N_44234,N_40937);
and U46906 (N_46906,N_42661,N_42760);
nor U46907 (N_46907,N_42862,N_42548);
and U46908 (N_46908,N_42003,N_43141);
nand U46909 (N_46909,N_40675,N_42237);
or U46910 (N_46910,N_40034,N_42061);
nand U46911 (N_46911,N_44694,N_43198);
nor U46912 (N_46912,N_41530,N_42407);
and U46913 (N_46913,N_44579,N_43614);
nor U46914 (N_46914,N_43493,N_42082);
nor U46915 (N_46915,N_40378,N_43743);
nor U46916 (N_46916,N_40566,N_41663);
and U46917 (N_46917,N_41939,N_42532);
xor U46918 (N_46918,N_43153,N_40212);
and U46919 (N_46919,N_42379,N_42393);
xor U46920 (N_46920,N_41629,N_42447);
or U46921 (N_46921,N_44943,N_41093);
or U46922 (N_46922,N_42320,N_42803);
or U46923 (N_46923,N_40953,N_41574);
and U46924 (N_46924,N_42929,N_40906);
nand U46925 (N_46925,N_43612,N_44077);
or U46926 (N_46926,N_44538,N_40534);
and U46927 (N_46927,N_41901,N_42800);
or U46928 (N_46928,N_42026,N_43439);
nand U46929 (N_46929,N_44039,N_42616);
nand U46930 (N_46930,N_42695,N_40854);
nand U46931 (N_46931,N_44634,N_41252);
xnor U46932 (N_46932,N_43698,N_42702);
and U46933 (N_46933,N_40140,N_41195);
and U46934 (N_46934,N_43821,N_41117);
xnor U46935 (N_46935,N_41029,N_43433);
and U46936 (N_46936,N_44198,N_43402);
nand U46937 (N_46937,N_42921,N_43782);
nor U46938 (N_46938,N_42383,N_42412);
xor U46939 (N_46939,N_44069,N_41022);
or U46940 (N_46940,N_40892,N_41517);
nand U46941 (N_46941,N_43412,N_41257);
nand U46942 (N_46942,N_40796,N_43078);
xor U46943 (N_46943,N_41217,N_42457);
and U46944 (N_46944,N_42493,N_42933);
nand U46945 (N_46945,N_41757,N_42323);
xor U46946 (N_46946,N_40808,N_44616);
or U46947 (N_46947,N_43603,N_43164);
and U46948 (N_46948,N_40352,N_41380);
and U46949 (N_46949,N_44233,N_40849);
nor U46950 (N_46950,N_43256,N_40121);
and U46951 (N_46951,N_44570,N_42806);
xnor U46952 (N_46952,N_43317,N_43112);
or U46953 (N_46953,N_44339,N_41212);
xnor U46954 (N_46954,N_42707,N_42221);
or U46955 (N_46955,N_42979,N_40802);
nor U46956 (N_46956,N_44152,N_41061);
and U46957 (N_46957,N_40828,N_41077);
or U46958 (N_46958,N_40035,N_41504);
and U46959 (N_46959,N_41373,N_44814);
and U46960 (N_46960,N_42736,N_42833);
and U46961 (N_46961,N_42408,N_42385);
or U46962 (N_46962,N_42319,N_42905);
and U46963 (N_46963,N_42498,N_43659);
nand U46964 (N_46964,N_44228,N_41761);
or U46965 (N_46965,N_41657,N_41915);
nor U46966 (N_46966,N_41101,N_44051);
nor U46967 (N_46967,N_40860,N_43326);
or U46968 (N_46968,N_44282,N_41130);
and U46969 (N_46969,N_41325,N_44932);
xor U46970 (N_46970,N_42015,N_40440);
or U46971 (N_46971,N_42352,N_40433);
nand U46972 (N_46972,N_42464,N_40115);
or U46973 (N_46973,N_41604,N_42875);
nor U46974 (N_46974,N_40473,N_41505);
nor U46975 (N_46975,N_44194,N_44510);
nand U46976 (N_46976,N_41540,N_43117);
nand U46977 (N_46977,N_43014,N_41324);
nand U46978 (N_46978,N_41345,N_43333);
or U46979 (N_46979,N_40656,N_43122);
nand U46980 (N_46980,N_40637,N_44320);
or U46981 (N_46981,N_41548,N_43555);
nor U46982 (N_46982,N_44546,N_41474);
or U46983 (N_46983,N_41690,N_41424);
or U46984 (N_46984,N_43487,N_40941);
and U46985 (N_46985,N_44793,N_43545);
nand U46986 (N_46986,N_44720,N_41569);
nor U46987 (N_46987,N_43234,N_41705);
xnor U46988 (N_46988,N_43480,N_43120);
nor U46989 (N_46989,N_43634,N_43021);
nand U46990 (N_46990,N_44509,N_42684);
or U46991 (N_46991,N_43973,N_44836);
xor U46992 (N_46992,N_43787,N_43550);
nor U46993 (N_46993,N_42676,N_41099);
nor U46994 (N_46994,N_40421,N_40655);
nor U46995 (N_46995,N_40002,N_41732);
or U46996 (N_46996,N_40939,N_40855);
xor U46997 (N_46997,N_43492,N_42169);
or U46998 (N_46998,N_41795,N_41546);
xnor U46999 (N_46999,N_41790,N_43362);
and U47000 (N_47000,N_42949,N_42983);
nor U47001 (N_47001,N_40830,N_41042);
or U47002 (N_47002,N_44594,N_42969);
or U47003 (N_47003,N_42285,N_42416);
nand U47004 (N_47004,N_43515,N_42038);
nor U47005 (N_47005,N_40073,N_43016);
nor U47006 (N_47006,N_41122,N_41846);
xor U47007 (N_47007,N_41818,N_43773);
nand U47008 (N_47008,N_43680,N_41376);
and U47009 (N_47009,N_42032,N_42887);
nand U47010 (N_47010,N_40801,N_44453);
nor U47011 (N_47011,N_43918,N_41026);
nand U47012 (N_47012,N_41819,N_43949);
or U47013 (N_47013,N_44327,N_44019);
nor U47014 (N_47014,N_44021,N_42603);
and U47015 (N_47015,N_44179,N_43886);
nand U47016 (N_47016,N_42350,N_44511);
or U47017 (N_47017,N_40009,N_40337);
or U47018 (N_47018,N_44686,N_42121);
or U47019 (N_47019,N_40718,N_42877);
nand U47020 (N_47020,N_43588,N_42400);
and U47021 (N_47021,N_41817,N_40447);
and U47022 (N_47022,N_41635,N_44224);
nor U47023 (N_47023,N_42626,N_41577);
xnor U47024 (N_47024,N_42530,N_41696);
and U47025 (N_47025,N_40144,N_41695);
or U47026 (N_47026,N_42718,N_41141);
nor U47027 (N_47027,N_41903,N_42749);
xnor U47028 (N_47028,N_44286,N_41425);
or U47029 (N_47029,N_41968,N_44551);
xnor U47030 (N_47030,N_41913,N_42841);
nor U47031 (N_47031,N_40918,N_40456);
and U47032 (N_47032,N_40547,N_40129);
nor U47033 (N_47033,N_41961,N_40304);
xnor U47034 (N_47034,N_44544,N_42176);
nor U47035 (N_47035,N_41133,N_42445);
xnor U47036 (N_47036,N_42612,N_44195);
xor U47037 (N_47037,N_43135,N_44528);
and U47038 (N_47038,N_44513,N_43088);
or U47039 (N_47039,N_40396,N_41489);
or U47040 (N_47040,N_41952,N_44708);
xnor U47041 (N_47041,N_43136,N_43580);
or U47042 (N_47042,N_40784,N_44772);
and U47043 (N_47043,N_43502,N_41336);
nor U47044 (N_47044,N_40942,N_43671);
nand U47045 (N_47045,N_43123,N_44807);
or U47046 (N_47046,N_43826,N_41056);
and U47047 (N_47047,N_42820,N_40174);
nand U47048 (N_47048,N_41573,N_42231);
xnor U47049 (N_47049,N_42682,N_44693);
nand U47050 (N_47050,N_41526,N_42781);
nand U47051 (N_47051,N_44749,N_40584);
xor U47052 (N_47052,N_43424,N_42109);
nand U47053 (N_47053,N_42673,N_41395);
nand U47054 (N_47054,N_43476,N_42166);
nor U47055 (N_47055,N_43804,N_41513);
or U47056 (N_47056,N_42838,N_40380);
nor U47057 (N_47057,N_43377,N_41935);
xor U47058 (N_47058,N_43450,N_42686);
nand U47059 (N_47059,N_43124,N_42780);
and U47060 (N_47060,N_40282,N_41118);
nand U47061 (N_47061,N_42962,N_44773);
xor U47062 (N_47062,N_41054,N_41809);
and U47063 (N_47063,N_44560,N_44832);
or U47064 (N_47064,N_43554,N_41488);
or U47065 (N_47065,N_41411,N_41683);
and U47066 (N_47066,N_42745,N_40251);
xor U47067 (N_47067,N_42423,N_42245);
nor U47068 (N_47068,N_44206,N_44554);
xnor U47069 (N_47069,N_41341,N_44175);
or U47070 (N_47070,N_41091,N_43159);
nor U47071 (N_47071,N_42575,N_42422);
and U47072 (N_47072,N_44104,N_44596);
nor U47073 (N_47073,N_41107,N_40990);
or U47074 (N_47074,N_41326,N_42547);
nor U47075 (N_47075,N_43316,N_42442);
nand U47076 (N_47076,N_40954,N_43637);
and U47077 (N_47077,N_44298,N_43387);
and U47078 (N_47078,N_44564,N_42236);
and U47079 (N_47079,N_42253,N_44082);
and U47080 (N_47080,N_41651,N_41062);
nor U47081 (N_47081,N_41235,N_40145);
and U47082 (N_47082,N_44358,N_41371);
or U47083 (N_47083,N_41407,N_41151);
nor U47084 (N_47084,N_40236,N_44130);
or U47085 (N_47085,N_43684,N_40551);
and U47086 (N_47086,N_44508,N_41164);
xnor U47087 (N_47087,N_40193,N_42823);
nand U47088 (N_47088,N_43532,N_40177);
nor U47089 (N_47089,N_42212,N_40645);
or U47090 (N_47090,N_44920,N_42327);
and U47091 (N_47091,N_42588,N_42961);
nand U47092 (N_47092,N_44717,N_42409);
and U47093 (N_47093,N_42507,N_41894);
xnor U47094 (N_47094,N_42599,N_41434);
and U47095 (N_47095,N_41645,N_44349);
and U47096 (N_47096,N_41372,N_43751);
xnor U47097 (N_47097,N_43209,N_43263);
nand U47098 (N_47098,N_42570,N_43481);
and U47099 (N_47099,N_41933,N_43577);
nor U47100 (N_47100,N_40136,N_43618);
nor U47101 (N_47101,N_42494,N_40059);
and U47102 (N_47102,N_42009,N_44356);
nor U47103 (N_47103,N_41538,N_43444);
nor U47104 (N_47104,N_44841,N_44813);
or U47105 (N_47105,N_44623,N_43761);
xnor U47106 (N_47106,N_40173,N_42022);
nor U47107 (N_47107,N_42081,N_41534);
xnor U47108 (N_47108,N_41312,N_40666);
nor U47109 (N_47109,N_41484,N_41008);
and U47110 (N_47110,N_41446,N_42277);
and U47111 (N_47111,N_41527,N_40707);
nand U47112 (N_47112,N_41665,N_44666);
xnor U47113 (N_47113,N_44771,N_42931);
nand U47114 (N_47114,N_44926,N_44332);
and U47115 (N_47115,N_42787,N_40809);
or U47116 (N_47116,N_41614,N_41930);
nand U47117 (N_47117,N_43038,N_41002);
or U47118 (N_47118,N_42973,N_40316);
or U47119 (N_47119,N_40690,N_41285);
nor U47120 (N_47120,N_40747,N_44440);
nand U47121 (N_47121,N_41612,N_41632);
xor U47122 (N_47122,N_42641,N_42858);
and U47123 (N_47123,N_43390,N_40646);
or U47124 (N_47124,N_40331,N_42964);
xor U47125 (N_47125,N_42545,N_43018);
xnor U47126 (N_47126,N_42276,N_44552);
or U47127 (N_47127,N_44937,N_44225);
nand U47128 (N_47128,N_41811,N_44084);
and U47129 (N_47129,N_42912,N_42337);
nor U47130 (N_47130,N_43987,N_44459);
xnor U47131 (N_47131,N_42357,N_40120);
or U47132 (N_47132,N_43488,N_40210);
and U47133 (N_47133,N_44330,N_43587);
xor U47134 (N_47134,N_41219,N_44923);
nor U47135 (N_47135,N_42092,N_44721);
and U47136 (N_47136,N_44115,N_43306);
xnor U47137 (N_47137,N_41849,N_42118);
xnor U47138 (N_47138,N_41972,N_43513);
and U47139 (N_47139,N_41670,N_42775);
and U47140 (N_47140,N_40895,N_42059);
nand U47141 (N_47141,N_42087,N_44809);
xnor U47142 (N_47142,N_40783,N_40462);
nor U47143 (N_47143,N_41932,N_40060);
and U47144 (N_47144,N_44426,N_44274);
nand U47145 (N_47145,N_44239,N_43610);
and U47146 (N_47146,N_41942,N_41271);
and U47147 (N_47147,N_42066,N_41329);
nand U47148 (N_47148,N_43996,N_40240);
xnor U47149 (N_47149,N_41402,N_42948);
nor U47150 (N_47150,N_42664,N_41382);
or U47151 (N_47151,N_40598,N_42935);
xnor U47152 (N_47152,N_44603,N_41821);
nand U47153 (N_47153,N_42436,N_42089);
or U47154 (N_47154,N_42976,N_43512);
or U47155 (N_47155,N_43935,N_43929);
xor U47156 (N_47156,N_44706,N_43157);
and U47157 (N_47157,N_43681,N_41814);
or U47158 (N_47158,N_40631,N_44652);
or U47159 (N_47159,N_41738,N_40041);
or U47160 (N_47160,N_42836,N_43113);
nor U47161 (N_47161,N_42853,N_44825);
or U47162 (N_47162,N_42986,N_41306);
xnor U47163 (N_47163,N_44080,N_41931);
or U47164 (N_47164,N_44992,N_42953);
xor U47165 (N_47165,N_42013,N_43222);
and U47166 (N_47166,N_40437,N_44765);
or U47167 (N_47167,N_43648,N_43218);
and U47168 (N_47168,N_44743,N_41985);
nand U47169 (N_47169,N_43672,N_42226);
xnor U47170 (N_47170,N_40033,N_42043);
nand U47171 (N_47171,N_44255,N_42175);
nand U47172 (N_47172,N_40244,N_43932);
xor U47173 (N_47173,N_43994,N_44955);
xnor U47174 (N_47174,N_44969,N_40665);
or U47175 (N_47175,N_40294,N_40279);
nor U47176 (N_47176,N_41875,N_41702);
and U47177 (N_47177,N_41980,N_44739);
nor U47178 (N_47178,N_41532,N_41789);
or U47179 (N_47179,N_42864,N_42214);
nor U47180 (N_47180,N_43299,N_42142);
nand U47181 (N_47181,N_40302,N_41406);
xnor U47182 (N_47182,N_41449,N_44609);
or U47183 (N_47183,N_40007,N_41774);
nor U47184 (N_47184,N_41824,N_44334);
nand U47185 (N_47185,N_41539,N_40143);
xor U47186 (N_47186,N_40272,N_42369);
nor U47187 (N_47187,N_43473,N_43505);
or U47188 (N_47188,N_40850,N_43963);
xor U47189 (N_47189,N_41121,N_43749);
xor U47190 (N_47190,N_43062,N_42818);
nand U47191 (N_47191,N_44968,N_40484);
and U47192 (N_47192,N_41428,N_42478);
xor U47193 (N_47193,N_43863,N_42651);
xnor U47194 (N_47194,N_44004,N_44472);
or U47195 (N_47195,N_41173,N_40743);
or U47196 (N_47196,N_43252,N_41417);
xor U47197 (N_47197,N_44798,N_43235);
nand U47198 (N_47198,N_44734,N_40761);
and U47199 (N_47199,N_44725,N_40329);
nand U47200 (N_47200,N_43184,N_44056);
xor U47201 (N_47201,N_40340,N_44410);
xor U47202 (N_47202,N_42403,N_43006);
nor U47203 (N_47203,N_40303,N_40438);
or U47204 (N_47204,N_43989,N_41340);
or U47205 (N_47205,N_41016,N_43762);
xor U47206 (N_47206,N_40327,N_44122);
xnor U47207 (N_47207,N_43410,N_41873);
nor U47208 (N_47208,N_42135,N_41564);
nand U47209 (N_47209,N_42571,N_42098);
or U47210 (N_47210,N_42293,N_41387);
nor U47211 (N_47211,N_40496,N_42579);
nand U47212 (N_47212,N_43539,N_44199);
nand U47213 (N_47213,N_41249,N_40558);
and U47214 (N_47214,N_44237,N_42488);
nand U47215 (N_47215,N_43964,N_41473);
or U47216 (N_47216,N_41912,N_43203);
and U47217 (N_47217,N_43666,N_42809);
xnor U47218 (N_47218,N_43849,N_44058);
and U47219 (N_47219,N_40722,N_41052);
xnor U47220 (N_47220,N_43593,N_44506);
or U47221 (N_47221,N_43985,N_41265);
nor U47222 (N_47222,N_42847,N_43307);
nor U47223 (N_47223,N_42741,N_41787);
xnor U47224 (N_47224,N_43131,N_43311);
or U47225 (N_47225,N_44517,N_42508);
and U47226 (N_47226,N_43434,N_40208);
nand U47227 (N_47227,N_43980,N_40464);
xor U47228 (N_47228,N_40758,N_44908);
xor U47229 (N_47229,N_41998,N_41547);
or U47230 (N_47230,N_43715,N_40928);
nand U47231 (N_47231,N_41698,N_40146);
or U47232 (N_47232,N_43093,N_41243);
xor U47233 (N_47233,N_40187,N_40346);
xor U47234 (N_47234,N_42576,N_42149);
xor U47235 (N_47235,N_44782,N_42339);
or U47236 (N_47236,N_43156,N_40163);
and U47237 (N_47237,N_44011,N_41720);
and U47238 (N_47238,N_40557,N_40907);
xor U47239 (N_47239,N_40427,N_42903);
or U47240 (N_47240,N_40845,N_44242);
nor U47241 (N_47241,N_43071,N_41227);
or U47242 (N_47242,N_44671,N_42914);
or U47243 (N_47243,N_43233,N_41295);
and U47244 (N_47244,N_41353,N_41001);
nor U47245 (N_47245,N_41020,N_42541);
nor U47246 (N_47246,N_42004,N_42269);
or U47247 (N_47247,N_43921,N_43650);
xor U47248 (N_47248,N_42314,N_41102);
or U47249 (N_47249,N_42814,N_43475);
or U47250 (N_47250,N_44157,N_44542);
or U47251 (N_47251,N_41859,N_42769);
nor U47252 (N_47252,N_42016,N_42433);
nor U47253 (N_47253,N_43406,N_42683);
or U47254 (N_47254,N_43706,N_42720);
xor U47255 (N_47255,N_41864,N_40650);
and U47256 (N_47256,N_42444,N_40817);
xor U47257 (N_47257,N_43840,N_42443);
nand U47258 (N_47258,N_42605,N_44532);
nand U47259 (N_47259,N_44653,N_42647);
nor U47260 (N_47260,N_41804,N_41438);
nand U47261 (N_47261,N_40138,N_41375);
nand U47262 (N_47262,N_41958,N_44331);
and U47263 (N_47263,N_42604,N_40276);
or U47264 (N_47264,N_40147,N_43432);
and U47265 (N_47265,N_44755,N_43442);
and U47266 (N_47266,N_44008,N_44834);
and U47267 (N_47267,N_43182,N_42917);
nor U47268 (N_47268,N_44523,N_40535);
nand U47269 (N_47269,N_43541,N_41247);
nand U47270 (N_47270,N_41511,N_41609);
nor U47271 (N_47271,N_43970,N_40218);
xor U47272 (N_47272,N_44308,N_41058);
or U47273 (N_47273,N_44500,N_40179);
or U47274 (N_47274,N_44303,N_44162);
or U47275 (N_47275,N_40871,N_44484);
nand U47276 (N_47276,N_44745,N_41854);
nand U47277 (N_47277,N_41178,N_44343);
xor U47278 (N_47278,N_41638,N_42658);
nand U47279 (N_47279,N_44441,N_41556);
nand U47280 (N_47280,N_41486,N_41725);
nand U47281 (N_47281,N_40803,N_43857);
nand U47282 (N_47282,N_44123,N_41095);
or U47283 (N_47283,N_40607,N_44941);
xnor U47284 (N_47284,N_44988,N_44512);
nand U47285 (N_47285,N_40230,N_40689);
and U47286 (N_47286,N_43163,N_43092);
xnor U47287 (N_47287,N_42913,N_44515);
nor U47288 (N_47288,N_41550,N_43143);
or U47289 (N_47289,N_43415,N_44578);
and U47290 (N_47290,N_41034,N_40394);
nand U47291 (N_47291,N_40794,N_42125);
nor U47292 (N_47292,N_44698,N_43564);
xor U47293 (N_47293,N_44724,N_40736);
xor U47294 (N_47294,N_44961,N_44811);
or U47295 (N_47295,N_43827,N_43365);
and U47296 (N_47296,N_44460,N_44990);
nor U47297 (N_47297,N_44770,N_42708);
or U47298 (N_47298,N_40565,N_43591);
nor U47299 (N_47299,N_42553,N_40411);
xnor U47300 (N_47300,N_43916,N_40948);
nand U47301 (N_47301,N_41900,N_42126);
or U47302 (N_47302,N_40362,N_42667);
nor U47303 (N_47303,N_43116,N_44788);
or U47304 (N_47304,N_44611,N_44141);
nor U47305 (N_47305,N_42282,N_41309);
and U47306 (N_47306,N_42455,N_40508);
or U47307 (N_47307,N_42863,N_43957);
and U47308 (N_47308,N_43904,N_44953);
nor U47309 (N_47309,N_40221,N_42067);
and U47310 (N_47310,N_40399,N_40814);
or U47311 (N_47311,N_43172,N_44812);
or U47312 (N_47312,N_40497,N_41637);
xor U47313 (N_47313,N_41128,N_44057);
nor U47314 (N_47314,N_44958,N_41003);
nand U47315 (N_47315,N_43615,N_44256);
nor U47316 (N_47316,N_42843,N_44819);
xor U47317 (N_47317,N_42474,N_40006);
nand U47318 (N_47318,N_43803,N_41870);
nand U47319 (N_47319,N_41863,N_40359);
xnor U47320 (N_47320,N_40869,N_44197);
xor U47321 (N_47321,N_43675,N_41867);
xnor U47322 (N_47322,N_44181,N_44548);
or U47323 (N_47323,N_40356,N_40628);
and U47324 (N_47324,N_42788,N_40372);
nor U47325 (N_47325,N_44140,N_40616);
or U47326 (N_47326,N_41724,N_40468);
and U47327 (N_47327,N_40663,N_43677);
nor U47328 (N_47328,N_44353,N_43342);
or U47329 (N_47329,N_41112,N_41711);
and U47330 (N_47330,N_43008,N_41766);
xor U47331 (N_47331,N_43426,N_44894);
and U47332 (N_47332,N_41923,N_41494);
nand U47333 (N_47333,N_44086,N_40206);
nand U47334 (N_47334,N_40422,N_42107);
nand U47335 (N_47335,N_41613,N_44142);
or U47336 (N_47336,N_44713,N_41157);
nor U47337 (N_47337,N_42909,N_40648);
nor U47338 (N_47338,N_42184,N_40585);
nor U47339 (N_47339,N_43035,N_40148);
xor U47340 (N_47340,N_44994,N_41633);
nor U47341 (N_47341,N_43391,N_43278);
nand U47342 (N_47342,N_42552,N_42928);
or U47343 (N_47343,N_43753,N_41189);
nor U47344 (N_47344,N_44640,N_42491);
xnor U47345 (N_47345,N_43206,N_41248);
and U47346 (N_47346,N_43730,N_41575);
xnor U47347 (N_47347,N_41241,N_43128);
nor U47348 (N_47348,N_42756,N_43097);
and U47349 (N_47349,N_43633,N_43552);
xnor U47350 (N_47350,N_40424,N_44887);
xor U47351 (N_47351,N_42215,N_42158);
or U47352 (N_47352,N_41466,N_41520);
or U47353 (N_47353,N_43308,N_42378);
and U47354 (N_47354,N_44354,N_43169);
nor U47355 (N_47355,N_43892,N_44964);
xor U47356 (N_47356,N_40102,N_44876);
nand U47357 (N_47357,N_43337,N_40092);
and U47358 (N_47358,N_44100,N_44723);
xor U47359 (N_47359,N_42275,N_44439);
or U47360 (N_47360,N_40326,N_41331);
xor U47361 (N_47361,N_44601,N_41275);
nor U47362 (N_47362,N_40130,N_43247);
nor U47363 (N_47363,N_42356,N_44840);
xnor U47364 (N_47364,N_44936,N_43643);
nor U47365 (N_47365,N_44705,N_40125);
nand U47366 (N_47366,N_42737,N_44848);
and U47367 (N_47367,N_42938,N_43622);
nand U47368 (N_47368,N_40410,N_44667);
xor U47369 (N_47369,N_43607,N_42974);
and U47370 (N_47370,N_43296,N_40930);
xor U47371 (N_47371,N_41256,N_41834);
nor U47372 (N_47372,N_44602,N_44520);
nor U47373 (N_47373,N_42244,N_42525);
xor U47374 (N_47374,N_41236,N_40629);
nand U47375 (N_47375,N_43229,N_41156);
nor U47376 (N_47376,N_42542,N_41926);
nand U47377 (N_47377,N_41799,N_41491);
xor U47378 (N_47378,N_40071,N_40412);
and U47379 (N_47379,N_42324,N_42533);
and U47380 (N_47380,N_42140,N_41640);
nor U47381 (N_47381,N_44900,N_44295);
nand U47382 (N_47382,N_41563,N_43036);
nor U47383 (N_47383,N_43847,N_41822);
or U47384 (N_47384,N_41350,N_43609);
and U47385 (N_47385,N_42888,N_40680);
nand U47386 (N_47386,N_41562,N_40719);
xnor U47387 (N_47387,N_41171,N_41983);
or U47388 (N_47388,N_44121,N_41076);
xor U47389 (N_47389,N_41358,N_43407);
xor U47390 (N_47390,N_42719,N_43869);
nor U47391 (N_47391,N_42006,N_44143);
or U47392 (N_47392,N_44912,N_41565);
or U47393 (N_47393,N_40657,N_41996);
and U47394 (N_47394,N_41242,N_40541);
nand U47395 (N_47395,N_40548,N_40103);
nor U47396 (N_47396,N_41519,N_43261);
or U47397 (N_47397,N_44401,N_41960);
nor U47398 (N_47398,N_42228,N_42648);
nand U47399 (N_47399,N_42366,N_44916);
or U47400 (N_47400,N_42703,N_42529);
xnor U47401 (N_47401,N_43004,N_41069);
nand U47402 (N_47402,N_43213,N_44661);
nor U47403 (N_47403,N_41416,N_44566);
xor U47404 (N_47404,N_40274,N_40788);
nor U47405 (N_47405,N_44730,N_43237);
nor U47406 (N_47406,N_40641,N_43259);
and U47407 (N_47407,N_42258,N_44824);
or U47408 (N_47408,N_42582,N_41772);
nor U47409 (N_47409,N_44543,N_43923);
xor U47410 (N_47410,N_43503,N_42951);
or U47411 (N_47411,N_42453,N_40111);
xor U47412 (N_47412,N_43997,N_42192);
or U47413 (N_47413,N_42074,N_40488);
or U47414 (N_47414,N_44468,N_40285);
and U47415 (N_47415,N_44350,N_43419);
nor U47416 (N_47416,N_41650,N_40406);
nand U47417 (N_47417,N_41860,N_40178);
or U47418 (N_47418,N_40931,N_43114);
nand U47419 (N_47419,N_42405,N_40777);
or U47420 (N_47420,N_43649,N_43028);
nand U47421 (N_47421,N_44949,N_42376);
xnor U47422 (N_47422,N_43499,N_44427);
nor U47423 (N_47423,N_40542,N_44040);
or U47424 (N_47424,N_42344,N_41047);
nor U47425 (N_47425,N_44888,N_42307);
nand U47426 (N_47426,N_43107,N_43223);
nand U47427 (N_47427,N_43685,N_40017);
and U47428 (N_47428,N_40956,N_44553);
and U47429 (N_47429,N_43000,N_42119);
or U47430 (N_47430,N_44780,N_40250);
or U47431 (N_47431,N_44196,N_40355);
and U47432 (N_47432,N_42211,N_43606);
nand U47433 (N_47433,N_43212,N_42281);
nand U47434 (N_47434,N_41908,N_40750);
nor U47435 (N_47435,N_41006,N_42890);
nor U47436 (N_47436,N_41823,N_41745);
nor U47437 (N_47437,N_42867,N_43583);
nor U47438 (N_47438,N_44481,N_42108);
nand U47439 (N_47439,N_42401,N_40591);
nor U47440 (N_47440,N_43400,N_40008);
nand U47441 (N_47441,N_44163,N_44978);
nand U47442 (N_47442,N_40141,N_44622);
or U47443 (N_47443,N_41793,N_43766);
nor U47444 (N_47444,N_44683,N_41465);
nor U47445 (N_47445,N_42475,N_42517);
nor U47446 (N_47446,N_40321,N_42578);
nand U47447 (N_47447,N_41925,N_42473);
or U47448 (N_47448,N_41159,N_43790);
or U47449 (N_47449,N_41500,N_40318);
nand U47450 (N_47450,N_44638,N_43868);
xnor U47451 (N_47451,N_44165,N_43249);
or U47452 (N_47452,N_42144,N_43535);
nor U47453 (N_47453,N_44637,N_43429);
or U47454 (N_47454,N_44259,N_42528);
nand U47455 (N_47455,N_40562,N_41397);
or U47456 (N_47456,N_43339,N_40963);
and U47457 (N_47457,N_42308,N_43207);
xnor U47458 (N_47458,N_44849,N_42312);
or U47459 (N_47459,N_44285,N_40420);
xnor U47460 (N_47460,N_44366,N_40833);
and U47461 (N_47461,N_41191,N_40154);
xor U47462 (N_47462,N_41750,N_44571);
nor U47463 (N_47463,N_42143,N_42997);
or U47464 (N_47464,N_41160,N_43525);
and U47465 (N_47465,N_42946,N_44018);
nand U47466 (N_47466,N_44582,N_44753);
and U47467 (N_47467,N_44752,N_44183);
and U47468 (N_47468,N_41481,N_42146);
nor U47469 (N_47469,N_44619,N_42609);
nand U47470 (N_47470,N_44351,N_41088);
or U47471 (N_47471,N_42073,N_42540);
nor U47472 (N_47472,N_40124,N_44129);
or U47473 (N_47473,N_44526,N_43779);
nand U47474 (N_47474,N_43495,N_44829);
xnor U47475 (N_47475,N_40728,N_43242);
and U47476 (N_47476,N_44556,N_40167);
xor U47477 (N_47477,N_42088,N_43500);
nand U47478 (N_47478,N_40981,N_41906);
and U47479 (N_47479,N_42375,N_42420);
or U47480 (N_47480,N_43472,N_43569);
and U47481 (N_47481,N_44761,N_44158);
nand U47482 (N_47482,N_40232,N_42959);
and U47483 (N_47483,N_41920,N_42342);
xnor U47484 (N_47484,N_43691,N_41092);
xnor U47485 (N_47485,N_43466,N_44700);
or U47486 (N_47486,N_43201,N_41116);
nor U47487 (N_47487,N_42213,N_44533);
or U47488 (N_47488,N_41842,N_42252);
and U47489 (N_47489,N_40539,N_41168);
nor U47490 (N_47490,N_43425,N_44696);
or U47491 (N_47491,N_44450,N_40003);
nor U47492 (N_47492,N_44685,N_43166);
nand U47493 (N_47493,N_43818,N_40806);
and U47494 (N_47494,N_42468,N_44485);
or U47495 (N_47495,N_41543,N_40888);
nor U47496 (N_47496,N_42001,N_44387);
or U47497 (N_47497,N_41584,N_44789);
or U47498 (N_47498,N_41015,N_43567);
xor U47499 (N_47499,N_43911,N_42848);
xnor U47500 (N_47500,N_44934,N_43039);
xnor U47501 (N_47501,N_42841,N_44401);
or U47502 (N_47502,N_41693,N_41353);
nor U47503 (N_47503,N_44003,N_44504);
xnor U47504 (N_47504,N_42917,N_40516);
nand U47505 (N_47505,N_40784,N_44375);
nor U47506 (N_47506,N_43544,N_41409);
or U47507 (N_47507,N_44955,N_44269);
xnor U47508 (N_47508,N_43544,N_43785);
and U47509 (N_47509,N_42758,N_40125);
xor U47510 (N_47510,N_40100,N_44500);
or U47511 (N_47511,N_44478,N_44017);
xnor U47512 (N_47512,N_44250,N_40229);
nand U47513 (N_47513,N_42496,N_41564);
nand U47514 (N_47514,N_44071,N_41948);
or U47515 (N_47515,N_41797,N_40520);
and U47516 (N_47516,N_41254,N_44310);
and U47517 (N_47517,N_44200,N_40519);
and U47518 (N_47518,N_43220,N_41600);
xnor U47519 (N_47519,N_40693,N_41678);
and U47520 (N_47520,N_42410,N_44073);
and U47521 (N_47521,N_41055,N_43946);
and U47522 (N_47522,N_44216,N_42409);
nor U47523 (N_47523,N_44763,N_43368);
xnor U47524 (N_47524,N_44225,N_40901);
and U47525 (N_47525,N_40577,N_40952);
xor U47526 (N_47526,N_44436,N_43383);
and U47527 (N_47527,N_41085,N_42831);
or U47528 (N_47528,N_42669,N_40582);
xnor U47529 (N_47529,N_40241,N_42650);
and U47530 (N_47530,N_41683,N_44206);
nand U47531 (N_47531,N_43320,N_40585);
and U47532 (N_47532,N_41785,N_43193);
or U47533 (N_47533,N_43762,N_43304);
and U47534 (N_47534,N_44012,N_44479);
or U47535 (N_47535,N_44067,N_41020);
nor U47536 (N_47536,N_40467,N_42950);
and U47537 (N_47537,N_40472,N_43206);
xnor U47538 (N_47538,N_42091,N_43230);
nor U47539 (N_47539,N_40886,N_41458);
or U47540 (N_47540,N_42403,N_42169);
nor U47541 (N_47541,N_40557,N_40213);
or U47542 (N_47542,N_42064,N_43687);
xor U47543 (N_47543,N_44703,N_42780);
nor U47544 (N_47544,N_41370,N_43265);
xor U47545 (N_47545,N_41004,N_44153);
or U47546 (N_47546,N_43721,N_41690);
nor U47547 (N_47547,N_41121,N_40057);
or U47548 (N_47548,N_40675,N_44424);
nand U47549 (N_47549,N_41172,N_43081);
or U47550 (N_47550,N_44503,N_40984);
nand U47551 (N_47551,N_42733,N_40071);
or U47552 (N_47552,N_42493,N_43204);
and U47553 (N_47553,N_43130,N_41035);
xor U47554 (N_47554,N_42244,N_41672);
nor U47555 (N_47555,N_42593,N_42209);
or U47556 (N_47556,N_40546,N_43828);
nand U47557 (N_47557,N_44994,N_40600);
xnor U47558 (N_47558,N_41686,N_44358);
nor U47559 (N_47559,N_42243,N_42678);
or U47560 (N_47560,N_40972,N_40881);
or U47561 (N_47561,N_42081,N_41873);
nor U47562 (N_47562,N_43601,N_40525);
nand U47563 (N_47563,N_44658,N_41122);
or U47564 (N_47564,N_41551,N_42952);
or U47565 (N_47565,N_42631,N_44302);
nand U47566 (N_47566,N_41850,N_43510);
or U47567 (N_47567,N_42379,N_41340);
or U47568 (N_47568,N_43136,N_43876);
and U47569 (N_47569,N_43519,N_43766);
and U47570 (N_47570,N_40676,N_44893);
xor U47571 (N_47571,N_44959,N_41218);
nor U47572 (N_47572,N_40052,N_43656);
nand U47573 (N_47573,N_43800,N_40537);
xnor U47574 (N_47574,N_40501,N_44599);
nand U47575 (N_47575,N_43009,N_42648);
xor U47576 (N_47576,N_43496,N_44345);
nor U47577 (N_47577,N_40901,N_40998);
and U47578 (N_47578,N_41211,N_40466);
and U47579 (N_47579,N_41518,N_43277);
or U47580 (N_47580,N_41581,N_42562);
xor U47581 (N_47581,N_44551,N_41695);
xor U47582 (N_47582,N_42718,N_42500);
or U47583 (N_47583,N_40312,N_43917);
nand U47584 (N_47584,N_40430,N_43055);
nor U47585 (N_47585,N_43065,N_43950);
and U47586 (N_47586,N_41035,N_43127);
and U47587 (N_47587,N_40621,N_41499);
nor U47588 (N_47588,N_42020,N_41392);
nand U47589 (N_47589,N_41309,N_44994);
xnor U47590 (N_47590,N_41764,N_44390);
or U47591 (N_47591,N_44856,N_40322);
or U47592 (N_47592,N_41267,N_44968);
xor U47593 (N_47593,N_44817,N_43348);
nand U47594 (N_47594,N_41966,N_43899);
or U47595 (N_47595,N_44130,N_41261);
nor U47596 (N_47596,N_40579,N_42024);
or U47597 (N_47597,N_41830,N_43338);
or U47598 (N_47598,N_42638,N_41118);
and U47599 (N_47599,N_40551,N_41899);
nand U47600 (N_47600,N_44831,N_40691);
or U47601 (N_47601,N_42151,N_41568);
xor U47602 (N_47602,N_44509,N_43793);
xnor U47603 (N_47603,N_44138,N_43394);
and U47604 (N_47604,N_44335,N_43762);
nor U47605 (N_47605,N_41271,N_42878);
and U47606 (N_47606,N_41812,N_40165);
nor U47607 (N_47607,N_41307,N_44584);
and U47608 (N_47608,N_43519,N_41396);
xor U47609 (N_47609,N_42298,N_40229);
xor U47610 (N_47610,N_41610,N_43154);
nor U47611 (N_47611,N_44544,N_42179);
nor U47612 (N_47612,N_43146,N_43207);
nand U47613 (N_47613,N_40661,N_42975);
nor U47614 (N_47614,N_40539,N_44268);
xnor U47615 (N_47615,N_43702,N_42806);
or U47616 (N_47616,N_44139,N_40529);
nor U47617 (N_47617,N_42957,N_44685);
nand U47618 (N_47618,N_42625,N_43579);
xnor U47619 (N_47619,N_41505,N_41466);
or U47620 (N_47620,N_41600,N_42409);
nand U47621 (N_47621,N_41811,N_44871);
or U47622 (N_47622,N_41914,N_44571);
nand U47623 (N_47623,N_43046,N_44792);
nor U47624 (N_47624,N_41084,N_44728);
nand U47625 (N_47625,N_41354,N_43495);
nand U47626 (N_47626,N_41856,N_44293);
or U47627 (N_47627,N_44418,N_40265);
xor U47628 (N_47628,N_41241,N_42992);
xnor U47629 (N_47629,N_41130,N_44735);
and U47630 (N_47630,N_40361,N_42853);
or U47631 (N_47631,N_40896,N_40639);
nand U47632 (N_47632,N_42119,N_43738);
or U47633 (N_47633,N_40701,N_42289);
nand U47634 (N_47634,N_43500,N_42666);
xnor U47635 (N_47635,N_41124,N_41965);
nand U47636 (N_47636,N_44231,N_43342);
xnor U47637 (N_47637,N_40424,N_41832);
nor U47638 (N_47638,N_42477,N_44522);
xor U47639 (N_47639,N_41836,N_42420);
xor U47640 (N_47640,N_44903,N_42305);
or U47641 (N_47641,N_41588,N_40081);
nand U47642 (N_47642,N_42471,N_41175);
nor U47643 (N_47643,N_40636,N_40054);
xnor U47644 (N_47644,N_41694,N_41185);
xnor U47645 (N_47645,N_42365,N_43521);
or U47646 (N_47646,N_43378,N_40366);
or U47647 (N_47647,N_41663,N_40598);
nor U47648 (N_47648,N_41003,N_44538);
or U47649 (N_47649,N_44934,N_42656);
xnor U47650 (N_47650,N_43034,N_44740);
xor U47651 (N_47651,N_44811,N_44137);
nand U47652 (N_47652,N_42446,N_42875);
or U47653 (N_47653,N_41640,N_43209);
xor U47654 (N_47654,N_42674,N_40245);
nand U47655 (N_47655,N_42392,N_42876);
nor U47656 (N_47656,N_43541,N_44785);
xnor U47657 (N_47657,N_40685,N_43172);
nor U47658 (N_47658,N_43326,N_40148);
nand U47659 (N_47659,N_41928,N_41888);
and U47660 (N_47660,N_41610,N_41193);
and U47661 (N_47661,N_41394,N_42128);
xnor U47662 (N_47662,N_42798,N_41403);
nor U47663 (N_47663,N_41977,N_44843);
nor U47664 (N_47664,N_44480,N_40433);
nor U47665 (N_47665,N_42657,N_43774);
and U47666 (N_47666,N_40591,N_40283);
nand U47667 (N_47667,N_42658,N_40936);
nand U47668 (N_47668,N_44056,N_40319);
xor U47669 (N_47669,N_44789,N_44403);
nand U47670 (N_47670,N_40428,N_44634);
or U47671 (N_47671,N_43620,N_40013);
xnor U47672 (N_47672,N_41152,N_44064);
xor U47673 (N_47673,N_42913,N_42193);
and U47674 (N_47674,N_41751,N_43553);
or U47675 (N_47675,N_44974,N_41129);
nor U47676 (N_47676,N_43917,N_44356);
nor U47677 (N_47677,N_43323,N_43913);
xnor U47678 (N_47678,N_43866,N_40340);
and U47679 (N_47679,N_40854,N_43941);
nor U47680 (N_47680,N_42525,N_44483);
or U47681 (N_47681,N_43222,N_43771);
and U47682 (N_47682,N_41229,N_40972);
nand U47683 (N_47683,N_44407,N_41397);
and U47684 (N_47684,N_40529,N_41686);
or U47685 (N_47685,N_43155,N_43024);
and U47686 (N_47686,N_41786,N_40521);
and U47687 (N_47687,N_44607,N_42040);
or U47688 (N_47688,N_40797,N_42216);
nor U47689 (N_47689,N_41196,N_40925);
nor U47690 (N_47690,N_41690,N_42674);
nand U47691 (N_47691,N_40200,N_43115);
or U47692 (N_47692,N_44931,N_41882);
nor U47693 (N_47693,N_44305,N_43598);
xnor U47694 (N_47694,N_40478,N_41561);
and U47695 (N_47695,N_41810,N_43003);
nand U47696 (N_47696,N_41140,N_42479);
or U47697 (N_47697,N_41674,N_42363);
nor U47698 (N_47698,N_42311,N_43529);
nand U47699 (N_47699,N_41687,N_43900);
nand U47700 (N_47700,N_42956,N_44703);
xor U47701 (N_47701,N_43885,N_42371);
nand U47702 (N_47702,N_40812,N_42756);
or U47703 (N_47703,N_44546,N_43367);
xnor U47704 (N_47704,N_41338,N_41503);
xnor U47705 (N_47705,N_44365,N_42544);
xor U47706 (N_47706,N_44438,N_41993);
or U47707 (N_47707,N_40916,N_40503);
nand U47708 (N_47708,N_41698,N_41058);
nand U47709 (N_47709,N_40372,N_40371);
nor U47710 (N_47710,N_42307,N_41829);
xnor U47711 (N_47711,N_41376,N_44405);
or U47712 (N_47712,N_44509,N_44014);
or U47713 (N_47713,N_41833,N_40387);
xor U47714 (N_47714,N_43081,N_44460);
or U47715 (N_47715,N_42586,N_40678);
xnor U47716 (N_47716,N_44078,N_40766);
nand U47717 (N_47717,N_40998,N_41992);
xor U47718 (N_47718,N_42570,N_42850);
nand U47719 (N_47719,N_42723,N_41480);
nand U47720 (N_47720,N_44999,N_44361);
nor U47721 (N_47721,N_43174,N_42381);
nor U47722 (N_47722,N_40145,N_44381);
or U47723 (N_47723,N_41229,N_44785);
nand U47724 (N_47724,N_41644,N_44177);
nor U47725 (N_47725,N_42085,N_41754);
nand U47726 (N_47726,N_42423,N_41170);
nor U47727 (N_47727,N_44893,N_43056);
and U47728 (N_47728,N_43753,N_44516);
or U47729 (N_47729,N_43560,N_43000);
and U47730 (N_47730,N_40047,N_44707);
xor U47731 (N_47731,N_42974,N_42599);
or U47732 (N_47732,N_42093,N_44051);
or U47733 (N_47733,N_41291,N_43808);
or U47734 (N_47734,N_44632,N_40715);
nor U47735 (N_47735,N_40573,N_40273);
and U47736 (N_47736,N_42730,N_40962);
nor U47737 (N_47737,N_42687,N_42127);
and U47738 (N_47738,N_42442,N_40340);
nand U47739 (N_47739,N_42395,N_43868);
xnor U47740 (N_47740,N_44312,N_43831);
xnor U47741 (N_47741,N_40985,N_42058);
and U47742 (N_47742,N_41653,N_43470);
or U47743 (N_47743,N_40054,N_43087);
nand U47744 (N_47744,N_42405,N_43916);
and U47745 (N_47745,N_42480,N_41355);
nand U47746 (N_47746,N_40886,N_44618);
nand U47747 (N_47747,N_44959,N_40219);
xnor U47748 (N_47748,N_41453,N_43298);
and U47749 (N_47749,N_43775,N_43289);
nand U47750 (N_47750,N_44930,N_42719);
and U47751 (N_47751,N_42918,N_40900);
nand U47752 (N_47752,N_44042,N_43138);
nand U47753 (N_47753,N_41766,N_41751);
nor U47754 (N_47754,N_40886,N_41939);
nand U47755 (N_47755,N_41825,N_42396);
or U47756 (N_47756,N_41644,N_42017);
nand U47757 (N_47757,N_41259,N_42453);
and U47758 (N_47758,N_43754,N_43355);
nor U47759 (N_47759,N_42447,N_44809);
nand U47760 (N_47760,N_40753,N_41873);
nor U47761 (N_47761,N_44711,N_40452);
or U47762 (N_47762,N_44762,N_42619);
or U47763 (N_47763,N_40621,N_41732);
nor U47764 (N_47764,N_44529,N_43656);
and U47765 (N_47765,N_42116,N_40332);
and U47766 (N_47766,N_40101,N_42558);
or U47767 (N_47767,N_40038,N_41678);
nor U47768 (N_47768,N_41592,N_41811);
or U47769 (N_47769,N_42269,N_44880);
and U47770 (N_47770,N_40898,N_41071);
and U47771 (N_47771,N_44884,N_41426);
or U47772 (N_47772,N_40898,N_44749);
nor U47773 (N_47773,N_44029,N_40525);
xor U47774 (N_47774,N_41493,N_44249);
nand U47775 (N_47775,N_42411,N_44961);
xor U47776 (N_47776,N_44073,N_42950);
xnor U47777 (N_47777,N_43677,N_41139);
xnor U47778 (N_47778,N_43972,N_41688);
or U47779 (N_47779,N_44041,N_40527);
nor U47780 (N_47780,N_41179,N_40323);
nand U47781 (N_47781,N_41582,N_43886);
xor U47782 (N_47782,N_42681,N_42075);
nand U47783 (N_47783,N_41938,N_41212);
or U47784 (N_47784,N_42779,N_40652);
nand U47785 (N_47785,N_42568,N_44916);
and U47786 (N_47786,N_43570,N_40733);
nor U47787 (N_47787,N_43129,N_42180);
nor U47788 (N_47788,N_44776,N_40262);
or U47789 (N_47789,N_42765,N_43963);
nand U47790 (N_47790,N_43524,N_40634);
and U47791 (N_47791,N_44909,N_43538);
nand U47792 (N_47792,N_40698,N_40011);
xnor U47793 (N_47793,N_42772,N_44358);
and U47794 (N_47794,N_44222,N_43745);
nand U47795 (N_47795,N_41146,N_41805);
xor U47796 (N_47796,N_44149,N_41421);
or U47797 (N_47797,N_43458,N_40697);
nor U47798 (N_47798,N_41830,N_40491);
nor U47799 (N_47799,N_44769,N_43664);
nor U47800 (N_47800,N_41560,N_42933);
nand U47801 (N_47801,N_43507,N_42620);
nand U47802 (N_47802,N_43364,N_44691);
or U47803 (N_47803,N_41702,N_41468);
nand U47804 (N_47804,N_42739,N_44399);
xor U47805 (N_47805,N_43752,N_42647);
or U47806 (N_47806,N_41523,N_43823);
or U47807 (N_47807,N_42980,N_41684);
nor U47808 (N_47808,N_43829,N_41187);
or U47809 (N_47809,N_44192,N_40305);
xor U47810 (N_47810,N_42374,N_40522);
nor U47811 (N_47811,N_44596,N_40112);
and U47812 (N_47812,N_42036,N_41768);
nand U47813 (N_47813,N_41244,N_42868);
and U47814 (N_47814,N_42887,N_44643);
or U47815 (N_47815,N_41432,N_44416);
or U47816 (N_47816,N_41020,N_44628);
nand U47817 (N_47817,N_43702,N_43672);
nand U47818 (N_47818,N_44390,N_44572);
xor U47819 (N_47819,N_43875,N_43438);
nand U47820 (N_47820,N_40529,N_41192);
or U47821 (N_47821,N_43155,N_44093);
or U47822 (N_47822,N_44953,N_42367);
nor U47823 (N_47823,N_41950,N_40760);
nor U47824 (N_47824,N_43847,N_40932);
or U47825 (N_47825,N_40398,N_40742);
nand U47826 (N_47826,N_42839,N_41225);
nor U47827 (N_47827,N_40806,N_41715);
nor U47828 (N_47828,N_44810,N_41139);
nand U47829 (N_47829,N_41452,N_40168);
and U47830 (N_47830,N_43537,N_40546);
or U47831 (N_47831,N_40350,N_40551);
or U47832 (N_47832,N_43150,N_40344);
xor U47833 (N_47833,N_40105,N_44996);
xnor U47834 (N_47834,N_43666,N_40402);
nand U47835 (N_47835,N_40537,N_43526);
nor U47836 (N_47836,N_42997,N_44152);
and U47837 (N_47837,N_41949,N_40880);
xnor U47838 (N_47838,N_40887,N_41025);
nand U47839 (N_47839,N_42833,N_44989);
or U47840 (N_47840,N_44740,N_43289);
nor U47841 (N_47841,N_44627,N_42536);
nand U47842 (N_47842,N_42397,N_44379);
xor U47843 (N_47843,N_40258,N_40153);
nand U47844 (N_47844,N_40060,N_42438);
or U47845 (N_47845,N_44020,N_43642);
and U47846 (N_47846,N_41399,N_43563);
xor U47847 (N_47847,N_41801,N_44661);
or U47848 (N_47848,N_43767,N_40959);
or U47849 (N_47849,N_42497,N_44204);
xnor U47850 (N_47850,N_44605,N_44866);
nand U47851 (N_47851,N_43727,N_44650);
xnor U47852 (N_47852,N_41017,N_41519);
xor U47853 (N_47853,N_44152,N_44300);
and U47854 (N_47854,N_40378,N_43178);
or U47855 (N_47855,N_40428,N_41878);
and U47856 (N_47856,N_42247,N_41230);
nand U47857 (N_47857,N_40297,N_44731);
or U47858 (N_47858,N_42863,N_41943);
xor U47859 (N_47859,N_42908,N_41027);
and U47860 (N_47860,N_42004,N_42719);
or U47861 (N_47861,N_41204,N_44975);
xor U47862 (N_47862,N_40570,N_43674);
xnor U47863 (N_47863,N_42604,N_42104);
nor U47864 (N_47864,N_44978,N_41838);
or U47865 (N_47865,N_41087,N_44864);
nand U47866 (N_47866,N_42557,N_43126);
nor U47867 (N_47867,N_44322,N_42553);
nor U47868 (N_47868,N_43666,N_42293);
nand U47869 (N_47869,N_40081,N_44344);
and U47870 (N_47870,N_44145,N_44911);
and U47871 (N_47871,N_44410,N_40895);
or U47872 (N_47872,N_40050,N_40525);
nor U47873 (N_47873,N_44447,N_44271);
nor U47874 (N_47874,N_44114,N_41306);
and U47875 (N_47875,N_44833,N_44334);
xnor U47876 (N_47876,N_42417,N_42924);
nor U47877 (N_47877,N_41458,N_42757);
nor U47878 (N_47878,N_44541,N_44515);
or U47879 (N_47879,N_42115,N_40775);
xor U47880 (N_47880,N_40456,N_43683);
or U47881 (N_47881,N_44454,N_43354);
nand U47882 (N_47882,N_44682,N_44621);
xor U47883 (N_47883,N_44872,N_41266);
or U47884 (N_47884,N_44899,N_41480);
and U47885 (N_47885,N_43563,N_41705);
nand U47886 (N_47886,N_43273,N_42710);
and U47887 (N_47887,N_40367,N_40341);
nand U47888 (N_47888,N_42374,N_40719);
nor U47889 (N_47889,N_42008,N_43507);
or U47890 (N_47890,N_44170,N_41136);
and U47891 (N_47891,N_40766,N_40043);
nand U47892 (N_47892,N_41605,N_41267);
or U47893 (N_47893,N_42182,N_43188);
nand U47894 (N_47894,N_40293,N_42640);
and U47895 (N_47895,N_43042,N_40816);
nand U47896 (N_47896,N_43460,N_43595);
or U47897 (N_47897,N_42797,N_42801);
or U47898 (N_47898,N_40210,N_40269);
nand U47899 (N_47899,N_42782,N_42021);
xor U47900 (N_47900,N_41394,N_42138);
nand U47901 (N_47901,N_41994,N_41081);
xor U47902 (N_47902,N_44228,N_44066);
nand U47903 (N_47903,N_42297,N_43306);
nor U47904 (N_47904,N_40575,N_40980);
nand U47905 (N_47905,N_43787,N_42130);
nand U47906 (N_47906,N_43284,N_41537);
xor U47907 (N_47907,N_40644,N_41039);
and U47908 (N_47908,N_43750,N_42057);
or U47909 (N_47909,N_41056,N_41739);
xor U47910 (N_47910,N_42757,N_40566);
xnor U47911 (N_47911,N_43095,N_43918);
nor U47912 (N_47912,N_43184,N_43821);
and U47913 (N_47913,N_42013,N_42885);
xor U47914 (N_47914,N_43955,N_44971);
or U47915 (N_47915,N_44656,N_43318);
or U47916 (N_47916,N_42905,N_42518);
xor U47917 (N_47917,N_43249,N_44881);
and U47918 (N_47918,N_42767,N_43921);
nor U47919 (N_47919,N_43852,N_43899);
nor U47920 (N_47920,N_41935,N_43794);
or U47921 (N_47921,N_44290,N_43627);
xnor U47922 (N_47922,N_41592,N_44759);
and U47923 (N_47923,N_40683,N_41780);
nand U47924 (N_47924,N_43924,N_41063);
xor U47925 (N_47925,N_44113,N_41642);
and U47926 (N_47926,N_40531,N_41871);
and U47927 (N_47927,N_40500,N_42122);
nor U47928 (N_47928,N_41491,N_40712);
or U47929 (N_47929,N_40920,N_41243);
and U47930 (N_47930,N_41061,N_42339);
and U47931 (N_47931,N_43151,N_41419);
xnor U47932 (N_47932,N_44410,N_40642);
and U47933 (N_47933,N_41622,N_40850);
nand U47934 (N_47934,N_44766,N_42136);
or U47935 (N_47935,N_42382,N_42868);
xnor U47936 (N_47936,N_44268,N_44821);
nor U47937 (N_47937,N_43866,N_43975);
nor U47938 (N_47938,N_40752,N_43178);
and U47939 (N_47939,N_44994,N_41804);
or U47940 (N_47940,N_43814,N_41006);
nand U47941 (N_47941,N_41417,N_41127);
nand U47942 (N_47942,N_40068,N_41966);
and U47943 (N_47943,N_42485,N_40270);
nor U47944 (N_47944,N_40354,N_41557);
and U47945 (N_47945,N_44661,N_43004);
and U47946 (N_47946,N_42100,N_44373);
nand U47947 (N_47947,N_44929,N_43271);
xnor U47948 (N_47948,N_42904,N_40535);
nor U47949 (N_47949,N_43233,N_40869);
and U47950 (N_47950,N_40460,N_40023);
and U47951 (N_47951,N_44450,N_40650);
or U47952 (N_47952,N_42635,N_42096);
or U47953 (N_47953,N_43205,N_44478);
or U47954 (N_47954,N_40937,N_42942);
nor U47955 (N_47955,N_44118,N_43135);
or U47956 (N_47956,N_44834,N_42784);
xnor U47957 (N_47957,N_41169,N_42983);
and U47958 (N_47958,N_43582,N_40988);
xnor U47959 (N_47959,N_43572,N_40107);
and U47960 (N_47960,N_44320,N_44701);
nand U47961 (N_47961,N_41741,N_43833);
and U47962 (N_47962,N_43536,N_43499);
or U47963 (N_47963,N_40740,N_43567);
nor U47964 (N_47964,N_42027,N_40135);
nor U47965 (N_47965,N_41242,N_40077);
nor U47966 (N_47966,N_43748,N_41771);
or U47967 (N_47967,N_42451,N_44375);
or U47968 (N_47968,N_42549,N_43319);
nand U47969 (N_47969,N_41959,N_40783);
nand U47970 (N_47970,N_41826,N_43377);
nor U47971 (N_47971,N_43288,N_43067);
xnor U47972 (N_47972,N_40104,N_43295);
nor U47973 (N_47973,N_41627,N_40130);
nor U47974 (N_47974,N_41493,N_41164);
nor U47975 (N_47975,N_42845,N_40032);
or U47976 (N_47976,N_42950,N_43670);
xor U47977 (N_47977,N_43635,N_43985);
nor U47978 (N_47978,N_43156,N_41101);
or U47979 (N_47979,N_40878,N_40766);
nand U47980 (N_47980,N_41282,N_43007);
or U47981 (N_47981,N_40563,N_41987);
and U47982 (N_47982,N_44935,N_44846);
and U47983 (N_47983,N_42845,N_43323);
xnor U47984 (N_47984,N_41869,N_40741);
and U47985 (N_47985,N_41622,N_41781);
and U47986 (N_47986,N_41483,N_42026);
xor U47987 (N_47987,N_43571,N_40442);
and U47988 (N_47988,N_40037,N_42086);
nand U47989 (N_47989,N_43751,N_44196);
and U47990 (N_47990,N_41839,N_44241);
nor U47991 (N_47991,N_42229,N_44440);
xor U47992 (N_47992,N_40754,N_44826);
or U47993 (N_47993,N_41169,N_43443);
or U47994 (N_47994,N_43047,N_43809);
xor U47995 (N_47995,N_43793,N_44862);
nand U47996 (N_47996,N_43865,N_43780);
nor U47997 (N_47997,N_41560,N_43838);
or U47998 (N_47998,N_41777,N_41223);
and U47999 (N_47999,N_44773,N_42649);
and U48000 (N_48000,N_41488,N_44826);
and U48001 (N_48001,N_40061,N_40795);
nand U48002 (N_48002,N_42865,N_43718);
and U48003 (N_48003,N_41979,N_41836);
nor U48004 (N_48004,N_42450,N_44304);
nand U48005 (N_48005,N_40548,N_43643);
and U48006 (N_48006,N_44809,N_44767);
nor U48007 (N_48007,N_41082,N_43605);
xor U48008 (N_48008,N_40326,N_40772);
or U48009 (N_48009,N_42667,N_40090);
or U48010 (N_48010,N_41126,N_40805);
nand U48011 (N_48011,N_40057,N_44444);
xnor U48012 (N_48012,N_41328,N_43397);
xnor U48013 (N_48013,N_44883,N_40173);
nor U48014 (N_48014,N_40906,N_41404);
nor U48015 (N_48015,N_44588,N_44372);
nand U48016 (N_48016,N_40809,N_44778);
or U48017 (N_48017,N_42010,N_42454);
nor U48018 (N_48018,N_44911,N_43924);
and U48019 (N_48019,N_44960,N_44765);
or U48020 (N_48020,N_43919,N_44462);
nand U48021 (N_48021,N_44670,N_41448);
nor U48022 (N_48022,N_41982,N_41426);
and U48023 (N_48023,N_42435,N_44981);
nand U48024 (N_48024,N_41399,N_44069);
xor U48025 (N_48025,N_40106,N_40250);
nor U48026 (N_48026,N_41541,N_40823);
xor U48027 (N_48027,N_44784,N_40502);
xnor U48028 (N_48028,N_41633,N_40105);
nor U48029 (N_48029,N_40022,N_44973);
and U48030 (N_48030,N_40161,N_42738);
and U48031 (N_48031,N_40423,N_43839);
or U48032 (N_48032,N_42564,N_41166);
nor U48033 (N_48033,N_40372,N_43719);
and U48034 (N_48034,N_42131,N_40478);
and U48035 (N_48035,N_42518,N_42520);
nand U48036 (N_48036,N_42870,N_40521);
nand U48037 (N_48037,N_42560,N_42984);
and U48038 (N_48038,N_40612,N_43628);
xnor U48039 (N_48039,N_44428,N_43803);
nand U48040 (N_48040,N_43514,N_44087);
nor U48041 (N_48041,N_40680,N_42645);
nand U48042 (N_48042,N_44713,N_44590);
nor U48043 (N_48043,N_43391,N_41434);
or U48044 (N_48044,N_40866,N_44526);
or U48045 (N_48045,N_44022,N_41515);
nand U48046 (N_48046,N_43195,N_42669);
and U48047 (N_48047,N_40671,N_44404);
xor U48048 (N_48048,N_44548,N_40652);
xnor U48049 (N_48049,N_44153,N_41092);
xnor U48050 (N_48050,N_40780,N_41859);
or U48051 (N_48051,N_44858,N_44387);
xor U48052 (N_48052,N_41431,N_40591);
and U48053 (N_48053,N_44791,N_41503);
xor U48054 (N_48054,N_42560,N_44606);
xnor U48055 (N_48055,N_42349,N_40791);
nand U48056 (N_48056,N_44645,N_41683);
or U48057 (N_48057,N_40157,N_44759);
nor U48058 (N_48058,N_40786,N_44003);
xnor U48059 (N_48059,N_42232,N_44877);
xor U48060 (N_48060,N_44366,N_43175);
nand U48061 (N_48061,N_40465,N_41000);
and U48062 (N_48062,N_43498,N_43669);
or U48063 (N_48063,N_44487,N_41148);
or U48064 (N_48064,N_40352,N_42030);
or U48065 (N_48065,N_44185,N_42197);
and U48066 (N_48066,N_41237,N_41286);
or U48067 (N_48067,N_42668,N_43486);
nor U48068 (N_48068,N_44649,N_42836);
nand U48069 (N_48069,N_43413,N_40459);
nand U48070 (N_48070,N_42430,N_42506);
or U48071 (N_48071,N_44895,N_44513);
and U48072 (N_48072,N_40010,N_41950);
or U48073 (N_48073,N_44992,N_40138);
nor U48074 (N_48074,N_42572,N_43260);
nand U48075 (N_48075,N_40694,N_43996);
nand U48076 (N_48076,N_40931,N_44767);
nor U48077 (N_48077,N_43838,N_42703);
nor U48078 (N_48078,N_43183,N_41046);
nor U48079 (N_48079,N_42541,N_43022);
or U48080 (N_48080,N_43097,N_41454);
xor U48081 (N_48081,N_43468,N_44554);
xnor U48082 (N_48082,N_40928,N_41387);
and U48083 (N_48083,N_41483,N_42320);
or U48084 (N_48084,N_42375,N_41069);
nor U48085 (N_48085,N_41514,N_41495);
nor U48086 (N_48086,N_41885,N_42728);
xor U48087 (N_48087,N_40297,N_43811);
and U48088 (N_48088,N_41526,N_43663);
xor U48089 (N_48089,N_43914,N_41638);
nor U48090 (N_48090,N_40921,N_40374);
and U48091 (N_48091,N_40487,N_43665);
or U48092 (N_48092,N_41722,N_43868);
and U48093 (N_48093,N_42422,N_43831);
xor U48094 (N_48094,N_44491,N_40380);
xor U48095 (N_48095,N_43485,N_43419);
nor U48096 (N_48096,N_40996,N_41607);
xnor U48097 (N_48097,N_42401,N_41383);
or U48098 (N_48098,N_44374,N_43503);
nand U48099 (N_48099,N_41603,N_40761);
xnor U48100 (N_48100,N_43343,N_44363);
or U48101 (N_48101,N_42775,N_40416);
nand U48102 (N_48102,N_43941,N_43917);
nand U48103 (N_48103,N_40511,N_42639);
nor U48104 (N_48104,N_40539,N_41855);
or U48105 (N_48105,N_41243,N_40007);
nand U48106 (N_48106,N_40337,N_44463);
nand U48107 (N_48107,N_44390,N_41795);
nor U48108 (N_48108,N_41743,N_44814);
nand U48109 (N_48109,N_43301,N_44121);
nand U48110 (N_48110,N_43886,N_42298);
nand U48111 (N_48111,N_41925,N_42547);
or U48112 (N_48112,N_40224,N_44505);
nor U48113 (N_48113,N_41638,N_42442);
or U48114 (N_48114,N_41302,N_40625);
nand U48115 (N_48115,N_40934,N_41078);
nand U48116 (N_48116,N_42914,N_42446);
nor U48117 (N_48117,N_44536,N_41474);
nor U48118 (N_48118,N_43684,N_43256);
nand U48119 (N_48119,N_40020,N_43553);
or U48120 (N_48120,N_41149,N_40874);
nand U48121 (N_48121,N_41609,N_42237);
or U48122 (N_48122,N_42221,N_43791);
or U48123 (N_48123,N_44589,N_43178);
xor U48124 (N_48124,N_44382,N_43030);
nand U48125 (N_48125,N_40535,N_41742);
xnor U48126 (N_48126,N_41543,N_42173);
xor U48127 (N_48127,N_40953,N_41183);
and U48128 (N_48128,N_44663,N_42483);
or U48129 (N_48129,N_42190,N_41341);
xnor U48130 (N_48130,N_42624,N_40781);
xor U48131 (N_48131,N_41473,N_42382);
or U48132 (N_48132,N_41029,N_40581);
nor U48133 (N_48133,N_41969,N_40750);
and U48134 (N_48134,N_42446,N_42772);
and U48135 (N_48135,N_43634,N_43768);
nor U48136 (N_48136,N_42508,N_40512);
xor U48137 (N_48137,N_41429,N_44256);
or U48138 (N_48138,N_43027,N_44791);
and U48139 (N_48139,N_41592,N_43237);
and U48140 (N_48140,N_41355,N_44183);
or U48141 (N_48141,N_41033,N_40639);
and U48142 (N_48142,N_40699,N_44969);
nor U48143 (N_48143,N_42341,N_43391);
and U48144 (N_48144,N_42532,N_44249);
nor U48145 (N_48145,N_40499,N_41475);
or U48146 (N_48146,N_41258,N_43116);
nand U48147 (N_48147,N_43388,N_42655);
nor U48148 (N_48148,N_41234,N_44727);
and U48149 (N_48149,N_44004,N_42382);
nor U48150 (N_48150,N_40911,N_42349);
and U48151 (N_48151,N_40318,N_43088);
and U48152 (N_48152,N_43853,N_41134);
nor U48153 (N_48153,N_43560,N_40626);
nor U48154 (N_48154,N_42107,N_41298);
and U48155 (N_48155,N_42479,N_41472);
xnor U48156 (N_48156,N_41927,N_41519);
nand U48157 (N_48157,N_43756,N_41562);
xnor U48158 (N_48158,N_40162,N_41035);
or U48159 (N_48159,N_41632,N_41376);
and U48160 (N_48160,N_44629,N_44489);
nor U48161 (N_48161,N_40873,N_42896);
xor U48162 (N_48162,N_41792,N_43691);
nand U48163 (N_48163,N_41938,N_44137);
and U48164 (N_48164,N_40917,N_41620);
nor U48165 (N_48165,N_41343,N_41539);
or U48166 (N_48166,N_40361,N_42491);
or U48167 (N_48167,N_44725,N_44102);
or U48168 (N_48168,N_40571,N_44153);
or U48169 (N_48169,N_40832,N_42144);
nand U48170 (N_48170,N_43013,N_41561);
or U48171 (N_48171,N_44158,N_44262);
and U48172 (N_48172,N_43576,N_42509);
nand U48173 (N_48173,N_44391,N_40679);
and U48174 (N_48174,N_44015,N_42025);
or U48175 (N_48175,N_40512,N_43735);
nor U48176 (N_48176,N_42971,N_44472);
xor U48177 (N_48177,N_43441,N_43941);
nand U48178 (N_48178,N_40015,N_41208);
xor U48179 (N_48179,N_41108,N_44010);
or U48180 (N_48180,N_42125,N_42993);
nor U48181 (N_48181,N_40752,N_42085);
nor U48182 (N_48182,N_43056,N_41399);
xor U48183 (N_48183,N_40569,N_41784);
xor U48184 (N_48184,N_41768,N_41013);
xor U48185 (N_48185,N_43468,N_43905);
and U48186 (N_48186,N_43281,N_43244);
nor U48187 (N_48187,N_43163,N_41313);
xnor U48188 (N_48188,N_42730,N_43072);
and U48189 (N_48189,N_43662,N_44391);
xnor U48190 (N_48190,N_42044,N_44324);
nor U48191 (N_48191,N_43420,N_41444);
nand U48192 (N_48192,N_42128,N_44257);
or U48193 (N_48193,N_43852,N_42715);
nor U48194 (N_48194,N_42572,N_44521);
nand U48195 (N_48195,N_44408,N_40257);
xor U48196 (N_48196,N_41639,N_42730);
xnor U48197 (N_48197,N_44855,N_42136);
nand U48198 (N_48198,N_43524,N_42984);
xor U48199 (N_48199,N_40171,N_43111);
or U48200 (N_48200,N_44410,N_41083);
xor U48201 (N_48201,N_44196,N_42624);
or U48202 (N_48202,N_41548,N_43046);
nor U48203 (N_48203,N_42035,N_41181);
and U48204 (N_48204,N_43936,N_42709);
and U48205 (N_48205,N_44791,N_41678);
nand U48206 (N_48206,N_43874,N_44344);
xor U48207 (N_48207,N_42178,N_41178);
or U48208 (N_48208,N_40900,N_44835);
nand U48209 (N_48209,N_44039,N_44097);
or U48210 (N_48210,N_44047,N_42259);
nand U48211 (N_48211,N_41459,N_40570);
nor U48212 (N_48212,N_44344,N_43077);
nor U48213 (N_48213,N_44870,N_42118);
and U48214 (N_48214,N_44564,N_40542);
xnor U48215 (N_48215,N_43359,N_41164);
nor U48216 (N_48216,N_40455,N_44649);
nand U48217 (N_48217,N_42427,N_44078);
nor U48218 (N_48218,N_40723,N_43390);
nand U48219 (N_48219,N_40791,N_43536);
nand U48220 (N_48220,N_40520,N_42955);
or U48221 (N_48221,N_42668,N_44332);
xnor U48222 (N_48222,N_40354,N_43997);
nor U48223 (N_48223,N_44855,N_43172);
xor U48224 (N_48224,N_40115,N_42556);
xor U48225 (N_48225,N_44746,N_44431);
and U48226 (N_48226,N_43686,N_43596);
and U48227 (N_48227,N_43802,N_42856);
nor U48228 (N_48228,N_41697,N_41080);
and U48229 (N_48229,N_43438,N_43226);
or U48230 (N_48230,N_44954,N_40835);
nor U48231 (N_48231,N_42518,N_41631);
or U48232 (N_48232,N_44223,N_41240);
nand U48233 (N_48233,N_44722,N_43959);
nor U48234 (N_48234,N_41222,N_44840);
and U48235 (N_48235,N_40696,N_42816);
or U48236 (N_48236,N_44545,N_41825);
nand U48237 (N_48237,N_40373,N_41074);
or U48238 (N_48238,N_42618,N_42048);
xor U48239 (N_48239,N_42413,N_40487);
nor U48240 (N_48240,N_41043,N_44469);
and U48241 (N_48241,N_42354,N_41415);
nand U48242 (N_48242,N_40693,N_40562);
or U48243 (N_48243,N_41975,N_40605);
or U48244 (N_48244,N_40940,N_40160);
or U48245 (N_48245,N_44595,N_41158);
nor U48246 (N_48246,N_41367,N_44073);
nand U48247 (N_48247,N_44034,N_41394);
nand U48248 (N_48248,N_44384,N_44402);
xor U48249 (N_48249,N_42692,N_43248);
and U48250 (N_48250,N_43379,N_41270);
and U48251 (N_48251,N_40647,N_41228);
nor U48252 (N_48252,N_43222,N_41961);
nor U48253 (N_48253,N_41076,N_41397);
or U48254 (N_48254,N_43897,N_40743);
nand U48255 (N_48255,N_44622,N_43400);
nand U48256 (N_48256,N_42639,N_44177);
and U48257 (N_48257,N_40299,N_41353);
nor U48258 (N_48258,N_44590,N_44229);
xnor U48259 (N_48259,N_42858,N_43363);
xor U48260 (N_48260,N_40443,N_41634);
xor U48261 (N_48261,N_41888,N_44011);
nand U48262 (N_48262,N_44015,N_44234);
nor U48263 (N_48263,N_40722,N_40981);
nand U48264 (N_48264,N_40790,N_41748);
and U48265 (N_48265,N_41475,N_41860);
nand U48266 (N_48266,N_44039,N_44022);
xor U48267 (N_48267,N_41478,N_43947);
and U48268 (N_48268,N_41201,N_41319);
nand U48269 (N_48269,N_43775,N_41608);
or U48270 (N_48270,N_40472,N_43705);
nor U48271 (N_48271,N_44384,N_44492);
nand U48272 (N_48272,N_43084,N_41273);
and U48273 (N_48273,N_43305,N_40563);
nor U48274 (N_48274,N_44999,N_42601);
xnor U48275 (N_48275,N_42522,N_44682);
and U48276 (N_48276,N_41849,N_44244);
or U48277 (N_48277,N_42104,N_40319);
nor U48278 (N_48278,N_41654,N_42087);
nand U48279 (N_48279,N_40379,N_40762);
xnor U48280 (N_48280,N_40333,N_42536);
or U48281 (N_48281,N_43505,N_41576);
and U48282 (N_48282,N_42361,N_43958);
nand U48283 (N_48283,N_42552,N_40145);
nand U48284 (N_48284,N_42454,N_41490);
nor U48285 (N_48285,N_43644,N_43879);
nand U48286 (N_48286,N_44068,N_44403);
xnor U48287 (N_48287,N_40909,N_44684);
xor U48288 (N_48288,N_41747,N_43706);
nand U48289 (N_48289,N_41650,N_40868);
and U48290 (N_48290,N_41338,N_40966);
xnor U48291 (N_48291,N_40473,N_44669);
and U48292 (N_48292,N_44323,N_41149);
xnor U48293 (N_48293,N_41142,N_43782);
or U48294 (N_48294,N_40585,N_42159);
xnor U48295 (N_48295,N_40519,N_44795);
xor U48296 (N_48296,N_44671,N_41383);
or U48297 (N_48297,N_40238,N_41780);
or U48298 (N_48298,N_40586,N_41625);
xor U48299 (N_48299,N_43380,N_40453);
or U48300 (N_48300,N_40171,N_43574);
nor U48301 (N_48301,N_43899,N_42131);
nand U48302 (N_48302,N_43257,N_41723);
and U48303 (N_48303,N_41811,N_44423);
nor U48304 (N_48304,N_44118,N_44207);
and U48305 (N_48305,N_42422,N_41129);
and U48306 (N_48306,N_42413,N_44867);
xnor U48307 (N_48307,N_43915,N_42478);
nand U48308 (N_48308,N_40790,N_40739);
and U48309 (N_48309,N_41866,N_40454);
xnor U48310 (N_48310,N_40127,N_43094);
xnor U48311 (N_48311,N_43387,N_43895);
nor U48312 (N_48312,N_41779,N_41383);
and U48313 (N_48313,N_40539,N_44753);
nand U48314 (N_48314,N_40442,N_42084);
and U48315 (N_48315,N_42626,N_43462);
xor U48316 (N_48316,N_41385,N_42431);
and U48317 (N_48317,N_44035,N_41951);
nand U48318 (N_48318,N_42131,N_44558);
nor U48319 (N_48319,N_41385,N_43046);
xor U48320 (N_48320,N_40900,N_40064);
xnor U48321 (N_48321,N_44901,N_40045);
and U48322 (N_48322,N_40691,N_41530);
nor U48323 (N_48323,N_40002,N_42755);
xor U48324 (N_48324,N_44057,N_42293);
nand U48325 (N_48325,N_40987,N_43269);
nor U48326 (N_48326,N_44848,N_44447);
xnor U48327 (N_48327,N_41064,N_44220);
or U48328 (N_48328,N_43799,N_44720);
nand U48329 (N_48329,N_40852,N_44652);
xnor U48330 (N_48330,N_40224,N_43787);
xor U48331 (N_48331,N_42126,N_42363);
nor U48332 (N_48332,N_41945,N_41032);
and U48333 (N_48333,N_43274,N_44992);
or U48334 (N_48334,N_43403,N_42057);
nor U48335 (N_48335,N_41000,N_43991);
xor U48336 (N_48336,N_40773,N_42232);
xnor U48337 (N_48337,N_42005,N_40897);
and U48338 (N_48338,N_42164,N_44565);
nor U48339 (N_48339,N_42755,N_40204);
nand U48340 (N_48340,N_40180,N_40902);
and U48341 (N_48341,N_41047,N_44722);
or U48342 (N_48342,N_43471,N_40866);
nand U48343 (N_48343,N_41113,N_40198);
and U48344 (N_48344,N_40323,N_40063);
and U48345 (N_48345,N_40562,N_41371);
nor U48346 (N_48346,N_40145,N_44667);
nor U48347 (N_48347,N_41151,N_42014);
nor U48348 (N_48348,N_43012,N_44052);
or U48349 (N_48349,N_40451,N_44841);
or U48350 (N_48350,N_42440,N_43593);
and U48351 (N_48351,N_40034,N_41234);
nand U48352 (N_48352,N_43931,N_40420);
nand U48353 (N_48353,N_42538,N_41191);
or U48354 (N_48354,N_44693,N_41253);
or U48355 (N_48355,N_43784,N_41494);
and U48356 (N_48356,N_41334,N_42561);
nand U48357 (N_48357,N_42512,N_41650);
nand U48358 (N_48358,N_41722,N_41493);
and U48359 (N_48359,N_43568,N_42192);
and U48360 (N_48360,N_44241,N_43277);
nand U48361 (N_48361,N_43146,N_43589);
and U48362 (N_48362,N_44042,N_40811);
or U48363 (N_48363,N_40184,N_40634);
and U48364 (N_48364,N_40651,N_43674);
nor U48365 (N_48365,N_44316,N_41453);
nor U48366 (N_48366,N_40148,N_40824);
nor U48367 (N_48367,N_44041,N_43394);
or U48368 (N_48368,N_44715,N_42360);
and U48369 (N_48369,N_41780,N_44212);
or U48370 (N_48370,N_40689,N_40901);
nand U48371 (N_48371,N_44020,N_42528);
or U48372 (N_48372,N_41483,N_40986);
and U48373 (N_48373,N_41418,N_41267);
or U48374 (N_48374,N_42398,N_43246);
or U48375 (N_48375,N_40119,N_43181);
or U48376 (N_48376,N_41727,N_43042);
xnor U48377 (N_48377,N_42149,N_40928);
or U48378 (N_48378,N_43837,N_41692);
nor U48379 (N_48379,N_42200,N_41939);
nand U48380 (N_48380,N_44419,N_42701);
xor U48381 (N_48381,N_43114,N_42777);
and U48382 (N_48382,N_43073,N_43806);
xnor U48383 (N_48383,N_43319,N_41682);
nand U48384 (N_48384,N_44452,N_40070);
and U48385 (N_48385,N_43518,N_44161);
nor U48386 (N_48386,N_41911,N_40996);
xnor U48387 (N_48387,N_43847,N_43260);
and U48388 (N_48388,N_43339,N_43366);
nand U48389 (N_48389,N_40149,N_43910);
nor U48390 (N_48390,N_40438,N_41571);
xor U48391 (N_48391,N_42020,N_41438);
nand U48392 (N_48392,N_44781,N_43466);
and U48393 (N_48393,N_44588,N_42637);
nand U48394 (N_48394,N_41158,N_41860);
nor U48395 (N_48395,N_41057,N_41924);
or U48396 (N_48396,N_43292,N_41573);
nor U48397 (N_48397,N_43200,N_44278);
and U48398 (N_48398,N_44552,N_44586);
nand U48399 (N_48399,N_42719,N_43663);
nor U48400 (N_48400,N_43567,N_41574);
xor U48401 (N_48401,N_42066,N_43928);
and U48402 (N_48402,N_44617,N_43183);
xor U48403 (N_48403,N_41337,N_42418);
or U48404 (N_48404,N_44035,N_40701);
nand U48405 (N_48405,N_43378,N_44292);
and U48406 (N_48406,N_40548,N_41852);
nor U48407 (N_48407,N_40896,N_40668);
or U48408 (N_48408,N_44552,N_40933);
xor U48409 (N_48409,N_40204,N_40975);
and U48410 (N_48410,N_40120,N_42372);
xnor U48411 (N_48411,N_43211,N_43939);
nand U48412 (N_48412,N_41520,N_41857);
and U48413 (N_48413,N_42586,N_43355);
xor U48414 (N_48414,N_44609,N_43696);
nor U48415 (N_48415,N_43825,N_40003);
and U48416 (N_48416,N_42790,N_43515);
and U48417 (N_48417,N_41263,N_40233);
or U48418 (N_48418,N_43659,N_40507);
nor U48419 (N_48419,N_43029,N_41095);
xnor U48420 (N_48420,N_43040,N_44788);
nand U48421 (N_48421,N_42392,N_44589);
nor U48422 (N_48422,N_42978,N_44122);
or U48423 (N_48423,N_40972,N_42247);
nand U48424 (N_48424,N_41839,N_40529);
and U48425 (N_48425,N_41220,N_42277);
nand U48426 (N_48426,N_42732,N_41089);
xor U48427 (N_48427,N_43972,N_43693);
nand U48428 (N_48428,N_43336,N_42412);
and U48429 (N_48429,N_42865,N_42639);
xor U48430 (N_48430,N_40301,N_44822);
nor U48431 (N_48431,N_43747,N_41934);
xor U48432 (N_48432,N_40930,N_44205);
xor U48433 (N_48433,N_43306,N_42629);
nor U48434 (N_48434,N_44266,N_41536);
and U48435 (N_48435,N_42813,N_42565);
and U48436 (N_48436,N_40250,N_44261);
nor U48437 (N_48437,N_43774,N_43476);
nand U48438 (N_48438,N_43745,N_40288);
or U48439 (N_48439,N_44550,N_42833);
and U48440 (N_48440,N_44268,N_44761);
nand U48441 (N_48441,N_43453,N_41185);
xnor U48442 (N_48442,N_44208,N_43633);
or U48443 (N_48443,N_40380,N_43454);
or U48444 (N_48444,N_43672,N_44333);
or U48445 (N_48445,N_44473,N_43005);
and U48446 (N_48446,N_42964,N_41727);
xor U48447 (N_48447,N_40183,N_40978);
or U48448 (N_48448,N_43653,N_43743);
and U48449 (N_48449,N_42441,N_43842);
and U48450 (N_48450,N_43477,N_40011);
or U48451 (N_48451,N_40087,N_41715);
nor U48452 (N_48452,N_42326,N_43780);
and U48453 (N_48453,N_40121,N_44888);
and U48454 (N_48454,N_42918,N_40898);
or U48455 (N_48455,N_44596,N_43055);
xor U48456 (N_48456,N_41525,N_41680);
and U48457 (N_48457,N_43745,N_43480);
nand U48458 (N_48458,N_44976,N_44293);
nor U48459 (N_48459,N_41162,N_40524);
and U48460 (N_48460,N_43566,N_41720);
nor U48461 (N_48461,N_41992,N_42631);
nor U48462 (N_48462,N_41512,N_40296);
and U48463 (N_48463,N_44817,N_43901);
and U48464 (N_48464,N_43234,N_44375);
and U48465 (N_48465,N_40979,N_44507);
or U48466 (N_48466,N_40479,N_40661);
nand U48467 (N_48467,N_42320,N_43792);
nand U48468 (N_48468,N_42046,N_41537);
or U48469 (N_48469,N_40290,N_43083);
xor U48470 (N_48470,N_40601,N_41228);
nor U48471 (N_48471,N_43350,N_42580);
nor U48472 (N_48472,N_43578,N_41241);
and U48473 (N_48473,N_43382,N_43016);
or U48474 (N_48474,N_43356,N_40566);
xnor U48475 (N_48475,N_40816,N_43944);
or U48476 (N_48476,N_43382,N_41094);
nor U48477 (N_48477,N_43404,N_44042);
xor U48478 (N_48478,N_42146,N_44434);
nand U48479 (N_48479,N_41699,N_43920);
nor U48480 (N_48480,N_40638,N_41802);
or U48481 (N_48481,N_44112,N_40174);
xor U48482 (N_48482,N_42542,N_41703);
nor U48483 (N_48483,N_43066,N_41573);
nor U48484 (N_48484,N_40802,N_41404);
nand U48485 (N_48485,N_42906,N_44333);
and U48486 (N_48486,N_44442,N_41549);
xor U48487 (N_48487,N_41439,N_42961);
nand U48488 (N_48488,N_44274,N_42272);
or U48489 (N_48489,N_44330,N_41918);
or U48490 (N_48490,N_40111,N_42669);
xnor U48491 (N_48491,N_41210,N_44750);
and U48492 (N_48492,N_40432,N_43978);
and U48493 (N_48493,N_44983,N_41057);
or U48494 (N_48494,N_44201,N_43917);
nand U48495 (N_48495,N_40744,N_43558);
xor U48496 (N_48496,N_42665,N_40575);
or U48497 (N_48497,N_40551,N_43082);
or U48498 (N_48498,N_42250,N_42954);
or U48499 (N_48499,N_43550,N_44091);
nand U48500 (N_48500,N_41971,N_41187);
xor U48501 (N_48501,N_41207,N_44689);
nor U48502 (N_48502,N_41617,N_43717);
or U48503 (N_48503,N_40618,N_44701);
nor U48504 (N_48504,N_42268,N_42609);
xnor U48505 (N_48505,N_44219,N_41275);
or U48506 (N_48506,N_40362,N_41328);
xor U48507 (N_48507,N_41083,N_40724);
or U48508 (N_48508,N_42693,N_42039);
nand U48509 (N_48509,N_43760,N_43888);
nor U48510 (N_48510,N_43804,N_42003);
or U48511 (N_48511,N_43260,N_42845);
nand U48512 (N_48512,N_40621,N_40856);
xor U48513 (N_48513,N_40013,N_42153);
nor U48514 (N_48514,N_43644,N_41114);
nand U48515 (N_48515,N_41387,N_43255);
nand U48516 (N_48516,N_44355,N_43227);
or U48517 (N_48517,N_40384,N_41194);
or U48518 (N_48518,N_44576,N_41315);
nor U48519 (N_48519,N_40303,N_42594);
nand U48520 (N_48520,N_41456,N_44240);
xnor U48521 (N_48521,N_44126,N_41542);
and U48522 (N_48522,N_42575,N_40999);
or U48523 (N_48523,N_43605,N_40773);
nor U48524 (N_48524,N_44058,N_42949);
nand U48525 (N_48525,N_43329,N_40952);
and U48526 (N_48526,N_43870,N_42511);
nand U48527 (N_48527,N_40443,N_41422);
nor U48528 (N_48528,N_41517,N_41445);
nand U48529 (N_48529,N_44161,N_41135);
and U48530 (N_48530,N_42282,N_44361);
or U48531 (N_48531,N_40861,N_41455);
or U48532 (N_48532,N_42283,N_40813);
and U48533 (N_48533,N_44009,N_41948);
xor U48534 (N_48534,N_43553,N_44207);
xor U48535 (N_48535,N_41048,N_40092);
or U48536 (N_48536,N_43778,N_40212);
nor U48537 (N_48537,N_43715,N_43915);
nand U48538 (N_48538,N_44839,N_44163);
xor U48539 (N_48539,N_41062,N_44599);
nand U48540 (N_48540,N_42196,N_40098);
nor U48541 (N_48541,N_43069,N_43666);
and U48542 (N_48542,N_42747,N_43214);
nor U48543 (N_48543,N_41185,N_43885);
nand U48544 (N_48544,N_40609,N_40912);
and U48545 (N_48545,N_43374,N_44734);
nand U48546 (N_48546,N_43990,N_40253);
xor U48547 (N_48547,N_40542,N_44773);
nor U48548 (N_48548,N_40722,N_41682);
nor U48549 (N_48549,N_40229,N_42681);
xor U48550 (N_48550,N_44272,N_43287);
nand U48551 (N_48551,N_43218,N_43299);
or U48552 (N_48552,N_43783,N_40634);
nor U48553 (N_48553,N_40147,N_41312);
nor U48554 (N_48554,N_41086,N_41632);
or U48555 (N_48555,N_43105,N_42169);
and U48556 (N_48556,N_40235,N_40224);
or U48557 (N_48557,N_44402,N_41004);
and U48558 (N_48558,N_40168,N_42764);
nor U48559 (N_48559,N_40302,N_41239);
nor U48560 (N_48560,N_44079,N_42055);
xor U48561 (N_48561,N_42793,N_42351);
nand U48562 (N_48562,N_44017,N_43830);
and U48563 (N_48563,N_42582,N_41079);
or U48564 (N_48564,N_40131,N_41989);
nor U48565 (N_48565,N_40229,N_44576);
nand U48566 (N_48566,N_40821,N_44505);
nor U48567 (N_48567,N_41409,N_42645);
or U48568 (N_48568,N_41111,N_40644);
nor U48569 (N_48569,N_42031,N_42446);
and U48570 (N_48570,N_41251,N_41280);
or U48571 (N_48571,N_42510,N_42883);
and U48572 (N_48572,N_44424,N_41944);
xnor U48573 (N_48573,N_42649,N_40088);
xor U48574 (N_48574,N_43347,N_44999);
nand U48575 (N_48575,N_44218,N_44102);
xor U48576 (N_48576,N_43072,N_44771);
nor U48577 (N_48577,N_42979,N_41383);
nor U48578 (N_48578,N_43831,N_44622);
xor U48579 (N_48579,N_42300,N_43095);
and U48580 (N_48580,N_43692,N_41240);
nand U48581 (N_48581,N_41962,N_41552);
nand U48582 (N_48582,N_42447,N_41826);
and U48583 (N_48583,N_44104,N_44225);
nor U48584 (N_48584,N_41395,N_43669);
xnor U48585 (N_48585,N_42813,N_41589);
or U48586 (N_48586,N_44902,N_40237);
or U48587 (N_48587,N_40833,N_44349);
xnor U48588 (N_48588,N_42152,N_44626);
xnor U48589 (N_48589,N_44922,N_42659);
xor U48590 (N_48590,N_44049,N_40505);
nand U48591 (N_48591,N_44545,N_43041);
or U48592 (N_48592,N_41528,N_44024);
nor U48593 (N_48593,N_42586,N_41045);
and U48594 (N_48594,N_42073,N_43705);
xnor U48595 (N_48595,N_41086,N_42852);
nand U48596 (N_48596,N_43052,N_42249);
nand U48597 (N_48597,N_43702,N_41804);
and U48598 (N_48598,N_42013,N_41250);
xor U48599 (N_48599,N_42765,N_40161);
xor U48600 (N_48600,N_42658,N_44837);
nor U48601 (N_48601,N_41753,N_44616);
nand U48602 (N_48602,N_40644,N_41839);
and U48603 (N_48603,N_41127,N_42549);
nand U48604 (N_48604,N_41565,N_40042);
or U48605 (N_48605,N_43129,N_44930);
and U48606 (N_48606,N_42255,N_41028);
nor U48607 (N_48607,N_42220,N_42945);
or U48608 (N_48608,N_44144,N_44201);
xnor U48609 (N_48609,N_44213,N_41819);
or U48610 (N_48610,N_40630,N_42556);
xnor U48611 (N_48611,N_41675,N_42879);
xor U48612 (N_48612,N_42916,N_44392);
nor U48613 (N_48613,N_41070,N_42457);
or U48614 (N_48614,N_44899,N_40282);
or U48615 (N_48615,N_43968,N_41307);
and U48616 (N_48616,N_44277,N_41864);
or U48617 (N_48617,N_43304,N_43062);
or U48618 (N_48618,N_40461,N_42249);
and U48619 (N_48619,N_42049,N_42746);
xor U48620 (N_48620,N_41864,N_40465);
or U48621 (N_48621,N_41569,N_42913);
or U48622 (N_48622,N_44701,N_41270);
xor U48623 (N_48623,N_44343,N_44461);
and U48624 (N_48624,N_44584,N_41300);
nand U48625 (N_48625,N_40087,N_42675);
and U48626 (N_48626,N_43890,N_42500);
nor U48627 (N_48627,N_40991,N_41137);
nand U48628 (N_48628,N_43485,N_41911);
xnor U48629 (N_48629,N_44769,N_44911);
nor U48630 (N_48630,N_43563,N_40240);
xor U48631 (N_48631,N_43611,N_44026);
nand U48632 (N_48632,N_44083,N_40699);
xnor U48633 (N_48633,N_42688,N_42473);
nor U48634 (N_48634,N_43312,N_42128);
or U48635 (N_48635,N_43416,N_44719);
and U48636 (N_48636,N_40321,N_44492);
nand U48637 (N_48637,N_43757,N_41120);
nand U48638 (N_48638,N_42710,N_44338);
xor U48639 (N_48639,N_41561,N_44164);
or U48640 (N_48640,N_44742,N_41560);
or U48641 (N_48641,N_43310,N_42848);
or U48642 (N_48642,N_41389,N_40897);
nor U48643 (N_48643,N_44723,N_40344);
or U48644 (N_48644,N_42003,N_44457);
nand U48645 (N_48645,N_44038,N_41489);
xor U48646 (N_48646,N_42196,N_44657);
or U48647 (N_48647,N_44944,N_40882);
and U48648 (N_48648,N_43681,N_41410);
nand U48649 (N_48649,N_41823,N_44508);
nand U48650 (N_48650,N_42991,N_44288);
xnor U48651 (N_48651,N_43488,N_43674);
or U48652 (N_48652,N_44030,N_42392);
or U48653 (N_48653,N_40589,N_40512);
nor U48654 (N_48654,N_41250,N_43303);
or U48655 (N_48655,N_40736,N_43278);
or U48656 (N_48656,N_40716,N_41933);
nand U48657 (N_48657,N_40786,N_40651);
xnor U48658 (N_48658,N_42168,N_40629);
nand U48659 (N_48659,N_40774,N_42730);
nor U48660 (N_48660,N_43878,N_43826);
nand U48661 (N_48661,N_40013,N_42084);
or U48662 (N_48662,N_40658,N_42888);
nor U48663 (N_48663,N_43483,N_44164);
or U48664 (N_48664,N_41175,N_43131);
nand U48665 (N_48665,N_44886,N_41650);
nand U48666 (N_48666,N_43505,N_42626);
nand U48667 (N_48667,N_40290,N_44019);
nand U48668 (N_48668,N_41654,N_42433);
nor U48669 (N_48669,N_41392,N_43756);
or U48670 (N_48670,N_42412,N_44839);
nand U48671 (N_48671,N_40449,N_43979);
nor U48672 (N_48672,N_41335,N_42149);
nor U48673 (N_48673,N_43320,N_42149);
xor U48674 (N_48674,N_40428,N_41424);
xor U48675 (N_48675,N_44744,N_43919);
nand U48676 (N_48676,N_41656,N_40405);
nand U48677 (N_48677,N_40603,N_40399);
xnor U48678 (N_48678,N_43782,N_41553);
xnor U48679 (N_48679,N_43231,N_42025);
nor U48680 (N_48680,N_40065,N_42891);
xnor U48681 (N_48681,N_44987,N_44960);
nand U48682 (N_48682,N_40161,N_43601);
and U48683 (N_48683,N_42574,N_40479);
nor U48684 (N_48684,N_43223,N_41167);
nand U48685 (N_48685,N_42365,N_40804);
and U48686 (N_48686,N_43159,N_41716);
nor U48687 (N_48687,N_43342,N_44197);
or U48688 (N_48688,N_40528,N_42286);
or U48689 (N_48689,N_44872,N_44904);
nand U48690 (N_48690,N_43127,N_42190);
and U48691 (N_48691,N_40955,N_42828);
and U48692 (N_48692,N_43133,N_44087);
nand U48693 (N_48693,N_40098,N_44638);
and U48694 (N_48694,N_42697,N_43033);
nand U48695 (N_48695,N_43167,N_44126);
or U48696 (N_48696,N_44164,N_42349);
or U48697 (N_48697,N_44774,N_42516);
nor U48698 (N_48698,N_41627,N_41448);
xnor U48699 (N_48699,N_42229,N_44633);
xnor U48700 (N_48700,N_43606,N_41972);
nor U48701 (N_48701,N_44573,N_44141);
and U48702 (N_48702,N_44939,N_42497);
xor U48703 (N_48703,N_42502,N_43286);
or U48704 (N_48704,N_42086,N_42928);
or U48705 (N_48705,N_44550,N_44415);
or U48706 (N_48706,N_41885,N_43669);
or U48707 (N_48707,N_42106,N_42903);
and U48708 (N_48708,N_41911,N_43142);
nand U48709 (N_48709,N_40059,N_40938);
and U48710 (N_48710,N_40000,N_41094);
nand U48711 (N_48711,N_42104,N_44151);
and U48712 (N_48712,N_44273,N_43563);
nand U48713 (N_48713,N_41320,N_40581);
or U48714 (N_48714,N_41910,N_40135);
nand U48715 (N_48715,N_41472,N_43546);
nand U48716 (N_48716,N_42372,N_40944);
nand U48717 (N_48717,N_42496,N_41780);
or U48718 (N_48718,N_40655,N_43871);
or U48719 (N_48719,N_42092,N_41034);
or U48720 (N_48720,N_43771,N_42482);
xnor U48721 (N_48721,N_44764,N_42320);
xor U48722 (N_48722,N_43551,N_44609);
and U48723 (N_48723,N_42435,N_44989);
and U48724 (N_48724,N_42429,N_42531);
or U48725 (N_48725,N_44250,N_42801);
nand U48726 (N_48726,N_43645,N_44910);
and U48727 (N_48727,N_44362,N_44974);
nand U48728 (N_48728,N_41688,N_43368);
or U48729 (N_48729,N_42872,N_41116);
nor U48730 (N_48730,N_42010,N_43270);
nand U48731 (N_48731,N_40889,N_40961);
nand U48732 (N_48732,N_41337,N_44704);
nand U48733 (N_48733,N_40997,N_41067);
or U48734 (N_48734,N_40370,N_42694);
and U48735 (N_48735,N_42185,N_41868);
or U48736 (N_48736,N_44555,N_41178);
and U48737 (N_48737,N_44763,N_41048);
nand U48738 (N_48738,N_42172,N_44009);
nor U48739 (N_48739,N_41257,N_41047);
and U48740 (N_48740,N_44007,N_43124);
and U48741 (N_48741,N_43704,N_42379);
nor U48742 (N_48742,N_41246,N_43770);
nand U48743 (N_48743,N_44149,N_41670);
xor U48744 (N_48744,N_41845,N_42677);
nand U48745 (N_48745,N_40014,N_40784);
or U48746 (N_48746,N_42169,N_44896);
xor U48747 (N_48747,N_44457,N_40212);
xnor U48748 (N_48748,N_43894,N_44728);
xor U48749 (N_48749,N_44051,N_40785);
and U48750 (N_48750,N_41426,N_44685);
and U48751 (N_48751,N_42389,N_40847);
nor U48752 (N_48752,N_43618,N_40844);
or U48753 (N_48753,N_44175,N_41769);
and U48754 (N_48754,N_43465,N_41609);
and U48755 (N_48755,N_44596,N_44878);
and U48756 (N_48756,N_43301,N_42537);
nand U48757 (N_48757,N_41323,N_40963);
or U48758 (N_48758,N_44229,N_43903);
xor U48759 (N_48759,N_41712,N_44964);
nor U48760 (N_48760,N_40023,N_43932);
and U48761 (N_48761,N_41137,N_43526);
nand U48762 (N_48762,N_41208,N_41115);
xnor U48763 (N_48763,N_42027,N_43124);
nor U48764 (N_48764,N_40076,N_40688);
xnor U48765 (N_48765,N_40296,N_43217);
xor U48766 (N_48766,N_43530,N_42017);
or U48767 (N_48767,N_40056,N_44381);
or U48768 (N_48768,N_43394,N_42695);
nor U48769 (N_48769,N_43799,N_40994);
xnor U48770 (N_48770,N_44474,N_43124);
xor U48771 (N_48771,N_42525,N_40853);
and U48772 (N_48772,N_43415,N_41937);
nand U48773 (N_48773,N_42941,N_44493);
and U48774 (N_48774,N_41209,N_43957);
xnor U48775 (N_48775,N_40287,N_42609);
and U48776 (N_48776,N_44597,N_42763);
or U48777 (N_48777,N_42677,N_42076);
nand U48778 (N_48778,N_42574,N_42885);
nand U48779 (N_48779,N_40698,N_44635);
and U48780 (N_48780,N_43669,N_44723);
and U48781 (N_48781,N_42672,N_40736);
and U48782 (N_48782,N_41485,N_42419);
nor U48783 (N_48783,N_42749,N_40344);
xor U48784 (N_48784,N_40988,N_44026);
or U48785 (N_48785,N_41766,N_41269);
and U48786 (N_48786,N_42177,N_41423);
nor U48787 (N_48787,N_42207,N_43708);
nor U48788 (N_48788,N_40633,N_43153);
xor U48789 (N_48789,N_40008,N_44503);
nand U48790 (N_48790,N_40911,N_43614);
xor U48791 (N_48791,N_44149,N_41235);
nor U48792 (N_48792,N_43277,N_40341);
xor U48793 (N_48793,N_43748,N_42206);
nor U48794 (N_48794,N_43472,N_40654);
nand U48795 (N_48795,N_44270,N_41263);
xnor U48796 (N_48796,N_43207,N_41927);
and U48797 (N_48797,N_41302,N_40070);
and U48798 (N_48798,N_44801,N_44019);
xnor U48799 (N_48799,N_40260,N_43442);
nor U48800 (N_48800,N_40455,N_40807);
nor U48801 (N_48801,N_42030,N_44811);
or U48802 (N_48802,N_40728,N_44162);
xnor U48803 (N_48803,N_43623,N_42996);
xor U48804 (N_48804,N_42588,N_40027);
nand U48805 (N_48805,N_40056,N_44588);
nand U48806 (N_48806,N_42680,N_42873);
nand U48807 (N_48807,N_43510,N_41187);
and U48808 (N_48808,N_41375,N_44714);
and U48809 (N_48809,N_42300,N_42723);
and U48810 (N_48810,N_42434,N_44308);
nand U48811 (N_48811,N_43763,N_42982);
nor U48812 (N_48812,N_41867,N_40310);
xor U48813 (N_48813,N_42502,N_43728);
and U48814 (N_48814,N_42449,N_43994);
xor U48815 (N_48815,N_42277,N_42622);
nand U48816 (N_48816,N_41934,N_40834);
and U48817 (N_48817,N_43863,N_42589);
nor U48818 (N_48818,N_41741,N_40988);
and U48819 (N_48819,N_44038,N_40718);
nor U48820 (N_48820,N_43845,N_40223);
nor U48821 (N_48821,N_42606,N_44717);
nand U48822 (N_48822,N_40281,N_43653);
and U48823 (N_48823,N_41036,N_42115);
nand U48824 (N_48824,N_44681,N_40313);
and U48825 (N_48825,N_41676,N_42872);
xor U48826 (N_48826,N_44451,N_41820);
nor U48827 (N_48827,N_42045,N_44757);
and U48828 (N_48828,N_40310,N_42420);
or U48829 (N_48829,N_41257,N_42023);
or U48830 (N_48830,N_44375,N_43028);
nor U48831 (N_48831,N_41576,N_42895);
nand U48832 (N_48832,N_40048,N_41130);
and U48833 (N_48833,N_41991,N_42153);
xnor U48834 (N_48834,N_43952,N_44094);
and U48835 (N_48835,N_40939,N_42559);
and U48836 (N_48836,N_42850,N_42275);
nor U48837 (N_48837,N_41533,N_42788);
nor U48838 (N_48838,N_40799,N_41907);
nand U48839 (N_48839,N_44993,N_43397);
nand U48840 (N_48840,N_40743,N_44078);
nor U48841 (N_48841,N_41826,N_40695);
and U48842 (N_48842,N_43331,N_44572);
or U48843 (N_48843,N_42960,N_42304);
nor U48844 (N_48844,N_42614,N_41414);
nor U48845 (N_48845,N_44455,N_43773);
nor U48846 (N_48846,N_43205,N_40656);
nand U48847 (N_48847,N_44301,N_44961);
and U48848 (N_48848,N_43245,N_40592);
and U48849 (N_48849,N_40693,N_42299);
nor U48850 (N_48850,N_41484,N_40976);
nor U48851 (N_48851,N_44098,N_42833);
or U48852 (N_48852,N_44310,N_40990);
and U48853 (N_48853,N_44818,N_40331);
xor U48854 (N_48854,N_43143,N_40229);
and U48855 (N_48855,N_43327,N_41825);
xor U48856 (N_48856,N_44240,N_42237);
xnor U48857 (N_48857,N_43423,N_40893);
xor U48858 (N_48858,N_43482,N_40249);
or U48859 (N_48859,N_42070,N_42156);
xor U48860 (N_48860,N_40584,N_40522);
nor U48861 (N_48861,N_41939,N_43579);
and U48862 (N_48862,N_44216,N_44671);
and U48863 (N_48863,N_43869,N_41324);
nor U48864 (N_48864,N_40309,N_44802);
xor U48865 (N_48865,N_42422,N_40804);
nor U48866 (N_48866,N_44596,N_41258);
nand U48867 (N_48867,N_40760,N_42644);
nor U48868 (N_48868,N_41904,N_43498);
xnor U48869 (N_48869,N_43953,N_44285);
xor U48870 (N_48870,N_43882,N_43873);
and U48871 (N_48871,N_41941,N_42206);
nor U48872 (N_48872,N_44277,N_40625);
and U48873 (N_48873,N_44771,N_40732);
nand U48874 (N_48874,N_44300,N_43971);
nor U48875 (N_48875,N_42061,N_41279);
nor U48876 (N_48876,N_40729,N_44244);
xor U48877 (N_48877,N_41179,N_43793);
and U48878 (N_48878,N_43767,N_40568);
nand U48879 (N_48879,N_43311,N_42286);
and U48880 (N_48880,N_44653,N_44161);
nand U48881 (N_48881,N_42646,N_42250);
or U48882 (N_48882,N_40992,N_42712);
and U48883 (N_48883,N_41793,N_41062);
xnor U48884 (N_48884,N_40418,N_44651);
and U48885 (N_48885,N_44459,N_44904);
nand U48886 (N_48886,N_44070,N_40961);
nand U48887 (N_48887,N_40310,N_42072);
or U48888 (N_48888,N_40114,N_44822);
xor U48889 (N_48889,N_42602,N_44006);
nand U48890 (N_48890,N_43731,N_41121);
and U48891 (N_48891,N_43829,N_41170);
nor U48892 (N_48892,N_44095,N_43755);
and U48893 (N_48893,N_44640,N_43515);
nor U48894 (N_48894,N_42368,N_44187);
nor U48895 (N_48895,N_42664,N_44838);
or U48896 (N_48896,N_43351,N_41746);
nand U48897 (N_48897,N_42195,N_42414);
nor U48898 (N_48898,N_40198,N_43554);
nand U48899 (N_48899,N_44372,N_40001);
or U48900 (N_48900,N_44076,N_44668);
nand U48901 (N_48901,N_40867,N_43458);
and U48902 (N_48902,N_41807,N_42413);
nand U48903 (N_48903,N_43728,N_40734);
xor U48904 (N_48904,N_42955,N_44040);
nand U48905 (N_48905,N_43216,N_40292);
and U48906 (N_48906,N_40969,N_44249);
nand U48907 (N_48907,N_44340,N_44032);
nor U48908 (N_48908,N_40474,N_40184);
and U48909 (N_48909,N_40725,N_41350);
nand U48910 (N_48910,N_41125,N_44422);
nor U48911 (N_48911,N_40104,N_44090);
or U48912 (N_48912,N_42160,N_40687);
and U48913 (N_48913,N_43537,N_41252);
or U48914 (N_48914,N_40158,N_44019);
and U48915 (N_48915,N_43718,N_44570);
nor U48916 (N_48916,N_43965,N_43328);
nand U48917 (N_48917,N_42241,N_44162);
and U48918 (N_48918,N_41753,N_43850);
nand U48919 (N_48919,N_43326,N_41771);
nand U48920 (N_48920,N_42927,N_43394);
nand U48921 (N_48921,N_44032,N_40906);
nand U48922 (N_48922,N_44212,N_41904);
xnor U48923 (N_48923,N_44354,N_42608);
nor U48924 (N_48924,N_41092,N_44129);
and U48925 (N_48925,N_42824,N_44213);
nand U48926 (N_48926,N_41051,N_41990);
or U48927 (N_48927,N_40620,N_43335);
nor U48928 (N_48928,N_41844,N_43637);
and U48929 (N_48929,N_42530,N_44717);
nor U48930 (N_48930,N_44309,N_41663);
and U48931 (N_48931,N_44090,N_42097);
nand U48932 (N_48932,N_40589,N_43078);
nand U48933 (N_48933,N_42089,N_42800);
nor U48934 (N_48934,N_43399,N_42861);
xor U48935 (N_48935,N_42764,N_42256);
or U48936 (N_48936,N_42165,N_40421);
nor U48937 (N_48937,N_43652,N_43297);
xor U48938 (N_48938,N_41944,N_43147);
xnor U48939 (N_48939,N_40204,N_41085);
nor U48940 (N_48940,N_43645,N_42659);
or U48941 (N_48941,N_43063,N_40864);
nor U48942 (N_48942,N_42468,N_40038);
xor U48943 (N_48943,N_42961,N_40292);
xor U48944 (N_48944,N_44634,N_40879);
or U48945 (N_48945,N_40527,N_43036);
and U48946 (N_48946,N_40792,N_44705);
nand U48947 (N_48947,N_42339,N_40171);
nand U48948 (N_48948,N_43684,N_41850);
and U48949 (N_48949,N_44997,N_41569);
and U48950 (N_48950,N_44679,N_40343);
nor U48951 (N_48951,N_41088,N_44727);
xor U48952 (N_48952,N_40319,N_42951);
nor U48953 (N_48953,N_42120,N_44981);
nor U48954 (N_48954,N_42007,N_43908);
xnor U48955 (N_48955,N_44117,N_40656);
nand U48956 (N_48956,N_44093,N_43060);
xor U48957 (N_48957,N_43612,N_41830);
and U48958 (N_48958,N_40849,N_40562);
or U48959 (N_48959,N_42964,N_41742);
nand U48960 (N_48960,N_42570,N_41063);
nor U48961 (N_48961,N_41799,N_42646);
or U48962 (N_48962,N_42980,N_41916);
or U48963 (N_48963,N_40610,N_40197);
or U48964 (N_48964,N_42247,N_42912);
and U48965 (N_48965,N_43505,N_40074);
nand U48966 (N_48966,N_41491,N_44565);
or U48967 (N_48967,N_40088,N_41480);
xor U48968 (N_48968,N_40012,N_40857);
and U48969 (N_48969,N_41851,N_44693);
nand U48970 (N_48970,N_44675,N_40319);
or U48971 (N_48971,N_41660,N_44276);
or U48972 (N_48972,N_41669,N_43644);
or U48973 (N_48973,N_44613,N_42658);
xor U48974 (N_48974,N_42951,N_42967);
nand U48975 (N_48975,N_41820,N_43754);
and U48976 (N_48976,N_44898,N_40769);
or U48977 (N_48977,N_41107,N_43222);
and U48978 (N_48978,N_44623,N_41396);
or U48979 (N_48979,N_42428,N_44422);
or U48980 (N_48980,N_43965,N_41728);
nand U48981 (N_48981,N_43026,N_40786);
and U48982 (N_48982,N_43309,N_44901);
xor U48983 (N_48983,N_41620,N_41374);
or U48984 (N_48984,N_42609,N_43254);
nand U48985 (N_48985,N_40571,N_42509);
or U48986 (N_48986,N_43757,N_44562);
or U48987 (N_48987,N_42456,N_41808);
or U48988 (N_48988,N_44980,N_43609);
or U48989 (N_48989,N_41874,N_44462);
xor U48990 (N_48990,N_40523,N_42531);
and U48991 (N_48991,N_41152,N_42509);
xor U48992 (N_48992,N_44935,N_41475);
nand U48993 (N_48993,N_43023,N_40634);
nor U48994 (N_48994,N_41568,N_42098);
nor U48995 (N_48995,N_40477,N_44690);
and U48996 (N_48996,N_44014,N_42664);
and U48997 (N_48997,N_44394,N_40029);
xor U48998 (N_48998,N_43537,N_42883);
xor U48999 (N_48999,N_40006,N_44397);
nor U49000 (N_49000,N_41297,N_42583);
or U49001 (N_49001,N_43021,N_41132);
or U49002 (N_49002,N_40678,N_42230);
or U49003 (N_49003,N_40627,N_43974);
nor U49004 (N_49004,N_43123,N_40201);
and U49005 (N_49005,N_42510,N_41554);
nor U49006 (N_49006,N_42061,N_41428);
nand U49007 (N_49007,N_42387,N_43682);
or U49008 (N_49008,N_43581,N_43949);
xnor U49009 (N_49009,N_41131,N_41333);
xor U49010 (N_49010,N_42430,N_43217);
nor U49011 (N_49011,N_44697,N_42312);
and U49012 (N_49012,N_42678,N_44252);
or U49013 (N_49013,N_44266,N_40893);
nand U49014 (N_49014,N_41510,N_40603);
nor U49015 (N_49015,N_43602,N_40241);
xnor U49016 (N_49016,N_41201,N_41250);
xnor U49017 (N_49017,N_41336,N_43048);
xnor U49018 (N_49018,N_42464,N_44317);
xor U49019 (N_49019,N_44446,N_40768);
nand U49020 (N_49020,N_44908,N_43042);
or U49021 (N_49021,N_42664,N_44804);
nor U49022 (N_49022,N_40860,N_41300);
nor U49023 (N_49023,N_41096,N_40561);
nor U49024 (N_49024,N_43572,N_44169);
and U49025 (N_49025,N_43590,N_43255);
nand U49026 (N_49026,N_43774,N_41666);
or U49027 (N_49027,N_40483,N_43839);
or U49028 (N_49028,N_44649,N_42409);
and U49029 (N_49029,N_42031,N_40899);
or U49030 (N_49030,N_41222,N_42055);
xor U49031 (N_49031,N_40147,N_44144);
or U49032 (N_49032,N_42090,N_40125);
or U49033 (N_49033,N_43723,N_44278);
nor U49034 (N_49034,N_43545,N_44341);
and U49035 (N_49035,N_43385,N_40452);
or U49036 (N_49036,N_40871,N_44478);
and U49037 (N_49037,N_43315,N_42037);
or U49038 (N_49038,N_42026,N_43352);
nand U49039 (N_49039,N_43079,N_41518);
xor U49040 (N_49040,N_44505,N_40013);
nand U49041 (N_49041,N_41067,N_43404);
nor U49042 (N_49042,N_42051,N_41736);
or U49043 (N_49043,N_44496,N_41364);
or U49044 (N_49044,N_43246,N_41002);
xor U49045 (N_49045,N_44615,N_41386);
nand U49046 (N_49046,N_40119,N_44704);
or U49047 (N_49047,N_44198,N_40711);
nor U49048 (N_49048,N_41678,N_42212);
or U49049 (N_49049,N_44716,N_44418);
nand U49050 (N_49050,N_42520,N_42692);
nor U49051 (N_49051,N_43848,N_41051);
and U49052 (N_49052,N_41914,N_42203);
and U49053 (N_49053,N_44374,N_44008);
xor U49054 (N_49054,N_42929,N_44872);
or U49055 (N_49055,N_43583,N_44260);
and U49056 (N_49056,N_44370,N_44910);
nor U49057 (N_49057,N_40390,N_41346);
or U49058 (N_49058,N_42967,N_40188);
xor U49059 (N_49059,N_43385,N_44817);
and U49060 (N_49060,N_42206,N_40590);
nor U49061 (N_49061,N_44545,N_43204);
xnor U49062 (N_49062,N_42814,N_44263);
xor U49063 (N_49063,N_43174,N_43027);
nor U49064 (N_49064,N_44928,N_43748);
and U49065 (N_49065,N_41025,N_40751);
or U49066 (N_49066,N_40029,N_41102);
or U49067 (N_49067,N_44753,N_43018);
xnor U49068 (N_49068,N_42930,N_40983);
nand U49069 (N_49069,N_40755,N_41042);
nor U49070 (N_49070,N_41002,N_40760);
or U49071 (N_49071,N_42582,N_42498);
xor U49072 (N_49072,N_41647,N_42275);
xor U49073 (N_49073,N_41881,N_42557);
or U49074 (N_49074,N_42678,N_40589);
nor U49075 (N_49075,N_40883,N_41877);
or U49076 (N_49076,N_43202,N_40330);
nand U49077 (N_49077,N_40716,N_43033);
xnor U49078 (N_49078,N_40752,N_42725);
and U49079 (N_49079,N_44599,N_43295);
nand U49080 (N_49080,N_40074,N_42310);
nand U49081 (N_49081,N_44617,N_41646);
nor U49082 (N_49082,N_44189,N_41366);
nand U49083 (N_49083,N_41196,N_40538);
xnor U49084 (N_49084,N_40286,N_44878);
and U49085 (N_49085,N_40092,N_41143);
or U49086 (N_49086,N_44923,N_40263);
and U49087 (N_49087,N_42755,N_43422);
nor U49088 (N_49088,N_44803,N_44485);
or U49089 (N_49089,N_41175,N_41177);
and U49090 (N_49090,N_44633,N_41840);
and U49091 (N_49091,N_40280,N_44108);
or U49092 (N_49092,N_40147,N_44552);
nand U49093 (N_49093,N_43106,N_43056);
and U49094 (N_49094,N_41674,N_41110);
xnor U49095 (N_49095,N_42924,N_44586);
xnor U49096 (N_49096,N_42133,N_42320);
nand U49097 (N_49097,N_42760,N_43276);
nand U49098 (N_49098,N_40925,N_41605);
xor U49099 (N_49099,N_40668,N_42055);
nor U49100 (N_49100,N_44946,N_42213);
nor U49101 (N_49101,N_43446,N_40588);
nor U49102 (N_49102,N_42167,N_43203);
nand U49103 (N_49103,N_43018,N_40527);
xor U49104 (N_49104,N_42303,N_43576);
nor U49105 (N_49105,N_43609,N_43604);
nand U49106 (N_49106,N_40731,N_42647);
nand U49107 (N_49107,N_43404,N_42178);
nor U49108 (N_49108,N_43557,N_40744);
nand U49109 (N_49109,N_44254,N_41121);
nor U49110 (N_49110,N_44949,N_43866);
nand U49111 (N_49111,N_43447,N_43370);
nor U49112 (N_49112,N_42009,N_42800);
nand U49113 (N_49113,N_41435,N_43491);
xor U49114 (N_49114,N_41566,N_40959);
nor U49115 (N_49115,N_40074,N_40933);
xnor U49116 (N_49116,N_40543,N_43099);
nor U49117 (N_49117,N_43798,N_40363);
and U49118 (N_49118,N_42069,N_43166);
or U49119 (N_49119,N_40618,N_41237);
or U49120 (N_49120,N_43720,N_44767);
nand U49121 (N_49121,N_41671,N_40524);
and U49122 (N_49122,N_42966,N_42993);
nor U49123 (N_49123,N_42917,N_43947);
nand U49124 (N_49124,N_42725,N_41987);
nand U49125 (N_49125,N_44304,N_42545);
nand U49126 (N_49126,N_40480,N_41582);
nor U49127 (N_49127,N_43592,N_43909);
nand U49128 (N_49128,N_42520,N_41816);
and U49129 (N_49129,N_41820,N_41126);
nor U49130 (N_49130,N_42425,N_43320);
xor U49131 (N_49131,N_44978,N_40897);
nor U49132 (N_49132,N_43754,N_44100);
xnor U49133 (N_49133,N_40058,N_42803);
or U49134 (N_49134,N_41139,N_42811);
nand U49135 (N_49135,N_43174,N_40117);
and U49136 (N_49136,N_42454,N_41270);
nor U49137 (N_49137,N_41445,N_42659);
and U49138 (N_49138,N_40796,N_44554);
nand U49139 (N_49139,N_43164,N_43240);
or U49140 (N_49140,N_44364,N_42203);
nor U49141 (N_49141,N_43661,N_44827);
nand U49142 (N_49142,N_44419,N_40711);
and U49143 (N_49143,N_40102,N_40981);
and U49144 (N_49144,N_40214,N_43236);
nor U49145 (N_49145,N_42956,N_40808);
or U49146 (N_49146,N_40399,N_42556);
and U49147 (N_49147,N_42884,N_42379);
xnor U49148 (N_49148,N_43550,N_41306);
xor U49149 (N_49149,N_43491,N_42905);
xor U49150 (N_49150,N_42877,N_44734);
and U49151 (N_49151,N_40585,N_44139);
nand U49152 (N_49152,N_41431,N_42140);
and U49153 (N_49153,N_44537,N_43558);
xnor U49154 (N_49154,N_40560,N_44529);
and U49155 (N_49155,N_40961,N_43323);
nand U49156 (N_49156,N_42218,N_41835);
and U49157 (N_49157,N_41959,N_44804);
or U49158 (N_49158,N_44984,N_44747);
nor U49159 (N_49159,N_42477,N_42341);
xor U49160 (N_49160,N_44816,N_40767);
and U49161 (N_49161,N_42807,N_42001);
nor U49162 (N_49162,N_41538,N_43608);
and U49163 (N_49163,N_43874,N_44892);
and U49164 (N_49164,N_40026,N_43540);
or U49165 (N_49165,N_40334,N_41753);
xnor U49166 (N_49166,N_41258,N_41867);
nor U49167 (N_49167,N_40012,N_44957);
or U49168 (N_49168,N_44265,N_42232);
or U49169 (N_49169,N_44710,N_41432);
xnor U49170 (N_49170,N_43568,N_41813);
and U49171 (N_49171,N_41853,N_44950);
nand U49172 (N_49172,N_42036,N_44809);
nor U49173 (N_49173,N_44280,N_40297);
or U49174 (N_49174,N_43266,N_43071);
nor U49175 (N_49175,N_43049,N_42639);
or U49176 (N_49176,N_40369,N_43202);
or U49177 (N_49177,N_41459,N_42321);
nand U49178 (N_49178,N_41167,N_40474);
or U49179 (N_49179,N_41482,N_41090);
and U49180 (N_49180,N_41659,N_43065);
nand U49181 (N_49181,N_43818,N_43927);
nor U49182 (N_49182,N_44239,N_41426);
and U49183 (N_49183,N_41954,N_41228);
nor U49184 (N_49184,N_41814,N_44008);
and U49185 (N_49185,N_40125,N_44341);
or U49186 (N_49186,N_42496,N_40609);
nor U49187 (N_49187,N_41607,N_42552);
nand U49188 (N_49188,N_44469,N_42836);
xor U49189 (N_49189,N_44380,N_43216);
xor U49190 (N_49190,N_44293,N_42799);
nor U49191 (N_49191,N_43810,N_44706);
xor U49192 (N_49192,N_42897,N_42637);
nor U49193 (N_49193,N_43256,N_42255);
and U49194 (N_49194,N_41225,N_41037);
nor U49195 (N_49195,N_44414,N_44036);
or U49196 (N_49196,N_41058,N_44837);
xor U49197 (N_49197,N_42185,N_44302);
xnor U49198 (N_49198,N_42804,N_44578);
nor U49199 (N_49199,N_41219,N_42230);
and U49200 (N_49200,N_42298,N_41249);
nand U49201 (N_49201,N_43285,N_43675);
nand U49202 (N_49202,N_43977,N_41561);
and U49203 (N_49203,N_42568,N_40459);
xor U49204 (N_49204,N_42881,N_43583);
nand U49205 (N_49205,N_43295,N_43185);
nand U49206 (N_49206,N_42970,N_43047);
xor U49207 (N_49207,N_44436,N_44292);
xor U49208 (N_49208,N_43157,N_42428);
xor U49209 (N_49209,N_44697,N_42320);
nor U49210 (N_49210,N_42084,N_44010);
nand U49211 (N_49211,N_40907,N_44074);
or U49212 (N_49212,N_42256,N_40609);
nand U49213 (N_49213,N_44848,N_40867);
or U49214 (N_49214,N_43749,N_40442);
and U49215 (N_49215,N_42370,N_42828);
or U49216 (N_49216,N_42925,N_42129);
xor U49217 (N_49217,N_44446,N_42701);
xnor U49218 (N_49218,N_40468,N_40860);
or U49219 (N_49219,N_40687,N_42099);
nand U49220 (N_49220,N_44788,N_40361);
and U49221 (N_49221,N_44430,N_42759);
nor U49222 (N_49222,N_41015,N_43659);
and U49223 (N_49223,N_42251,N_41430);
xnor U49224 (N_49224,N_42440,N_41316);
and U49225 (N_49225,N_42740,N_44404);
and U49226 (N_49226,N_43854,N_44938);
and U49227 (N_49227,N_44242,N_44185);
or U49228 (N_49228,N_44760,N_42466);
and U49229 (N_49229,N_44668,N_41684);
or U49230 (N_49230,N_44582,N_42852);
xor U49231 (N_49231,N_40604,N_41933);
or U49232 (N_49232,N_42808,N_40096);
xor U49233 (N_49233,N_40569,N_41818);
or U49234 (N_49234,N_44652,N_42335);
nand U49235 (N_49235,N_42994,N_40753);
and U49236 (N_49236,N_41841,N_41351);
or U49237 (N_49237,N_43534,N_41697);
nor U49238 (N_49238,N_40299,N_40877);
xnor U49239 (N_49239,N_44685,N_41362);
or U49240 (N_49240,N_44816,N_42910);
nor U49241 (N_49241,N_43157,N_44409);
nand U49242 (N_49242,N_44037,N_42097);
nor U49243 (N_49243,N_41412,N_44053);
or U49244 (N_49244,N_42065,N_40599);
nand U49245 (N_49245,N_44855,N_41097);
xnor U49246 (N_49246,N_41944,N_42337);
and U49247 (N_49247,N_41161,N_41467);
nor U49248 (N_49248,N_41164,N_41438);
nand U49249 (N_49249,N_40327,N_40049);
xnor U49250 (N_49250,N_41959,N_41464);
xor U49251 (N_49251,N_44255,N_44935);
nand U49252 (N_49252,N_41054,N_42187);
and U49253 (N_49253,N_40496,N_40775);
nand U49254 (N_49254,N_44253,N_43166);
nor U49255 (N_49255,N_41289,N_44372);
xnor U49256 (N_49256,N_40917,N_43780);
nor U49257 (N_49257,N_44943,N_42821);
nor U49258 (N_49258,N_42753,N_42757);
or U49259 (N_49259,N_40350,N_41376);
nand U49260 (N_49260,N_43152,N_43147);
nand U49261 (N_49261,N_42408,N_43694);
nand U49262 (N_49262,N_43894,N_41757);
xnor U49263 (N_49263,N_40893,N_44907);
or U49264 (N_49264,N_40241,N_42162);
nor U49265 (N_49265,N_44033,N_44414);
xnor U49266 (N_49266,N_41331,N_42768);
xor U49267 (N_49267,N_41222,N_40374);
nand U49268 (N_49268,N_44915,N_41652);
or U49269 (N_49269,N_41376,N_43816);
nor U49270 (N_49270,N_43565,N_40889);
nand U49271 (N_49271,N_42777,N_43446);
nor U49272 (N_49272,N_44719,N_43024);
or U49273 (N_49273,N_42827,N_41421);
or U49274 (N_49274,N_41573,N_41524);
nor U49275 (N_49275,N_42715,N_41186);
xor U49276 (N_49276,N_42516,N_44863);
or U49277 (N_49277,N_44986,N_44304);
nor U49278 (N_49278,N_43561,N_42847);
xor U49279 (N_49279,N_40474,N_41027);
nand U49280 (N_49280,N_43305,N_42042);
nor U49281 (N_49281,N_41049,N_42426);
nor U49282 (N_49282,N_43528,N_41801);
and U49283 (N_49283,N_41559,N_40670);
nor U49284 (N_49284,N_42121,N_41868);
nand U49285 (N_49285,N_44342,N_42614);
or U49286 (N_49286,N_42478,N_41599);
xnor U49287 (N_49287,N_43890,N_42758);
xor U49288 (N_49288,N_40344,N_42566);
xor U49289 (N_49289,N_43780,N_41785);
xnor U49290 (N_49290,N_43173,N_41673);
or U49291 (N_49291,N_43744,N_41758);
xnor U49292 (N_49292,N_43340,N_43231);
and U49293 (N_49293,N_43019,N_40797);
and U49294 (N_49294,N_43975,N_44844);
or U49295 (N_49295,N_44228,N_43863);
and U49296 (N_49296,N_40175,N_44012);
or U49297 (N_49297,N_40156,N_42740);
or U49298 (N_49298,N_44469,N_42493);
and U49299 (N_49299,N_42856,N_41830);
nand U49300 (N_49300,N_41818,N_41544);
xnor U49301 (N_49301,N_42156,N_44024);
and U49302 (N_49302,N_41240,N_41981);
and U49303 (N_49303,N_43546,N_42712);
nor U49304 (N_49304,N_41299,N_40087);
nor U49305 (N_49305,N_44977,N_43709);
nand U49306 (N_49306,N_42272,N_40560);
and U49307 (N_49307,N_40706,N_41882);
nand U49308 (N_49308,N_43096,N_44995);
xor U49309 (N_49309,N_42274,N_44464);
nor U49310 (N_49310,N_40841,N_40603);
or U49311 (N_49311,N_40941,N_43440);
nor U49312 (N_49312,N_40724,N_42657);
xnor U49313 (N_49313,N_44566,N_41413);
or U49314 (N_49314,N_44843,N_43408);
nor U49315 (N_49315,N_43818,N_40507);
nor U49316 (N_49316,N_43211,N_40972);
xnor U49317 (N_49317,N_44687,N_40879);
nand U49318 (N_49318,N_41721,N_40345);
and U49319 (N_49319,N_44979,N_44946);
nand U49320 (N_49320,N_43439,N_44379);
nand U49321 (N_49321,N_41221,N_40031);
or U49322 (N_49322,N_43783,N_42565);
and U49323 (N_49323,N_41305,N_44143);
nand U49324 (N_49324,N_43833,N_44475);
nor U49325 (N_49325,N_41282,N_40809);
and U49326 (N_49326,N_41755,N_40436);
and U49327 (N_49327,N_44875,N_44011);
xnor U49328 (N_49328,N_44485,N_42259);
nand U49329 (N_49329,N_44114,N_44833);
or U49330 (N_49330,N_41293,N_40823);
nor U49331 (N_49331,N_41981,N_43078);
xor U49332 (N_49332,N_40891,N_44243);
nor U49333 (N_49333,N_40172,N_40414);
xor U49334 (N_49334,N_40352,N_41289);
and U49335 (N_49335,N_42351,N_42905);
nand U49336 (N_49336,N_42089,N_40351);
and U49337 (N_49337,N_43977,N_41830);
or U49338 (N_49338,N_42324,N_43234);
xor U49339 (N_49339,N_40703,N_40538);
and U49340 (N_49340,N_41159,N_43035);
or U49341 (N_49341,N_41807,N_40401);
nand U49342 (N_49342,N_44918,N_40153);
nand U49343 (N_49343,N_42129,N_40512);
nor U49344 (N_49344,N_40320,N_41399);
nor U49345 (N_49345,N_43016,N_40227);
or U49346 (N_49346,N_44703,N_42072);
and U49347 (N_49347,N_42779,N_42962);
nand U49348 (N_49348,N_44438,N_42921);
and U49349 (N_49349,N_44674,N_43415);
and U49350 (N_49350,N_41152,N_44628);
xor U49351 (N_49351,N_40449,N_42754);
or U49352 (N_49352,N_42061,N_43744);
nor U49353 (N_49353,N_40467,N_42238);
nor U49354 (N_49354,N_43553,N_41376);
or U49355 (N_49355,N_42861,N_42542);
nand U49356 (N_49356,N_42858,N_42885);
and U49357 (N_49357,N_40263,N_43776);
or U49358 (N_49358,N_44696,N_44013);
or U49359 (N_49359,N_43316,N_44136);
or U49360 (N_49360,N_41507,N_42506);
xnor U49361 (N_49361,N_41089,N_42099);
and U49362 (N_49362,N_41954,N_42681);
xnor U49363 (N_49363,N_41913,N_40549);
and U49364 (N_49364,N_43323,N_41793);
nand U49365 (N_49365,N_42005,N_40969);
nand U49366 (N_49366,N_42633,N_42851);
xor U49367 (N_49367,N_40096,N_42875);
nand U49368 (N_49368,N_42351,N_44414);
nand U49369 (N_49369,N_40349,N_40337);
and U49370 (N_49370,N_44628,N_44395);
or U49371 (N_49371,N_43547,N_41443);
and U49372 (N_49372,N_40906,N_44921);
nor U49373 (N_49373,N_41099,N_43292);
or U49374 (N_49374,N_44734,N_43117);
xor U49375 (N_49375,N_42196,N_40808);
or U49376 (N_49376,N_44696,N_40100);
and U49377 (N_49377,N_44542,N_40493);
nand U49378 (N_49378,N_43396,N_40548);
nor U49379 (N_49379,N_43902,N_44197);
nor U49380 (N_49380,N_41903,N_41283);
or U49381 (N_49381,N_42541,N_40791);
and U49382 (N_49382,N_42432,N_42335);
nand U49383 (N_49383,N_41841,N_43174);
or U49384 (N_49384,N_44853,N_44673);
nor U49385 (N_49385,N_41803,N_41560);
and U49386 (N_49386,N_43705,N_44081);
nand U49387 (N_49387,N_41459,N_42480);
xor U49388 (N_49388,N_44080,N_40633);
and U49389 (N_49389,N_42202,N_42999);
nand U49390 (N_49390,N_41895,N_41489);
and U49391 (N_49391,N_43307,N_42299);
and U49392 (N_49392,N_43636,N_41585);
nor U49393 (N_49393,N_40905,N_42566);
xnor U49394 (N_49394,N_44301,N_40375);
and U49395 (N_49395,N_44394,N_41641);
xor U49396 (N_49396,N_43628,N_41348);
or U49397 (N_49397,N_42970,N_40037);
or U49398 (N_49398,N_42322,N_41739);
nand U49399 (N_49399,N_44201,N_43564);
and U49400 (N_49400,N_40783,N_43542);
or U49401 (N_49401,N_41370,N_43855);
xor U49402 (N_49402,N_40224,N_42272);
nor U49403 (N_49403,N_43768,N_40188);
nor U49404 (N_49404,N_40926,N_42734);
or U49405 (N_49405,N_44191,N_44900);
xnor U49406 (N_49406,N_40199,N_40695);
nor U49407 (N_49407,N_41400,N_44298);
or U49408 (N_49408,N_41338,N_43664);
xnor U49409 (N_49409,N_43431,N_40431);
or U49410 (N_49410,N_41404,N_42844);
and U49411 (N_49411,N_41530,N_44899);
xnor U49412 (N_49412,N_43511,N_41754);
and U49413 (N_49413,N_40735,N_43400);
or U49414 (N_49414,N_44365,N_44471);
nand U49415 (N_49415,N_44361,N_43634);
or U49416 (N_49416,N_40364,N_40575);
or U49417 (N_49417,N_40020,N_40933);
nor U49418 (N_49418,N_41135,N_40620);
nor U49419 (N_49419,N_41459,N_42487);
nand U49420 (N_49420,N_43047,N_40924);
or U49421 (N_49421,N_43251,N_42208);
nand U49422 (N_49422,N_40522,N_40088);
nor U49423 (N_49423,N_43431,N_43289);
xnor U49424 (N_49424,N_40953,N_42431);
xor U49425 (N_49425,N_41777,N_40301);
xnor U49426 (N_49426,N_44592,N_40250);
nand U49427 (N_49427,N_44058,N_44730);
or U49428 (N_49428,N_40595,N_44278);
xor U49429 (N_49429,N_44055,N_41566);
or U49430 (N_49430,N_40865,N_40467);
and U49431 (N_49431,N_40814,N_44063);
nand U49432 (N_49432,N_42319,N_42539);
or U49433 (N_49433,N_40063,N_42098);
nor U49434 (N_49434,N_41094,N_44437);
and U49435 (N_49435,N_42138,N_40463);
nand U49436 (N_49436,N_42709,N_40778);
or U49437 (N_49437,N_43786,N_44589);
and U49438 (N_49438,N_42128,N_43621);
xor U49439 (N_49439,N_42557,N_43760);
or U49440 (N_49440,N_44534,N_44370);
nand U49441 (N_49441,N_44212,N_42718);
xnor U49442 (N_49442,N_40803,N_40746);
nor U49443 (N_49443,N_42207,N_43929);
nand U49444 (N_49444,N_42114,N_44315);
or U49445 (N_49445,N_41429,N_43341);
xor U49446 (N_49446,N_44974,N_42805);
or U49447 (N_49447,N_40015,N_40082);
and U49448 (N_49448,N_43119,N_41202);
and U49449 (N_49449,N_41337,N_43352);
and U49450 (N_49450,N_42484,N_44865);
and U49451 (N_49451,N_43278,N_43123);
xnor U49452 (N_49452,N_44409,N_40460);
or U49453 (N_49453,N_43048,N_41065);
nand U49454 (N_49454,N_43279,N_42805);
xor U49455 (N_49455,N_42405,N_44089);
xor U49456 (N_49456,N_42283,N_43704);
nor U49457 (N_49457,N_42989,N_41606);
nand U49458 (N_49458,N_42071,N_42816);
and U49459 (N_49459,N_41998,N_41001);
nor U49460 (N_49460,N_40162,N_42971);
xor U49461 (N_49461,N_40848,N_42285);
nor U49462 (N_49462,N_40949,N_44267);
and U49463 (N_49463,N_41738,N_42799);
xor U49464 (N_49464,N_44627,N_40278);
nand U49465 (N_49465,N_44018,N_42870);
and U49466 (N_49466,N_41729,N_44647);
xnor U49467 (N_49467,N_43973,N_43526);
and U49468 (N_49468,N_42579,N_42173);
nor U49469 (N_49469,N_41220,N_43797);
nor U49470 (N_49470,N_43383,N_42059);
xnor U49471 (N_49471,N_43686,N_44867);
xor U49472 (N_49472,N_44103,N_42978);
and U49473 (N_49473,N_43461,N_40426);
and U49474 (N_49474,N_41628,N_42305);
or U49475 (N_49475,N_40028,N_44614);
and U49476 (N_49476,N_42583,N_44912);
or U49477 (N_49477,N_40728,N_43925);
xor U49478 (N_49478,N_41936,N_43679);
nand U49479 (N_49479,N_44512,N_42026);
and U49480 (N_49480,N_41711,N_44317);
and U49481 (N_49481,N_42444,N_40420);
nand U49482 (N_49482,N_44642,N_40417);
and U49483 (N_49483,N_40197,N_42270);
nand U49484 (N_49484,N_40945,N_40292);
nor U49485 (N_49485,N_43631,N_44574);
and U49486 (N_49486,N_41665,N_40499);
xnor U49487 (N_49487,N_40650,N_41486);
or U49488 (N_49488,N_40807,N_41733);
xor U49489 (N_49489,N_40069,N_42121);
nand U49490 (N_49490,N_42786,N_40974);
nand U49491 (N_49491,N_43549,N_42972);
xnor U49492 (N_49492,N_43429,N_40629);
nand U49493 (N_49493,N_42341,N_41668);
or U49494 (N_49494,N_41048,N_40489);
xnor U49495 (N_49495,N_42542,N_42851);
nand U49496 (N_49496,N_40869,N_41291);
nor U49497 (N_49497,N_42768,N_43788);
or U49498 (N_49498,N_44966,N_44768);
xnor U49499 (N_49499,N_42311,N_44100);
xnor U49500 (N_49500,N_40145,N_44808);
nand U49501 (N_49501,N_44904,N_41001);
and U49502 (N_49502,N_44781,N_44790);
or U49503 (N_49503,N_41371,N_42811);
and U49504 (N_49504,N_41346,N_44464);
or U49505 (N_49505,N_41914,N_43344);
or U49506 (N_49506,N_43747,N_40185);
xor U49507 (N_49507,N_42588,N_41629);
xor U49508 (N_49508,N_43935,N_41378);
nand U49509 (N_49509,N_44087,N_40473);
nand U49510 (N_49510,N_43568,N_43886);
xor U49511 (N_49511,N_42490,N_42424);
xnor U49512 (N_49512,N_44302,N_41424);
nand U49513 (N_49513,N_40087,N_41389);
or U49514 (N_49514,N_40664,N_43394);
nor U49515 (N_49515,N_43023,N_42913);
xnor U49516 (N_49516,N_43904,N_40497);
or U49517 (N_49517,N_40334,N_43111);
xnor U49518 (N_49518,N_44325,N_44542);
and U49519 (N_49519,N_41278,N_44474);
or U49520 (N_49520,N_40741,N_44798);
nand U49521 (N_49521,N_44244,N_41140);
xnor U49522 (N_49522,N_42076,N_44823);
or U49523 (N_49523,N_42121,N_43726);
nor U49524 (N_49524,N_44812,N_41416);
xor U49525 (N_49525,N_44024,N_43305);
or U49526 (N_49526,N_42164,N_44998);
xnor U49527 (N_49527,N_40715,N_41541);
nor U49528 (N_49528,N_43986,N_41120);
or U49529 (N_49529,N_40664,N_41040);
nand U49530 (N_49530,N_43991,N_41445);
or U49531 (N_49531,N_40854,N_43400);
nand U49532 (N_49532,N_42592,N_44274);
and U49533 (N_49533,N_42360,N_40342);
nor U49534 (N_49534,N_44966,N_42806);
and U49535 (N_49535,N_44829,N_40335);
nor U49536 (N_49536,N_43782,N_44687);
and U49537 (N_49537,N_44407,N_44995);
xor U49538 (N_49538,N_40820,N_43580);
or U49539 (N_49539,N_42858,N_43570);
nand U49540 (N_49540,N_44032,N_44921);
nor U49541 (N_49541,N_40894,N_41469);
nand U49542 (N_49542,N_44675,N_43868);
xnor U49543 (N_49543,N_44628,N_40241);
nand U49544 (N_49544,N_44744,N_40218);
xor U49545 (N_49545,N_44867,N_40511);
nand U49546 (N_49546,N_42852,N_42466);
or U49547 (N_49547,N_41636,N_44546);
xnor U49548 (N_49548,N_43304,N_44266);
nor U49549 (N_49549,N_42498,N_43574);
xnor U49550 (N_49550,N_44812,N_41591);
or U49551 (N_49551,N_44485,N_42018);
or U49552 (N_49552,N_43275,N_44123);
and U49553 (N_49553,N_41037,N_43883);
nor U49554 (N_49554,N_43437,N_42233);
or U49555 (N_49555,N_44088,N_41771);
or U49556 (N_49556,N_42671,N_42484);
xor U49557 (N_49557,N_41469,N_40076);
nand U49558 (N_49558,N_43120,N_41625);
xnor U49559 (N_49559,N_44252,N_41714);
xor U49560 (N_49560,N_40254,N_40985);
xnor U49561 (N_49561,N_41516,N_43698);
or U49562 (N_49562,N_40680,N_42186);
and U49563 (N_49563,N_42818,N_43335);
and U49564 (N_49564,N_43822,N_43367);
nor U49565 (N_49565,N_42808,N_40742);
and U49566 (N_49566,N_42790,N_44213);
nor U49567 (N_49567,N_41146,N_43010);
nand U49568 (N_49568,N_42800,N_44085);
nand U49569 (N_49569,N_41053,N_41250);
nand U49570 (N_49570,N_43606,N_44433);
and U49571 (N_49571,N_40931,N_42250);
xnor U49572 (N_49572,N_40245,N_43982);
xor U49573 (N_49573,N_40331,N_42131);
or U49574 (N_49574,N_40766,N_43821);
nand U49575 (N_49575,N_41216,N_43267);
nor U49576 (N_49576,N_40835,N_44063);
or U49577 (N_49577,N_41793,N_41457);
nand U49578 (N_49578,N_40488,N_42523);
and U49579 (N_49579,N_40629,N_42452);
xnor U49580 (N_49580,N_44621,N_42513);
nor U49581 (N_49581,N_41881,N_41424);
and U49582 (N_49582,N_44659,N_40643);
nand U49583 (N_49583,N_40690,N_41441);
or U49584 (N_49584,N_43869,N_43961);
and U49585 (N_49585,N_42944,N_43916);
xor U49586 (N_49586,N_40424,N_43868);
or U49587 (N_49587,N_40866,N_44466);
or U49588 (N_49588,N_40853,N_41505);
nand U49589 (N_49589,N_42533,N_42621);
nor U49590 (N_49590,N_44631,N_43537);
nor U49591 (N_49591,N_43479,N_44491);
and U49592 (N_49592,N_44145,N_42595);
or U49593 (N_49593,N_44018,N_42509);
xor U49594 (N_49594,N_43940,N_44420);
nor U49595 (N_49595,N_42791,N_43180);
xor U49596 (N_49596,N_43525,N_41458);
nor U49597 (N_49597,N_44358,N_42221);
and U49598 (N_49598,N_42891,N_42764);
xnor U49599 (N_49599,N_41820,N_43753);
nor U49600 (N_49600,N_41247,N_42313);
nand U49601 (N_49601,N_42598,N_41261);
and U49602 (N_49602,N_40692,N_40084);
and U49603 (N_49603,N_44075,N_43388);
xnor U49604 (N_49604,N_41734,N_43219);
and U49605 (N_49605,N_43157,N_44588);
and U49606 (N_49606,N_41658,N_41398);
nor U49607 (N_49607,N_44155,N_42518);
xnor U49608 (N_49608,N_44485,N_40925);
xor U49609 (N_49609,N_40939,N_43206);
nor U49610 (N_49610,N_40260,N_43469);
xor U49611 (N_49611,N_41657,N_40918);
nor U49612 (N_49612,N_44451,N_41456);
xnor U49613 (N_49613,N_40472,N_40459);
or U49614 (N_49614,N_40536,N_44832);
nor U49615 (N_49615,N_43850,N_43767);
xor U49616 (N_49616,N_44684,N_43112);
and U49617 (N_49617,N_43394,N_43822);
and U49618 (N_49618,N_42836,N_40263);
nand U49619 (N_49619,N_40120,N_42885);
xnor U49620 (N_49620,N_42114,N_41135);
or U49621 (N_49621,N_41441,N_40249);
and U49622 (N_49622,N_43241,N_41540);
xor U49623 (N_49623,N_43862,N_40287);
nor U49624 (N_49624,N_43352,N_44955);
nor U49625 (N_49625,N_42953,N_44884);
nand U49626 (N_49626,N_43565,N_40815);
xnor U49627 (N_49627,N_40454,N_43153);
xor U49628 (N_49628,N_40194,N_41111);
nand U49629 (N_49629,N_42567,N_41544);
nor U49630 (N_49630,N_40371,N_41569);
and U49631 (N_49631,N_40897,N_44362);
xor U49632 (N_49632,N_42715,N_43744);
or U49633 (N_49633,N_43714,N_41411);
and U49634 (N_49634,N_44066,N_42316);
nor U49635 (N_49635,N_44631,N_44835);
xor U49636 (N_49636,N_42137,N_40075);
xnor U49637 (N_49637,N_42032,N_42522);
and U49638 (N_49638,N_41829,N_40749);
or U49639 (N_49639,N_41024,N_41416);
nand U49640 (N_49640,N_41556,N_40752);
xnor U49641 (N_49641,N_42336,N_42539);
nor U49642 (N_49642,N_44605,N_44353);
nand U49643 (N_49643,N_40715,N_41680);
and U49644 (N_49644,N_43538,N_43635);
nand U49645 (N_49645,N_41422,N_42078);
nor U49646 (N_49646,N_44806,N_41644);
or U49647 (N_49647,N_42096,N_43198);
nor U49648 (N_49648,N_43247,N_43508);
nand U49649 (N_49649,N_42880,N_40505);
xor U49650 (N_49650,N_44942,N_43895);
xor U49651 (N_49651,N_40982,N_40640);
or U49652 (N_49652,N_43382,N_43534);
nor U49653 (N_49653,N_40375,N_40776);
and U49654 (N_49654,N_44759,N_43597);
and U49655 (N_49655,N_40557,N_44918);
xor U49656 (N_49656,N_41797,N_44817);
and U49657 (N_49657,N_42742,N_43752);
nand U49658 (N_49658,N_40075,N_43109);
nor U49659 (N_49659,N_44201,N_44962);
or U49660 (N_49660,N_44659,N_42661);
nand U49661 (N_49661,N_41040,N_40246);
and U49662 (N_49662,N_44798,N_40373);
and U49663 (N_49663,N_44172,N_40930);
nand U49664 (N_49664,N_41129,N_41430);
and U49665 (N_49665,N_41430,N_43602);
and U49666 (N_49666,N_42151,N_44489);
nor U49667 (N_49667,N_43902,N_44490);
xnor U49668 (N_49668,N_42234,N_43603);
xor U49669 (N_49669,N_43373,N_42108);
and U49670 (N_49670,N_42407,N_41468);
or U49671 (N_49671,N_43144,N_44388);
and U49672 (N_49672,N_41147,N_42134);
and U49673 (N_49673,N_44459,N_42819);
nand U49674 (N_49674,N_42107,N_44817);
nor U49675 (N_49675,N_40665,N_41917);
xnor U49676 (N_49676,N_40588,N_42538);
nand U49677 (N_49677,N_40580,N_44539);
or U49678 (N_49678,N_40528,N_44071);
or U49679 (N_49679,N_44535,N_43702);
or U49680 (N_49680,N_44080,N_40691);
or U49681 (N_49681,N_44154,N_40172);
nand U49682 (N_49682,N_41627,N_41923);
and U49683 (N_49683,N_43892,N_41370);
xnor U49684 (N_49684,N_40105,N_43689);
and U49685 (N_49685,N_43746,N_43443);
and U49686 (N_49686,N_44341,N_44710);
xor U49687 (N_49687,N_44048,N_42794);
xor U49688 (N_49688,N_43397,N_43813);
or U49689 (N_49689,N_43390,N_40684);
nor U49690 (N_49690,N_42639,N_41333);
and U49691 (N_49691,N_43934,N_43429);
or U49692 (N_49692,N_40314,N_40183);
and U49693 (N_49693,N_41612,N_43655);
nand U49694 (N_49694,N_44773,N_44590);
and U49695 (N_49695,N_41118,N_42582);
or U49696 (N_49696,N_41165,N_43675);
xor U49697 (N_49697,N_40796,N_41917);
or U49698 (N_49698,N_40438,N_41648);
nand U49699 (N_49699,N_44276,N_40608);
and U49700 (N_49700,N_44097,N_40564);
or U49701 (N_49701,N_43757,N_42418);
nor U49702 (N_49702,N_44579,N_41917);
or U49703 (N_49703,N_42158,N_40731);
nor U49704 (N_49704,N_41677,N_44055);
and U49705 (N_49705,N_41555,N_42686);
nor U49706 (N_49706,N_40110,N_41106);
and U49707 (N_49707,N_41673,N_40011);
xor U49708 (N_49708,N_42784,N_42316);
or U49709 (N_49709,N_42664,N_41965);
and U49710 (N_49710,N_43141,N_41128);
and U49711 (N_49711,N_43409,N_44388);
nor U49712 (N_49712,N_42879,N_43417);
nand U49713 (N_49713,N_43014,N_44380);
nand U49714 (N_49714,N_43982,N_42501);
nand U49715 (N_49715,N_42540,N_41759);
xnor U49716 (N_49716,N_43008,N_44116);
and U49717 (N_49717,N_43975,N_44711);
and U49718 (N_49718,N_44293,N_42443);
and U49719 (N_49719,N_44023,N_41906);
xor U49720 (N_49720,N_44287,N_42322);
and U49721 (N_49721,N_44585,N_43908);
xor U49722 (N_49722,N_44670,N_42711);
nor U49723 (N_49723,N_42953,N_44525);
nand U49724 (N_49724,N_42928,N_41028);
and U49725 (N_49725,N_40624,N_40201);
nor U49726 (N_49726,N_42354,N_41271);
nand U49727 (N_49727,N_44760,N_43056);
nand U49728 (N_49728,N_41759,N_44364);
and U49729 (N_49729,N_43243,N_42025);
nand U49730 (N_49730,N_41712,N_40576);
and U49731 (N_49731,N_40260,N_40283);
nand U49732 (N_49732,N_40250,N_40850);
and U49733 (N_49733,N_41542,N_40372);
nor U49734 (N_49734,N_44386,N_44493);
nor U49735 (N_49735,N_44027,N_43615);
xor U49736 (N_49736,N_41200,N_43558);
xor U49737 (N_49737,N_42539,N_44144);
and U49738 (N_49738,N_41171,N_42982);
nand U49739 (N_49739,N_43776,N_44512);
nor U49740 (N_49740,N_44275,N_44449);
and U49741 (N_49741,N_40377,N_40286);
nor U49742 (N_49742,N_41596,N_41208);
xnor U49743 (N_49743,N_41200,N_44539);
and U49744 (N_49744,N_41431,N_41540);
nor U49745 (N_49745,N_41796,N_44047);
or U49746 (N_49746,N_43120,N_43755);
nand U49747 (N_49747,N_44137,N_40970);
nand U49748 (N_49748,N_42152,N_40279);
nand U49749 (N_49749,N_42398,N_43008);
or U49750 (N_49750,N_42950,N_40832);
and U49751 (N_49751,N_42406,N_43298);
or U49752 (N_49752,N_40097,N_42326);
nand U49753 (N_49753,N_43345,N_44210);
xor U49754 (N_49754,N_42916,N_40018);
and U49755 (N_49755,N_41867,N_42523);
nor U49756 (N_49756,N_40336,N_41062);
nand U49757 (N_49757,N_42519,N_44770);
and U49758 (N_49758,N_42060,N_43179);
nor U49759 (N_49759,N_42235,N_41373);
or U49760 (N_49760,N_41384,N_42736);
and U49761 (N_49761,N_44549,N_43853);
nand U49762 (N_49762,N_41157,N_41639);
and U49763 (N_49763,N_40944,N_44894);
and U49764 (N_49764,N_44819,N_42671);
or U49765 (N_49765,N_42913,N_42746);
and U49766 (N_49766,N_42109,N_42176);
nand U49767 (N_49767,N_43084,N_43236);
or U49768 (N_49768,N_42272,N_43398);
nor U49769 (N_49769,N_43128,N_42310);
xnor U49770 (N_49770,N_44109,N_44087);
nor U49771 (N_49771,N_44994,N_43684);
or U49772 (N_49772,N_43130,N_44177);
and U49773 (N_49773,N_43849,N_43225);
nor U49774 (N_49774,N_40886,N_41579);
xnor U49775 (N_49775,N_42416,N_44195);
nor U49776 (N_49776,N_44268,N_41028);
nand U49777 (N_49777,N_43568,N_44139);
nand U49778 (N_49778,N_41811,N_40061);
xnor U49779 (N_49779,N_42951,N_44008);
xor U49780 (N_49780,N_43097,N_40860);
xor U49781 (N_49781,N_44356,N_40857);
nor U49782 (N_49782,N_41065,N_41020);
xnor U49783 (N_49783,N_44218,N_42547);
and U49784 (N_49784,N_44009,N_40412);
nand U49785 (N_49785,N_41834,N_44511);
nor U49786 (N_49786,N_43116,N_43670);
and U49787 (N_49787,N_44491,N_40245);
nand U49788 (N_49788,N_42498,N_44040);
nand U49789 (N_49789,N_40832,N_43235);
and U49790 (N_49790,N_41355,N_42501);
xnor U49791 (N_49791,N_43045,N_40397);
and U49792 (N_49792,N_40498,N_40557);
and U49793 (N_49793,N_42998,N_43314);
nor U49794 (N_49794,N_41628,N_40119);
xnor U49795 (N_49795,N_44941,N_41515);
nor U49796 (N_49796,N_43766,N_40663);
or U49797 (N_49797,N_40673,N_44468);
nor U49798 (N_49798,N_40837,N_40059);
or U49799 (N_49799,N_41200,N_42384);
and U49800 (N_49800,N_43959,N_42315);
xnor U49801 (N_49801,N_42400,N_44809);
xnor U49802 (N_49802,N_42902,N_42643);
or U49803 (N_49803,N_42214,N_42264);
and U49804 (N_49804,N_44090,N_43866);
nand U49805 (N_49805,N_40499,N_44436);
xnor U49806 (N_49806,N_42968,N_41315);
nor U49807 (N_49807,N_42691,N_41799);
nand U49808 (N_49808,N_43153,N_40232);
or U49809 (N_49809,N_43636,N_42812);
and U49810 (N_49810,N_43297,N_41415);
nor U49811 (N_49811,N_42909,N_42753);
or U49812 (N_49812,N_42648,N_41214);
and U49813 (N_49813,N_42040,N_44483);
xnor U49814 (N_49814,N_41776,N_43346);
and U49815 (N_49815,N_43646,N_42549);
xor U49816 (N_49816,N_40603,N_44888);
or U49817 (N_49817,N_44530,N_44268);
xnor U49818 (N_49818,N_44501,N_43953);
xor U49819 (N_49819,N_43945,N_42111);
and U49820 (N_49820,N_44208,N_40494);
nand U49821 (N_49821,N_43956,N_41493);
nor U49822 (N_49822,N_42999,N_44829);
nor U49823 (N_49823,N_40096,N_40213);
and U49824 (N_49824,N_44958,N_43799);
xor U49825 (N_49825,N_43738,N_40886);
nor U49826 (N_49826,N_44406,N_42269);
or U49827 (N_49827,N_43782,N_42366);
and U49828 (N_49828,N_41696,N_41152);
nand U49829 (N_49829,N_44964,N_44723);
and U49830 (N_49830,N_43977,N_44382);
or U49831 (N_49831,N_40304,N_42929);
nor U49832 (N_49832,N_41741,N_40645);
nor U49833 (N_49833,N_41828,N_40632);
or U49834 (N_49834,N_41046,N_43453);
nand U49835 (N_49835,N_44784,N_44608);
and U49836 (N_49836,N_43214,N_41440);
or U49837 (N_49837,N_40165,N_40222);
nor U49838 (N_49838,N_43906,N_44863);
nand U49839 (N_49839,N_43009,N_42025);
and U49840 (N_49840,N_40621,N_40272);
xor U49841 (N_49841,N_43364,N_42807);
and U49842 (N_49842,N_42978,N_44955);
nor U49843 (N_49843,N_44692,N_44950);
and U49844 (N_49844,N_43643,N_41448);
xnor U49845 (N_49845,N_42444,N_42451);
or U49846 (N_49846,N_41954,N_41595);
and U49847 (N_49847,N_43003,N_44315);
xnor U49848 (N_49848,N_43944,N_41494);
and U49849 (N_49849,N_40717,N_40751);
or U49850 (N_49850,N_41533,N_43322);
nor U49851 (N_49851,N_43015,N_40592);
or U49852 (N_49852,N_41237,N_42751);
or U49853 (N_49853,N_43724,N_44845);
and U49854 (N_49854,N_44713,N_41152);
nor U49855 (N_49855,N_44445,N_43363);
and U49856 (N_49856,N_40700,N_42984);
nand U49857 (N_49857,N_42139,N_43674);
and U49858 (N_49858,N_44820,N_40815);
or U49859 (N_49859,N_40112,N_44628);
or U49860 (N_49860,N_43548,N_40241);
nand U49861 (N_49861,N_42695,N_42375);
or U49862 (N_49862,N_44847,N_41542);
and U49863 (N_49863,N_42977,N_40232);
and U49864 (N_49864,N_41585,N_40343);
nor U49865 (N_49865,N_41134,N_44996);
nor U49866 (N_49866,N_43496,N_40397);
nand U49867 (N_49867,N_40840,N_43241);
xor U49868 (N_49868,N_41583,N_40487);
and U49869 (N_49869,N_44192,N_40251);
xnor U49870 (N_49870,N_42849,N_41463);
xor U49871 (N_49871,N_42098,N_40565);
or U49872 (N_49872,N_43779,N_42387);
nand U49873 (N_49873,N_44487,N_40453);
nand U49874 (N_49874,N_43643,N_43657);
nor U49875 (N_49875,N_40134,N_44150);
nor U49876 (N_49876,N_41382,N_40023);
nor U49877 (N_49877,N_44820,N_43730);
and U49878 (N_49878,N_41873,N_44509);
nor U49879 (N_49879,N_43021,N_43815);
or U49880 (N_49880,N_41539,N_41563);
nand U49881 (N_49881,N_44648,N_42561);
or U49882 (N_49882,N_44735,N_44169);
nand U49883 (N_49883,N_40540,N_42689);
nand U49884 (N_49884,N_40758,N_40485);
xor U49885 (N_49885,N_42377,N_41807);
nand U49886 (N_49886,N_42443,N_41229);
nor U49887 (N_49887,N_43338,N_42730);
and U49888 (N_49888,N_42934,N_43954);
nor U49889 (N_49889,N_43022,N_44193);
or U49890 (N_49890,N_43075,N_42176);
xnor U49891 (N_49891,N_43670,N_42464);
or U49892 (N_49892,N_40640,N_44625);
nand U49893 (N_49893,N_41707,N_42751);
nand U49894 (N_49894,N_43406,N_42156);
nor U49895 (N_49895,N_43106,N_41557);
xnor U49896 (N_49896,N_41794,N_44584);
nor U49897 (N_49897,N_42434,N_40755);
nand U49898 (N_49898,N_42333,N_43472);
nor U49899 (N_49899,N_43159,N_44902);
xnor U49900 (N_49900,N_43510,N_40397);
nor U49901 (N_49901,N_42201,N_42040);
or U49902 (N_49902,N_42144,N_44494);
nand U49903 (N_49903,N_40194,N_42581);
and U49904 (N_49904,N_42121,N_42415);
and U49905 (N_49905,N_42126,N_42551);
and U49906 (N_49906,N_43331,N_42951);
nand U49907 (N_49907,N_44032,N_43773);
nor U49908 (N_49908,N_41187,N_41518);
nor U49909 (N_49909,N_42466,N_42906);
or U49910 (N_49910,N_42320,N_42247);
or U49911 (N_49911,N_44577,N_40967);
xor U49912 (N_49912,N_43962,N_41136);
and U49913 (N_49913,N_43218,N_40853);
xor U49914 (N_49914,N_41821,N_43621);
nor U49915 (N_49915,N_40576,N_44125);
and U49916 (N_49916,N_40297,N_40375);
nand U49917 (N_49917,N_43373,N_41654);
or U49918 (N_49918,N_44239,N_42954);
xnor U49919 (N_49919,N_42067,N_42750);
and U49920 (N_49920,N_44817,N_41279);
and U49921 (N_49921,N_40984,N_40502);
or U49922 (N_49922,N_40836,N_40753);
or U49923 (N_49923,N_42950,N_44563);
nand U49924 (N_49924,N_44465,N_42892);
xnor U49925 (N_49925,N_42755,N_43156);
and U49926 (N_49926,N_42597,N_44441);
xnor U49927 (N_49927,N_40657,N_40168);
and U49928 (N_49928,N_40919,N_40479);
xor U49929 (N_49929,N_42544,N_42539);
xor U49930 (N_49930,N_42185,N_41143);
nand U49931 (N_49931,N_42914,N_42281);
nand U49932 (N_49932,N_41331,N_42316);
nand U49933 (N_49933,N_43004,N_43482);
nor U49934 (N_49934,N_42179,N_44164);
and U49935 (N_49935,N_44124,N_44458);
nand U49936 (N_49936,N_44063,N_44447);
or U49937 (N_49937,N_40962,N_41876);
or U49938 (N_49938,N_43893,N_44410);
nor U49939 (N_49939,N_41434,N_43900);
nand U49940 (N_49940,N_40436,N_44855);
xnor U49941 (N_49941,N_43525,N_40217);
and U49942 (N_49942,N_40392,N_43170);
xnor U49943 (N_49943,N_41750,N_41464);
xnor U49944 (N_49944,N_41884,N_42635);
and U49945 (N_49945,N_42063,N_41496);
nand U49946 (N_49946,N_44624,N_43136);
nand U49947 (N_49947,N_41366,N_42647);
and U49948 (N_49948,N_43862,N_40676);
nand U49949 (N_49949,N_44808,N_41644);
or U49950 (N_49950,N_43739,N_41251);
nand U49951 (N_49951,N_41553,N_41652);
and U49952 (N_49952,N_42098,N_41218);
xor U49953 (N_49953,N_41119,N_44864);
nor U49954 (N_49954,N_42209,N_44836);
nor U49955 (N_49955,N_44293,N_42872);
xor U49956 (N_49956,N_44701,N_42147);
or U49957 (N_49957,N_43320,N_44773);
and U49958 (N_49958,N_40560,N_44020);
and U49959 (N_49959,N_40662,N_41033);
nand U49960 (N_49960,N_42667,N_40576);
xor U49961 (N_49961,N_41447,N_43359);
xor U49962 (N_49962,N_42119,N_42040);
nand U49963 (N_49963,N_43312,N_43768);
and U49964 (N_49964,N_41366,N_41019);
nor U49965 (N_49965,N_41450,N_40814);
and U49966 (N_49966,N_44784,N_44057);
xor U49967 (N_49967,N_41305,N_43757);
xnor U49968 (N_49968,N_40729,N_44784);
nand U49969 (N_49969,N_44089,N_43221);
or U49970 (N_49970,N_42511,N_41366);
nor U49971 (N_49971,N_40415,N_43386);
and U49972 (N_49972,N_42733,N_43211);
and U49973 (N_49973,N_43700,N_41870);
nand U49974 (N_49974,N_40264,N_40266);
nand U49975 (N_49975,N_44281,N_41309);
and U49976 (N_49976,N_40762,N_40652);
and U49977 (N_49977,N_44889,N_43957);
or U49978 (N_49978,N_40041,N_41391);
xor U49979 (N_49979,N_44584,N_43771);
nand U49980 (N_49980,N_42111,N_44027);
nand U49981 (N_49981,N_42518,N_42105);
or U49982 (N_49982,N_40459,N_42296);
nor U49983 (N_49983,N_43084,N_43056);
or U49984 (N_49984,N_42566,N_42122);
nor U49985 (N_49985,N_43702,N_40248);
and U49986 (N_49986,N_43584,N_42163);
nor U49987 (N_49987,N_44992,N_44743);
nand U49988 (N_49988,N_44035,N_40655);
nor U49989 (N_49989,N_41065,N_40897);
nand U49990 (N_49990,N_40363,N_41372);
nand U49991 (N_49991,N_44047,N_44615);
nand U49992 (N_49992,N_40594,N_40841);
nor U49993 (N_49993,N_40675,N_43772);
or U49994 (N_49994,N_41336,N_41058);
nor U49995 (N_49995,N_42640,N_44656);
nand U49996 (N_49996,N_44335,N_42660);
nand U49997 (N_49997,N_44857,N_41188);
nor U49998 (N_49998,N_41962,N_44022);
or U49999 (N_49999,N_41288,N_40246);
xnor UO_0 (O_0,N_49572,N_46339);
and UO_1 (O_1,N_49795,N_46842);
or UO_2 (O_2,N_49944,N_45229);
and UO_3 (O_3,N_48664,N_45035);
nor UO_4 (O_4,N_49831,N_47552);
and UO_5 (O_5,N_49450,N_46840);
nand UO_6 (O_6,N_48514,N_46082);
or UO_7 (O_7,N_48677,N_45353);
or UO_8 (O_8,N_47622,N_49123);
nand UO_9 (O_9,N_48265,N_46252);
nor UO_10 (O_10,N_48117,N_45961);
xnor UO_11 (O_11,N_45940,N_46578);
nand UO_12 (O_12,N_49136,N_49401);
nor UO_13 (O_13,N_49183,N_47952);
or UO_14 (O_14,N_45547,N_48856);
and UO_15 (O_15,N_47838,N_49232);
nor UO_16 (O_16,N_45232,N_47741);
or UO_17 (O_17,N_47508,N_47750);
and UO_18 (O_18,N_49162,N_47253);
and UO_19 (O_19,N_49967,N_49928);
nand UO_20 (O_20,N_45589,N_49905);
and UO_21 (O_21,N_46924,N_47491);
nor UO_22 (O_22,N_46378,N_48651);
and UO_23 (O_23,N_47836,N_47537);
or UO_24 (O_24,N_48272,N_49823);
and UO_25 (O_25,N_46529,N_48018);
nor UO_26 (O_26,N_49835,N_47662);
xor UO_27 (O_27,N_49644,N_48137);
nor UO_28 (O_28,N_47281,N_46572);
nand UO_29 (O_29,N_48735,N_47794);
nand UO_30 (O_30,N_47874,N_46060);
xnor UO_31 (O_31,N_46332,N_45455);
and UO_32 (O_32,N_49268,N_47489);
xor UO_33 (O_33,N_46386,N_48756);
and UO_34 (O_34,N_46870,N_46308);
or UO_35 (O_35,N_48177,N_49314);
xor UO_36 (O_36,N_49921,N_45731);
xnor UO_37 (O_37,N_45134,N_45064);
nor UO_38 (O_38,N_46912,N_49796);
and UO_39 (O_39,N_47638,N_45632);
nand UO_40 (O_40,N_45457,N_46949);
nand UO_41 (O_41,N_45877,N_47008);
xnor UO_42 (O_42,N_45833,N_47873);
or UO_43 (O_43,N_46732,N_46625);
xor UO_44 (O_44,N_47585,N_47151);
or UO_45 (O_45,N_49470,N_45079);
nor UO_46 (O_46,N_49022,N_45803);
or UO_47 (O_47,N_49850,N_45549);
nand UO_48 (O_48,N_49651,N_49742);
xor UO_49 (O_49,N_45490,N_45849);
and UO_50 (O_50,N_49545,N_45146);
nor UO_51 (O_51,N_46017,N_49141);
or UO_52 (O_52,N_49008,N_45850);
nor UO_53 (O_53,N_49784,N_45659);
nand UO_54 (O_54,N_45984,N_47311);
or UO_55 (O_55,N_49191,N_48928);
or UO_56 (O_56,N_47887,N_48899);
nand UO_57 (O_57,N_45373,N_45913);
and UO_58 (O_58,N_47995,N_47130);
and UO_59 (O_59,N_48919,N_47528);
xor UO_60 (O_60,N_49167,N_45751);
or UO_61 (O_61,N_46177,N_47204);
nand UO_62 (O_62,N_49629,N_49280);
and UO_63 (O_63,N_46963,N_47513);
nor UO_64 (O_64,N_45969,N_46504);
nand UO_65 (O_65,N_45464,N_45186);
xnor UO_66 (O_66,N_45652,N_48698);
or UO_67 (O_67,N_45591,N_47796);
nand UO_68 (O_68,N_46793,N_47372);
nand UO_69 (O_69,N_46834,N_45109);
xor UO_70 (O_70,N_49716,N_48446);
and UO_71 (O_71,N_48325,N_45418);
xor UO_72 (O_72,N_49297,N_47682);
and UO_73 (O_73,N_49101,N_46629);
xor UO_74 (O_74,N_45805,N_47527);
nand UO_75 (O_75,N_48162,N_49005);
and UO_76 (O_76,N_48381,N_47553);
nor UO_77 (O_77,N_45218,N_48705);
nor UO_78 (O_78,N_49212,N_47230);
or UO_79 (O_79,N_46894,N_48387);
nand UO_80 (O_80,N_46087,N_49529);
xnor UO_81 (O_81,N_47855,N_47381);
xnor UO_82 (O_82,N_46026,N_47573);
nor UO_83 (O_83,N_45511,N_49275);
nor UO_84 (O_84,N_47065,N_48057);
nand UO_85 (O_85,N_45949,N_48666);
xor UO_86 (O_86,N_46491,N_49128);
and UO_87 (O_87,N_47283,N_47548);
or UO_88 (O_88,N_48992,N_46762);
xnor UO_89 (O_89,N_46123,N_48227);
or UO_90 (O_90,N_47704,N_45931);
and UO_91 (O_91,N_48744,N_46190);
xor UO_92 (O_92,N_45107,N_45008);
or UO_93 (O_93,N_47824,N_45136);
nand UO_94 (O_94,N_48947,N_46575);
nand UO_95 (O_95,N_48816,N_45978);
and UO_96 (O_96,N_47900,N_49900);
or UO_97 (O_97,N_47007,N_46598);
nor UO_98 (O_98,N_48260,N_45370);
xnor UO_99 (O_99,N_45611,N_45785);
and UO_100 (O_100,N_48089,N_49233);
and UO_101 (O_101,N_46228,N_48077);
nor UO_102 (O_102,N_48598,N_45838);
xor UO_103 (O_103,N_47772,N_46658);
nand UO_104 (O_104,N_47726,N_45286);
or UO_105 (O_105,N_47771,N_45205);
or UO_106 (O_106,N_46558,N_46846);
or UO_107 (O_107,N_49947,N_45879);
and UO_108 (O_108,N_48893,N_49257);
or UO_109 (O_109,N_46914,N_48726);
and UO_110 (O_110,N_46365,N_47308);
xor UO_111 (O_111,N_45648,N_47068);
xor UO_112 (O_112,N_45513,N_49664);
nor UO_113 (O_113,N_47785,N_48670);
xor UO_114 (O_114,N_45571,N_45974);
and UO_115 (O_115,N_46954,N_48024);
and UO_116 (O_116,N_46305,N_47298);
and UO_117 (O_117,N_46774,N_45859);
nand UO_118 (O_118,N_46107,N_45635);
xor UO_119 (O_119,N_47962,N_45120);
or UO_120 (O_120,N_45830,N_49279);
nand UO_121 (O_121,N_45679,N_49412);
and UO_122 (O_122,N_49107,N_49695);
xor UO_123 (O_123,N_45482,N_45819);
and UO_124 (O_124,N_46248,N_45098);
or UO_125 (O_125,N_48640,N_47781);
and UO_126 (O_126,N_49993,N_48034);
xor UO_127 (O_127,N_47577,N_46229);
and UO_128 (O_128,N_46582,N_48920);
nor UO_129 (O_129,N_47484,N_45090);
or UO_130 (O_130,N_48659,N_48786);
or UO_131 (O_131,N_49806,N_46302);
or UO_132 (O_132,N_45665,N_48292);
and UO_133 (O_133,N_48013,N_47498);
nor UO_134 (O_134,N_48541,N_47437);
nand UO_135 (O_135,N_46257,N_49499);
nand UO_136 (O_136,N_45856,N_46376);
and UO_137 (O_137,N_46896,N_45620);
or UO_138 (O_138,N_46351,N_47276);
nor UO_139 (O_139,N_48793,N_49498);
nor UO_140 (O_140,N_49869,N_48217);
nand UO_141 (O_141,N_49326,N_48451);
or UO_142 (O_142,N_47054,N_45282);
or UO_143 (O_143,N_48654,N_47334);
or UO_144 (O_144,N_47877,N_47757);
nor UO_145 (O_145,N_45980,N_45788);
or UO_146 (O_146,N_47574,N_45223);
nand UO_147 (O_147,N_47713,N_45020);
or UO_148 (O_148,N_46668,N_49030);
or UO_149 (O_149,N_45553,N_49096);
nor UO_150 (O_150,N_49339,N_46715);
nand UO_151 (O_151,N_45963,N_47401);
nor UO_152 (O_152,N_46819,N_49408);
nor UO_153 (O_153,N_48620,N_48282);
or UO_154 (O_154,N_46489,N_48969);
or UO_155 (O_155,N_46643,N_46208);
nor UO_156 (O_156,N_45349,N_49604);
and UO_157 (O_157,N_46324,N_47270);
and UO_158 (O_158,N_49840,N_45734);
or UO_159 (O_159,N_47284,N_47324);
nand UO_160 (O_160,N_49345,N_45432);
nand UO_161 (O_161,N_48403,N_45394);
nor UO_162 (O_162,N_46084,N_47249);
or UO_163 (O_163,N_48220,N_48909);
and UO_164 (O_164,N_47199,N_49732);
xor UO_165 (O_165,N_46016,N_49100);
nor UO_166 (O_166,N_47086,N_46903);
or UO_167 (O_167,N_49559,N_46534);
xnor UO_168 (O_168,N_49991,N_49042);
xor UO_169 (O_169,N_46772,N_47612);
or UO_170 (O_170,N_47997,N_47338);
or UO_171 (O_171,N_46950,N_49636);
or UO_172 (O_172,N_46266,N_48110);
nand UO_173 (O_173,N_48968,N_48875);
and UO_174 (O_174,N_45621,N_48005);
and UO_175 (O_175,N_47031,N_49773);
and UO_176 (O_176,N_48836,N_48722);
nand UO_177 (O_177,N_48810,N_49495);
xor UO_178 (O_178,N_48393,N_46277);
nor UO_179 (O_179,N_48248,N_45973);
nor UO_180 (O_180,N_46057,N_45874);
nor UO_181 (O_181,N_45427,N_46313);
xnor UO_182 (O_182,N_45826,N_47184);
xnor UO_183 (O_183,N_47393,N_45161);
nor UO_184 (O_184,N_45654,N_49067);
and UO_185 (O_185,N_46085,N_45255);
and UO_186 (O_186,N_46995,N_49676);
and UO_187 (O_187,N_45616,N_46663);
or UO_188 (O_188,N_46756,N_47686);
and UO_189 (O_189,N_49709,N_47705);
or UO_190 (O_190,N_45791,N_46158);
nor UO_191 (O_191,N_47210,N_45463);
nor UO_192 (O_192,N_45633,N_47170);
nor UO_193 (O_193,N_46580,N_47187);
xnor UO_194 (O_194,N_45461,N_45899);
nand UO_195 (O_195,N_45031,N_45933);
or UO_196 (O_196,N_48916,N_45853);
nand UO_197 (O_197,N_48399,N_47155);
nor UO_198 (O_198,N_47636,N_45124);
xor UO_199 (O_199,N_45770,N_48210);
and UO_200 (O_200,N_46259,N_48789);
xnor UO_201 (O_201,N_48055,N_48849);
xor UO_202 (O_202,N_48501,N_49674);
nand UO_203 (O_203,N_48475,N_49848);
or UO_204 (O_204,N_45097,N_47992);
xnor UO_205 (O_205,N_46556,N_46074);
nand UO_206 (O_206,N_47278,N_48589);
and UO_207 (O_207,N_46839,N_49447);
or UO_208 (O_208,N_49429,N_49739);
xor UO_209 (O_209,N_49622,N_49414);
and UO_210 (O_210,N_45559,N_46695);
nand UO_211 (O_211,N_47522,N_46510);
nor UO_212 (O_212,N_49700,N_49769);
and UO_213 (O_213,N_48287,N_46258);
nand UO_214 (O_214,N_47434,N_46826);
nand UO_215 (O_215,N_49290,N_45638);
or UO_216 (O_216,N_48745,N_47132);
nand UO_217 (O_217,N_46059,N_47212);
nor UO_218 (O_218,N_45092,N_46350);
xor UO_219 (O_219,N_48846,N_46019);
and UO_220 (O_220,N_45171,N_48635);
nand UO_221 (O_221,N_45944,N_49810);
nand UO_222 (O_222,N_45947,N_48578);
nor UO_223 (O_223,N_46642,N_45225);
nand UO_224 (O_224,N_48888,N_48095);
and UO_225 (O_225,N_49288,N_47179);
nor UO_226 (O_226,N_49938,N_45011);
or UO_227 (O_227,N_45604,N_48045);
or UO_228 (O_228,N_49815,N_47304);
nor UO_229 (O_229,N_47268,N_46620);
nand UO_230 (O_230,N_48761,N_46486);
or UO_231 (O_231,N_47349,N_47493);
xor UO_232 (O_232,N_46564,N_48533);
nor UO_233 (O_233,N_45637,N_49770);
or UO_234 (O_234,N_46614,N_45564);
nand UO_235 (O_235,N_45668,N_45884);
xor UO_236 (O_236,N_46735,N_48588);
xnor UO_237 (O_237,N_48225,N_46434);
nand UO_238 (O_238,N_47206,N_46079);
nor UO_239 (O_239,N_46563,N_47412);
or UO_240 (O_240,N_48648,N_47378);
or UO_241 (O_241,N_48092,N_45000);
nand UO_242 (O_242,N_46552,N_47057);
nor UO_243 (O_243,N_46783,N_47764);
xnor UO_244 (O_244,N_45548,N_47517);
nand UO_245 (O_245,N_47219,N_49047);
and UO_246 (O_246,N_47748,N_47398);
nand UO_247 (O_247,N_49449,N_49758);
or UO_248 (O_248,N_47663,N_45608);
and UO_249 (O_249,N_46526,N_48555);
and UO_250 (O_250,N_47858,N_45708);
and UO_251 (O_251,N_48763,N_45300);
nand UO_252 (O_252,N_46942,N_49502);
xor UO_253 (O_253,N_47465,N_49983);
nor UO_254 (O_254,N_46962,N_48870);
and UO_255 (O_255,N_47989,N_46922);
or UO_256 (O_256,N_45673,N_45509);
or UO_257 (O_257,N_48794,N_48736);
or UO_258 (O_258,N_49509,N_47941);
nand UO_259 (O_259,N_46430,N_49415);
nand UO_260 (O_260,N_46586,N_46784);
nor UO_261 (O_261,N_49469,N_49175);
or UO_262 (O_262,N_48646,N_47703);
and UO_263 (O_263,N_47728,N_45821);
xor UO_264 (O_264,N_49369,N_47791);
xor UO_265 (O_265,N_45917,N_45368);
or UO_266 (O_266,N_47605,N_47911);
nor UO_267 (O_267,N_47455,N_46519);
nand UO_268 (O_268,N_48583,N_48731);
nor UO_269 (O_269,N_49431,N_48021);
xor UO_270 (O_270,N_45858,N_49109);
and UO_271 (O_271,N_45515,N_49289);
and UO_272 (O_272,N_49619,N_48837);
or UO_273 (O_273,N_45752,N_46303);
and UO_274 (O_274,N_47407,N_47943);
or UO_275 (O_275,N_45934,N_45082);
xor UO_276 (O_276,N_47492,N_47603);
nor UO_277 (O_277,N_47937,N_45982);
nor UO_278 (O_278,N_45878,N_48884);
nor UO_279 (O_279,N_48285,N_48702);
or UO_280 (O_280,N_47377,N_49276);
nand UO_281 (O_281,N_45975,N_49321);
xnor UO_282 (O_282,N_48079,N_46346);
xnor UO_283 (O_283,N_47441,N_47743);
nor UO_284 (O_284,N_48516,N_45240);
nor UO_285 (O_285,N_47606,N_47649);
xnor UO_286 (O_286,N_45898,N_49176);
or UO_287 (O_287,N_45471,N_48324);
nor UO_288 (O_288,N_47096,N_49218);
xnor UO_289 (O_289,N_45063,N_45308);
xor UO_290 (O_290,N_48511,N_48804);
xor UO_291 (O_291,N_45842,N_49072);
nor UO_292 (O_292,N_49421,N_45721);
xnor UO_293 (O_293,N_46559,N_47673);
xnor UO_294 (O_294,N_49007,N_46130);
nor UO_295 (O_295,N_47217,N_48070);
xnor UO_296 (O_296,N_45643,N_46408);
xor UO_297 (O_297,N_47134,N_46724);
and UO_298 (O_298,N_48781,N_47314);
and UO_299 (O_299,N_49645,N_49519);
nand UO_300 (O_300,N_49968,N_49922);
xor UO_301 (O_301,N_45603,N_47352);
xor UO_302 (O_302,N_49076,N_46712);
xnor UO_303 (O_303,N_48610,N_47263);
nand UO_304 (O_304,N_46103,N_48823);
nor UO_305 (O_305,N_48703,N_48112);
xnor UO_306 (O_306,N_49975,N_45410);
xnor UO_307 (O_307,N_48412,N_46230);
nor UO_308 (O_308,N_45759,N_46247);
xnor UO_309 (O_309,N_46731,N_48988);
and UO_310 (O_310,N_48085,N_48560);
nand UO_311 (O_311,N_48867,N_48831);
xor UO_312 (O_312,N_47301,N_46980);
nor UO_313 (O_313,N_48518,N_48910);
and UO_314 (O_314,N_48022,N_49256);
nand UO_315 (O_315,N_48007,N_45622);
and UO_316 (O_316,N_45657,N_46566);
or UO_317 (O_317,N_49272,N_47156);
and UO_318 (O_318,N_46565,N_48760);
and UO_319 (O_319,N_46484,N_48774);
or UO_320 (O_320,N_49740,N_49735);
xnor UO_321 (O_321,N_45269,N_47018);
xnor UO_322 (O_322,N_46897,N_49605);
nor UO_323 (O_323,N_47812,N_46382);
and UO_324 (O_324,N_48345,N_49597);
and UO_325 (O_325,N_48949,N_46210);
xnor UO_326 (O_326,N_49426,N_48604);
or UO_327 (O_327,N_49507,N_48615);
nor UO_328 (O_328,N_47222,N_46627);
xor UO_329 (O_329,N_45967,N_47614);
xnor UO_330 (O_330,N_48936,N_49747);
xor UO_331 (O_331,N_49265,N_46075);
xor UO_332 (O_332,N_47256,N_45028);
or UO_333 (O_333,N_45854,N_46527);
xnor UO_334 (O_334,N_49749,N_46776);
and UO_335 (O_335,N_48003,N_47464);
and UO_336 (O_336,N_49755,N_49374);
xor UO_337 (O_337,N_45755,N_47424);
or UO_338 (O_338,N_46108,N_49878);
nand UO_339 (O_339,N_47925,N_45609);
nand UO_340 (O_340,N_47415,N_46058);
or UO_341 (O_341,N_45615,N_47266);
and UO_342 (O_342,N_47981,N_46866);
xor UO_343 (O_343,N_45623,N_45243);
or UO_344 (O_344,N_49195,N_48987);
or UO_345 (O_345,N_45324,N_46213);
xnor UO_346 (O_346,N_47336,N_48618);
or UO_347 (O_347,N_45377,N_45529);
and UO_348 (O_348,N_48842,N_47584);
nand UO_349 (O_349,N_46162,N_48682);
nand UO_350 (O_350,N_45474,N_46116);
or UO_351 (O_351,N_48950,N_48540);
nor UO_352 (O_352,N_47113,N_46166);
and UO_353 (O_353,N_49767,N_45906);
and UO_354 (O_354,N_47879,N_48914);
xnor UO_355 (O_355,N_45188,N_48241);
or UO_356 (O_356,N_49788,N_47734);
nand UO_357 (O_357,N_49106,N_46759);
and UO_358 (O_358,N_45383,N_47312);
and UO_359 (O_359,N_45437,N_49880);
or UO_360 (O_360,N_46699,N_49309);
and UO_361 (O_361,N_48565,N_45211);
or UO_362 (O_362,N_46992,N_49253);
nand UO_363 (O_363,N_48985,N_46164);
xnor UO_364 (O_364,N_47845,N_45217);
xor UO_365 (O_365,N_46876,N_47665);
nor UO_366 (O_366,N_49771,N_48155);
and UO_367 (O_367,N_49908,N_48141);
nand UO_368 (O_368,N_45159,N_47055);
xor UO_369 (O_369,N_48840,N_48890);
nand UO_370 (O_370,N_47938,N_48554);
nand UO_371 (O_371,N_49164,N_47837);
xnor UO_372 (O_372,N_45142,N_45627);
xnor UO_373 (O_373,N_49649,N_46173);
or UO_374 (O_374,N_45288,N_47092);
nand UO_375 (O_375,N_45185,N_45670);
xnor UO_376 (O_376,N_48386,N_47379);
or UO_377 (O_377,N_45742,N_49384);
or UO_378 (O_378,N_45417,N_49871);
xor UO_379 (O_379,N_46803,N_47882);
nand UO_380 (O_380,N_49440,N_47466);
or UO_381 (O_381,N_49221,N_49066);
nor UO_382 (O_382,N_49686,N_46825);
nand UO_383 (O_383,N_47642,N_48882);
xnor UO_384 (O_384,N_48198,N_48359);
nor UO_385 (O_385,N_47000,N_49002);
xor UO_386 (O_386,N_47708,N_47546);
and UO_387 (O_387,N_46716,N_46102);
nor UO_388 (O_388,N_48941,N_48746);
nor UO_389 (O_389,N_46220,N_49443);
and UO_390 (O_390,N_48373,N_49508);
nand UO_391 (O_391,N_47017,N_47979);
or UO_392 (O_392,N_48379,N_45572);
or UO_393 (O_393,N_48036,N_45104);
and UO_394 (O_394,N_49786,N_48959);
or UO_395 (O_395,N_48796,N_48256);
or UO_396 (O_396,N_45409,N_48060);
or UO_397 (O_397,N_45034,N_45954);
nor UO_398 (O_398,N_46573,N_48841);
or UO_399 (O_399,N_46684,N_45449);
or UO_400 (O_400,N_48181,N_46231);
nor UO_401 (O_401,N_48401,N_47329);
xor UO_402 (O_402,N_49293,N_48035);
xor UO_403 (O_403,N_48172,N_49228);
xnor UO_404 (O_404,N_46574,N_47045);
xor UO_405 (O_405,N_47817,N_48099);
and UO_406 (O_406,N_48558,N_46795);
and UO_407 (O_407,N_47689,N_47860);
xnor UO_408 (O_408,N_48952,N_48607);
or UO_409 (O_409,N_47602,N_46387);
nand UO_410 (O_410,N_45002,N_45153);
nand UO_411 (O_411,N_48215,N_49521);
nor UO_412 (O_412,N_47236,N_48608);
nor UO_413 (O_413,N_46416,N_49360);
nand UO_414 (O_414,N_47869,N_46284);
nor UO_415 (O_415,N_49235,N_49791);
or UO_416 (O_416,N_49040,N_48298);
nor UO_417 (O_417,N_47878,N_49160);
or UO_418 (O_418,N_47174,N_49018);
and UO_419 (O_419,N_49154,N_45653);
nand UO_420 (O_420,N_45279,N_47296);
or UO_421 (O_421,N_48297,N_47145);
xor UO_422 (O_422,N_48996,N_45492);
or UO_423 (O_423,N_49438,N_49949);
or UO_424 (O_424,N_45045,N_45908);
or UO_425 (O_425,N_46850,N_49575);
nor UO_426 (O_426,N_46348,N_48074);
xnor UO_427 (O_427,N_47262,N_49399);
xnor UO_428 (O_428,N_46971,N_46283);
and UO_429 (O_429,N_48688,N_47255);
nand UO_430 (O_430,N_45013,N_45506);
nand UO_431 (O_431,N_48738,N_46734);
nand UO_432 (O_432,N_46518,N_46422);
nand UO_433 (O_433,N_49019,N_46030);
xor UO_434 (O_434,N_48829,N_46607);
xnor UO_435 (O_435,N_46369,N_45520);
xnor UO_436 (O_436,N_46122,N_46862);
nor UO_437 (O_437,N_47910,N_45369);
or UO_438 (O_438,N_45009,N_45691);
nor UO_439 (O_439,N_47637,N_49574);
nor UO_440 (O_440,N_47477,N_45724);
and UO_441 (O_441,N_47084,N_49504);
nor UO_442 (O_442,N_45254,N_48832);
and UO_443 (O_443,N_45361,N_46708);
nor UO_444 (O_444,N_49668,N_48127);
nor UO_445 (O_445,N_47913,N_47813);
or UO_446 (O_446,N_45903,N_46701);
xor UO_447 (O_447,N_47406,N_47893);
or UO_448 (O_448,N_47062,N_47423);
and UO_449 (O_449,N_45600,N_48064);
nand UO_450 (O_450,N_48417,N_49316);
nand UO_451 (O_451,N_45663,N_45544);
nand UO_452 (O_452,N_49017,N_46462);
nand UO_453 (O_453,N_46847,N_46520);
xnor UO_454 (O_454,N_46101,N_47368);
and UO_455 (O_455,N_47929,N_48335);
xnor UO_456 (O_456,N_48844,N_45113);
nor UO_457 (O_457,N_49188,N_49540);
nand UO_458 (O_458,N_49303,N_48951);
and UO_459 (O_459,N_45429,N_46179);
nor UO_460 (O_460,N_49048,N_47659);
or UO_461 (O_461,N_45351,N_49992);
and UO_462 (O_462,N_49790,N_48649);
xor UO_463 (O_463,N_48869,N_49208);
or UO_464 (O_464,N_47361,N_47056);
and UO_465 (O_465,N_47322,N_49573);
or UO_466 (O_466,N_47557,N_45184);
xnor UO_467 (O_467,N_46150,N_47690);
and UO_468 (O_468,N_48924,N_46070);
and UO_469 (O_469,N_47157,N_49801);
nand UO_470 (O_470,N_46909,N_48130);
nand UO_471 (O_471,N_46316,N_47207);
and UO_472 (O_472,N_47500,N_45845);
xnor UO_473 (O_473,N_46021,N_49051);
nand UO_474 (O_474,N_48425,N_47438);
nor UO_475 (O_475,N_48176,N_48404);
nor UO_476 (O_476,N_47560,N_49904);
or UO_477 (O_477,N_47403,N_45386);
nand UO_478 (O_478,N_45263,N_48480);
nor UO_479 (O_479,N_48208,N_48000);
or UO_480 (O_480,N_45326,N_45613);
nand UO_481 (O_481,N_48319,N_45340);
or UO_482 (O_482,N_48984,N_46679);
and UO_483 (O_483,N_47272,N_49859);
and UO_484 (O_484,N_45890,N_47698);
xor UO_485 (O_485,N_47966,N_47725);
xnor UO_486 (O_486,N_46691,N_49643);
nor UO_487 (O_487,N_46488,N_48246);
nand UO_488 (O_488,N_47205,N_48101);
nand UO_489 (O_489,N_47535,N_48073);
and UO_490 (O_490,N_45952,N_46341);
and UO_491 (O_491,N_45556,N_46038);
and UO_492 (O_492,N_45403,N_49127);
nand UO_493 (O_493,N_49385,N_45767);
and UO_494 (O_494,N_45840,N_47216);
xnor UO_495 (O_495,N_46304,N_49915);
nand UO_496 (O_496,N_46856,N_49170);
nor UO_497 (O_497,N_46402,N_47829);
nor UO_498 (O_498,N_47416,N_45998);
nand UO_499 (O_499,N_48068,N_49957);
or UO_500 (O_500,N_47760,N_47835);
nand UO_501 (O_501,N_47936,N_49746);
or UO_502 (O_502,N_46094,N_47999);
or UO_503 (O_503,N_49407,N_46739);
xnor UO_504 (O_504,N_46569,N_46192);
nand UO_505 (O_505,N_47758,N_48204);
and UO_506 (O_506,N_45631,N_48033);
nor UO_507 (O_507,N_47857,N_46623);
nor UO_508 (O_508,N_47529,N_45182);
nand UO_509 (O_509,N_46923,N_49225);
nor UO_510 (O_510,N_45685,N_47971);
nor UO_511 (O_511,N_48859,N_49491);
or UO_512 (O_512,N_46718,N_48190);
and UO_513 (O_513,N_47515,N_45360);
or UO_514 (O_514,N_48792,N_49737);
nor UO_515 (O_515,N_48268,N_45156);
nand UO_516 (O_516,N_45111,N_48510);
or UO_517 (O_517,N_48502,N_47119);
xnor UO_518 (O_518,N_47462,N_47797);
or UO_519 (O_519,N_47861,N_46852);
nand UO_520 (O_520,N_46243,N_47425);
nand UO_521 (O_521,N_49341,N_48413);
and UO_522 (O_522,N_48779,N_47946);
or UO_523 (O_523,N_48430,N_47384);
and UO_524 (O_524,N_46721,N_45162);
and UO_525 (O_525,N_47683,N_48491);
and UO_526 (O_526,N_47976,N_48805);
or UO_527 (O_527,N_45454,N_46503);
or UO_528 (O_528,N_48903,N_47258);
nor UO_529 (O_529,N_46612,N_48328);
and UO_530 (O_530,N_45715,N_47731);
nor UO_531 (O_531,N_45181,N_46859);
and UO_532 (O_532,N_46297,N_47834);
xnor UO_533 (O_533,N_49568,N_46737);
or UO_534 (O_534,N_45711,N_45817);
nor UO_535 (O_535,N_46212,N_47892);
nor UO_536 (O_536,N_45929,N_46638);
or UO_537 (O_537,N_49889,N_46149);
or UO_538 (O_538,N_47196,N_47386);
xnor UO_539 (O_539,N_46851,N_49547);
and UO_540 (O_540,N_49219,N_45504);
xnor UO_541 (O_541,N_48531,N_45246);
nand UO_542 (O_542,N_46384,N_49623);
xor UO_543 (O_543,N_46292,N_47536);
and UO_544 (O_544,N_49198,N_45839);
xor UO_545 (O_545,N_47819,N_48029);
and UO_546 (O_546,N_45970,N_47654);
or UO_547 (O_547,N_46336,N_46831);
and UO_548 (O_548,N_47138,N_49163);
or UO_549 (O_549,N_48308,N_48693);
and UO_550 (O_550,N_45450,N_49893);
nor UO_551 (O_551,N_48866,N_47480);
and UO_552 (O_552,N_46298,N_48752);
xor UO_553 (O_553,N_46861,N_49972);
nand UO_554 (O_554,N_48183,N_45178);
nand UO_555 (O_555,N_48463,N_47956);
nor UO_556 (O_556,N_48093,N_48126);
and UO_557 (O_557,N_45552,N_47419);
nor UO_558 (O_558,N_46993,N_49792);
xor UO_559 (O_559,N_49750,N_47111);
or UO_560 (O_560,N_47444,N_48314);
nand UO_561 (O_561,N_45499,N_47467);
and UO_562 (O_562,N_45004,N_47078);
or UO_563 (O_563,N_47099,N_48264);
or UO_564 (O_564,N_45810,N_47635);
nand UO_565 (O_565,N_49406,N_48323);
xor UO_566 (O_566,N_45707,N_49380);
and UO_567 (O_567,N_46945,N_48833);
or UO_568 (O_568,N_47970,N_46282);
nor UO_569 (O_569,N_49624,N_48685);
nor UO_570 (O_570,N_49378,N_45389);
or UO_571 (O_571,N_47295,N_48537);
xor UO_572 (O_572,N_48907,N_45605);
and UO_573 (O_573,N_48020,N_46632);
xor UO_574 (O_574,N_48114,N_45362);
xor UO_575 (O_575,N_48242,N_46245);
and UO_576 (O_576,N_45909,N_45396);
nor UO_577 (O_577,N_47209,N_48590);
and UO_578 (O_578,N_47234,N_45466);
xnor UO_579 (O_579,N_45539,N_46940);
xor UO_580 (O_580,N_45010,N_48768);
xnor UO_581 (O_581,N_45398,N_47594);
nand UO_582 (O_582,N_45816,N_47744);
xor UO_583 (O_583,N_45078,N_45048);
nand UO_584 (O_584,N_45210,N_46736);
xor UO_585 (O_585,N_49836,N_45741);
nand UO_586 (O_586,N_48562,N_48506);
nor UO_587 (O_587,N_49255,N_47944);
nor UO_588 (O_588,N_47090,N_46595);
nor UO_589 (O_589,N_49650,N_45425);
or UO_590 (O_590,N_47317,N_49069);
xnor UO_591 (O_591,N_48926,N_45230);
nor UO_592 (O_592,N_46933,N_45047);
xnor UO_593 (O_593,N_45214,N_45451);
or UO_594 (O_594,N_48863,N_46991);
or UO_595 (O_595,N_46329,N_46807);
or UO_596 (O_596,N_49652,N_48732);
and UO_597 (O_597,N_45640,N_49362);
and UO_598 (O_598,N_46399,N_47718);
and UO_599 (O_599,N_48713,N_48053);
or UO_600 (O_600,N_49787,N_48499);
xor UO_601 (O_601,N_47142,N_46978);
and UO_602 (O_602,N_47626,N_45175);
xnor UO_603 (O_603,N_49673,N_48709);
nand UO_604 (O_604,N_49594,N_46487);
nand UO_605 (O_605,N_45789,N_45328);
and UO_606 (O_606,N_45695,N_45441);
nor UO_607 (O_607,N_45498,N_49876);
or UO_608 (O_608,N_47122,N_46674);
nand UO_609 (O_609,N_46507,N_48906);
or UO_610 (O_610,N_46692,N_49860);
xor UO_611 (O_611,N_46749,N_46468);
nand UO_612 (O_612,N_48019,N_48770);
xor UO_613 (O_613,N_46990,N_48032);
nand UO_614 (O_614,N_48690,N_46033);
and UO_615 (O_615,N_48358,N_46185);
nand UO_616 (O_616,N_45997,N_45199);
and UO_617 (O_617,N_47618,N_49989);
xor UO_618 (O_618,N_47735,N_49238);
nor UO_619 (O_619,N_45928,N_48908);
xor UO_620 (O_620,N_47061,N_45139);
nor UO_621 (O_621,N_49906,N_48119);
and UO_622 (O_622,N_46802,N_48637);
xor UO_623 (O_623,N_47211,N_48147);
nor UO_624 (O_624,N_47509,N_49593);
and UO_625 (O_625,N_48639,N_46889);
and UO_626 (O_626,N_47319,N_48150);
nor UO_627 (O_627,N_47676,N_45042);
or UO_628 (O_628,N_47148,N_45968);
nand UO_629 (O_629,N_48739,N_49684);
nand UO_630 (O_630,N_49531,N_48179);
xnor UO_631 (O_631,N_49418,N_47485);
xnor UO_632 (O_632,N_49999,N_45157);
and UO_633 (O_633,N_46134,N_46524);
and UO_634 (O_634,N_48466,N_46659);
nor UO_635 (O_635,N_47414,N_48365);
and UO_636 (O_636,N_45675,N_47027);
nand UO_637 (O_637,N_47024,N_45702);
xnor UO_638 (O_638,N_49681,N_48497);
xor UO_639 (O_639,N_45710,N_45091);
and UO_640 (O_640,N_46646,N_47564);
or UO_641 (O_641,N_46505,N_46309);
and UO_642 (O_642,N_48253,N_46240);
nor UO_643 (O_643,N_49515,N_47589);
nand UO_644 (O_644,N_49173,N_46467);
nor UO_645 (O_645,N_45639,N_48933);
nand UO_646 (O_646,N_48440,N_49775);
or UO_647 (O_647,N_46250,N_48168);
or UO_648 (O_648,N_49059,N_47083);
xor UO_649 (O_649,N_49435,N_47647);
and UO_650 (O_650,N_49201,N_48585);
nand UO_651 (O_651,N_45535,N_48507);
nand UO_652 (O_652,N_48647,N_47820);
and UO_653 (O_653,N_46886,N_49931);
xor UO_654 (O_654,N_46136,N_48825);
nand UO_655 (O_655,N_49958,N_49004);
nor UO_656 (O_656,N_47215,N_45683);
and UO_657 (O_657,N_47942,N_49896);
xnor UO_658 (O_658,N_45372,N_49063);
and UO_659 (O_659,N_45804,N_49299);
nand UO_660 (O_660,N_47783,N_47275);
or UO_661 (O_661,N_46694,N_45776);
nand UO_662 (O_662,N_46901,N_45080);
or UO_663 (O_663,N_46045,N_46567);
nand UO_664 (O_664,N_48998,N_49982);
or UO_665 (O_665,N_46409,N_47816);
xnor UO_666 (O_666,N_46126,N_48676);
nand UO_667 (O_667,N_47998,N_48433);
or UO_668 (O_668,N_48009,N_48187);
or UO_669 (O_669,N_45187,N_48228);
xnor UO_670 (O_670,N_46235,N_49112);
nor UO_671 (O_671,N_48843,N_48124);
nand UO_672 (O_672,N_46478,N_46048);
or UO_673 (O_673,N_45280,N_46454);
and UO_674 (O_674,N_49659,N_48629);
or UO_675 (O_675,N_46171,N_47044);
nand UO_676 (O_676,N_47043,N_47389);
or UO_677 (O_677,N_48938,N_46601);
and UO_678 (O_678,N_46472,N_49184);
xnor UO_679 (O_679,N_46453,N_47669);
xnor UO_680 (O_680,N_48508,N_46407);
nand UO_681 (O_681,N_47050,N_47190);
nor UO_682 (O_682,N_46455,N_46343);
nor UO_683 (O_683,N_48729,N_47141);
xnor UO_684 (O_684,N_45145,N_45988);
or UO_685 (O_685,N_46159,N_48609);
or UO_686 (O_686,N_48571,N_48409);
xor UO_687 (O_687,N_46725,N_47749);
xor UO_688 (O_688,N_45256,N_48930);
nand UO_689 (O_689,N_45761,N_46077);
and UO_690 (O_690,N_48790,N_45407);
xnor UO_691 (O_691,N_49093,N_46360);
nand UO_692 (O_692,N_47933,N_46746);
or UO_693 (O_693,N_46010,N_46687);
nor UO_694 (O_694,N_46480,N_46090);
and UO_695 (O_695,N_46466,N_47339);
xor UO_696 (O_696,N_48678,N_49245);
or UO_697 (O_697,N_45158,N_48223);
nor UO_698 (O_698,N_49655,N_46198);
xnor UO_699 (O_699,N_48456,N_47843);
or UO_700 (O_700,N_47201,N_47098);
or UO_701 (O_701,N_47456,N_46191);
or UO_702 (O_702,N_45160,N_47779);
or UO_703 (O_703,N_47526,N_46804);
nor UO_704 (O_704,N_46860,N_45018);
xor UO_705 (O_705,N_47175,N_46279);
nor UO_706 (O_706,N_48492,N_48965);
and UO_707 (O_707,N_48939,N_46738);
and UO_708 (O_708,N_47897,N_48313);
and UO_709 (O_709,N_45397,N_48730);
xnor UO_710 (O_710,N_46670,N_45177);
nand UO_711 (O_711,N_49111,N_46758);
xor UO_712 (O_712,N_48132,N_47644);
xnor UO_713 (O_713,N_48717,N_47445);
and UO_714 (O_714,N_48470,N_48632);
nor UO_715 (O_715,N_46628,N_45445);
nor UO_716 (O_716,N_48809,N_47409);
xnor UO_717 (O_717,N_45335,N_45517);
nand UO_718 (O_718,N_45918,N_47666);
and UO_719 (O_719,N_47439,N_45778);
xor UO_720 (O_720,N_45075,N_46895);
or UO_721 (O_721,N_47627,N_46875);
nor UO_722 (O_722,N_47405,N_45697);
nand UO_723 (O_723,N_47291,N_45626);
xnor UO_724 (O_724,N_45130,N_49772);
nand UO_725 (O_725,N_49844,N_45392);
nand UO_726 (O_726,N_45236,N_45179);
xnor UO_727 (O_727,N_46542,N_47582);
xor UO_728 (O_728,N_45486,N_47488);
or UO_729 (O_729,N_46988,N_49522);
xor UO_730 (O_730,N_49554,N_49082);
or UO_731 (O_731,N_47006,N_46456);
or UO_732 (O_732,N_46633,N_48694);
or UO_733 (O_733,N_46854,N_45439);
or UO_734 (O_734,N_45337,N_45775);
xor UO_735 (O_735,N_48415,N_49205);
nand UO_736 (O_736,N_49578,N_45222);
and UO_737 (O_737,N_47294,N_47901);
nand UO_738 (O_738,N_48390,N_47067);
xnor UO_739 (O_739,N_46379,N_49666);
and UO_740 (O_740,N_48605,N_47241);
or UO_741 (O_741,N_49872,N_47506);
or UO_742 (O_742,N_45768,N_47073);
or UO_743 (O_743,N_47335,N_48205);
nand UO_744 (O_744,N_46723,N_46215);
nand UO_745 (O_745,N_47575,N_48234);
and UO_746 (O_746,N_46743,N_48336);
nor UO_747 (O_747,N_47239,N_45847);
xor UO_748 (O_748,N_46610,N_47029);
nand UO_749 (O_749,N_48166,N_49482);
nor UO_750 (O_750,N_49660,N_46093);
xor UO_751 (O_751,N_47802,N_46072);
nand UO_752 (O_752,N_45641,N_45001);
nor UO_753 (O_753,N_48971,N_48991);
nor UO_754 (O_754,N_49424,N_49672);
nand UO_755 (O_755,N_47344,N_47013);
xnor UO_756 (O_756,N_48953,N_45272);
or UO_757 (O_757,N_48817,N_49079);
or UO_758 (O_758,N_46441,N_49320);
or UO_759 (O_759,N_45190,N_48370);
and UO_760 (O_760,N_49138,N_47833);
nand UO_761 (O_761,N_45072,N_45876);
xnor UO_762 (O_762,N_47960,N_46106);
and UO_763 (O_763,N_46673,N_45945);
nor UO_764 (O_764,N_45312,N_46865);
or UO_765 (O_765,N_49145,N_46929);
and UO_766 (O_766,N_48304,N_45215);
nor UO_767 (O_767,N_49156,N_49284);
or UO_768 (O_768,N_46727,N_45102);
nand UO_769 (O_769,N_46280,N_45066);
nor UO_770 (O_770,N_47809,N_46651);
nor UO_771 (O_771,N_45069,N_45579);
nor UO_772 (O_772,N_48750,N_47060);
and UO_773 (O_773,N_47035,N_46681);
nand UO_774 (O_774,N_48154,N_49441);
or UO_775 (O_775,N_49778,N_45213);
xnor UO_776 (O_776,N_48069,N_47070);
xor UO_777 (O_777,N_48262,N_48599);
nand UO_778 (O_778,N_45780,N_48490);
or UO_779 (O_779,N_47105,N_49566);
or UO_780 (O_780,N_47611,N_46286);
and UO_781 (O_781,N_45592,N_45039);
nand UO_782 (O_782,N_47002,N_46608);
and UO_783 (O_783,N_47950,N_45669);
nor UO_784 (O_784,N_46741,N_48286);
xnor UO_785 (O_785,N_47367,N_49861);
and UO_786 (O_786,N_48273,N_49661);
nand UO_787 (O_787,N_49064,N_49444);
and UO_788 (O_788,N_45472,N_47351);
and UO_789 (O_789,N_47140,N_45743);
nor UO_790 (O_790,N_48641,N_45524);
xnor UO_791 (O_791,N_46869,N_45376);
and UO_792 (O_792,N_46984,N_47316);
or UO_793 (O_793,N_46906,N_49016);
xor UO_794 (O_794,N_48881,N_46311);
xor UO_795 (O_795,N_47590,N_46028);
and UO_796 (O_796,N_48973,N_45131);
nand UO_797 (O_797,N_45607,N_48580);
and UO_798 (O_798,N_45251,N_49960);
nand UO_799 (O_799,N_46237,N_49372);
or UO_800 (O_800,N_48734,N_47126);
and UO_801 (O_801,N_47350,N_49337);
nor UO_802 (O_802,N_45910,N_46761);
or UO_803 (O_803,N_48538,N_47667);
nand UO_804 (O_804,N_45204,N_48476);
nor UO_805 (O_805,N_46449,N_45647);
and UO_806 (O_806,N_47332,N_46704);
or UO_807 (O_807,N_49727,N_49553);
or UO_808 (O_808,N_48199,N_47124);
and UO_809 (O_809,N_46448,N_48174);
xor UO_810 (O_810,N_49977,N_46385);
or UO_811 (O_811,N_45478,N_47830);
or UO_812 (O_812,N_45321,N_49129);
xnor UO_813 (O_813,N_47650,N_48125);
nor UO_814 (O_814,N_47089,N_47046);
and UO_815 (O_815,N_47458,N_49322);
or UO_816 (O_816,N_49058,N_46535);
xnor UO_817 (O_817,N_45095,N_46540);
nand UO_818 (O_818,N_48724,N_48041);
xnor UO_819 (O_819,N_47136,N_48934);
xnor UO_820 (O_820,N_45393,N_46345);
or UO_821 (O_821,N_47623,N_47213);
xor UO_822 (O_822,N_49834,N_48288);
nand UO_823 (O_823,N_49114,N_48600);
or UO_824 (O_824,N_47227,N_47022);
or UO_825 (O_825,N_47366,N_46916);
or UO_826 (O_826,N_48146,N_47282);
or UO_827 (O_827,N_46947,N_49535);
nor UO_828 (O_828,N_45844,N_47476);
nand UO_829 (O_829,N_48338,N_45196);
or UO_830 (O_830,N_49021,N_45822);
and UO_831 (O_831,N_48230,N_45950);
nand UO_832 (O_832,N_48989,N_48261);
nor UO_833 (O_833,N_47987,N_46098);
and UO_834 (O_834,N_47115,N_45875);
nand UO_835 (O_835,N_49980,N_46799);
or UO_836 (O_836,N_47766,N_45739);
and UO_837 (O_837,N_46446,N_47009);
xor UO_838 (O_838,N_45200,N_47395);
and UO_839 (O_839,N_45802,N_49994);
and UO_840 (O_840,N_49886,N_48536);
nand UO_841 (O_841,N_49635,N_49379);
xnor UO_842 (O_842,N_46710,N_46757);
xor UO_843 (O_843,N_48353,N_49663);
nand UO_844 (O_844,N_47531,N_49413);
xor UO_845 (O_845,N_48361,N_45901);
or UO_846 (O_846,N_46513,N_47171);
nor UO_847 (O_847,N_49315,N_49607);
xnor UO_848 (O_848,N_49382,N_48428);
nand UO_849 (O_849,N_46766,N_47082);
or UO_850 (O_850,N_48001,N_47259);
nand UO_851 (O_851,N_45883,N_47544);
nor UO_852 (O_852,N_47864,N_45430);
nand UO_853 (O_853,N_48317,N_47639);
nor UO_854 (O_854,N_48294,N_47630);
nand UO_855 (O_855,N_46686,N_45976);
nor UO_856 (O_856,N_45525,N_49135);
xor UO_857 (O_857,N_49270,N_47871);
nand UO_858 (O_858,N_48046,N_49862);
and UO_859 (O_859,N_49446,N_48927);
nor UO_860 (O_860,N_47737,N_45566);
or UO_861 (O_861,N_49817,N_47680);
nor UO_862 (O_862,N_48447,N_48207);
or UO_863 (O_863,N_46624,N_45658);
and UO_864 (O_864,N_49598,N_46095);
nor UO_865 (O_865,N_46403,N_49962);
nand UO_866 (O_866,N_45629,N_47965);
nor UO_867 (O_867,N_46848,N_45966);
xor UO_868 (O_868,N_48755,N_45495);
xor UO_869 (O_869,N_48798,N_45325);
and UO_870 (O_870,N_47158,N_45646);
nor UO_871 (O_871,N_47714,N_48251);
nand UO_872 (O_872,N_48026,N_46671);
nor UO_873 (O_873,N_49979,N_48081);
nor UO_874 (O_874,N_49899,N_49855);
nand UO_875 (O_875,N_48303,N_45044);
nor UO_876 (O_876,N_45596,N_46000);
or UO_877 (O_877,N_46015,N_46157);
xor UO_878 (O_878,N_47396,N_48544);
xor UO_879 (O_879,N_48331,N_48281);
and UO_880 (O_880,N_45103,N_47841);
xor UO_881 (O_881,N_48695,N_47354);
nand UO_882 (O_882,N_46153,N_45434);
and UO_883 (O_883,N_45404,N_47102);
xnor UO_884 (O_884,N_45718,N_46374);
nand UO_885 (O_885,N_49330,N_48439);
and UO_886 (O_886,N_48917,N_46227);
nand UO_887 (O_887,N_47761,N_48202);
and UO_888 (O_888,N_45234,N_46593);
xnor UO_889 (O_889,N_48616,N_46012);
nand UO_890 (O_890,N_49483,N_49157);
and UO_891 (O_891,N_48037,N_48240);
xor UO_892 (O_892,N_49698,N_47767);
and UO_893 (O_893,N_45485,N_45007);
xnor UO_894 (O_894,N_45891,N_46055);
xnor UO_895 (O_895,N_47340,N_45421);
nand UO_896 (O_896,N_45671,N_46111);
nand UO_897 (O_897,N_49196,N_48467);
nand UO_898 (O_898,N_47427,N_45634);
nand UO_899 (O_899,N_49202,N_48877);
or UO_900 (O_900,N_49174,N_47889);
or UO_901 (O_901,N_45872,N_47991);
xor UO_902 (O_902,N_47549,N_49582);
nor UO_903 (O_903,N_49526,N_49756);
or UO_904 (O_904,N_47313,N_46160);
xor UO_905 (O_905,N_45419,N_46200);
nand UO_906 (O_906,N_49744,N_45773);
nand UO_907 (O_907,N_47185,N_47246);
or UO_908 (O_908,N_49359,N_46867);
and UO_909 (O_909,N_47421,N_48944);
xnor UO_910 (O_910,N_49278,N_45593);
xnor UO_911 (O_911,N_48556,N_46698);
and UO_912 (O_912,N_48681,N_46244);
or UO_913 (O_913,N_46473,N_48096);
xor UO_914 (O_914,N_49344,N_45835);
xnor UO_915 (O_915,N_48023,N_49990);
nor UO_916 (O_916,N_45391,N_47631);
nor UO_917 (O_917,N_48103,N_47152);
nand UO_918 (O_918,N_46356,N_47279);
nor UO_919 (O_919,N_48098,N_46844);
nand UO_920 (O_920,N_47495,N_48769);
nor UO_921 (O_921,N_46068,N_47643);
nor UO_922 (O_922,N_47240,N_47195);
nand UO_923 (O_923,N_47675,N_46970);
and UO_924 (O_924,N_45195,N_46481);
xnor UO_925 (O_925,N_46667,N_49615);
xor UO_926 (O_926,N_48151,N_46423);
nor UO_927 (O_927,N_45194,N_46855);
nor UO_928 (O_928,N_49302,N_45598);
or UO_929 (O_929,N_45828,N_48574);
or UO_930 (O_930,N_48010,N_46004);
nor UO_931 (O_931,N_48532,N_45061);
and UO_932 (O_932,N_45748,N_45895);
xor UO_933 (O_933,N_46251,N_47243);
nand UO_934 (O_934,N_47047,N_46312);
xnor UO_935 (O_935,N_47011,N_47810);
or UO_936 (O_936,N_48716,N_48889);
nor UO_937 (O_937,N_49015,N_46533);
and UO_938 (O_938,N_46530,N_45526);
nand UO_939 (O_939,N_49503,N_47208);
nor UO_940 (O_940,N_46868,N_49095);
nand UO_941 (O_941,N_47733,N_45612);
nor UO_942 (O_942,N_47144,N_48674);
nor UO_943 (O_943,N_49394,N_45758);
xor UO_944 (O_944,N_46926,N_47839);
nand UO_945 (O_945,N_47568,N_45367);
and UO_946 (O_946,N_49995,N_46706);
and UO_947 (O_947,N_46944,N_45355);
or UO_948 (O_948,N_48721,N_45431);
and UO_949 (O_949,N_47375,N_48429);
or UO_950 (O_950,N_45088,N_47595);
nor UO_951 (O_951,N_45123,N_47327);
or UO_952 (O_952,N_45003,N_47473);
xnor UO_953 (O_953,N_46863,N_46680);
xnor UO_954 (O_954,N_48344,N_46392);
nand UO_955 (O_955,N_49776,N_47727);
nand UO_956 (O_956,N_45022,N_45505);
nor UO_957 (O_957,N_45174,N_45354);
nor UO_958 (O_958,N_45806,N_46433);
and UO_959 (O_959,N_46830,N_48612);
and UO_960 (O_960,N_49743,N_46833);
nand UO_961 (O_961,N_45698,N_46644);
and UO_962 (O_962,N_48534,N_48707);
and UO_963 (O_963,N_47969,N_47374);
xnor UO_964 (O_964,N_45528,N_46500);
or UO_965 (O_965,N_46105,N_48797);
nor UO_966 (O_966,N_48535,N_48818);
xnor UO_967 (O_967,N_46129,N_45220);
nor UO_968 (O_968,N_49794,N_48008);
nand UO_969 (O_969,N_46415,N_48921);
and UO_970 (O_970,N_48627,N_45678);
xnor UO_971 (O_971,N_46675,N_45041);
and UO_972 (O_972,N_45264,N_45693);
nand UO_973 (O_973,N_45165,N_47472);
xor UO_974 (O_974,N_45764,N_49116);
or UO_975 (O_975,N_45996,N_46648);
and UO_976 (O_976,N_47133,N_45414);
and UO_977 (O_977,N_48025,N_47440);
or UO_978 (O_978,N_49696,N_45105);
xnor UO_979 (O_979,N_49722,N_46114);
xnor UO_980 (O_980,N_48249,N_46935);
or UO_981 (O_981,N_45774,N_45480);
nand UO_982 (O_982,N_48961,N_48725);
xnor UO_983 (O_983,N_46435,N_47678);
nor UO_984 (O_984,N_47165,N_47709);
and UO_985 (O_985,N_48657,N_46354);
or UO_986 (O_986,N_47135,N_49094);
xor UO_987 (O_987,N_45387,N_46952);
nor UO_988 (O_988,N_49139,N_47719);
or UO_989 (O_989,N_49356,N_49765);
and UO_990 (O_990,N_49287,N_46275);
or UO_991 (O_991,N_45690,N_47963);
or UO_992 (O_992,N_49713,N_47450);
nor UO_993 (O_993,N_49555,N_46662);
and UO_994 (O_994,N_47565,N_45568);
or UO_995 (O_995,N_45907,N_48728);
nand UO_996 (O_996,N_48613,N_47117);
nor UO_997 (O_997,N_46688,N_49909);
or UO_998 (O_998,N_49455,N_46241);
xnor UO_999 (O_999,N_45163,N_48667);
and UO_1000 (O_1000,N_45846,N_47499);
nand UO_1001 (O_1001,N_46063,N_45363);
and UO_1002 (O_1002,N_48878,N_48845);
xnor UO_1003 (O_1003,N_48185,N_45644);
nor UO_1004 (O_1004,N_46334,N_48479);
or UO_1005 (O_1005,N_48795,N_47765);
nand UO_1006 (O_1006,N_48071,N_45762);
xnor UO_1007 (O_1007,N_45424,N_45197);
or UO_1008 (O_1008,N_45892,N_45994);
nand UO_1009 (O_1009,N_49172,N_49825);
nor UO_1010 (O_1010,N_48911,N_49080);
nand UO_1011 (O_1011,N_48318,N_46172);
nand UO_1012 (O_1012,N_45676,N_49620);
or UO_1013 (O_1013,N_45831,N_45036);
xor UO_1014 (O_1014,N_48300,N_48134);
nand UO_1015 (O_1015,N_45905,N_46451);
or UO_1016 (O_1016,N_49169,N_45807);
and UO_1017 (O_1017,N_46352,N_45812);
and UO_1018 (O_1018,N_49028,N_45346);
or UO_1019 (O_1019,N_45293,N_47578);
nor UO_1020 (O_1020,N_49313,N_49974);
xor UO_1021 (O_1021,N_47930,N_46450);
and UO_1022 (O_1022,N_46665,N_47831);
nor UO_1023 (O_1023,N_48787,N_46545);
or UO_1024 (O_1024,N_47826,N_49389);
xnor UO_1025 (O_1025,N_49318,N_47903);
nor UO_1026 (O_1026,N_47840,N_49403);
nor UO_1027 (O_1027,N_47928,N_45244);
and UO_1028 (O_1028,N_48250,N_46857);
xnor UO_1029 (O_1029,N_45959,N_47988);
nor UO_1030 (O_1030,N_49951,N_49300);
and UO_1031 (O_1031,N_46616,N_47621);
and UO_1032 (O_1032,N_49124,N_49966);
or UO_1033 (O_1033,N_49728,N_49588);
nor UO_1034 (O_1034,N_48193,N_45025);
nand UO_1035 (O_1035,N_46619,N_45296);
nand UO_1036 (O_1036,N_49295,N_47524);
xnor UO_1037 (O_1037,N_47547,N_46274);
nand UO_1038 (O_1038,N_47261,N_49774);
nand UO_1039 (O_1039,N_45467,N_46713);
nor UO_1040 (O_1040,N_47945,N_46890);
nand UO_1041 (O_1041,N_45541,N_45787);
or UO_1042 (O_1042,N_46204,N_49428);
nand UO_1043 (O_1043,N_46398,N_47487);
nand UO_1044 (O_1044,N_46800,N_49430);
and UO_1045 (O_1045,N_47562,N_46653);
or UO_1046 (O_1046,N_49032,N_45680);
and UO_1047 (O_1047,N_48500,N_49587);
nor UO_1048 (O_1048,N_46056,N_48235);
nand UO_1049 (O_1049,N_45057,N_46307);
or UO_1050 (O_1050,N_45307,N_45227);
nand UO_1051 (O_1051,N_49550,N_48421);
nor UO_1052 (O_1052,N_49658,N_46777);
nor UO_1053 (O_1053,N_49849,N_48658);
xor UO_1054 (O_1054,N_46957,N_48293);
nor UO_1055 (O_1055,N_47411,N_46985);
xnor UO_1056 (O_1056,N_48683,N_46104);
or UO_1057 (O_1057,N_49736,N_45460);
xnor UO_1058 (O_1058,N_47402,N_45226);
and UO_1059 (O_1059,N_46823,N_46790);
xnor UO_1060 (O_1060,N_47523,N_48873);
nand UO_1061 (O_1061,N_47645,N_46765);
nor UO_1062 (O_1062,N_46490,N_47715);
nand UO_1063 (O_1063,N_45965,N_45333);
and UO_1064 (O_1064,N_46246,N_47701);
xnor UO_1065 (O_1065,N_47883,N_49286);
nor UO_1066 (O_1066,N_48834,N_48762);
or UO_1067 (O_1067,N_47982,N_46268);
or UO_1068 (O_1068,N_49911,N_47567);
xor UO_1069 (O_1069,N_49230,N_49062);
or UO_1070 (O_1070,N_49381,N_49485);
or UO_1071 (O_1071,N_45099,N_48054);
xor UO_1072 (O_1072,N_48394,N_49711);
and UO_1073 (O_1073,N_47688,N_46583);
nor UO_1074 (O_1074,N_47914,N_48624);
xnor UO_1075 (O_1075,N_48956,N_47619);
and UO_1076 (O_1076,N_46592,N_46040);
nor UO_1077 (O_1077,N_45521,N_48445);
nand UO_1078 (O_1078,N_49070,N_47020);
nand UO_1079 (O_1079,N_45385,N_46613);
xor UO_1080 (O_1080,N_47640,N_46042);
or UO_1081 (O_1081,N_49025,N_47410);
or UO_1082 (O_1082,N_49442,N_45473);
nand UO_1083 (O_1083,N_49667,N_47964);
and UO_1084 (O_1084,N_49340,N_47571);
and UO_1085 (O_1085,N_47583,N_47400);
nor UO_1086 (O_1086,N_48879,N_46050);
nor UO_1087 (O_1087,N_45580,N_45448);
nand UO_1088 (O_1088,N_48048,N_48047);
nand UO_1089 (O_1089,N_45247,N_45935);
nand UO_1090 (O_1090,N_45503,N_48237);
xnor UO_1091 (O_1091,N_49950,N_48209);
or UO_1092 (O_1092,N_45692,N_46714);
nand UO_1093 (O_1093,N_45888,N_47881);
and UO_1094 (O_1094,N_49946,N_47346);
nand UO_1095 (O_1095,N_47699,N_48113);
nor UO_1096 (O_1096,N_48858,N_46969);
nor UO_1097 (O_1097,N_45141,N_45413);
xor UO_1098 (O_1098,N_47116,N_45006);
nand UO_1099 (O_1099,N_48570,N_47248);
xnor UO_1100 (O_1100,N_45757,N_46666);
xor UO_1101 (O_1101,N_48782,N_49366);
xor UO_1102 (O_1102,N_49687,N_47822);
or UO_1103 (O_1103,N_47042,N_47862);
nand UO_1104 (O_1104,N_47265,N_45666);
nor UO_1105 (O_1105,N_46281,N_47475);
and UO_1106 (O_1106,N_45560,N_46269);
nor UO_1107 (O_1107,N_49131,N_46438);
or UO_1108 (O_1108,N_45729,N_48523);
nor UO_1109 (O_1109,N_47127,N_45574);
nor UO_1110 (O_1110,N_45259,N_49158);
and UO_1111 (O_1111,N_48857,N_49549);
or UO_1112 (O_1112,N_46330,N_48329);
nand UO_1113 (O_1113,N_45765,N_45800);
nand UO_1114 (O_1114,N_46314,N_47554);
nand UO_1115 (O_1115,N_48316,N_49346);
nand UO_1116 (O_1116,N_46233,N_48120);
nor UO_1117 (O_1117,N_46989,N_48775);
nand UO_1118 (O_1118,N_49602,N_46693);
xor UO_1119 (O_1119,N_46789,N_46318);
nand UO_1120 (O_1120,N_46635,N_47580);
nor UO_1121 (O_1121,N_45290,N_46609);
and UO_1122 (O_1122,N_46813,N_49692);
xnor UO_1123 (O_1123,N_45170,N_48104);
and UO_1124 (O_1124,N_47696,N_48121);
or UO_1125 (O_1125,N_47778,N_49847);
nand UO_1126 (O_1126,N_45399,N_48967);
xor UO_1127 (O_1127,N_45677,N_49608);
or UO_1128 (O_1128,N_46025,N_46994);
xor UO_1129 (O_1129,N_47461,N_45100);
or UO_1130 (O_1130,N_49866,N_46444);
nor UO_1131 (O_1131,N_45534,N_46596);
and UO_1132 (O_1132,N_48226,N_49383);
nand UO_1133 (O_1133,N_45149,N_47848);
xnor UO_1134 (O_1134,N_49614,N_45584);
nand UO_1135 (O_1135,N_46689,N_46887);
or UO_1136 (O_1136,N_46412,N_45051);
nand UO_1137 (O_1137,N_48673,N_48385);
nor UO_1138 (O_1138,N_47428,N_48975);
and UO_1139 (O_1139,N_48090,N_46238);
and UO_1140 (O_1140,N_48771,N_46645);
xor UO_1141 (O_1141,N_49479,N_47069);
and UO_1142 (O_1142,N_48310,N_47203);
and UO_1143 (O_1143,N_47660,N_49586);
nand UO_1144 (O_1144,N_46373,N_45848);
and UO_1145 (O_1145,N_47355,N_46788);
nand UO_1146 (O_1146,N_46432,N_46930);
or UO_1147 (O_1147,N_47866,N_49596);
nor UO_1148 (O_1148,N_48592,N_45555);
xor UO_1149 (O_1149,N_46096,N_45017);
and UO_1150 (O_1150,N_47091,N_47934);
nand UO_1151 (O_1151,N_46537,N_48660);
or UO_1152 (O_1152,N_49867,N_49953);
nor UO_1153 (O_1153,N_45043,N_49818);
xor UO_1154 (O_1154,N_48206,N_45712);
and UO_1155 (O_1155,N_47653,N_46333);
nand UO_1156 (O_1156,N_49068,N_45636);
or UO_1157 (O_1157,N_49764,N_49912);
nor UO_1158 (O_1158,N_45977,N_46657);
and UO_1159 (O_1159,N_46522,N_47443);
or UO_1160 (O_1160,N_46141,N_45297);
nand UO_1161 (O_1161,N_48896,N_48549);
and UO_1162 (O_1162,N_46951,N_48509);
or UO_1163 (O_1163,N_49334,N_46218);
nand UO_1164 (O_1164,N_48448,N_47154);
nor UO_1165 (O_1165,N_46769,N_49451);
nor UO_1166 (O_1166,N_46331,N_49653);
nand UO_1167 (O_1167,N_48999,N_49013);
xor UO_1168 (O_1168,N_49998,N_49603);
xor UO_1169 (O_1169,N_47109,N_46827);
xor UO_1170 (O_1170,N_49273,N_49464);
and UO_1171 (O_1171,N_47376,N_48195);
and UO_1172 (O_1172,N_49352,N_49186);
nor UO_1173 (O_1173,N_47657,N_45416);
and UO_1174 (O_1174,N_49718,N_46109);
or UO_1175 (O_1175,N_46395,N_47729);
xor UO_1176 (O_1176,N_48411,N_45597);
nor UO_1177 (O_1177,N_49471,N_46301);
or UO_1178 (O_1178,N_46587,N_46836);
or UO_1179 (O_1179,N_47921,N_46660);
or UO_1180 (O_1180,N_46753,N_47538);
nor UO_1181 (O_1181,N_45999,N_47579);
nor UO_1182 (O_1182,N_46647,N_46300);
nand UO_1183 (O_1183,N_48252,N_46594);
nor UO_1184 (O_1184,N_47103,N_48550);
and UO_1185 (O_1185,N_47519,N_46707);
or UO_1186 (O_1186,N_45575,N_48280);
nor UO_1187 (O_1187,N_48259,N_49488);
or UO_1188 (O_1188,N_47967,N_45446);
xor UO_1189 (O_1189,N_46576,N_45684);
and UO_1190 (O_1190,N_47948,N_48567);
nand UO_1191 (O_1191,N_46020,N_46262);
nand UO_1192 (O_1192,N_45681,N_49725);
nand UO_1193 (O_1193,N_48420,N_45749);
nand UO_1194 (O_1194,N_49561,N_46219);
or UO_1195 (O_1195,N_48389,N_48799);
nor UO_1196 (O_1196,N_49961,N_47632);
nand UO_1197 (O_1197,N_49258,N_49146);
xnor UO_1198 (O_1198,N_48065,N_47514);
nor UO_1199 (O_1199,N_49956,N_49486);
or UO_1200 (O_1200,N_47033,N_48852);
and UO_1201 (O_1201,N_45305,N_47383);
xor UO_1202 (O_1202,N_46871,N_49045);
nor UO_1203 (O_1203,N_49475,N_47616);
nand UO_1204 (O_1204,N_49182,N_49926);
or UO_1205 (O_1205,N_47408,N_49358);
and UO_1206 (O_1206,N_48123,N_49611);
xor UO_1207 (O_1207,N_47418,N_47915);
or UO_1208 (O_1208,N_49811,N_45242);
xor UO_1209 (O_1209,N_48116,N_47919);
nor UO_1210 (O_1210,N_46872,N_45985);
nor UO_1211 (O_1211,N_48348,N_47094);
and UO_1212 (O_1212,N_48351,N_49864);
nand UO_1213 (O_1213,N_48970,N_46405);
nand UO_1214 (O_1214,N_49884,N_46733);
and UO_1215 (O_1215,N_49031,N_48360);
xnor UO_1216 (O_1216,N_45442,N_49704);
xor UO_1217 (O_1217,N_49854,N_47167);
nand UO_1218 (O_1218,N_45938,N_45302);
nor UO_1219 (O_1219,N_49304,N_47832);
nor UO_1220 (O_1220,N_45329,N_47909);
and UO_1221 (O_1221,N_46521,N_48216);
and UO_1222 (O_1222,N_46810,N_47177);
nand UO_1223 (O_1223,N_45939,N_49707);
nor UO_1224 (O_1224,N_47823,N_48083);
xnor UO_1225 (O_1225,N_48980,N_46340);
and UO_1226 (O_1226,N_45023,N_48573);
and UO_1227 (O_1227,N_49073,N_48747);
nand UO_1228 (O_1228,N_47710,N_48767);
nor UO_1229 (O_1229,N_46146,N_49422);
nand UO_1230 (O_1230,N_49216,N_48027);
nor UO_1231 (O_1231,N_46965,N_47811);
and UO_1232 (O_1232,N_45056,N_49932);
and UO_1233 (O_1233,N_48801,N_47847);
or UO_1234 (O_1234,N_45140,N_45049);
nand UO_1235 (O_1235,N_47712,N_45144);
nand UO_1236 (O_1236,N_45694,N_48274);
nand UO_1237 (O_1237,N_49193,N_46429);
nor UO_1238 (O_1238,N_45557,N_45268);
and UO_1239 (O_1239,N_45323,N_48940);
nand UO_1240 (O_1240,N_46782,N_46196);
xor UO_1241 (O_1241,N_48231,N_47559);
and UO_1242 (O_1242,N_48645,N_46905);
or UO_1243 (O_1243,N_48471,N_48672);
and UO_1244 (O_1244,N_45599,N_45189);
nand UO_1245 (O_1245,N_47016,N_46849);
or UO_1246 (O_1246,N_46132,N_49266);
nor UO_1247 (O_1247,N_48221,N_48106);
nand UO_1248 (O_1248,N_48751,N_47596);
nor UO_1249 (O_1249,N_49074,N_46742);
and UO_1250 (O_1250,N_48979,N_48056);
nor UO_1251 (O_1251,N_46367,N_46005);
nand UO_1252 (O_1252,N_49452,N_46442);
and UO_1253 (O_1253,N_49925,N_45811);
nor UO_1254 (O_1254,N_48559,N_46911);
or UO_1255 (O_1255,N_45512,N_47746);
nor UO_1256 (O_1256,N_49458,N_47274);
nand UO_1257 (O_1257,N_48449,N_47231);
or UO_1258 (O_1258,N_45719,N_48321);
and UO_1259 (O_1259,N_48758,N_48061);
nor UO_1260 (O_1260,N_48464,N_46447);
or UO_1261 (O_1261,N_49567,N_46602);
or UO_1262 (O_1262,N_49845,N_48108);
nand UO_1263 (O_1263,N_49803,N_45026);
nor UO_1264 (O_1264,N_49978,N_49647);
nor UO_1265 (O_1265,N_45922,N_45958);
xnor UO_1266 (O_1266,N_49077,N_49263);
and UO_1267 (O_1267,N_47162,N_49416);
nor UO_1268 (O_1268,N_46703,N_46013);
or UO_1269 (O_1269,N_47482,N_47471);
nor UO_1270 (O_1270,N_47747,N_47805);
or UO_1271 (O_1271,N_48255,N_49056);
nor UO_1272 (O_1272,N_49534,N_47610);
nand UO_1273 (O_1273,N_46502,N_49281);
nor UO_1274 (O_1274,N_47080,N_47194);
xnor UO_1275 (O_1275,N_45880,N_49606);
or UO_1276 (O_1276,N_48197,N_46672);
nor UO_1277 (O_1277,N_47147,N_47609);
xor UO_1278 (O_1278,N_47740,N_48652);
xnor UO_1279 (O_1279,N_49789,N_45357);
xor UO_1280 (O_1280,N_46966,N_49821);
nand UO_1281 (O_1281,N_47906,N_49955);
nand UO_1282 (O_1282,N_45469,N_47214);
nand UO_1283 (O_1283,N_48572,N_46956);
xnor UO_1284 (O_1284,N_47570,N_46417);
nand UO_1285 (O_1285,N_48194,N_49349);
or UO_1286 (O_1286,N_45651,N_48239);
nor UO_1287 (O_1287,N_45682,N_46568);
and UO_1288 (O_1288,N_47260,N_46760);
and UO_1289 (O_1289,N_47539,N_48016);
nor UO_1290 (O_1290,N_49677,N_45920);
nand UO_1291 (O_1291,N_46603,N_45824);
nor UO_1292 (O_1292,N_46163,N_49536);
and UO_1293 (O_1293,N_47202,N_47394);
xnor UO_1294 (O_1294,N_49306,N_46900);
nand UO_1295 (O_1295,N_45481,N_46821);
or UO_1296 (O_1296,N_48133,N_48701);
and UO_1297 (O_1297,N_48462,N_48143);
xnor UO_1298 (O_1298,N_49510,N_45852);
nand UO_1299 (O_1299,N_47711,N_49152);
nor UO_1300 (O_1300,N_47218,N_47671);
and UO_1301 (O_1301,N_47100,N_49113);
and UO_1302 (O_1302,N_47875,N_49558);
nor UO_1303 (O_1303,N_46463,N_48489);
and UO_1304 (O_1304,N_48165,N_45497);
or UO_1305 (O_1305,N_47188,N_46630);
nor UO_1306 (O_1306,N_48913,N_45070);
or UO_1307 (O_1307,N_47363,N_48102);
nor UO_1308 (O_1308,N_47059,N_48808);
nand UO_1309 (O_1309,N_49613,N_46941);
nor UO_1310 (O_1310,N_48457,N_49542);
xnor UO_1311 (O_1311,N_46029,N_45106);
xor UO_1312 (O_1312,N_45772,N_48017);
nor UO_1313 (O_1313,N_45384,N_45313);
xnor UO_1314 (O_1314,N_45382,N_47163);
nand UO_1315 (O_1315,N_47429,N_45582);
xor UO_1316 (O_1316,N_47814,N_49920);
and UO_1317 (O_1317,N_46054,N_48277);
nand UO_1318 (O_1318,N_46528,N_45338);
xor UO_1319 (O_1319,N_45202,N_49357);
and UO_1320 (O_1320,N_48791,N_47288);
nor UO_1321 (O_1321,N_46722,N_49552);
nor UO_1322 (O_1322,N_47774,N_46877);
or UO_1323 (O_1323,N_45792,N_47867);
nor UO_1324 (O_1324,N_46719,N_46726);
or UO_1325 (O_1325,N_49189,N_45015);
and UO_1326 (O_1326,N_45366,N_47131);
nor UO_1327 (O_1327,N_49759,N_49437);
or UO_1328 (O_1328,N_46626,N_49192);
nor UO_1329 (O_1329,N_46427,N_47181);
and UO_1330 (O_1330,N_46349,N_46032);
xnor UO_1331 (O_1331,N_49217,N_48886);
nand UO_1332 (O_1332,N_46167,N_46256);
nand UO_1333 (O_1333,N_47545,N_48800);
or UO_1334 (O_1334,N_47773,N_49377);
nor UO_1335 (O_1335,N_46987,N_49639);
or UO_1336 (O_1336,N_49234,N_47591);
nand UO_1337 (O_1337,N_46549,N_47380);
nor UO_1338 (O_1338,N_49292,N_48397);
and UO_1339 (O_1339,N_46364,N_48838);
or UO_1340 (O_1340,N_48144,N_46203);
xor UO_1341 (O_1341,N_45065,N_48689);
and UO_1342 (O_1342,N_46357,N_47899);
nor UO_1343 (O_1343,N_45991,N_48545);
and UO_1344 (O_1344,N_47432,N_48634);
and UO_1345 (O_1345,N_49490,N_47169);
or UO_1346 (O_1346,N_45271,N_49548);
and UO_1347 (O_1347,N_48958,N_46234);
nand UO_1348 (O_1348,N_49147,N_49506);
and UO_1349 (O_1349,N_48566,N_47468);
xnor UO_1350 (O_1350,N_46805,N_49798);
xnor UO_1351 (O_1351,N_46426,N_46193);
nor UO_1352 (O_1352,N_47232,N_49985);
and UO_1353 (O_1353,N_49190,N_45122);
and UO_1354 (O_1354,N_47128,N_46064);
xor UO_1355 (O_1355,N_47039,N_47001);
nor UO_1356 (O_1356,N_49410,N_48295);
and UO_1357 (O_1357,N_47088,N_47828);
and UO_1358 (O_1358,N_46370,N_45304);
xnor UO_1359 (O_1359,N_47153,N_49477);
xor UO_1360 (O_1360,N_45085,N_48525);
xor UO_1361 (O_1361,N_48711,N_45860);
or UO_1362 (O_1362,N_48052,N_48291);
nor UO_1363 (O_1363,N_49738,N_47996);
xor UO_1364 (O_1364,N_49473,N_48785);
nor UO_1365 (O_1365,N_49678,N_48434);
xor UO_1366 (O_1366,N_47173,N_49863);
or UO_1367 (O_1367,N_45946,N_45459);
nand UO_1368 (O_1368,N_49050,N_49797);
or UO_1369 (O_1369,N_46511,N_46683);
or UO_1370 (O_1370,N_45687,N_49748);
xor UO_1371 (O_1371,N_47815,N_48169);
and UO_1372 (O_1372,N_45135,N_46018);
xnor UO_1373 (O_1373,N_45453,N_49213);
xor UO_1374 (O_1374,N_49325,N_49583);
and UO_1375 (O_1375,N_48929,N_46979);
nand UO_1376 (O_1376,N_48883,N_48186);
xnor UO_1377 (O_1377,N_49103,N_46812);
xnor UO_1378 (O_1378,N_48278,N_46785);
or UO_1379 (O_1379,N_48826,N_45030);
xor UO_1380 (O_1380,N_49853,N_45531);
nand UO_1381 (O_1381,N_49682,N_49327);
xnor UO_1382 (O_1382,N_47125,N_49528);
or UO_1383 (O_1383,N_45904,N_45456);
nor UO_1384 (O_1384,N_46543,N_49242);
xnor UO_1385 (O_1385,N_47668,N_48986);
xor UO_1386 (O_1386,N_48332,N_45016);
xnor UO_1387 (O_1387,N_46600,N_45164);
or UO_1388 (O_1388,N_48957,N_47808);
nand UO_1389 (O_1389,N_49044,N_48232);
or UO_1390 (O_1390,N_48229,N_47483);
nand UO_1391 (O_1391,N_45316,N_49630);
nor UO_1392 (O_1392,N_49500,N_45730);
nor UO_1393 (O_1393,N_46073,N_45198);
nand UO_1394 (O_1394,N_45960,N_46325);
xnor UO_1395 (O_1395,N_46031,N_46086);
and UO_1396 (O_1396,N_47318,N_49563);
nand UO_1397 (O_1397,N_46289,N_45532);
or UO_1398 (O_1398,N_46047,N_47121);
nor UO_1399 (O_1399,N_45794,N_46967);
and UO_1400 (O_1400,N_45201,N_48539);
xor UO_1401 (O_1401,N_48031,N_49291);
or UO_1402 (O_1402,N_48269,N_48139);
or UO_1403 (O_1403,N_47923,N_45930);
nor UO_1404 (O_1404,N_46561,N_46483);
or UO_1405 (O_1405,N_47721,N_45277);
xnor UO_1406 (O_1406,N_47692,N_49637);
xnor UO_1407 (O_1407,N_46711,N_49913);
nand UO_1408 (O_1408,N_48371,N_45203);
and UO_1409 (O_1409,N_47370,N_45502);
nor UO_1410 (O_1410,N_48718,N_47983);
or UO_1411 (O_1411,N_45809,N_45262);
nor UO_1412 (O_1412,N_47732,N_45740);
xor UO_1413 (O_1413,N_48862,N_45422);
xor UO_1414 (O_1414,N_47896,N_45793);
and UO_1415 (O_1415,N_47357,N_45561);
or UO_1416 (O_1416,N_46217,N_45628);
xnor UO_1417 (O_1417,N_47072,N_45400);
xor UO_1418 (O_1418,N_47670,N_48011);
nor UO_1419 (O_1419,N_48352,N_49981);
or UO_1420 (O_1420,N_48925,N_48306);
nor UO_1421 (O_1421,N_47700,N_48158);
nand UO_1422 (O_1422,N_46768,N_46960);
and UO_1423 (O_1423,N_49248,N_49240);
and UO_1424 (O_1424,N_48898,N_47369);
nor UO_1425 (O_1425,N_47333,N_45554);
nand UO_1426 (O_1426,N_46509,N_49099);
or UO_1427 (O_1427,N_49580,N_47385);
or UO_1428 (O_1428,N_45343,N_47237);
xor UO_1429 (O_1429,N_48244,N_45336);
and UO_1430 (O_1430,N_49020,N_48742);
nor UO_1431 (O_1431,N_48173,N_49376);
or UO_1432 (O_1432,N_47328,N_48163);
xor UO_1433 (O_1433,N_49719,N_48312);
or UO_1434 (O_1434,N_45119,N_47777);
nor UO_1435 (O_1435,N_45265,N_45315);
and UO_1436 (O_1436,N_48213,N_46089);
nor UO_1437 (O_1437,N_48340,N_49084);
and UO_1438 (O_1438,N_47191,N_45115);
or UO_1439 (O_1439,N_45726,N_49969);
xor UO_1440 (O_1440,N_49541,N_48431);
nor UO_1441 (O_1441,N_48636,N_49075);
or UO_1442 (O_1442,N_48484,N_47993);
and UO_1443 (O_1443,N_47005,N_48459);
nor UO_1444 (O_1444,N_47353,N_47321);
or UO_1445 (O_1445,N_45114,N_48777);
or UO_1446 (O_1446,N_48097,N_46236);
nor UO_1447 (O_1447,N_46548,N_45086);
nor UO_1448 (O_1448,N_49035,N_47599);
nand UO_1449 (O_1449,N_47801,N_46049);
and UO_1450 (O_1450,N_49691,N_46977);
nand UO_1451 (O_1451,N_48643,N_49907);
or UO_1452 (O_1452,N_46183,N_45808);
and UO_1453 (O_1453,N_46997,N_49006);
xnor UO_1454 (O_1454,N_49701,N_48043);
xnor UO_1455 (O_1455,N_49807,N_45252);
xnor UO_1456 (O_1456,N_47325,N_49814);
and UO_1457 (O_1457,N_46361,N_47752);
nand UO_1458 (O_1458,N_49984,N_49768);
nor UO_1459 (O_1459,N_45581,N_49215);
or UO_1460 (O_1460,N_46982,N_45745);
nand UO_1461 (O_1461,N_46655,N_47694);
nor UO_1462 (O_1462,N_45058,N_49329);
nand UO_1463 (O_1463,N_45818,N_45458);
and UO_1464 (O_1464,N_45483,N_45167);
or UO_1465 (O_1465,N_49714,N_47245);
nor UO_1466 (O_1466,N_47474,N_46506);
nor UO_1467 (O_1467,N_45868,N_49875);
or UO_1468 (O_1468,N_48628,N_47844);
nand UO_1469 (O_1469,N_47252,N_47789);
nand UO_1470 (O_1470,N_46410,N_48118);
or UO_1471 (O_1471,N_49168,N_45301);
nand UO_1472 (O_1472,N_48974,N_45763);
or UO_1473 (O_1473,N_49496,N_47244);
nor UO_1474 (O_1474,N_48486,N_49827);
nand UO_1475 (O_1475,N_48377,N_46763);
nand UO_1476 (O_1476,N_48727,N_46792);
nand UO_1477 (O_1477,N_47345,N_47371);
and UO_1478 (O_1478,N_46337,N_47798);
xnor UO_1479 (O_1479,N_48290,N_46907);
nand UO_1480 (O_1480,N_48175,N_49285);
nor UO_1481 (O_1481,N_45779,N_47868);
nor UO_1482 (O_1482,N_46338,N_47360);
nor UO_1483 (O_1483,N_47388,N_48284);
or UO_1484 (O_1484,N_47452,N_48978);
nand UO_1485 (O_1485,N_48679,N_45911);
nand UO_1486 (O_1486,N_48894,N_48042);
and UO_1487 (O_1487,N_47242,N_47891);
or UO_1488 (O_1488,N_46904,N_47189);
nor UO_1489 (O_1489,N_49102,N_46263);
or UO_1490 (O_1490,N_47182,N_49104);
nand UO_1491 (O_1491,N_48577,N_46794);
nand UO_1492 (O_1492,N_48778,N_46959);
or UO_1493 (O_1493,N_46539,N_45530);
nand UO_1494 (O_1494,N_46091,N_46260);
and UO_1495 (O_1495,N_46754,N_48078);
or UO_1496 (O_1496,N_49513,N_49948);
xnor UO_1497 (O_1497,N_48655,N_46288);
xor UO_1498 (O_1498,N_49757,N_46879);
nor UO_1499 (O_1499,N_46750,N_45813);
and UO_1500 (O_1500,N_45374,N_46188);
and UO_1501 (O_1501,N_45732,N_47977);
or UO_1502 (O_1502,N_49919,N_45180);
xor UO_1503 (O_1503,N_45083,N_49354);
xor UO_1504 (O_1504,N_49390,N_48650);
nor UO_1505 (O_1505,N_48822,N_49670);
or UO_1506 (O_1506,N_49976,N_47931);
xor UO_1507 (O_1507,N_46808,N_47343);
nor UO_1508 (O_1508,N_46700,N_46326);
nand UO_1509 (O_1509,N_47504,N_49065);
and UO_1510 (O_1510,N_49936,N_48851);
nand UO_1511 (O_1511,N_48485,N_48153);
or UO_1512 (O_1512,N_49467,N_48802);
nor UO_1513 (O_1513,N_48653,N_45408);
and UO_1514 (O_1514,N_49328,N_45402);
xor UO_1515 (O_1515,N_48611,N_45550);
and UO_1516 (O_1516,N_45055,N_45864);
nand UO_1517 (O_1517,N_49918,N_49445);
nor UO_1518 (O_1518,N_45067,N_46880);
or UO_1519 (O_1519,N_45736,N_45438);
nor UO_1520 (O_1520,N_46161,N_49143);
or UO_1521 (O_1521,N_47435,N_46682);
xor UO_1522 (O_1522,N_47114,N_48247);
nor UO_1523 (O_1523,N_49487,N_49231);
or UO_1524 (O_1524,N_47722,N_48824);
nor UO_1525 (O_1525,N_49963,N_48861);
nand UO_1526 (O_1526,N_48700,N_47974);
and UO_1527 (O_1527,N_46437,N_49873);
nand UO_1528 (O_1528,N_46791,N_48341);
and UO_1529 (O_1529,N_49901,N_45558);
xor UO_1530 (O_1530,N_45420,N_47512);
xnor UO_1531 (O_1531,N_48167,N_47818);
and UO_1532 (O_1532,N_45112,N_47320);
nor UO_1533 (O_1533,N_46133,N_49133);
xor UO_1534 (O_1534,N_45583,N_47220);
nand UO_1535 (O_1535,N_47884,N_49694);
nor UO_1536 (O_1536,N_45815,N_45972);
and UO_1537 (O_1537,N_47661,N_47034);
nor UO_1538 (O_1538,N_47706,N_47927);
xor UO_1539 (O_1539,N_45068,N_49556);
or UO_1540 (O_1540,N_45237,N_45832);
nand UO_1541 (O_1541,N_48473,N_47555);
nor UO_1542 (O_1542,N_47664,N_46581);
nand UO_1543 (O_1543,N_45889,N_48432);
and UO_1544 (O_1544,N_48772,N_49715);
nand UO_1545 (O_1545,N_49780,N_46272);
xor UO_1546 (O_1546,N_45465,N_49155);
nor UO_1547 (O_1547,N_49222,N_47516);
nand UO_1548 (O_1548,N_48644,N_47876);
nor UO_1549 (O_1549,N_45121,N_45405);
nand UO_1550 (O_1550,N_49517,N_47037);
nor UO_1551 (O_1551,N_45444,N_46401);
xor UO_1552 (O_1552,N_46536,N_48584);
or UO_1553 (O_1553,N_46770,N_48408);
nor UO_1554 (O_1554,N_48482,N_49283);
and UO_1555 (O_1555,N_46606,N_49331);
xnor UO_1556 (O_1556,N_47064,N_47807);
nor UO_1557 (O_1557,N_48355,N_46796);
or UO_1558 (O_1558,N_48885,N_46071);
xnor UO_1559 (O_1559,N_45287,N_45235);
or UO_1560 (O_1560,N_49126,N_49842);
xnor UO_1561 (O_1561,N_48807,N_46143);
nor UO_1562 (O_1562,N_46182,N_48603);
nand UO_1563 (O_1563,N_49462,N_45914);
or UO_1564 (O_1564,N_47079,N_49577);
xor UO_1565 (O_1565,N_49837,N_48712);
xor UO_1566 (O_1566,N_46465,N_48900);
nand UO_1567 (O_1567,N_46135,N_48519);
nand UO_1568 (O_1568,N_48596,N_48977);
and UO_1569 (O_1569,N_46801,N_49841);
or UO_1570 (O_1570,N_48923,N_45475);
or UO_1571 (O_1571,N_49891,N_48441);
nor UO_1572 (O_1572,N_46065,N_46319);
nand UO_1573 (O_1573,N_49456,N_48362);
or UO_1574 (O_1574,N_46062,N_46420);
or UO_1575 (O_1575,N_47066,N_46216);
xnor UO_1576 (O_1576,N_45129,N_47561);
and UO_1577 (O_1577,N_46751,N_49052);
xor UO_1578 (O_1578,N_45900,N_47026);
xnor UO_1579 (O_1579,N_45971,N_49375);
nor UO_1580 (O_1580,N_45401,N_45881);
or UO_1581 (O_1581,N_49436,N_49527);
nor UO_1582 (O_1582,N_45133,N_45193);
or UO_1583 (O_1583,N_48733,N_45380);
nor UO_1584 (O_1584,N_47192,N_48301);
nor UO_1585 (O_1585,N_47453,N_45320);
or UO_1586 (O_1586,N_46523,N_47716);
nor UO_1587 (O_1587,N_48754,N_48749);
nand UO_1588 (O_1588,N_49941,N_45209);
nor UO_1589 (O_1589,N_49902,N_49874);
nor UO_1590 (O_1590,N_47551,N_47223);
nand UO_1591 (O_1591,N_45295,N_47137);
nand UO_1592 (O_1592,N_49119,N_49324);
and UO_1593 (O_1593,N_49478,N_46131);
or UO_1594 (O_1594,N_46406,N_46615);
xor UO_1595 (O_1595,N_45661,N_49493);
and UO_1596 (O_1596,N_45339,N_47853);
nand UO_1597 (O_1597,N_49599,N_45143);
or UO_1598 (O_1598,N_45038,N_47918);
nand UO_1599 (O_1599,N_49120,N_46242);
and UO_1600 (O_1600,N_45585,N_46069);
or UO_1601 (O_1601,N_45703,N_48191);
and UO_1602 (O_1602,N_47112,N_49551);
or UO_1603 (O_1603,N_48395,N_48461);
or UO_1604 (O_1604,N_45390,N_47095);
xnor UO_1605 (O_1605,N_48568,N_49730);
and UO_1606 (O_1606,N_47040,N_48963);
nor UO_1607 (O_1607,N_49633,N_48481);
nor UO_1608 (O_1608,N_45551,N_45299);
and UO_1609 (O_1609,N_48902,N_45518);
nand UO_1610 (O_1610,N_45019,N_48521);
xnor UO_1611 (O_1611,N_46938,N_49165);
xor UO_1612 (O_1612,N_46696,N_45278);
nor UO_1613 (O_1613,N_49819,N_45117);
nand UO_1614 (O_1614,N_49544,N_49524);
nand UO_1615 (O_1615,N_49537,N_46577);
nand UO_1616 (O_1616,N_48960,N_49785);
xor UO_1617 (O_1617,N_49914,N_48238);
and UO_1618 (O_1618,N_45292,N_49618);
nand UO_1619 (O_1619,N_45562,N_48157);
xnor UO_1620 (O_1620,N_46176,N_49338);
and UO_1621 (O_1621,N_49332,N_47958);
xnor UO_1622 (O_1622,N_46814,N_46428);
nor UO_1623 (O_1623,N_46022,N_46043);
nor UO_1624 (O_1624,N_46881,N_48211);
and UO_1625 (O_1625,N_48942,N_46389);
nand UO_1626 (O_1626,N_47289,N_47063);
or UO_1627 (O_1627,N_49463,N_45126);
and UO_1628 (O_1628,N_48710,N_47922);
or UO_1629 (O_1629,N_45667,N_47762);
xor UO_1630 (O_1630,N_46747,N_48160);
nor UO_1631 (O_1631,N_46589,N_49027);
xor UO_1632 (O_1632,N_45358,N_45923);
or UO_1633 (O_1633,N_48478,N_48391);
nand UO_1634 (O_1634,N_49538,N_46621);
or UO_1635 (O_1635,N_49965,N_49934);
and UO_1636 (O_1636,N_47107,N_47285);
nand UO_1637 (O_1637,N_45601,N_45138);
nor UO_1638 (O_1638,N_48582,N_49484);
nand UO_1639 (O_1639,N_46214,N_47870);
nor UO_1640 (O_1640,N_48400,N_47856);
and UO_1641 (O_1641,N_46902,N_45101);
xor UO_1642 (O_1642,N_49439,N_47542);
nor UO_1643 (O_1643,N_47615,N_46253);
and UO_1644 (O_1644,N_48245,N_48171);
or UO_1645 (O_1645,N_47655,N_45426);
xnor UO_1646 (O_1646,N_46474,N_49824);
nand UO_1647 (O_1647,N_46744,N_48815);
nor UO_1648 (O_1648,N_48922,N_45624);
and UO_1649 (O_1649,N_46493,N_48551);
nand UO_1650 (O_1650,N_45415,N_49179);
nand UO_1651 (O_1651,N_46986,N_49301);
nand UO_1652 (O_1652,N_49274,N_49363);
and UO_1653 (O_1653,N_47038,N_46515);
and UO_1654 (O_1654,N_46117,N_45093);
xor UO_1655 (O_1655,N_47397,N_46740);
nor UO_1656 (O_1656,N_47058,N_49868);
xnor UO_1657 (O_1657,N_48504,N_46127);
or UO_1658 (O_1658,N_46838,N_45169);
xnor UO_1659 (O_1659,N_45688,N_46893);
or UO_1660 (O_1660,N_48422,N_49916);
nor UO_1661 (O_1661,N_49480,N_46458);
xnor UO_1662 (O_1662,N_45893,N_47041);
xor UO_1663 (O_1663,N_48814,N_47093);
or UO_1664 (O_1664,N_45350,N_48122);
nand UO_1665 (O_1665,N_45250,N_47724);
xnor UO_1666 (O_1666,N_47087,N_49134);
nand UO_1667 (O_1667,N_45606,N_48955);
nor UO_1668 (O_1668,N_47390,N_45926);
xor UO_1669 (O_1669,N_46205,N_45737);
or UO_1670 (O_1670,N_48587,N_47634);
xor UO_1671 (O_1671,N_48416,N_49361);
or UO_1672 (O_1672,N_49856,N_49453);
xnor UO_1673 (O_1673,N_46265,N_47940);
and UO_1674 (O_1674,N_48602,N_48993);
or UO_1675 (O_1675,N_49425,N_48995);
nand UO_1676 (O_1676,N_46585,N_49628);
and UO_1677 (O_1677,N_48082,N_46380);
or UO_1678 (O_1678,N_45722,N_48563);
nand UO_1679 (O_1679,N_47932,N_46202);
nand UO_1680 (O_1680,N_45132,N_46878);
xor UO_1681 (O_1681,N_45650,N_46936);
xor UO_1682 (O_1682,N_45625,N_49461);
xor UO_1683 (O_1683,N_49090,N_46910);
nor UO_1684 (O_1684,N_48188,N_48575);
and UO_1685 (O_1685,N_49616,N_46328);
xor UO_1686 (O_1686,N_45266,N_49569);
nor UO_1687 (O_1687,N_46709,N_46973);
and UO_1688 (O_1688,N_46983,N_45941);
xor UO_1689 (O_1689,N_47224,N_46180);
nand UO_1690 (O_1690,N_46291,N_48623);
or UO_1691 (O_1691,N_48895,N_47417);
nor UO_1692 (O_1692,N_45796,N_49779);
xnor UO_1693 (O_1693,N_45942,N_46974);
nor UO_1694 (O_1694,N_47233,N_49923);
xor UO_1695 (O_1695,N_49259,N_46046);
or UO_1696 (O_1696,N_49247,N_45241);
nor UO_1697 (O_1697,N_46181,N_45309);
nand UO_1698 (O_1698,N_45701,N_46306);
nand UO_1699 (O_1699,N_48349,N_45253);
nand UO_1700 (O_1700,N_48438,N_45238);
or UO_1701 (O_1701,N_49933,N_45040);
and UO_1702 (O_1702,N_49432,N_46113);
nand UO_1703 (O_1703,N_45375,N_49335);
and UO_1704 (O_1704,N_48138,N_48347);
xor UO_1705 (O_1705,N_45989,N_45871);
nor UO_1706 (O_1706,N_49036,N_46080);
nor UO_1707 (O_1707,N_48773,N_46377);
nand UO_1708 (O_1708,N_47486,N_49585);
or UO_1709 (O_1709,N_46174,N_47129);
nor UO_1710 (O_1710,N_46781,N_46934);
nand UO_1711 (O_1711,N_48820,N_46170);
nand UO_1712 (O_1712,N_49150,N_49505);
and UO_1713 (O_1713,N_49685,N_49296);
nor UO_1714 (O_1714,N_45219,N_49612);
nand UO_1715 (O_1715,N_45771,N_45081);
and UO_1716 (O_1716,N_46139,N_46664);
or UO_1717 (O_1717,N_49937,N_47633);
xor UO_1718 (O_1718,N_46811,N_47648);
nor UO_1719 (O_1719,N_49117,N_48591);
nor UO_1720 (O_1720,N_47566,N_49197);
or UO_1721 (O_1721,N_47225,N_47160);
xor UO_1722 (O_1722,N_49110,N_47957);
xor UO_1723 (O_1723,N_47250,N_47908);
and UO_1724 (O_1724,N_49812,N_46100);
and UO_1725 (O_1725,N_48905,N_48715);
xnor UO_1726 (O_1726,N_46928,N_48855);
and UO_1727 (O_1727,N_47293,N_48051);
nand UO_1728 (O_1728,N_45152,N_49433);
and UO_1729 (O_1729,N_45310,N_48661);
or UO_1730 (O_1730,N_46271,N_48436);
nor UO_1731 (O_1731,N_45797,N_45894);
and UO_1732 (O_1732,N_45447,N_46485);
and UO_1733 (O_1733,N_48964,N_48780);
or UO_1734 (O_1734,N_45912,N_49041);
nand UO_1735 (O_1735,N_45754,N_47292);
nand UO_1736 (O_1736,N_48982,N_47198);
or UO_1737 (O_1737,N_47315,N_48363);
xnor UO_1738 (O_1738,N_49881,N_48579);
and UO_1739 (O_1739,N_45932,N_45381);
nor UO_1740 (O_1740,N_49351,N_45943);
nor UO_1741 (O_1741,N_48788,N_47799);
and UO_1742 (O_1742,N_46832,N_49669);
xor UO_1743 (O_1743,N_49149,N_45602);
xor UO_1744 (O_1744,N_48267,N_49870);
xor UO_1745 (O_1745,N_46837,N_45686);
nand UO_1746 (O_1746,N_46261,N_46702);
or UO_1747 (O_1747,N_46027,N_48135);
nor UO_1748 (O_1748,N_48443,N_49858);
xnor UO_1749 (O_1749,N_47717,N_47532);
or UO_1750 (O_1750,N_48622,N_49766);
nand UO_1751 (O_1751,N_47681,N_48593);
and UO_1752 (O_1752,N_47905,N_46035);
nor UO_1753 (O_1753,N_47850,N_48435);
or UO_1754 (O_1754,N_46209,N_45897);
xnor UO_1755 (O_1755,N_49753,N_47012);
xor UO_1756 (O_1756,N_48299,N_47792);
nor UO_1757 (O_1757,N_49419,N_46296);
or UO_1758 (O_1758,N_45500,N_47470);
or UO_1759 (O_1759,N_47920,N_49688);
or UO_1760 (O_1760,N_48212,N_48493);
nand UO_1761 (O_1761,N_45867,N_49092);
and UO_1762 (O_1762,N_49800,N_48044);
and UO_1763 (O_1763,N_48614,N_49634);
or UO_1764 (O_1764,N_48128,N_47825);
nand UO_1765 (O_1765,N_45610,N_49083);
nand UO_1766 (O_1766,N_47540,N_47770);
xor UO_1767 (O_1767,N_48219,N_45948);
xnor UO_1768 (O_1768,N_45108,N_45054);
nand UO_1769 (O_1769,N_47955,N_45992);
and UO_1770 (O_1770,N_46884,N_46891);
nor UO_1771 (O_1771,N_49533,N_48458);
nand UO_1772 (O_1772,N_45825,N_48576);
or UO_1773 (O_1773,N_48737,N_45014);
or UO_1774 (O_1774,N_49822,N_47356);
and UO_1775 (O_1775,N_47821,N_46882);
or UO_1776 (O_1776,N_49805,N_47307);
nor UO_1777 (O_1777,N_47431,N_49368);
nand UO_1778 (O_1778,N_48990,N_47077);
xnor UO_1779 (O_1779,N_45352,N_48469);
nor UO_1780 (O_1780,N_48233,N_46948);
xor UO_1781 (O_1781,N_47030,N_49319);
or UO_1782 (O_1782,N_48398,N_49829);
or UO_1783 (O_1783,N_47166,N_48561);
xnor UO_1784 (O_1784,N_48743,N_46014);
or UO_1785 (O_1785,N_45700,N_46457);
xnor UO_1786 (O_1786,N_47947,N_48418);
xnor UO_1787 (O_1787,N_46211,N_45291);
xnor UO_1788 (O_1788,N_49060,N_47793);
and UO_1789 (O_1789,N_47071,N_49125);
or UO_1790 (O_1790,N_49355,N_49122);
nor UO_1791 (O_1791,N_45725,N_45576);
xor UO_1792 (O_1792,N_48236,N_46932);
nor UO_1793 (O_1793,N_48748,N_49883);
xnor UO_1794 (O_1794,N_49472,N_46381);
nand UO_1795 (O_1795,N_46036,N_45151);
xnor UO_1796 (O_1796,N_49252,N_48159);
nor UO_1797 (O_1797,N_47382,N_47685);
nand UO_1798 (O_1798,N_48388,N_45062);
nor UO_1799 (O_1799,N_49996,N_46285);
or UO_1800 (O_1800,N_47048,N_47890);
nand UO_1801 (O_1801,N_47912,N_49745);
nor UO_1802 (O_1802,N_49543,N_46584);
xnor UO_1803 (O_1803,N_48305,N_49720);
and UO_1804 (O_1804,N_47442,N_48904);
nand UO_1805 (O_1805,N_49350,N_48954);
and UO_1806 (O_1806,N_45261,N_49514);
or UO_1807 (O_1807,N_49370,N_47652);
nor UO_1808 (O_1808,N_45183,N_47101);
or UO_1809 (O_1809,N_49210,N_48378);
and UO_1810 (O_1810,N_46151,N_47028);
nor UO_1811 (O_1811,N_49365,N_47804);
nand UO_1812 (O_1812,N_49220,N_48784);
nand UO_1813 (O_1813,N_46154,N_46550);
and UO_1814 (O_1814,N_46516,N_48513);
nand UO_1815 (O_1815,N_47730,N_47362);
nand UO_1816 (O_1816,N_47021,N_49648);
xor UO_1817 (O_1817,N_46396,N_48178);
xor UO_1818 (O_1818,N_47803,N_48617);
or UO_1819 (O_1819,N_46322,N_45656);
and UO_1820 (O_1820,N_46061,N_48066);
nor UO_1821 (O_1821,N_46443,N_48871);
or UO_1822 (O_1822,N_49323,N_45257);
xor UO_1823 (O_1823,N_49391,N_45191);
or UO_1824 (O_1824,N_47951,N_48145);
and UO_1825 (O_1825,N_49808,N_46998);
nand UO_1826 (O_1826,N_49001,N_49640);
and UO_1827 (O_1827,N_48283,N_45443);
or UO_1828 (O_1828,N_46553,N_49395);
and UO_1829 (O_1829,N_45705,N_46186);
or UO_1830 (O_1830,N_49409,N_45590);
nand UO_1831 (O_1831,N_46254,N_49802);
nand UO_1832 (O_1832,N_49986,N_48049);
nand UO_1833 (O_1833,N_46767,N_48839);
nor UO_1834 (O_1834,N_48369,N_45128);
nand UO_1835 (O_1835,N_47769,N_49294);
nor UO_1836 (O_1836,N_49733,N_47501);
nand UO_1837 (O_1837,N_45260,N_48115);
nand UO_1838 (O_1838,N_48320,N_46195);
xor UO_1839 (O_1839,N_49702,N_45322);
xnor UO_1840 (O_1840,N_48932,N_49177);
nand UO_1841 (O_1841,N_48757,N_45829);
and UO_1842 (O_1842,N_47854,N_49251);
xor UO_1843 (O_1843,N_47558,N_48868);
or UO_1844 (O_1844,N_48380,N_48819);
nor UO_1845 (O_1845,N_48266,N_48419);
xnor UO_1846 (O_1846,N_46083,N_49269);
or UO_1847 (O_1847,N_48218,N_45777);
nor UO_1848 (O_1848,N_48943,N_46355);
or UO_1849 (O_1849,N_48072,N_49298);
and UO_1850 (O_1850,N_49940,N_48581);
or UO_1851 (O_1851,N_49929,N_48483);
nor UO_1852 (O_1852,N_47502,N_45096);
or UO_1853 (O_1853,N_46797,N_46512);
and UO_1854 (O_1854,N_45630,N_49731);
xor UO_1855 (O_1855,N_48263,N_49055);
xor UO_1856 (O_1856,N_49010,N_46044);
xor UO_1857 (O_1857,N_47511,N_47788);
or UO_1858 (O_1858,N_45784,N_45173);
and UO_1859 (O_1859,N_48675,N_45327);
xor UO_1860 (O_1860,N_45798,N_47961);
xor UO_1861 (O_1861,N_47586,N_47697);
or UO_1862 (O_1862,N_48496,N_48686);
and UO_1863 (O_1863,N_45388,N_45709);
xnor UO_1864 (O_1864,N_49689,N_47494);
and UO_1865 (O_1865,N_49964,N_49782);
or UO_1866 (O_1866,N_49890,N_49843);
and UO_1867 (O_1867,N_47479,N_48642);
and UO_1868 (O_1868,N_49166,N_46824);
xor UO_1869 (O_1869,N_46397,N_47695);
xor UO_1870 (O_1870,N_48201,N_49518);
xnor UO_1871 (O_1871,N_49236,N_45334);
nand UO_1872 (O_1872,N_45689,N_47986);
nand UO_1873 (O_1873,N_45378,N_48865);
and UO_1874 (O_1874,N_46393,N_45127);
xnor UO_1875 (O_1875,N_48601,N_47885);
nor UO_1876 (O_1876,N_47608,N_48548);
xnor UO_1877 (O_1877,N_49576,N_47980);
nor UO_1878 (O_1878,N_48699,N_47110);
xnor UO_1879 (O_1879,N_45990,N_45843);
or UO_1880 (O_1880,N_46943,N_45258);
nand UO_1881 (O_1881,N_46469,N_47898);
nor UO_1882 (O_1882,N_47180,N_45440);
xor UO_1883 (O_1883,N_49565,N_46184);
nand UO_1884 (O_1884,N_45594,N_48058);
nor UO_1885 (O_1885,N_45921,N_47341);
or UO_1886 (O_1886,N_49011,N_49427);
nor UO_1887 (O_1887,N_47413,N_45713);
nor UO_1888 (O_1888,N_46439,N_46915);
nor UO_1889 (O_1889,N_47457,N_46051);
xor UO_1890 (O_1890,N_46806,N_48302);
nor UO_1891 (O_1891,N_49033,N_45342);
nor UO_1892 (O_1892,N_47264,N_47533);
xnor UO_1893 (O_1893,N_46591,N_49148);
nor UO_1894 (O_1894,N_48595,N_46579);
xnor UO_1895 (O_1895,N_47939,N_49943);
xnor UO_1896 (O_1896,N_46517,N_48275);
xnor UO_1897 (O_1897,N_45747,N_49516);
xnor UO_1898 (O_1898,N_46999,N_46501);
nand UO_1899 (O_1899,N_46147,N_45750);
xnor UO_1900 (O_1900,N_48131,N_46347);
nand UO_1901 (O_1901,N_49882,N_47306);
nand UO_1902 (O_1902,N_49140,N_46482);
or UO_1903 (O_1903,N_49348,N_48912);
xor UO_1904 (O_1904,N_46400,N_45827);
or UO_1905 (O_1905,N_48196,N_46310);
xnor UO_1906 (O_1906,N_48630,N_45735);
nand UO_1907 (O_1907,N_45862,N_47597);
or UO_1908 (O_1908,N_45050,N_45510);
nand UO_1909 (O_1909,N_49087,N_45986);
xnor UO_1910 (O_1910,N_48706,N_45172);
nor UO_1911 (O_1911,N_45331,N_45533);
and UO_1912 (O_1912,N_48853,N_49917);
or UO_1913 (O_1913,N_48383,N_48901);
or UO_1914 (O_1914,N_49310,N_48356);
nor UO_1915 (O_1915,N_45866,N_46006);
nor UO_1916 (O_1916,N_45823,N_45674);
or UO_1917 (O_1917,N_47723,N_46295);
or UO_1918 (O_1918,N_46008,N_47739);
xor UO_1919 (O_1919,N_49159,N_47392);
and UO_1920 (O_1920,N_46835,N_45470);
nor UO_1921 (O_1921,N_49665,N_49830);
or UO_1922 (O_1922,N_47310,N_47448);
xnor UO_1923 (O_1923,N_49741,N_47651);
xnor UO_1924 (O_1924,N_46088,N_47541);
xnor UO_1925 (O_1925,N_47975,N_45046);
and UO_1926 (O_1926,N_46368,N_45228);
or UO_1927 (O_1927,N_49180,N_48405);
nor UO_1928 (O_1928,N_48631,N_48966);
or UO_1929 (O_1929,N_48444,N_49153);
xor UO_1930 (O_1930,N_49204,N_45484);
nor UO_1931 (O_1931,N_46538,N_48004);
xor UO_1932 (O_1932,N_49262,N_49397);
xnor UO_1933 (O_1933,N_46419,N_49367);
nor UO_1934 (O_1934,N_49364,N_48142);
and UO_1935 (O_1935,N_45865,N_49987);
and UO_1936 (O_1936,N_45728,N_45543);
nor UO_1937 (O_1937,N_49024,N_45614);
or UO_1938 (O_1938,N_48526,N_46541);
xnor UO_1939 (O_1939,N_45837,N_46745);
nor UO_1940 (O_1940,N_45546,N_47865);
xor UO_1941 (O_1941,N_49879,N_46597);
nand UO_1942 (O_1942,N_48528,N_46676);
nor UO_1943 (O_1943,N_48468,N_45412);
xnor UO_1944 (O_1944,N_47572,N_48342);
nor UO_1945 (O_1945,N_46634,N_49229);
nand UO_1946 (O_1946,N_47305,N_49511);
or UO_1947 (O_1947,N_47926,N_48270);
xor UO_1948 (O_1948,N_45094,N_48437);
nor UO_1949 (O_1949,N_47968,N_46560);
and UO_1950 (O_1950,N_47592,N_49892);
nor UO_1951 (O_1951,N_45569,N_49254);
and UO_1952 (O_1952,N_48662,N_48557);
and UO_1953 (O_1953,N_47449,N_46414);
nand UO_1954 (O_1954,N_48243,N_45987);
nand UO_1955 (O_1955,N_49089,N_46120);
xor UO_1956 (O_1956,N_45507,N_47139);
and UO_1957 (O_1957,N_49617,N_45820);
or UO_1958 (O_1958,N_49246,N_48530);
or UO_1959 (O_1959,N_48854,N_45995);
or UO_1960 (O_1960,N_49959,N_48050);
xor UO_1961 (O_1961,N_49012,N_49721);
xnor UO_1962 (O_1962,N_46773,N_47290);
nor UO_1963 (O_1963,N_45723,N_48759);
nor UO_1964 (O_1964,N_46496,N_45231);
or UO_1965 (O_1965,N_46508,N_46276);
and UO_1966 (O_1966,N_45118,N_49207);
or UO_1967 (O_1967,N_45206,N_49584);
xnor UO_1968 (O_1968,N_49752,N_46076);
xor UO_1969 (O_1969,N_49417,N_45289);
xor UO_1970 (O_1970,N_45270,N_45964);
nor UO_1971 (O_1971,N_48945,N_46728);
and UO_1972 (O_1972,N_45344,N_47387);
nand UO_1973 (O_1973,N_48148,N_46067);
and UO_1974 (O_1974,N_49865,N_49046);
and UO_1975 (O_1975,N_45887,N_45962);
xnor UO_1976 (O_1976,N_47521,N_46669);
nor UO_1977 (O_1977,N_45012,N_46786);
nor UO_1978 (O_1978,N_45148,N_47496);
nand UO_1979 (O_1979,N_49839,N_45937);
xor UO_1980 (O_1980,N_46148,N_45283);
xnor UO_1981 (O_1981,N_47674,N_49271);
and UO_1982 (O_1982,N_46961,N_45577);
xor UO_1983 (O_1983,N_45662,N_45916);
nand UO_1984 (O_1984,N_47399,N_49061);
xnor UO_1985 (O_1985,N_47200,N_46551);
and UO_1986 (O_1986,N_46003,N_49405);
nor UO_1987 (O_1987,N_45790,N_47587);
nor UO_1988 (O_1988,N_45479,N_48354);
xor UO_1989 (O_1989,N_49305,N_45514);
nor UO_1990 (O_1990,N_49512,N_48372);
and UO_1991 (O_1991,N_49734,N_49579);
nand UO_1992 (O_1992,N_48935,N_45294);
nand UO_1993 (O_1993,N_49371,N_49034);
and UO_1994 (O_1994,N_46344,N_47164);
nor UO_1995 (O_1995,N_47365,N_46729);
nand UO_1996 (O_1996,N_48680,N_49420);
and UO_1997 (O_1997,N_48830,N_45345);
xnor UO_1998 (O_1998,N_46958,N_48812);
or UO_1999 (O_1999,N_49942,N_46828);
and UO_2000 (O_2000,N_48427,N_49454);
and UO_2001 (O_2001,N_46097,N_49690);
nand UO_2002 (O_2002,N_49557,N_48876);
or UO_2003 (O_2003,N_49703,N_47197);
or UO_2004 (O_2004,N_46752,N_48753);
nand UO_2005 (O_2005,N_49751,N_46363);
or UO_2006 (O_2006,N_46820,N_49121);
nor UO_2007 (O_2007,N_47273,N_47984);
xor UO_2008 (O_2008,N_49457,N_45462);
nor UO_2009 (O_2009,N_49589,N_46843);
nand UO_2010 (O_2010,N_48850,N_49038);
xor UO_2011 (O_2011,N_48028,N_45208);
and UO_2012 (O_2012,N_47019,N_49029);
and UO_2013 (O_2013,N_48765,N_47679);
xor UO_2014 (O_2014,N_45727,N_49562);
or UO_2015 (O_2015,N_46656,N_47490);
and UO_2016 (O_2016,N_47852,N_49465);
xor UO_2017 (O_2017,N_47081,N_47753);
nor UO_2018 (O_2018,N_47613,N_49211);
or UO_2019 (O_2019,N_47656,N_49970);
or UO_2020 (O_2020,N_49161,N_45216);
xor UO_2021 (O_2021,N_48828,N_47014);
xnor UO_2022 (O_2022,N_47569,N_47049);
nor UO_2023 (O_2023,N_46755,N_48915);
nor UO_2024 (O_2024,N_46557,N_48891);
and UO_2025 (O_2025,N_49224,N_47895);
and UO_2026 (O_2026,N_49476,N_46787);
or UO_2027 (O_2027,N_46829,N_46037);
nor UO_2028 (O_2028,N_49828,N_46152);
and UO_2029 (O_2029,N_46461,N_46815);
and UO_2030 (O_2030,N_46475,N_49877);
nor UO_2031 (O_2031,N_47229,N_48619);
xor UO_2032 (O_2032,N_47097,N_49132);
or UO_2033 (O_2033,N_49638,N_48776);
nor UO_2034 (O_2034,N_47759,N_48375);
nand UO_2035 (O_2035,N_46617,N_46052);
and UO_2036 (O_2036,N_47556,N_46547);
nand UO_2037 (O_2037,N_45084,N_47404);
nor UO_2038 (O_2038,N_49171,N_48357);
and UO_2039 (O_2039,N_49699,N_46918);
xnor UO_2040 (O_2040,N_46267,N_46996);
or UO_2041 (O_2041,N_48063,N_45089);
or UO_2042 (O_2042,N_46497,N_47985);
xnor UO_2043 (O_2043,N_48343,N_49085);
or UO_2044 (O_2044,N_48012,N_45319);
nor UO_2045 (O_2045,N_46221,N_49404);
and UO_2046 (O_2046,N_49474,N_46460);
nand UO_2047 (O_2047,N_46809,N_45927);
or UO_2048 (O_2048,N_48626,N_48783);
nand UO_2049 (O_2049,N_47738,N_46418);
xor UO_2050 (O_2050,N_46817,N_47326);
or UO_2051 (O_2051,N_45538,N_46921);
xor UO_2052 (O_2052,N_49023,N_46128);
or UO_2053 (O_2053,N_47120,N_45704);
or UO_2054 (O_2054,N_48687,N_48088);
and UO_2055 (O_2055,N_47108,N_49997);
nand UO_2056 (O_2056,N_48552,N_46436);
nor UO_2057 (O_2057,N_49656,N_47004);
xnor UO_2058 (O_2058,N_49105,N_48309);
nor UO_2059 (O_2059,N_48334,N_45523);
and UO_2060 (O_2060,N_48972,N_48367);
nor UO_2061 (O_2061,N_47786,N_46946);
nor UO_2062 (O_2062,N_46372,N_48708);
xnor UO_2063 (O_2063,N_48946,N_45760);
nor UO_2064 (O_2064,N_47023,N_49973);
nand UO_2065 (O_2065,N_45406,N_46404);
and UO_2066 (O_2066,N_46748,N_45332);
or UO_2067 (O_2067,N_46383,N_46499);
or UO_2068 (O_2068,N_47280,N_48091);
xor UO_2069 (O_2069,N_47953,N_48182);
nand UO_2070 (O_2070,N_46431,N_47863);
and UO_2071 (O_2071,N_47420,N_49353);
nor UO_2072 (O_2072,N_48442,N_49894);
or UO_2073 (O_2073,N_46294,N_47534);
xnor UO_2074 (O_2074,N_45477,N_45869);
nor UO_2075 (O_2075,N_49209,N_48606);
or UO_2076 (O_2076,N_47451,N_45873);
or UO_2077 (O_2077,N_46937,N_47600);
or UO_2078 (O_2078,N_48553,N_45487);
xnor UO_2079 (O_2079,N_49343,N_46640);
nand UO_2080 (O_2080,N_49387,N_49249);
and UO_2081 (O_2081,N_46730,N_46818);
or UO_2082 (O_2082,N_49546,N_48410);
and UO_2083 (O_2083,N_45249,N_47851);
nor UO_2084 (O_2084,N_46165,N_49601);
or UO_2085 (O_2085,N_49264,N_47620);
or UO_2086 (O_2086,N_46359,N_49799);
xnor UO_2087 (O_2087,N_45248,N_47348);
nor UO_2088 (O_2088,N_45595,N_46413);
nor UO_2089 (O_2089,N_46290,N_47782);
nand UO_2090 (O_2090,N_46925,N_49466);
nand UO_2091 (O_2091,N_49760,N_48547);
and UO_2092 (O_2092,N_49777,N_46920);
xor UO_2093 (O_2093,N_46335,N_48140);
and UO_2094 (O_2094,N_46264,N_46864);
or UO_2095 (O_2095,N_46287,N_49762);
and UO_2096 (O_2096,N_48200,N_46690);
and UO_2097 (O_2097,N_47085,N_46099);
xor UO_2098 (O_2098,N_46845,N_49952);
nand UO_2099 (O_2099,N_46362,N_48524);
and UO_2100 (O_2100,N_49267,N_46464);
xnor UO_2101 (O_2101,N_46187,N_48813);
xnor UO_2102 (O_2102,N_49434,N_46494);
and UO_2103 (O_2103,N_46555,N_47426);
and UO_2104 (O_2104,N_45032,N_47702);
and UO_2105 (O_2105,N_48214,N_48723);
nor UO_2106 (O_2106,N_49097,N_46053);
nor UO_2107 (O_2107,N_49523,N_49857);
xor UO_2108 (O_2108,N_47271,N_47894);
nand UO_2109 (O_2109,N_45706,N_48976);
xnor UO_2110 (O_2110,N_49118,N_47624);
or UO_2111 (O_2111,N_48597,N_47768);
xor UO_2112 (O_2112,N_48529,N_49935);
and UO_2113 (O_2113,N_46661,N_45060);
nor UO_2114 (O_2114,N_45395,N_47795);
nor UO_2115 (O_2115,N_47601,N_48638);
or UO_2116 (O_2116,N_48346,N_49626);
nor UO_2117 (O_2117,N_45150,N_46424);
or UO_2118 (O_2118,N_47846,N_46498);
nor UO_2119 (O_2119,N_47481,N_45645);
nand UO_2120 (O_2120,N_48656,N_47463);
nor UO_2121 (O_2121,N_46939,N_49130);
xnor UO_2122 (O_2122,N_47364,N_46639);
nand UO_2123 (O_2123,N_49239,N_45330);
nor UO_2124 (O_2124,N_49250,N_45660);
nand UO_2125 (O_2125,N_49396,N_45029);
nand UO_2126 (O_2126,N_47247,N_45902);
xor UO_2127 (O_2127,N_46371,N_46390);
or UO_2128 (O_2128,N_48384,N_45087);
or UO_2129 (O_2129,N_47503,N_46888);
xor UO_2130 (O_2130,N_47973,N_45245);
nor UO_2131 (O_2131,N_47254,N_46178);
nand UO_2132 (O_2132,N_46720,N_48224);
or UO_2133 (O_2133,N_48586,N_45649);
xor UO_2134 (O_2134,N_49833,N_48505);
nand UO_2135 (O_2135,N_47143,N_47790);
and UO_2136 (O_2136,N_45221,N_47904);
nor UO_2137 (O_2137,N_47010,N_48322);
and UO_2138 (O_2138,N_49804,N_48803);
xor UO_2139 (O_2139,N_46001,N_48364);
nand UO_2140 (O_2140,N_49520,N_48714);
or UO_2141 (O_2141,N_45273,N_47015);
xnor UO_2142 (O_2142,N_46972,N_48180);
xor UO_2143 (O_2143,N_46194,N_47787);
xnor UO_2144 (O_2144,N_46189,N_48376);
and UO_2145 (O_2145,N_49988,N_47193);
and UO_2146 (O_2146,N_48860,N_46841);
nor UO_2147 (O_2147,N_45542,N_47629);
nand UO_2148 (O_2148,N_48543,N_47228);
or UO_2149 (O_2149,N_48931,N_48189);
and UO_2150 (O_2150,N_48488,N_49468);
or UO_2151 (O_2151,N_49481,N_49631);
nand UO_2152 (O_2152,N_48569,N_47658);
nand UO_2153 (O_2153,N_45545,N_47924);
xnor UO_2154 (O_2154,N_46225,N_46388);
nand UO_2155 (O_2155,N_46618,N_46239);
nor UO_2156 (O_2156,N_48669,N_45955);
nand UO_2157 (O_2157,N_47330,N_49081);
or UO_2158 (O_2158,N_46908,N_46471);
nand UO_2159 (O_2159,N_47235,N_45311);
xor UO_2160 (O_2160,N_47447,N_46636);
and UO_2161 (O_2161,N_49459,N_47150);
or UO_2162 (O_2162,N_46124,N_49662);
xor UO_2163 (O_2163,N_47505,N_45224);
nor UO_2164 (O_2164,N_45664,N_45801);
nand UO_2165 (O_2165,N_45981,N_45433);
or UO_2166 (O_2166,N_48542,N_47238);
and UO_2167 (O_2167,N_46156,N_49539);
nor UO_2168 (O_2168,N_48149,N_46169);
nand UO_2169 (O_2169,N_48821,N_49492);
nor UO_2170 (O_2170,N_49591,N_47459);
and UO_2171 (O_2171,N_46041,N_47604);
xnor UO_2172 (O_2172,N_47358,N_45356);
nand UO_2173 (O_2173,N_48203,N_47800);
nand UO_2174 (O_2174,N_45371,N_45005);
nor UO_2175 (O_2175,N_48170,N_45347);
or UO_2176 (O_2176,N_48704,N_49530);
nand UO_2177 (O_2177,N_45496,N_46118);
xnor UO_2178 (O_2178,N_46697,N_49642);
and UO_2179 (O_2179,N_46544,N_49333);
and UO_2180 (O_2180,N_46222,N_46981);
nor UO_2181 (O_2181,N_49609,N_46142);
xor UO_2182 (O_2182,N_46270,N_49494);
nor UO_2183 (O_2183,N_45076,N_46853);
and UO_2184 (O_2184,N_45274,N_48455);
or UO_2185 (O_2185,N_47520,N_49625);
and UO_2186 (O_2186,N_45619,N_46599);
nor UO_2187 (O_2187,N_47625,N_48847);
or UO_2188 (O_2188,N_47776,N_45110);
nand UO_2189 (O_2189,N_47257,N_47359);
nand UO_2190 (O_2190,N_49088,N_46654);
or UO_2191 (O_2191,N_46226,N_48040);
and UO_2192 (O_2192,N_47226,N_46327);
xor UO_2193 (O_2193,N_45435,N_47576);
nand UO_2194 (O_2194,N_48015,N_46562);
or UO_2195 (O_2195,N_47994,N_48452);
nand UO_2196 (O_2196,N_46039,N_47269);
and UO_2197 (O_2197,N_46223,N_47581);
nand UO_2198 (O_2198,N_49181,N_48424);
xnor UO_2199 (O_2199,N_48407,N_46366);
and UO_2200 (O_2200,N_49888,N_48522);
and UO_2201 (O_2201,N_47342,N_47025);
or UO_2202 (O_2202,N_45746,N_47745);
xnor UO_2203 (O_2203,N_45834,N_45672);
or UO_2204 (O_2204,N_46778,N_45870);
xor UO_2205 (O_2205,N_49595,N_45053);
or UO_2206 (O_2206,N_45781,N_46798);
nand UO_2207 (O_2207,N_48086,N_48156);
nor UO_2208 (O_2208,N_45863,N_45814);
or UO_2209 (O_2209,N_45567,N_48720);
or UO_2210 (O_2210,N_47607,N_45468);
and UO_2211 (O_2211,N_45786,N_46299);
and UO_2212 (O_2212,N_45925,N_48997);
and UO_2213 (O_2213,N_49307,N_48564);
nand UO_2214 (O_2214,N_48164,N_45147);
nor UO_2215 (O_2215,N_46931,N_48080);
and UO_2216 (O_2216,N_45993,N_48254);
nand UO_2217 (O_2217,N_46976,N_45519);
nand UO_2218 (O_2218,N_47159,N_49680);
and UO_2219 (O_2219,N_45168,N_48684);
nor UO_2220 (O_2220,N_49783,N_49761);
or UO_2221 (O_2221,N_46023,N_48892);
xor UO_2222 (O_2222,N_48474,N_48872);
xor UO_2223 (O_2223,N_47972,N_46590);
and UO_2224 (O_2224,N_49185,N_46964);
xor UO_2225 (O_2225,N_46780,N_45716);
nand UO_2226 (O_2226,N_48423,N_45565);
and UO_2227 (O_2227,N_45782,N_45071);
nor UO_2228 (O_2228,N_46873,N_45359);
nor UO_2229 (O_2229,N_46919,N_49532);
or UO_2230 (O_2230,N_46115,N_46899);
nand UO_2231 (O_2231,N_49627,N_47337);
nand UO_2232 (O_2232,N_45855,N_46353);
xor UO_2233 (O_2233,N_49838,N_47806);
and UO_2234 (O_2234,N_47677,N_45501);
xor UO_2235 (O_2235,N_45699,N_49227);
nor UO_2236 (O_2236,N_46249,N_49910);
and UO_2237 (O_2237,N_48366,N_48406);
nand UO_2238 (O_2238,N_46394,N_48094);
or UO_2239 (O_2239,N_46605,N_47687);
and UO_2240 (O_2240,N_49646,N_48874);
nor UO_2241 (O_2241,N_45696,N_46898);
xnor UO_2242 (O_2242,N_47598,N_49708);
nand UO_2243 (O_2243,N_48671,N_47720);
nor UO_2244 (O_2244,N_45073,N_49654);
xnor UO_2245 (O_2245,N_49054,N_49311);
and UO_2246 (O_2246,N_47051,N_47172);
or UO_2247 (O_2247,N_45341,N_49729);
or UO_2248 (O_2248,N_48527,N_49726);
or UO_2249 (O_2249,N_49423,N_45116);
nor UO_2250 (O_2250,N_46411,N_48498);
and UO_2251 (O_2251,N_47251,N_49388);
and UO_2252 (O_2252,N_45522,N_46421);
nand UO_2253 (O_2253,N_46197,N_45491);
nand UO_2254 (O_2254,N_47309,N_47267);
nor UO_2255 (O_2255,N_48594,N_46315);
xnor UO_2256 (O_2256,N_46532,N_46206);
and UO_2257 (O_2257,N_48465,N_48392);
and UO_2258 (O_2258,N_47780,N_46477);
nand UO_2259 (O_2259,N_45488,N_46955);
nor UO_2260 (O_2260,N_49003,N_47146);
and UO_2261 (O_2261,N_45570,N_47286);
or UO_2262 (O_2262,N_46571,N_45212);
or UO_2263 (O_2263,N_49763,N_46138);
and UO_2264 (O_2264,N_48494,N_46144);
or UO_2265 (O_2265,N_45795,N_47628);
nand UO_2266 (O_2266,N_45365,N_46514);
nand UO_2267 (O_2267,N_49402,N_49336);
nand UO_2268 (O_2268,N_48311,N_47221);
nor UO_2269 (O_2269,N_45125,N_46110);
or UO_2270 (O_2270,N_48897,N_48741);
nand UO_2271 (O_2271,N_49852,N_49223);
and UO_2272 (O_2272,N_47755,N_47104);
xor UO_2273 (O_2273,N_45537,N_45281);
nand UO_2274 (O_2274,N_49226,N_48002);
nor UO_2275 (O_2275,N_46232,N_45516);
nor UO_2276 (O_2276,N_49671,N_46323);
nor UO_2277 (O_2277,N_47436,N_45137);
nand UO_2278 (O_2278,N_45720,N_47277);
nand UO_2279 (O_2279,N_49851,N_46892);
nor UO_2280 (O_2280,N_49194,N_47888);
or UO_2281 (O_2281,N_48084,N_48453);
xnor UO_2282 (O_2282,N_48129,N_45436);
or UO_2283 (O_2283,N_48472,N_46440);
nor UO_2284 (O_2284,N_48512,N_49693);
nand UO_2285 (O_2285,N_48330,N_49971);
and UO_2286 (O_2286,N_48503,N_46009);
and UO_2287 (O_2287,N_46677,N_46717);
xor UO_2288 (O_2288,N_49571,N_45411);
or UO_2289 (O_2289,N_49898,N_49039);
nand UO_2290 (O_2290,N_49460,N_45769);
and UO_2291 (O_2291,N_47872,N_47859);
or UO_2292 (O_2292,N_46975,N_45586);
and UO_2293 (O_2293,N_45799,N_48396);
nor UO_2294 (O_2294,N_47563,N_46913);
and UO_2295 (O_2295,N_48806,N_48006);
nand UO_2296 (O_2296,N_46459,N_49813);
xor UO_2297 (O_2297,N_48621,N_45239);
nand UO_2298 (O_2298,N_45233,N_47880);
nor UO_2299 (O_2299,N_48257,N_49260);
and UO_2300 (O_2300,N_49793,N_49706);
xor UO_2301 (O_2301,N_47756,N_45493);
nand UO_2302 (O_2302,N_45536,N_47075);
or UO_2303 (O_2303,N_49026,N_47183);
and UO_2304 (O_2304,N_49091,N_49723);
nor UO_2305 (O_2305,N_46495,N_45155);
nor UO_2306 (O_2306,N_49717,N_49214);
and UO_2307 (O_2307,N_48692,N_49009);
nor UO_2308 (O_2308,N_49897,N_45924);
and UO_2309 (O_2309,N_48402,N_46531);
xnor UO_2310 (O_2310,N_47300,N_47588);
xor UO_2311 (O_2311,N_47297,N_47935);
and UO_2312 (O_2312,N_46858,N_46953);
nand UO_2313 (O_2313,N_49610,N_47842);
and UO_2314 (O_2314,N_47684,N_48414);
or UO_2315 (O_2315,N_45753,N_45033);
or UO_2316 (O_2316,N_49108,N_47550);
nand UO_2317 (O_2317,N_48811,N_49809);
nor UO_2318 (O_2318,N_45021,N_47303);
nor UO_2319 (O_2319,N_47106,N_46273);
or UO_2320 (O_2320,N_47391,N_46011);
nor UO_2321 (O_2321,N_49781,N_49237);
and UO_2322 (O_2322,N_49581,N_45655);
and UO_2323 (O_2323,N_49137,N_45956);
nor UO_2324 (O_2324,N_47886,N_46358);
or UO_2325 (O_2325,N_48515,N_49000);
and UO_2326 (O_2326,N_48740,N_49675);
xor UO_2327 (O_2327,N_47446,N_45348);
nor UO_2328 (O_2328,N_47907,N_49820);
or UO_2329 (O_2329,N_48948,N_47347);
or UO_2330 (O_2330,N_46078,N_48059);
or UO_2331 (O_2331,N_46445,N_47299);
xor UO_2332 (O_2332,N_45573,N_46391);
and UO_2333 (O_2333,N_46024,N_48192);
nand UO_2334 (O_2334,N_46705,N_49705);
xnor UO_2335 (O_2335,N_48136,N_48038);
nand UO_2336 (O_2336,N_48887,N_48697);
and UO_2337 (O_2337,N_45896,N_48520);
xnor UO_2338 (O_2338,N_49373,N_45077);
xor UO_2339 (O_2339,N_48258,N_46207);
xor UO_2340 (O_2340,N_47422,N_48517);
nand UO_2341 (O_2341,N_45841,N_47742);
nand UO_2342 (O_2342,N_45037,N_45176);
nand UO_2343 (O_2343,N_49826,N_48276);
nand UO_2344 (O_2344,N_49078,N_49187);
or UO_2345 (O_2345,N_46375,N_48111);
and UO_2346 (O_2346,N_46145,N_45936);
nor UO_2347 (O_2347,N_46168,N_49398);
or UO_2348 (O_2348,N_45618,N_45885);
and UO_2349 (O_2349,N_49393,N_48835);
and UO_2350 (O_2350,N_45024,N_46554);
or UO_2351 (O_2351,N_48546,N_49086);
or UO_2352 (O_2352,N_48105,N_46293);
nor UO_2353 (O_2353,N_47978,N_49683);
xnor UO_2354 (O_2354,N_48337,N_46140);
and UO_2355 (O_2355,N_48665,N_47691);
nor UO_2356 (O_2356,N_47707,N_48296);
or UO_2357 (O_2357,N_49712,N_49400);
xor UO_2358 (O_2358,N_46652,N_47149);
and UO_2359 (O_2359,N_49241,N_46137);
nor UO_2360 (O_2360,N_47460,N_45783);
and UO_2361 (O_2361,N_47186,N_46874);
nand UO_2362 (O_2362,N_46775,N_45267);
nand UO_2363 (O_2363,N_46611,N_47454);
and UO_2364 (O_2364,N_48477,N_49724);
or UO_2365 (O_2365,N_45857,N_47323);
or UO_2366 (O_2366,N_49098,N_47161);
or UO_2367 (O_2367,N_47751,N_48184);
nor UO_2368 (O_2368,N_45851,N_48918);
nand UO_2369 (O_2369,N_48696,N_49679);
nand UO_2370 (O_2370,N_49057,N_47902);
xnor UO_2371 (O_2371,N_47646,N_46470);
xnor UO_2372 (O_2372,N_46649,N_49203);
and UO_2373 (O_2373,N_46034,N_45298);
and UO_2374 (O_2374,N_48109,N_45861);
nor UO_2375 (O_2375,N_45318,N_45953);
nor UO_2376 (O_2376,N_48460,N_48937);
and UO_2377 (O_2377,N_48981,N_47775);
nand UO_2378 (O_2378,N_49308,N_47917);
nand UO_2379 (O_2379,N_47990,N_46278);
and UO_2380 (O_2380,N_46155,N_46321);
nand UO_2381 (O_2381,N_49142,N_45476);
nand UO_2382 (O_2382,N_49392,N_49144);
xnor UO_2383 (O_2383,N_45192,N_47525);
or UO_2384 (O_2384,N_48327,N_45423);
nand UO_2385 (O_2385,N_47076,N_46546);
nand UO_2386 (O_2386,N_47373,N_48368);
or UO_2387 (O_2387,N_47784,N_48848);
or UO_2388 (O_2388,N_45756,N_45494);
nor UO_2389 (O_2389,N_45052,N_45508);
nand UO_2390 (O_2390,N_45489,N_49037);
or UO_2391 (O_2391,N_46425,N_45983);
and UO_2392 (O_2392,N_49347,N_45617);
nand UO_2393 (O_2393,N_45428,N_46479);
nand UO_2394 (O_2394,N_48487,N_46968);
or UO_2395 (O_2395,N_46081,N_45527);
xor UO_2396 (O_2396,N_49386,N_49816);
or UO_2397 (O_2397,N_49261,N_48374);
and UO_2398 (O_2398,N_48075,N_48271);
nand UO_2399 (O_2399,N_45587,N_49049);
nor UO_2400 (O_2400,N_49282,N_45285);
xor UO_2401 (O_2401,N_45915,N_48161);
nor UO_2402 (O_2402,N_48030,N_46007);
and UO_2403 (O_2403,N_47954,N_45379);
xor UO_2404 (O_2404,N_47469,N_49895);
nand UO_2405 (O_2405,N_45882,N_48766);
or UO_2406 (O_2406,N_47736,N_49497);
or UO_2407 (O_2407,N_46779,N_46764);
xnor UO_2408 (O_2408,N_46121,N_49954);
or UO_2409 (O_2409,N_47959,N_49525);
xnor UO_2410 (O_2410,N_47593,N_48339);
nand UO_2411 (O_2411,N_49887,N_45766);
or UO_2412 (O_2412,N_45452,N_46002);
and UO_2413 (O_2413,N_46883,N_48107);
or UO_2414 (O_2414,N_47118,N_46641);
and UO_2415 (O_2415,N_45540,N_49277);
xor UO_2416 (O_2416,N_49564,N_45836);
nor UO_2417 (O_2417,N_46476,N_46604);
nand UO_2418 (O_2418,N_45303,N_46320);
and UO_2419 (O_2419,N_45314,N_49885);
nand UO_2420 (O_2420,N_48880,N_46199);
and UO_2421 (O_2421,N_46492,N_49014);
and UO_2422 (O_2422,N_49903,N_47497);
nor UO_2423 (O_2423,N_45207,N_46119);
or UO_2424 (O_2424,N_47617,N_46255);
nand UO_2425 (O_2425,N_49930,N_45276);
or UO_2426 (O_2426,N_48289,N_45717);
xnor UO_2427 (O_2427,N_49592,N_49832);
nor UO_2428 (O_2428,N_48382,N_49927);
nor UO_2429 (O_2429,N_46927,N_46125);
xnor UO_2430 (O_2430,N_45275,N_48100);
nand UO_2431 (O_2431,N_45027,N_46452);
or UO_2432 (O_2432,N_46637,N_48994);
or UO_2433 (O_2433,N_47641,N_47003);
and UO_2434 (O_2434,N_48076,N_49697);
or UO_2435 (O_2435,N_47053,N_48067);
xnor UO_2436 (O_2436,N_49244,N_47430);
nand UO_2437 (O_2437,N_49053,N_46342);
nor UO_2438 (O_2438,N_45059,N_49945);
nor UO_2439 (O_2439,N_48983,N_49657);
xor UO_2440 (O_2440,N_45284,N_49924);
nand UO_2441 (O_2441,N_48633,N_49621);
or UO_2442 (O_2442,N_46650,N_46822);
nand UO_2443 (O_2443,N_45317,N_46631);
and UO_2444 (O_2444,N_48764,N_45744);
nor UO_2445 (O_2445,N_48062,N_47949);
nand UO_2446 (O_2446,N_48279,N_47763);
or UO_2447 (O_2447,N_45951,N_49178);
nor UO_2448 (O_2448,N_46201,N_47510);
nand UO_2449 (O_2449,N_48495,N_48014);
or UO_2450 (O_2450,N_46317,N_49312);
xor UO_2451 (O_2451,N_48087,N_47478);
nor UO_2452 (O_2452,N_47507,N_46066);
or UO_2453 (O_2453,N_48719,N_47543);
nor UO_2454 (O_2454,N_45886,N_45074);
nand UO_2455 (O_2455,N_48222,N_47754);
or UO_2456 (O_2456,N_49939,N_48333);
xor UO_2457 (O_2457,N_48307,N_48326);
nand UO_2458 (O_2458,N_46525,N_45979);
or UO_2459 (O_2459,N_46885,N_45738);
nand UO_2460 (O_2460,N_48625,N_46685);
xor UO_2461 (O_2461,N_45588,N_47168);
nand UO_2462 (O_2462,N_49043,N_47123);
xnor UO_2463 (O_2463,N_45563,N_46224);
nand UO_2464 (O_2464,N_48450,N_49846);
or UO_2465 (O_2465,N_49243,N_47693);
nand UO_2466 (O_2466,N_49317,N_48152);
nor UO_2467 (O_2467,N_46175,N_45306);
xnor UO_2468 (O_2468,N_49590,N_47433);
xor UO_2469 (O_2469,N_48315,N_49200);
xor UO_2470 (O_2470,N_47827,N_48668);
xnor UO_2471 (O_2471,N_48864,N_48827);
and UO_2472 (O_2472,N_48426,N_48962);
and UO_2473 (O_2473,N_49570,N_47518);
nand UO_2474 (O_2474,N_49600,N_49501);
or UO_2475 (O_2475,N_49489,N_46570);
and UO_2476 (O_2476,N_47916,N_49115);
nor UO_2477 (O_2477,N_49710,N_47176);
nor UO_2478 (O_2478,N_49411,N_46588);
nor UO_2479 (O_2479,N_47672,N_46771);
nor UO_2480 (O_2480,N_49632,N_48691);
nor UO_2481 (O_2481,N_49448,N_48350);
or UO_2482 (O_2482,N_47849,N_46112);
nor UO_2483 (O_2483,N_49641,N_47530);
nand UO_2484 (O_2484,N_48663,N_47331);
or UO_2485 (O_2485,N_49560,N_47074);
nor UO_2486 (O_2486,N_45957,N_45733);
nor UO_2487 (O_2487,N_49199,N_45578);
or UO_2488 (O_2488,N_46622,N_47052);
xnor UO_2489 (O_2489,N_46917,N_46092);
or UO_2490 (O_2490,N_49071,N_45919);
or UO_2491 (O_2491,N_45364,N_48039);
xnor UO_2492 (O_2492,N_45642,N_47287);
nand UO_2493 (O_2493,N_48454,N_47032);
or UO_2494 (O_2494,N_49151,N_49342);
nor UO_2495 (O_2495,N_46678,N_47178);
or UO_2496 (O_2496,N_47036,N_49206);
nor UO_2497 (O_2497,N_45166,N_49754);
or UO_2498 (O_2498,N_47302,N_45714);
or UO_2499 (O_2499,N_46816,N_45154);
nand UO_2500 (O_2500,N_49878,N_45049);
and UO_2501 (O_2501,N_45101,N_49447);
or UO_2502 (O_2502,N_46168,N_45494);
or UO_2503 (O_2503,N_47013,N_46768);
and UO_2504 (O_2504,N_45732,N_45221);
nand UO_2505 (O_2505,N_48676,N_47256);
nor UO_2506 (O_2506,N_46523,N_48177);
nand UO_2507 (O_2507,N_46876,N_46954);
and UO_2508 (O_2508,N_48307,N_47577);
or UO_2509 (O_2509,N_45119,N_49512);
or UO_2510 (O_2510,N_48031,N_46200);
and UO_2511 (O_2511,N_46356,N_45487);
and UO_2512 (O_2512,N_46442,N_48619);
nor UO_2513 (O_2513,N_45421,N_45816);
xor UO_2514 (O_2514,N_46109,N_47990);
nor UO_2515 (O_2515,N_48488,N_47949);
or UO_2516 (O_2516,N_45928,N_46393);
and UO_2517 (O_2517,N_45894,N_46142);
nor UO_2518 (O_2518,N_46299,N_48985);
xnor UO_2519 (O_2519,N_47479,N_45589);
or UO_2520 (O_2520,N_46398,N_49411);
and UO_2521 (O_2521,N_46604,N_47471);
and UO_2522 (O_2522,N_46158,N_45940);
xnor UO_2523 (O_2523,N_49538,N_49618);
xor UO_2524 (O_2524,N_47111,N_47630);
nand UO_2525 (O_2525,N_47998,N_45113);
nand UO_2526 (O_2526,N_46931,N_47312);
and UO_2527 (O_2527,N_47332,N_45766);
and UO_2528 (O_2528,N_48222,N_49593);
nand UO_2529 (O_2529,N_47056,N_46052);
nor UO_2530 (O_2530,N_45349,N_45889);
or UO_2531 (O_2531,N_49869,N_45547);
and UO_2532 (O_2532,N_47210,N_48713);
and UO_2533 (O_2533,N_46508,N_45969);
or UO_2534 (O_2534,N_49025,N_49106);
xnor UO_2535 (O_2535,N_48841,N_48958);
and UO_2536 (O_2536,N_45585,N_45786);
nor UO_2537 (O_2537,N_47277,N_45790);
xnor UO_2538 (O_2538,N_45385,N_49466);
xnor UO_2539 (O_2539,N_48325,N_47607);
nor UO_2540 (O_2540,N_45099,N_48944);
nor UO_2541 (O_2541,N_47157,N_45809);
nand UO_2542 (O_2542,N_49330,N_46685);
nor UO_2543 (O_2543,N_49486,N_48265);
nor UO_2544 (O_2544,N_47330,N_46053);
xor UO_2545 (O_2545,N_48337,N_45913);
or UO_2546 (O_2546,N_46366,N_46834);
xnor UO_2547 (O_2547,N_45160,N_45159);
xnor UO_2548 (O_2548,N_45296,N_47408);
nand UO_2549 (O_2549,N_48350,N_45570);
nand UO_2550 (O_2550,N_47949,N_48808);
nor UO_2551 (O_2551,N_49242,N_47965);
nand UO_2552 (O_2552,N_49082,N_48665);
nand UO_2553 (O_2553,N_48329,N_48672);
nor UO_2554 (O_2554,N_48448,N_45579);
or UO_2555 (O_2555,N_45805,N_45426);
or UO_2556 (O_2556,N_48293,N_47936);
nor UO_2557 (O_2557,N_47025,N_45169);
xor UO_2558 (O_2558,N_45135,N_48220);
or UO_2559 (O_2559,N_49775,N_46839);
nand UO_2560 (O_2560,N_48273,N_46016);
nor UO_2561 (O_2561,N_46424,N_49221);
nand UO_2562 (O_2562,N_48340,N_49374);
and UO_2563 (O_2563,N_46581,N_48643);
nand UO_2564 (O_2564,N_47062,N_49737);
nand UO_2565 (O_2565,N_47713,N_46073);
nor UO_2566 (O_2566,N_47701,N_49437);
nand UO_2567 (O_2567,N_48018,N_47541);
or UO_2568 (O_2568,N_47709,N_45127);
nor UO_2569 (O_2569,N_46387,N_46312);
nor UO_2570 (O_2570,N_48287,N_45833);
xor UO_2571 (O_2571,N_47586,N_45716);
xor UO_2572 (O_2572,N_49491,N_46672);
and UO_2573 (O_2573,N_48206,N_49393);
or UO_2574 (O_2574,N_47721,N_46810);
and UO_2575 (O_2575,N_46641,N_47201);
nor UO_2576 (O_2576,N_46613,N_47075);
and UO_2577 (O_2577,N_46568,N_48563);
nor UO_2578 (O_2578,N_47075,N_45753);
nor UO_2579 (O_2579,N_46145,N_49448);
or UO_2580 (O_2580,N_47599,N_49851);
xor UO_2581 (O_2581,N_45943,N_49530);
and UO_2582 (O_2582,N_46355,N_49076);
nand UO_2583 (O_2583,N_49951,N_47723);
and UO_2584 (O_2584,N_46853,N_47102);
or UO_2585 (O_2585,N_46346,N_49126);
and UO_2586 (O_2586,N_49118,N_49984);
or UO_2587 (O_2587,N_48357,N_48999);
or UO_2588 (O_2588,N_49570,N_46339);
and UO_2589 (O_2589,N_49361,N_47809);
and UO_2590 (O_2590,N_46066,N_49395);
xnor UO_2591 (O_2591,N_47471,N_46598);
nor UO_2592 (O_2592,N_47783,N_47698);
or UO_2593 (O_2593,N_47895,N_49361);
nor UO_2594 (O_2594,N_48142,N_48438);
or UO_2595 (O_2595,N_48689,N_46108);
nand UO_2596 (O_2596,N_45185,N_48081);
nand UO_2597 (O_2597,N_48156,N_45437);
and UO_2598 (O_2598,N_46513,N_45677);
nand UO_2599 (O_2599,N_49547,N_49264);
xnor UO_2600 (O_2600,N_48175,N_47423);
nor UO_2601 (O_2601,N_45975,N_47200);
or UO_2602 (O_2602,N_48684,N_45516);
nor UO_2603 (O_2603,N_46972,N_49887);
xor UO_2604 (O_2604,N_47955,N_46726);
nand UO_2605 (O_2605,N_46188,N_46752);
nor UO_2606 (O_2606,N_48042,N_49686);
and UO_2607 (O_2607,N_46685,N_45437);
and UO_2608 (O_2608,N_49503,N_45166);
and UO_2609 (O_2609,N_49033,N_45509);
and UO_2610 (O_2610,N_46038,N_46570);
nand UO_2611 (O_2611,N_45146,N_47217);
nand UO_2612 (O_2612,N_45035,N_48825);
nand UO_2613 (O_2613,N_48407,N_49353);
nand UO_2614 (O_2614,N_45903,N_49938);
and UO_2615 (O_2615,N_48196,N_47425);
nor UO_2616 (O_2616,N_48653,N_47157);
and UO_2617 (O_2617,N_45938,N_47431);
xnor UO_2618 (O_2618,N_49566,N_47453);
and UO_2619 (O_2619,N_47060,N_49958);
and UO_2620 (O_2620,N_45543,N_47543);
xor UO_2621 (O_2621,N_45003,N_45886);
xor UO_2622 (O_2622,N_45681,N_46826);
or UO_2623 (O_2623,N_48779,N_47360);
or UO_2624 (O_2624,N_47892,N_46699);
xor UO_2625 (O_2625,N_47153,N_45802);
or UO_2626 (O_2626,N_48139,N_48677);
or UO_2627 (O_2627,N_48304,N_48669);
or UO_2628 (O_2628,N_48000,N_48990);
nand UO_2629 (O_2629,N_47603,N_46475);
and UO_2630 (O_2630,N_48260,N_49572);
nand UO_2631 (O_2631,N_46037,N_46931);
or UO_2632 (O_2632,N_49753,N_49506);
and UO_2633 (O_2633,N_49485,N_49636);
nand UO_2634 (O_2634,N_46920,N_49493);
nor UO_2635 (O_2635,N_49994,N_47242);
or UO_2636 (O_2636,N_46617,N_45105);
nand UO_2637 (O_2637,N_48350,N_49998);
and UO_2638 (O_2638,N_49025,N_47343);
xor UO_2639 (O_2639,N_47353,N_45261);
or UO_2640 (O_2640,N_49802,N_46004);
and UO_2641 (O_2641,N_47008,N_47133);
xnor UO_2642 (O_2642,N_49900,N_48210);
xnor UO_2643 (O_2643,N_49050,N_49991);
and UO_2644 (O_2644,N_49861,N_49499);
nand UO_2645 (O_2645,N_48767,N_49410);
and UO_2646 (O_2646,N_47419,N_45394);
nand UO_2647 (O_2647,N_48179,N_47020);
nor UO_2648 (O_2648,N_49096,N_47237);
nand UO_2649 (O_2649,N_48045,N_46996);
nand UO_2650 (O_2650,N_48794,N_46100);
or UO_2651 (O_2651,N_49518,N_49069);
nand UO_2652 (O_2652,N_47008,N_47619);
or UO_2653 (O_2653,N_47398,N_46445);
nor UO_2654 (O_2654,N_45798,N_49971);
nor UO_2655 (O_2655,N_47054,N_47287);
nand UO_2656 (O_2656,N_47359,N_46814);
or UO_2657 (O_2657,N_46027,N_45654);
xnor UO_2658 (O_2658,N_47362,N_46896);
nand UO_2659 (O_2659,N_48503,N_46797);
and UO_2660 (O_2660,N_48498,N_48887);
or UO_2661 (O_2661,N_45096,N_45290);
or UO_2662 (O_2662,N_47447,N_45673);
or UO_2663 (O_2663,N_48761,N_45608);
and UO_2664 (O_2664,N_47020,N_46622);
nand UO_2665 (O_2665,N_47794,N_45226);
or UO_2666 (O_2666,N_48798,N_45373);
and UO_2667 (O_2667,N_47124,N_48424);
nand UO_2668 (O_2668,N_48190,N_49470);
or UO_2669 (O_2669,N_45968,N_48064);
or UO_2670 (O_2670,N_48950,N_47930);
nand UO_2671 (O_2671,N_48824,N_46846);
and UO_2672 (O_2672,N_45599,N_49977);
xor UO_2673 (O_2673,N_45291,N_45922);
nor UO_2674 (O_2674,N_45115,N_48139);
or UO_2675 (O_2675,N_45715,N_45537);
and UO_2676 (O_2676,N_48588,N_49785);
or UO_2677 (O_2677,N_46532,N_49246);
nor UO_2678 (O_2678,N_45021,N_49711);
and UO_2679 (O_2679,N_47051,N_48277);
and UO_2680 (O_2680,N_46526,N_48986);
and UO_2681 (O_2681,N_47714,N_47994);
nor UO_2682 (O_2682,N_48193,N_49781);
and UO_2683 (O_2683,N_48197,N_47178);
xor UO_2684 (O_2684,N_49758,N_47712);
nand UO_2685 (O_2685,N_46451,N_47642);
nand UO_2686 (O_2686,N_48478,N_46128);
nor UO_2687 (O_2687,N_45339,N_46763);
xor UO_2688 (O_2688,N_47370,N_49660);
or UO_2689 (O_2689,N_45251,N_45278);
or UO_2690 (O_2690,N_46836,N_49633);
and UO_2691 (O_2691,N_49758,N_47079);
nand UO_2692 (O_2692,N_45056,N_46729);
and UO_2693 (O_2693,N_48969,N_48185);
nand UO_2694 (O_2694,N_47577,N_49449);
nor UO_2695 (O_2695,N_47957,N_47590);
nor UO_2696 (O_2696,N_45532,N_48866);
nor UO_2697 (O_2697,N_49292,N_46843);
nand UO_2698 (O_2698,N_48023,N_45279);
and UO_2699 (O_2699,N_49008,N_49564);
or UO_2700 (O_2700,N_45940,N_48328);
nand UO_2701 (O_2701,N_46243,N_46583);
and UO_2702 (O_2702,N_49216,N_46154);
nor UO_2703 (O_2703,N_48494,N_49796);
and UO_2704 (O_2704,N_46074,N_46227);
nand UO_2705 (O_2705,N_45416,N_45288);
nand UO_2706 (O_2706,N_49621,N_47364);
nand UO_2707 (O_2707,N_47784,N_48949);
xnor UO_2708 (O_2708,N_45746,N_49236);
and UO_2709 (O_2709,N_45528,N_48285);
nand UO_2710 (O_2710,N_49006,N_48124);
xnor UO_2711 (O_2711,N_48421,N_46902);
nor UO_2712 (O_2712,N_48000,N_45946);
nand UO_2713 (O_2713,N_47308,N_47708);
nor UO_2714 (O_2714,N_46833,N_46330);
or UO_2715 (O_2715,N_45829,N_49999);
or UO_2716 (O_2716,N_45794,N_49187);
nor UO_2717 (O_2717,N_47217,N_46755);
nor UO_2718 (O_2718,N_45832,N_48851);
xnor UO_2719 (O_2719,N_48511,N_47430);
or UO_2720 (O_2720,N_48914,N_47984);
nor UO_2721 (O_2721,N_48448,N_46980);
nand UO_2722 (O_2722,N_47590,N_48702);
nand UO_2723 (O_2723,N_49109,N_45466);
nor UO_2724 (O_2724,N_48346,N_48736);
nand UO_2725 (O_2725,N_48156,N_46846);
and UO_2726 (O_2726,N_47114,N_49026);
nor UO_2727 (O_2727,N_47289,N_47820);
and UO_2728 (O_2728,N_46088,N_45703);
nand UO_2729 (O_2729,N_49894,N_48193);
or UO_2730 (O_2730,N_46340,N_47810);
and UO_2731 (O_2731,N_49404,N_47045);
or UO_2732 (O_2732,N_49513,N_49853);
nand UO_2733 (O_2733,N_47526,N_48041);
nor UO_2734 (O_2734,N_49566,N_46556);
or UO_2735 (O_2735,N_48129,N_46519);
and UO_2736 (O_2736,N_48529,N_48711);
nor UO_2737 (O_2737,N_46371,N_49832);
nand UO_2738 (O_2738,N_46501,N_47613);
nand UO_2739 (O_2739,N_48029,N_46745);
nor UO_2740 (O_2740,N_46628,N_46056);
nor UO_2741 (O_2741,N_45171,N_49761);
xnor UO_2742 (O_2742,N_48861,N_46880);
or UO_2743 (O_2743,N_46677,N_47485);
or UO_2744 (O_2744,N_48808,N_49879);
or UO_2745 (O_2745,N_45801,N_45106);
xor UO_2746 (O_2746,N_46189,N_45857);
nand UO_2747 (O_2747,N_48675,N_49279);
nand UO_2748 (O_2748,N_45672,N_48089);
xor UO_2749 (O_2749,N_45266,N_47046);
and UO_2750 (O_2750,N_45747,N_45279);
or UO_2751 (O_2751,N_47568,N_47159);
nand UO_2752 (O_2752,N_46983,N_47847);
or UO_2753 (O_2753,N_48804,N_45639);
and UO_2754 (O_2754,N_46944,N_46534);
nor UO_2755 (O_2755,N_48556,N_47554);
nor UO_2756 (O_2756,N_45405,N_46237);
xor UO_2757 (O_2757,N_47740,N_47753);
and UO_2758 (O_2758,N_47114,N_45177);
or UO_2759 (O_2759,N_48750,N_48210);
xnor UO_2760 (O_2760,N_45860,N_47240);
and UO_2761 (O_2761,N_45345,N_47640);
nor UO_2762 (O_2762,N_48502,N_47496);
xor UO_2763 (O_2763,N_47859,N_45581);
or UO_2764 (O_2764,N_49404,N_47549);
or UO_2765 (O_2765,N_46419,N_49208);
or UO_2766 (O_2766,N_47207,N_45145);
and UO_2767 (O_2767,N_49595,N_47335);
nor UO_2768 (O_2768,N_48727,N_47359);
xor UO_2769 (O_2769,N_48238,N_46171);
xnor UO_2770 (O_2770,N_45551,N_46286);
nand UO_2771 (O_2771,N_45303,N_46258);
or UO_2772 (O_2772,N_48326,N_46034);
and UO_2773 (O_2773,N_47226,N_46032);
xor UO_2774 (O_2774,N_48087,N_46530);
nor UO_2775 (O_2775,N_49950,N_49283);
nand UO_2776 (O_2776,N_48706,N_47908);
nand UO_2777 (O_2777,N_49003,N_48617);
or UO_2778 (O_2778,N_48805,N_45550);
xor UO_2779 (O_2779,N_45807,N_47199);
and UO_2780 (O_2780,N_49769,N_48266);
xnor UO_2781 (O_2781,N_46834,N_46286);
nor UO_2782 (O_2782,N_48420,N_47085);
and UO_2783 (O_2783,N_49959,N_48819);
nor UO_2784 (O_2784,N_46333,N_46511);
and UO_2785 (O_2785,N_45548,N_47804);
nand UO_2786 (O_2786,N_47770,N_49011);
xnor UO_2787 (O_2787,N_49667,N_45382);
and UO_2788 (O_2788,N_48641,N_48378);
or UO_2789 (O_2789,N_49547,N_48004);
nand UO_2790 (O_2790,N_49127,N_45755);
nand UO_2791 (O_2791,N_45333,N_45258);
or UO_2792 (O_2792,N_48833,N_49943);
or UO_2793 (O_2793,N_45838,N_47777);
nor UO_2794 (O_2794,N_48097,N_45910);
nor UO_2795 (O_2795,N_45833,N_47470);
nor UO_2796 (O_2796,N_47515,N_49805);
xnor UO_2797 (O_2797,N_45490,N_49011);
xor UO_2798 (O_2798,N_47802,N_47481);
nand UO_2799 (O_2799,N_46412,N_47425);
xnor UO_2800 (O_2800,N_46685,N_46380);
or UO_2801 (O_2801,N_49449,N_47946);
nor UO_2802 (O_2802,N_47077,N_46496);
or UO_2803 (O_2803,N_45972,N_46191);
nand UO_2804 (O_2804,N_47539,N_47289);
nand UO_2805 (O_2805,N_45756,N_48498);
xnor UO_2806 (O_2806,N_45478,N_49488);
or UO_2807 (O_2807,N_49197,N_46642);
nand UO_2808 (O_2808,N_47557,N_45893);
nand UO_2809 (O_2809,N_47899,N_46364);
nor UO_2810 (O_2810,N_48969,N_46230);
and UO_2811 (O_2811,N_45972,N_47917);
and UO_2812 (O_2812,N_46230,N_45657);
or UO_2813 (O_2813,N_45407,N_47100);
or UO_2814 (O_2814,N_46809,N_46680);
nor UO_2815 (O_2815,N_46821,N_45873);
or UO_2816 (O_2816,N_48964,N_45606);
or UO_2817 (O_2817,N_47017,N_45713);
nand UO_2818 (O_2818,N_48118,N_45747);
and UO_2819 (O_2819,N_48115,N_48275);
or UO_2820 (O_2820,N_45607,N_49372);
nand UO_2821 (O_2821,N_47156,N_45463);
and UO_2822 (O_2822,N_45291,N_47738);
nand UO_2823 (O_2823,N_45003,N_45509);
or UO_2824 (O_2824,N_49939,N_47718);
nor UO_2825 (O_2825,N_48795,N_48726);
and UO_2826 (O_2826,N_45975,N_45193);
xor UO_2827 (O_2827,N_48798,N_45415);
nor UO_2828 (O_2828,N_48447,N_49726);
and UO_2829 (O_2829,N_46713,N_47062);
nand UO_2830 (O_2830,N_47491,N_45702);
or UO_2831 (O_2831,N_48373,N_45839);
xnor UO_2832 (O_2832,N_46938,N_48493);
and UO_2833 (O_2833,N_46264,N_47515);
nand UO_2834 (O_2834,N_49204,N_48685);
and UO_2835 (O_2835,N_45237,N_47044);
and UO_2836 (O_2836,N_48872,N_47096);
or UO_2837 (O_2837,N_48848,N_47365);
xnor UO_2838 (O_2838,N_47528,N_47016);
xnor UO_2839 (O_2839,N_48966,N_47959);
nand UO_2840 (O_2840,N_48087,N_46439);
xor UO_2841 (O_2841,N_48263,N_45024);
or UO_2842 (O_2842,N_46889,N_45321);
xnor UO_2843 (O_2843,N_46203,N_46385);
or UO_2844 (O_2844,N_49018,N_46914);
or UO_2845 (O_2845,N_49834,N_46398);
nor UO_2846 (O_2846,N_47018,N_47831);
nor UO_2847 (O_2847,N_49163,N_46694);
nand UO_2848 (O_2848,N_49708,N_47399);
xnor UO_2849 (O_2849,N_47411,N_49255);
and UO_2850 (O_2850,N_48629,N_48082);
nor UO_2851 (O_2851,N_49989,N_47557);
xor UO_2852 (O_2852,N_45982,N_49122);
nor UO_2853 (O_2853,N_48314,N_47661);
and UO_2854 (O_2854,N_48328,N_48797);
xor UO_2855 (O_2855,N_45828,N_45502);
nand UO_2856 (O_2856,N_47316,N_47837);
nand UO_2857 (O_2857,N_45105,N_48459);
or UO_2858 (O_2858,N_48476,N_49835);
nand UO_2859 (O_2859,N_47471,N_48141);
nand UO_2860 (O_2860,N_47341,N_47222);
nand UO_2861 (O_2861,N_46138,N_49256);
nand UO_2862 (O_2862,N_47088,N_46760);
or UO_2863 (O_2863,N_49819,N_47571);
xor UO_2864 (O_2864,N_47993,N_46717);
or UO_2865 (O_2865,N_47256,N_49776);
nand UO_2866 (O_2866,N_45381,N_48664);
and UO_2867 (O_2867,N_46039,N_45741);
nor UO_2868 (O_2868,N_45107,N_45235);
or UO_2869 (O_2869,N_46079,N_47111);
and UO_2870 (O_2870,N_48286,N_45239);
nand UO_2871 (O_2871,N_47062,N_48973);
or UO_2872 (O_2872,N_47606,N_46249);
and UO_2873 (O_2873,N_47744,N_47416);
and UO_2874 (O_2874,N_49162,N_48317);
nand UO_2875 (O_2875,N_45961,N_48673);
or UO_2876 (O_2876,N_49018,N_48750);
nand UO_2877 (O_2877,N_47728,N_49794);
nor UO_2878 (O_2878,N_48576,N_47603);
and UO_2879 (O_2879,N_45866,N_45711);
nor UO_2880 (O_2880,N_49155,N_45563);
nor UO_2881 (O_2881,N_47182,N_49915);
nor UO_2882 (O_2882,N_45367,N_49979);
and UO_2883 (O_2883,N_48669,N_45002);
and UO_2884 (O_2884,N_48487,N_46033);
or UO_2885 (O_2885,N_46737,N_47849);
xor UO_2886 (O_2886,N_49156,N_45050);
and UO_2887 (O_2887,N_45997,N_45974);
nor UO_2888 (O_2888,N_48531,N_49561);
or UO_2889 (O_2889,N_46219,N_45354);
nand UO_2890 (O_2890,N_48751,N_49671);
or UO_2891 (O_2891,N_48766,N_49405);
nand UO_2892 (O_2892,N_47597,N_46261);
or UO_2893 (O_2893,N_47088,N_45100);
or UO_2894 (O_2894,N_46244,N_48269);
nor UO_2895 (O_2895,N_48598,N_47690);
nor UO_2896 (O_2896,N_46798,N_45117);
or UO_2897 (O_2897,N_48134,N_47844);
nand UO_2898 (O_2898,N_46983,N_48578);
xor UO_2899 (O_2899,N_46433,N_49268);
nand UO_2900 (O_2900,N_48487,N_46370);
and UO_2901 (O_2901,N_48761,N_46239);
nor UO_2902 (O_2902,N_45336,N_49386);
nor UO_2903 (O_2903,N_46349,N_45629);
xor UO_2904 (O_2904,N_48537,N_46635);
xnor UO_2905 (O_2905,N_47367,N_48972);
and UO_2906 (O_2906,N_46286,N_48233);
nand UO_2907 (O_2907,N_45572,N_48912);
xor UO_2908 (O_2908,N_45953,N_47145);
xor UO_2909 (O_2909,N_46279,N_48924);
or UO_2910 (O_2910,N_45055,N_46543);
or UO_2911 (O_2911,N_49396,N_46686);
xor UO_2912 (O_2912,N_46978,N_49718);
nor UO_2913 (O_2913,N_49961,N_46763);
and UO_2914 (O_2914,N_45201,N_47622);
and UO_2915 (O_2915,N_49396,N_45571);
and UO_2916 (O_2916,N_46085,N_47577);
or UO_2917 (O_2917,N_48735,N_45473);
nand UO_2918 (O_2918,N_48983,N_45889);
xnor UO_2919 (O_2919,N_45601,N_48800);
or UO_2920 (O_2920,N_47669,N_46491);
or UO_2921 (O_2921,N_45033,N_48251);
and UO_2922 (O_2922,N_46788,N_47931);
nand UO_2923 (O_2923,N_45806,N_46387);
and UO_2924 (O_2924,N_46428,N_45350);
nand UO_2925 (O_2925,N_49942,N_45115);
nand UO_2926 (O_2926,N_48296,N_45762);
or UO_2927 (O_2927,N_47762,N_45779);
nand UO_2928 (O_2928,N_47647,N_45100);
or UO_2929 (O_2929,N_46433,N_46138);
nor UO_2930 (O_2930,N_46985,N_45283);
and UO_2931 (O_2931,N_47362,N_45201);
nor UO_2932 (O_2932,N_46181,N_48882);
xnor UO_2933 (O_2933,N_48320,N_47524);
nand UO_2934 (O_2934,N_49388,N_46327);
and UO_2935 (O_2935,N_48899,N_48789);
nor UO_2936 (O_2936,N_48494,N_46625);
nand UO_2937 (O_2937,N_49493,N_48917);
nor UO_2938 (O_2938,N_48950,N_48817);
or UO_2939 (O_2939,N_49908,N_48184);
nor UO_2940 (O_2940,N_45976,N_48428);
xor UO_2941 (O_2941,N_48755,N_46634);
and UO_2942 (O_2942,N_49285,N_47534);
or UO_2943 (O_2943,N_48594,N_47420);
and UO_2944 (O_2944,N_47468,N_45338);
and UO_2945 (O_2945,N_47981,N_45540);
or UO_2946 (O_2946,N_49954,N_49403);
nor UO_2947 (O_2947,N_49618,N_47352);
and UO_2948 (O_2948,N_49013,N_46210);
xnor UO_2949 (O_2949,N_47081,N_47426);
nor UO_2950 (O_2950,N_48325,N_47783);
nor UO_2951 (O_2951,N_47752,N_47867);
xnor UO_2952 (O_2952,N_45103,N_45751);
nor UO_2953 (O_2953,N_45712,N_49498);
nand UO_2954 (O_2954,N_45911,N_46916);
or UO_2955 (O_2955,N_45590,N_47484);
or UO_2956 (O_2956,N_45461,N_48728);
nor UO_2957 (O_2957,N_46240,N_48159);
nand UO_2958 (O_2958,N_47756,N_49366);
xnor UO_2959 (O_2959,N_46255,N_45903);
and UO_2960 (O_2960,N_48351,N_47689);
or UO_2961 (O_2961,N_47823,N_48422);
and UO_2962 (O_2962,N_48056,N_49821);
or UO_2963 (O_2963,N_46824,N_47532);
xor UO_2964 (O_2964,N_49786,N_45236);
nor UO_2965 (O_2965,N_46355,N_49951);
nand UO_2966 (O_2966,N_47583,N_49852);
nand UO_2967 (O_2967,N_46475,N_46660);
and UO_2968 (O_2968,N_46970,N_45816);
nand UO_2969 (O_2969,N_49156,N_48725);
or UO_2970 (O_2970,N_46889,N_49793);
nand UO_2971 (O_2971,N_48118,N_49786);
or UO_2972 (O_2972,N_47272,N_49045);
and UO_2973 (O_2973,N_46583,N_48990);
nand UO_2974 (O_2974,N_49464,N_45021);
nand UO_2975 (O_2975,N_49897,N_48312);
or UO_2976 (O_2976,N_45631,N_49206);
xnor UO_2977 (O_2977,N_48690,N_47340);
and UO_2978 (O_2978,N_47091,N_45784);
or UO_2979 (O_2979,N_48514,N_48766);
nand UO_2980 (O_2980,N_46318,N_47929);
nor UO_2981 (O_2981,N_45975,N_49440);
xnor UO_2982 (O_2982,N_46592,N_47407);
or UO_2983 (O_2983,N_47613,N_45178);
nor UO_2984 (O_2984,N_46892,N_48245);
xor UO_2985 (O_2985,N_46187,N_45544);
nor UO_2986 (O_2986,N_46751,N_46592);
nor UO_2987 (O_2987,N_49426,N_48865);
or UO_2988 (O_2988,N_45421,N_49321);
and UO_2989 (O_2989,N_45221,N_47382);
nand UO_2990 (O_2990,N_49464,N_49774);
xnor UO_2991 (O_2991,N_48923,N_47822);
or UO_2992 (O_2992,N_47403,N_48982);
nand UO_2993 (O_2993,N_47859,N_46207);
or UO_2994 (O_2994,N_48304,N_49274);
xor UO_2995 (O_2995,N_46097,N_48010);
nand UO_2996 (O_2996,N_46833,N_46143);
nor UO_2997 (O_2997,N_45139,N_49448);
and UO_2998 (O_2998,N_47131,N_45015);
and UO_2999 (O_2999,N_49957,N_45996);
nand UO_3000 (O_3000,N_48130,N_48921);
and UO_3001 (O_3001,N_48910,N_49932);
and UO_3002 (O_3002,N_47299,N_48321);
or UO_3003 (O_3003,N_47397,N_48360);
and UO_3004 (O_3004,N_45508,N_46098);
nor UO_3005 (O_3005,N_49347,N_47213);
and UO_3006 (O_3006,N_47975,N_46223);
nand UO_3007 (O_3007,N_45459,N_46585);
or UO_3008 (O_3008,N_48297,N_49969);
xor UO_3009 (O_3009,N_45681,N_46045);
xor UO_3010 (O_3010,N_46460,N_47448);
and UO_3011 (O_3011,N_49895,N_47433);
nor UO_3012 (O_3012,N_49107,N_48471);
nand UO_3013 (O_3013,N_46409,N_47870);
nand UO_3014 (O_3014,N_45532,N_49106);
nand UO_3015 (O_3015,N_49595,N_48581);
nand UO_3016 (O_3016,N_47280,N_47483);
xnor UO_3017 (O_3017,N_48163,N_47708);
xor UO_3018 (O_3018,N_49371,N_45943);
nor UO_3019 (O_3019,N_48933,N_47649);
or UO_3020 (O_3020,N_45907,N_45736);
xnor UO_3021 (O_3021,N_45581,N_49965);
nor UO_3022 (O_3022,N_48373,N_47543);
nor UO_3023 (O_3023,N_49750,N_49048);
nor UO_3024 (O_3024,N_45306,N_47172);
nand UO_3025 (O_3025,N_48689,N_47387);
and UO_3026 (O_3026,N_46206,N_46115);
and UO_3027 (O_3027,N_47757,N_47824);
and UO_3028 (O_3028,N_47176,N_47649);
nor UO_3029 (O_3029,N_46647,N_48640);
nor UO_3030 (O_3030,N_47973,N_48516);
nor UO_3031 (O_3031,N_49460,N_45657);
or UO_3032 (O_3032,N_46453,N_49577);
and UO_3033 (O_3033,N_46468,N_48273);
xnor UO_3034 (O_3034,N_45300,N_46652);
nand UO_3035 (O_3035,N_48628,N_47267);
nor UO_3036 (O_3036,N_47799,N_48699);
xnor UO_3037 (O_3037,N_47763,N_49002);
nor UO_3038 (O_3038,N_48413,N_45060);
and UO_3039 (O_3039,N_47718,N_48591);
nand UO_3040 (O_3040,N_46131,N_49508);
nor UO_3041 (O_3041,N_45832,N_47531);
xnor UO_3042 (O_3042,N_47162,N_49124);
or UO_3043 (O_3043,N_47253,N_45380);
nor UO_3044 (O_3044,N_45614,N_48558);
xnor UO_3045 (O_3045,N_49718,N_45262);
nor UO_3046 (O_3046,N_48818,N_48206);
and UO_3047 (O_3047,N_48591,N_48267);
nand UO_3048 (O_3048,N_49259,N_47822);
nand UO_3049 (O_3049,N_47264,N_47544);
or UO_3050 (O_3050,N_47657,N_47580);
nor UO_3051 (O_3051,N_45583,N_46278);
and UO_3052 (O_3052,N_45314,N_47856);
nand UO_3053 (O_3053,N_45650,N_47924);
and UO_3054 (O_3054,N_46748,N_47024);
or UO_3055 (O_3055,N_47499,N_46562);
nor UO_3056 (O_3056,N_46649,N_47799);
nor UO_3057 (O_3057,N_46949,N_47516);
or UO_3058 (O_3058,N_46633,N_45812);
xor UO_3059 (O_3059,N_47087,N_46889);
nor UO_3060 (O_3060,N_45906,N_49945);
xnor UO_3061 (O_3061,N_47808,N_48141);
and UO_3062 (O_3062,N_48375,N_48182);
nand UO_3063 (O_3063,N_48864,N_47283);
or UO_3064 (O_3064,N_46359,N_48022);
and UO_3065 (O_3065,N_46947,N_46586);
nand UO_3066 (O_3066,N_48433,N_49364);
nor UO_3067 (O_3067,N_46015,N_48570);
and UO_3068 (O_3068,N_46540,N_49510);
and UO_3069 (O_3069,N_46279,N_48362);
nand UO_3070 (O_3070,N_47996,N_47871);
xnor UO_3071 (O_3071,N_48843,N_47619);
or UO_3072 (O_3072,N_47465,N_49603);
nand UO_3073 (O_3073,N_48163,N_49747);
and UO_3074 (O_3074,N_49125,N_45504);
nand UO_3075 (O_3075,N_45826,N_47237);
or UO_3076 (O_3076,N_48989,N_48066);
xor UO_3077 (O_3077,N_46579,N_49639);
nor UO_3078 (O_3078,N_48805,N_48347);
and UO_3079 (O_3079,N_47651,N_48077);
nor UO_3080 (O_3080,N_46974,N_45621);
or UO_3081 (O_3081,N_47621,N_49237);
xor UO_3082 (O_3082,N_47605,N_45382);
nor UO_3083 (O_3083,N_49928,N_45315);
nor UO_3084 (O_3084,N_48453,N_47627);
or UO_3085 (O_3085,N_47392,N_45281);
or UO_3086 (O_3086,N_45859,N_47111);
xor UO_3087 (O_3087,N_48126,N_49528);
nand UO_3088 (O_3088,N_46061,N_45778);
nand UO_3089 (O_3089,N_46049,N_48020);
nor UO_3090 (O_3090,N_49328,N_46460);
or UO_3091 (O_3091,N_45691,N_48618);
xor UO_3092 (O_3092,N_47409,N_46357);
and UO_3093 (O_3093,N_46777,N_45507);
nand UO_3094 (O_3094,N_47478,N_47455);
and UO_3095 (O_3095,N_48940,N_46402);
and UO_3096 (O_3096,N_48966,N_47428);
or UO_3097 (O_3097,N_49698,N_47468);
nor UO_3098 (O_3098,N_46681,N_49970);
xor UO_3099 (O_3099,N_45720,N_49617);
or UO_3100 (O_3100,N_47379,N_45692);
nand UO_3101 (O_3101,N_49737,N_46732);
nor UO_3102 (O_3102,N_47742,N_47094);
or UO_3103 (O_3103,N_49529,N_49189);
xnor UO_3104 (O_3104,N_45004,N_49223);
or UO_3105 (O_3105,N_49684,N_46517);
xnor UO_3106 (O_3106,N_45085,N_47956);
xnor UO_3107 (O_3107,N_45903,N_49017);
or UO_3108 (O_3108,N_45239,N_49094);
nor UO_3109 (O_3109,N_48582,N_48779);
nand UO_3110 (O_3110,N_48094,N_45963);
xnor UO_3111 (O_3111,N_46781,N_45956);
nor UO_3112 (O_3112,N_48688,N_49903);
and UO_3113 (O_3113,N_45298,N_45773);
or UO_3114 (O_3114,N_47989,N_45731);
nor UO_3115 (O_3115,N_49033,N_46720);
xnor UO_3116 (O_3116,N_46180,N_48741);
xor UO_3117 (O_3117,N_49089,N_49829);
or UO_3118 (O_3118,N_46854,N_45705);
xnor UO_3119 (O_3119,N_47094,N_48044);
xor UO_3120 (O_3120,N_48567,N_48159);
nor UO_3121 (O_3121,N_48420,N_48100);
and UO_3122 (O_3122,N_49788,N_45549);
and UO_3123 (O_3123,N_46681,N_49358);
and UO_3124 (O_3124,N_47376,N_49965);
nand UO_3125 (O_3125,N_46445,N_48113);
or UO_3126 (O_3126,N_47497,N_45901);
nor UO_3127 (O_3127,N_47547,N_47062);
or UO_3128 (O_3128,N_46838,N_48595);
and UO_3129 (O_3129,N_49308,N_49871);
and UO_3130 (O_3130,N_46200,N_47066);
nand UO_3131 (O_3131,N_46330,N_49999);
nand UO_3132 (O_3132,N_48336,N_48450);
or UO_3133 (O_3133,N_48888,N_45925);
and UO_3134 (O_3134,N_47486,N_47769);
and UO_3135 (O_3135,N_49459,N_49833);
nand UO_3136 (O_3136,N_47721,N_48126);
nor UO_3137 (O_3137,N_45885,N_46024);
nor UO_3138 (O_3138,N_47142,N_47711);
xnor UO_3139 (O_3139,N_46775,N_47527);
nor UO_3140 (O_3140,N_49985,N_46724);
nor UO_3141 (O_3141,N_47870,N_45502);
or UO_3142 (O_3142,N_45423,N_47118);
and UO_3143 (O_3143,N_46993,N_46238);
and UO_3144 (O_3144,N_48739,N_46075);
or UO_3145 (O_3145,N_46728,N_46227);
or UO_3146 (O_3146,N_46926,N_45141);
xnor UO_3147 (O_3147,N_48319,N_46007);
and UO_3148 (O_3148,N_48922,N_48370);
and UO_3149 (O_3149,N_45374,N_45764);
and UO_3150 (O_3150,N_49136,N_47346);
xnor UO_3151 (O_3151,N_46699,N_48059);
xnor UO_3152 (O_3152,N_47777,N_48637);
nand UO_3153 (O_3153,N_47524,N_46889);
nor UO_3154 (O_3154,N_46436,N_45277);
nor UO_3155 (O_3155,N_48994,N_48840);
nor UO_3156 (O_3156,N_48360,N_47761);
and UO_3157 (O_3157,N_47535,N_49258);
xnor UO_3158 (O_3158,N_48180,N_46107);
or UO_3159 (O_3159,N_45561,N_45470);
nor UO_3160 (O_3160,N_48360,N_48539);
and UO_3161 (O_3161,N_47790,N_49954);
and UO_3162 (O_3162,N_48085,N_48402);
and UO_3163 (O_3163,N_49597,N_48849);
nand UO_3164 (O_3164,N_47129,N_45717);
nor UO_3165 (O_3165,N_46813,N_47921);
and UO_3166 (O_3166,N_47412,N_49331);
nand UO_3167 (O_3167,N_49090,N_49964);
nor UO_3168 (O_3168,N_46145,N_45851);
nor UO_3169 (O_3169,N_45815,N_48029);
and UO_3170 (O_3170,N_45369,N_49658);
and UO_3171 (O_3171,N_49598,N_49555);
xor UO_3172 (O_3172,N_48717,N_47158);
or UO_3173 (O_3173,N_48016,N_48937);
nor UO_3174 (O_3174,N_47297,N_45674);
xnor UO_3175 (O_3175,N_48084,N_49840);
xor UO_3176 (O_3176,N_45300,N_49282);
nor UO_3177 (O_3177,N_48149,N_48545);
xnor UO_3178 (O_3178,N_46173,N_49115);
nor UO_3179 (O_3179,N_45007,N_45762);
nand UO_3180 (O_3180,N_45412,N_46426);
and UO_3181 (O_3181,N_45218,N_47838);
nor UO_3182 (O_3182,N_47589,N_45012);
xnor UO_3183 (O_3183,N_47171,N_46258);
or UO_3184 (O_3184,N_48232,N_46457);
or UO_3185 (O_3185,N_48921,N_48009);
nor UO_3186 (O_3186,N_46041,N_49358);
nand UO_3187 (O_3187,N_49315,N_48436);
nor UO_3188 (O_3188,N_45747,N_49129);
nor UO_3189 (O_3189,N_46661,N_48519);
nand UO_3190 (O_3190,N_49422,N_46839);
and UO_3191 (O_3191,N_47417,N_45567);
or UO_3192 (O_3192,N_46191,N_49602);
nor UO_3193 (O_3193,N_46078,N_46805);
nand UO_3194 (O_3194,N_45536,N_45651);
or UO_3195 (O_3195,N_46971,N_49749);
or UO_3196 (O_3196,N_46523,N_49783);
or UO_3197 (O_3197,N_46740,N_47090);
nor UO_3198 (O_3198,N_46259,N_49298);
nor UO_3199 (O_3199,N_48575,N_48708);
or UO_3200 (O_3200,N_48772,N_47612);
or UO_3201 (O_3201,N_47127,N_46795);
nand UO_3202 (O_3202,N_45871,N_47759);
xnor UO_3203 (O_3203,N_46347,N_46912);
or UO_3204 (O_3204,N_48180,N_48116);
xnor UO_3205 (O_3205,N_45410,N_49852);
xnor UO_3206 (O_3206,N_46796,N_47853);
xnor UO_3207 (O_3207,N_46503,N_45652);
or UO_3208 (O_3208,N_49850,N_48931);
nand UO_3209 (O_3209,N_48924,N_46199);
nor UO_3210 (O_3210,N_46833,N_48251);
or UO_3211 (O_3211,N_46773,N_46061);
nor UO_3212 (O_3212,N_49481,N_45886);
and UO_3213 (O_3213,N_45435,N_46054);
xor UO_3214 (O_3214,N_46919,N_46230);
nand UO_3215 (O_3215,N_47995,N_47979);
nor UO_3216 (O_3216,N_46194,N_49067);
or UO_3217 (O_3217,N_45959,N_45334);
xnor UO_3218 (O_3218,N_48875,N_47481);
or UO_3219 (O_3219,N_49453,N_48780);
nor UO_3220 (O_3220,N_47295,N_49865);
or UO_3221 (O_3221,N_48552,N_46045);
xnor UO_3222 (O_3222,N_49625,N_48475);
xnor UO_3223 (O_3223,N_47328,N_45026);
nand UO_3224 (O_3224,N_46541,N_47857);
or UO_3225 (O_3225,N_48042,N_49585);
xor UO_3226 (O_3226,N_49615,N_49136);
nor UO_3227 (O_3227,N_46705,N_46848);
nand UO_3228 (O_3228,N_47459,N_47294);
xor UO_3229 (O_3229,N_45350,N_47012);
or UO_3230 (O_3230,N_46133,N_46561);
or UO_3231 (O_3231,N_46478,N_48539);
nand UO_3232 (O_3232,N_48842,N_49872);
nand UO_3233 (O_3233,N_47573,N_46911);
xor UO_3234 (O_3234,N_47518,N_48246);
or UO_3235 (O_3235,N_49620,N_45946);
nand UO_3236 (O_3236,N_46419,N_48287);
and UO_3237 (O_3237,N_48925,N_47923);
nand UO_3238 (O_3238,N_45114,N_49358);
xor UO_3239 (O_3239,N_49617,N_49214);
or UO_3240 (O_3240,N_49247,N_48585);
nor UO_3241 (O_3241,N_47172,N_47374);
nand UO_3242 (O_3242,N_48233,N_48487);
xor UO_3243 (O_3243,N_45898,N_47805);
and UO_3244 (O_3244,N_47312,N_47498);
and UO_3245 (O_3245,N_49613,N_45895);
xnor UO_3246 (O_3246,N_49581,N_49092);
and UO_3247 (O_3247,N_45923,N_49624);
or UO_3248 (O_3248,N_47839,N_45438);
xnor UO_3249 (O_3249,N_45378,N_48778);
xor UO_3250 (O_3250,N_48884,N_45978);
or UO_3251 (O_3251,N_48772,N_49004);
nor UO_3252 (O_3252,N_47414,N_47754);
and UO_3253 (O_3253,N_48056,N_46387);
nand UO_3254 (O_3254,N_47731,N_47060);
and UO_3255 (O_3255,N_48703,N_46089);
and UO_3256 (O_3256,N_46278,N_48799);
xnor UO_3257 (O_3257,N_47988,N_47220);
nor UO_3258 (O_3258,N_47269,N_45471);
nand UO_3259 (O_3259,N_48116,N_47587);
xnor UO_3260 (O_3260,N_49695,N_48926);
nor UO_3261 (O_3261,N_45942,N_45529);
xor UO_3262 (O_3262,N_45769,N_48927);
nor UO_3263 (O_3263,N_47049,N_47710);
xnor UO_3264 (O_3264,N_45943,N_49764);
nor UO_3265 (O_3265,N_49119,N_49758);
or UO_3266 (O_3266,N_47702,N_46465);
and UO_3267 (O_3267,N_46128,N_45831);
nand UO_3268 (O_3268,N_45966,N_48554);
nor UO_3269 (O_3269,N_45156,N_46499);
nand UO_3270 (O_3270,N_48459,N_49492);
or UO_3271 (O_3271,N_49789,N_48991);
nand UO_3272 (O_3272,N_49664,N_49191);
nand UO_3273 (O_3273,N_45281,N_49774);
nand UO_3274 (O_3274,N_46319,N_45985);
or UO_3275 (O_3275,N_45108,N_48029);
nand UO_3276 (O_3276,N_49944,N_45048);
or UO_3277 (O_3277,N_45965,N_46283);
and UO_3278 (O_3278,N_47416,N_49900);
nand UO_3279 (O_3279,N_49283,N_45041);
xnor UO_3280 (O_3280,N_48951,N_46698);
nand UO_3281 (O_3281,N_48906,N_47070);
nand UO_3282 (O_3282,N_49939,N_49690);
or UO_3283 (O_3283,N_46237,N_49616);
nor UO_3284 (O_3284,N_49514,N_49254);
and UO_3285 (O_3285,N_46264,N_49878);
and UO_3286 (O_3286,N_45446,N_49193);
or UO_3287 (O_3287,N_46897,N_49879);
or UO_3288 (O_3288,N_46571,N_49747);
nor UO_3289 (O_3289,N_49966,N_45258);
and UO_3290 (O_3290,N_47750,N_45846);
and UO_3291 (O_3291,N_46579,N_45780);
xor UO_3292 (O_3292,N_47935,N_46592);
and UO_3293 (O_3293,N_45252,N_45045);
nor UO_3294 (O_3294,N_46655,N_49942);
and UO_3295 (O_3295,N_49996,N_46766);
or UO_3296 (O_3296,N_49423,N_46356);
nand UO_3297 (O_3297,N_48869,N_47318);
nand UO_3298 (O_3298,N_49480,N_49566);
nor UO_3299 (O_3299,N_48467,N_48125);
and UO_3300 (O_3300,N_49315,N_48187);
and UO_3301 (O_3301,N_46567,N_49990);
or UO_3302 (O_3302,N_46577,N_46239);
xor UO_3303 (O_3303,N_46907,N_46606);
xor UO_3304 (O_3304,N_46752,N_45836);
or UO_3305 (O_3305,N_49216,N_48149);
or UO_3306 (O_3306,N_48284,N_48122);
xor UO_3307 (O_3307,N_45515,N_49625);
and UO_3308 (O_3308,N_46907,N_46883);
or UO_3309 (O_3309,N_49463,N_45465);
and UO_3310 (O_3310,N_46339,N_45603);
and UO_3311 (O_3311,N_45842,N_49291);
or UO_3312 (O_3312,N_48182,N_45904);
and UO_3313 (O_3313,N_46598,N_48713);
and UO_3314 (O_3314,N_47171,N_46787);
and UO_3315 (O_3315,N_47081,N_48196);
and UO_3316 (O_3316,N_46527,N_47415);
xor UO_3317 (O_3317,N_47125,N_48849);
nand UO_3318 (O_3318,N_46824,N_48871);
nor UO_3319 (O_3319,N_46538,N_46518);
or UO_3320 (O_3320,N_48939,N_47074);
and UO_3321 (O_3321,N_45372,N_48787);
nor UO_3322 (O_3322,N_46653,N_47599);
nor UO_3323 (O_3323,N_47179,N_45958);
and UO_3324 (O_3324,N_49173,N_45521);
or UO_3325 (O_3325,N_47749,N_47563);
nand UO_3326 (O_3326,N_49109,N_49747);
nor UO_3327 (O_3327,N_47194,N_48778);
xnor UO_3328 (O_3328,N_49261,N_48796);
nand UO_3329 (O_3329,N_49329,N_47619);
nor UO_3330 (O_3330,N_45541,N_47381);
nor UO_3331 (O_3331,N_45005,N_46025);
xnor UO_3332 (O_3332,N_45735,N_48718);
xor UO_3333 (O_3333,N_49139,N_48703);
or UO_3334 (O_3334,N_46772,N_49178);
and UO_3335 (O_3335,N_45050,N_49658);
or UO_3336 (O_3336,N_48048,N_48785);
nand UO_3337 (O_3337,N_47772,N_45571);
and UO_3338 (O_3338,N_48786,N_49240);
nor UO_3339 (O_3339,N_46758,N_46221);
xnor UO_3340 (O_3340,N_49858,N_47299);
xor UO_3341 (O_3341,N_47411,N_46117);
nand UO_3342 (O_3342,N_48016,N_48439);
xnor UO_3343 (O_3343,N_49595,N_46974);
nand UO_3344 (O_3344,N_48483,N_49441);
nand UO_3345 (O_3345,N_45366,N_45514);
nor UO_3346 (O_3346,N_47284,N_48393);
nand UO_3347 (O_3347,N_45163,N_46803);
nor UO_3348 (O_3348,N_48101,N_45663);
nand UO_3349 (O_3349,N_49462,N_49697);
and UO_3350 (O_3350,N_46259,N_48548);
or UO_3351 (O_3351,N_47418,N_45311);
or UO_3352 (O_3352,N_48764,N_46946);
or UO_3353 (O_3353,N_45287,N_49088);
nor UO_3354 (O_3354,N_46429,N_47455);
nand UO_3355 (O_3355,N_48241,N_46339);
xnor UO_3356 (O_3356,N_45758,N_48599);
and UO_3357 (O_3357,N_46057,N_47720);
or UO_3358 (O_3358,N_47982,N_47849);
nor UO_3359 (O_3359,N_49424,N_46383);
and UO_3360 (O_3360,N_48508,N_46211);
xnor UO_3361 (O_3361,N_47260,N_47208);
and UO_3362 (O_3362,N_49597,N_45626);
and UO_3363 (O_3363,N_47656,N_46271);
xor UO_3364 (O_3364,N_47974,N_49316);
or UO_3365 (O_3365,N_46522,N_49801);
xor UO_3366 (O_3366,N_47095,N_47447);
xor UO_3367 (O_3367,N_46972,N_49376);
nor UO_3368 (O_3368,N_45059,N_46531);
and UO_3369 (O_3369,N_45881,N_46836);
xor UO_3370 (O_3370,N_49993,N_48371);
or UO_3371 (O_3371,N_45767,N_45977);
nor UO_3372 (O_3372,N_45776,N_47624);
nor UO_3373 (O_3373,N_48122,N_45248);
xnor UO_3374 (O_3374,N_46755,N_49328);
xnor UO_3375 (O_3375,N_47576,N_45973);
nand UO_3376 (O_3376,N_48041,N_47120);
or UO_3377 (O_3377,N_49871,N_46876);
xnor UO_3378 (O_3378,N_46862,N_47606);
nor UO_3379 (O_3379,N_48064,N_46018);
and UO_3380 (O_3380,N_49731,N_46785);
nor UO_3381 (O_3381,N_47243,N_49033);
xor UO_3382 (O_3382,N_49125,N_46953);
xnor UO_3383 (O_3383,N_45371,N_46947);
nand UO_3384 (O_3384,N_49430,N_46247);
nor UO_3385 (O_3385,N_47056,N_47028);
and UO_3386 (O_3386,N_47641,N_48404);
and UO_3387 (O_3387,N_47291,N_49612);
nand UO_3388 (O_3388,N_49330,N_49375);
nand UO_3389 (O_3389,N_49184,N_46889);
or UO_3390 (O_3390,N_49076,N_47693);
xnor UO_3391 (O_3391,N_49393,N_49500);
xnor UO_3392 (O_3392,N_48158,N_45435);
nor UO_3393 (O_3393,N_47955,N_49404);
nand UO_3394 (O_3394,N_49713,N_46237);
nand UO_3395 (O_3395,N_45813,N_45676);
nand UO_3396 (O_3396,N_46779,N_46605);
xor UO_3397 (O_3397,N_45247,N_48194);
nor UO_3398 (O_3398,N_45513,N_45011);
xor UO_3399 (O_3399,N_46200,N_46392);
nand UO_3400 (O_3400,N_48800,N_47729);
nand UO_3401 (O_3401,N_48286,N_45733);
nand UO_3402 (O_3402,N_47939,N_46126);
xnor UO_3403 (O_3403,N_47008,N_48584);
and UO_3404 (O_3404,N_46764,N_48927);
xnor UO_3405 (O_3405,N_49105,N_47863);
nand UO_3406 (O_3406,N_45739,N_48239);
nor UO_3407 (O_3407,N_46717,N_47245);
xnor UO_3408 (O_3408,N_46171,N_46814);
and UO_3409 (O_3409,N_46460,N_47223);
nor UO_3410 (O_3410,N_45745,N_46331);
xor UO_3411 (O_3411,N_49333,N_47608);
and UO_3412 (O_3412,N_48889,N_49085);
xnor UO_3413 (O_3413,N_47155,N_45322);
xor UO_3414 (O_3414,N_47864,N_46338);
and UO_3415 (O_3415,N_45862,N_47593);
nand UO_3416 (O_3416,N_48405,N_49913);
or UO_3417 (O_3417,N_49404,N_49106);
nand UO_3418 (O_3418,N_47460,N_48592);
xor UO_3419 (O_3419,N_49816,N_45716);
and UO_3420 (O_3420,N_48266,N_47113);
nand UO_3421 (O_3421,N_48574,N_45327);
and UO_3422 (O_3422,N_45776,N_45701);
nand UO_3423 (O_3423,N_48186,N_47772);
or UO_3424 (O_3424,N_45356,N_45361);
and UO_3425 (O_3425,N_47938,N_47661);
and UO_3426 (O_3426,N_45879,N_49395);
nor UO_3427 (O_3427,N_47611,N_49294);
and UO_3428 (O_3428,N_46569,N_47106);
nor UO_3429 (O_3429,N_48980,N_47435);
or UO_3430 (O_3430,N_48569,N_48709);
xnor UO_3431 (O_3431,N_46068,N_45559);
and UO_3432 (O_3432,N_46607,N_49485);
and UO_3433 (O_3433,N_45573,N_45501);
or UO_3434 (O_3434,N_48664,N_48034);
or UO_3435 (O_3435,N_45255,N_46698);
nand UO_3436 (O_3436,N_46077,N_46744);
or UO_3437 (O_3437,N_45732,N_47290);
or UO_3438 (O_3438,N_49683,N_49743);
or UO_3439 (O_3439,N_46509,N_49535);
and UO_3440 (O_3440,N_47464,N_45323);
and UO_3441 (O_3441,N_46670,N_47207);
nor UO_3442 (O_3442,N_48868,N_45874);
or UO_3443 (O_3443,N_45992,N_47486);
nor UO_3444 (O_3444,N_48258,N_47518);
xor UO_3445 (O_3445,N_46216,N_47087);
xnor UO_3446 (O_3446,N_47887,N_45997);
and UO_3447 (O_3447,N_49894,N_45837);
nor UO_3448 (O_3448,N_46376,N_48351);
or UO_3449 (O_3449,N_47852,N_45729);
xnor UO_3450 (O_3450,N_47736,N_48417);
xor UO_3451 (O_3451,N_49310,N_45050);
xnor UO_3452 (O_3452,N_47397,N_47708);
or UO_3453 (O_3453,N_49334,N_48919);
or UO_3454 (O_3454,N_45819,N_49253);
nand UO_3455 (O_3455,N_45274,N_47265);
nand UO_3456 (O_3456,N_47622,N_46484);
nor UO_3457 (O_3457,N_48511,N_47106);
nor UO_3458 (O_3458,N_47069,N_45355);
nand UO_3459 (O_3459,N_45427,N_48393);
nor UO_3460 (O_3460,N_47880,N_49308);
nor UO_3461 (O_3461,N_45744,N_46807);
nor UO_3462 (O_3462,N_46614,N_49447);
nand UO_3463 (O_3463,N_49839,N_49323);
and UO_3464 (O_3464,N_49397,N_49567);
nor UO_3465 (O_3465,N_47036,N_49774);
nand UO_3466 (O_3466,N_45263,N_46432);
or UO_3467 (O_3467,N_46721,N_45190);
nor UO_3468 (O_3468,N_48223,N_47105);
or UO_3469 (O_3469,N_47622,N_49880);
or UO_3470 (O_3470,N_49075,N_49679);
or UO_3471 (O_3471,N_46172,N_48795);
and UO_3472 (O_3472,N_47042,N_49981);
xor UO_3473 (O_3473,N_49400,N_47962);
and UO_3474 (O_3474,N_45716,N_47399);
nand UO_3475 (O_3475,N_47127,N_46401);
nand UO_3476 (O_3476,N_46832,N_46863);
and UO_3477 (O_3477,N_45916,N_48191);
nor UO_3478 (O_3478,N_46890,N_47198);
nor UO_3479 (O_3479,N_47014,N_46277);
or UO_3480 (O_3480,N_47481,N_46391);
and UO_3481 (O_3481,N_47784,N_46330);
xnor UO_3482 (O_3482,N_49666,N_49845);
or UO_3483 (O_3483,N_47382,N_46227);
xnor UO_3484 (O_3484,N_48356,N_49614);
or UO_3485 (O_3485,N_45571,N_45530);
or UO_3486 (O_3486,N_48580,N_45982);
or UO_3487 (O_3487,N_48606,N_46033);
nor UO_3488 (O_3488,N_46341,N_48963);
nor UO_3489 (O_3489,N_49928,N_46700);
nand UO_3490 (O_3490,N_48419,N_48155);
and UO_3491 (O_3491,N_45261,N_47073);
xor UO_3492 (O_3492,N_46862,N_46701);
nand UO_3493 (O_3493,N_49159,N_47934);
nand UO_3494 (O_3494,N_45423,N_45242);
or UO_3495 (O_3495,N_49386,N_48469);
xnor UO_3496 (O_3496,N_48887,N_49199);
nand UO_3497 (O_3497,N_46000,N_49561);
or UO_3498 (O_3498,N_45784,N_48303);
xor UO_3499 (O_3499,N_48014,N_49469);
and UO_3500 (O_3500,N_46802,N_45220);
and UO_3501 (O_3501,N_47426,N_49430);
nand UO_3502 (O_3502,N_45165,N_49865);
xor UO_3503 (O_3503,N_49198,N_47202);
and UO_3504 (O_3504,N_48605,N_47748);
nor UO_3505 (O_3505,N_46099,N_45771);
nor UO_3506 (O_3506,N_45649,N_47559);
or UO_3507 (O_3507,N_45807,N_45593);
xor UO_3508 (O_3508,N_49344,N_46223);
and UO_3509 (O_3509,N_46805,N_46112);
xnor UO_3510 (O_3510,N_47858,N_48836);
nor UO_3511 (O_3511,N_47638,N_48171);
or UO_3512 (O_3512,N_49241,N_46743);
nand UO_3513 (O_3513,N_48942,N_48897);
nor UO_3514 (O_3514,N_45453,N_47211);
nor UO_3515 (O_3515,N_45302,N_45619);
or UO_3516 (O_3516,N_49643,N_48217);
or UO_3517 (O_3517,N_45151,N_45410);
or UO_3518 (O_3518,N_47465,N_49144);
xnor UO_3519 (O_3519,N_49426,N_49875);
xor UO_3520 (O_3520,N_49336,N_49820);
xor UO_3521 (O_3521,N_49628,N_45395);
nand UO_3522 (O_3522,N_45868,N_45874);
nand UO_3523 (O_3523,N_46550,N_47371);
nand UO_3524 (O_3524,N_48622,N_49999);
and UO_3525 (O_3525,N_49962,N_45050);
and UO_3526 (O_3526,N_47322,N_49853);
nand UO_3527 (O_3527,N_45241,N_49467);
or UO_3528 (O_3528,N_48829,N_45305);
nand UO_3529 (O_3529,N_45035,N_47384);
or UO_3530 (O_3530,N_46115,N_48625);
nor UO_3531 (O_3531,N_46337,N_49280);
nand UO_3532 (O_3532,N_45919,N_49212);
or UO_3533 (O_3533,N_46626,N_48203);
nor UO_3534 (O_3534,N_48701,N_49978);
nor UO_3535 (O_3535,N_46230,N_46611);
xnor UO_3536 (O_3536,N_48259,N_48012);
nor UO_3537 (O_3537,N_47386,N_46915);
nand UO_3538 (O_3538,N_49226,N_45901);
and UO_3539 (O_3539,N_45092,N_49616);
nand UO_3540 (O_3540,N_47040,N_48725);
nor UO_3541 (O_3541,N_47704,N_45227);
nor UO_3542 (O_3542,N_48528,N_48263);
nand UO_3543 (O_3543,N_45159,N_49681);
or UO_3544 (O_3544,N_45107,N_47913);
nand UO_3545 (O_3545,N_47257,N_47302);
and UO_3546 (O_3546,N_49410,N_47371);
and UO_3547 (O_3547,N_48053,N_48132);
xnor UO_3548 (O_3548,N_45128,N_49518);
or UO_3549 (O_3549,N_46436,N_47864);
or UO_3550 (O_3550,N_48331,N_45074);
and UO_3551 (O_3551,N_47016,N_49228);
nor UO_3552 (O_3552,N_49667,N_49682);
nand UO_3553 (O_3553,N_47501,N_48298);
and UO_3554 (O_3554,N_46497,N_48663);
nor UO_3555 (O_3555,N_49955,N_45081);
or UO_3556 (O_3556,N_46500,N_46680);
nor UO_3557 (O_3557,N_47629,N_45112);
nor UO_3558 (O_3558,N_48093,N_46026);
and UO_3559 (O_3559,N_45420,N_45343);
nor UO_3560 (O_3560,N_47379,N_48277);
nand UO_3561 (O_3561,N_47914,N_45734);
nor UO_3562 (O_3562,N_47192,N_49729);
nand UO_3563 (O_3563,N_47939,N_49193);
and UO_3564 (O_3564,N_47721,N_46850);
and UO_3565 (O_3565,N_48463,N_45371);
xnor UO_3566 (O_3566,N_46711,N_47275);
and UO_3567 (O_3567,N_48747,N_46108);
and UO_3568 (O_3568,N_49454,N_45959);
xor UO_3569 (O_3569,N_46479,N_49963);
nor UO_3570 (O_3570,N_45993,N_45706);
xnor UO_3571 (O_3571,N_48763,N_47383);
nor UO_3572 (O_3572,N_49770,N_47789);
nand UO_3573 (O_3573,N_48059,N_49719);
or UO_3574 (O_3574,N_47256,N_46518);
nor UO_3575 (O_3575,N_48982,N_47249);
xnor UO_3576 (O_3576,N_47104,N_48232);
nor UO_3577 (O_3577,N_49741,N_48825);
and UO_3578 (O_3578,N_45264,N_49972);
or UO_3579 (O_3579,N_47675,N_45579);
and UO_3580 (O_3580,N_46607,N_48596);
and UO_3581 (O_3581,N_47815,N_47880);
nor UO_3582 (O_3582,N_45604,N_47629);
nor UO_3583 (O_3583,N_46333,N_46706);
nor UO_3584 (O_3584,N_48845,N_46068);
nand UO_3585 (O_3585,N_46425,N_46630);
and UO_3586 (O_3586,N_45787,N_45199);
and UO_3587 (O_3587,N_48698,N_46581);
nor UO_3588 (O_3588,N_48014,N_48755);
nand UO_3589 (O_3589,N_48634,N_47294);
or UO_3590 (O_3590,N_46018,N_49105);
nand UO_3591 (O_3591,N_49911,N_46200);
nor UO_3592 (O_3592,N_49232,N_47355);
or UO_3593 (O_3593,N_47407,N_48145);
or UO_3594 (O_3594,N_45149,N_47726);
xor UO_3595 (O_3595,N_46345,N_45485);
nand UO_3596 (O_3596,N_47345,N_46875);
or UO_3597 (O_3597,N_45996,N_45260);
and UO_3598 (O_3598,N_49310,N_47710);
nor UO_3599 (O_3599,N_47672,N_47948);
nor UO_3600 (O_3600,N_45990,N_45543);
xnor UO_3601 (O_3601,N_45817,N_46789);
and UO_3602 (O_3602,N_47273,N_45191);
nand UO_3603 (O_3603,N_49354,N_48058);
nand UO_3604 (O_3604,N_47518,N_47047);
nand UO_3605 (O_3605,N_45094,N_45002);
or UO_3606 (O_3606,N_47157,N_47286);
or UO_3607 (O_3607,N_45795,N_45841);
nor UO_3608 (O_3608,N_47267,N_47994);
nand UO_3609 (O_3609,N_46642,N_45892);
nand UO_3610 (O_3610,N_48015,N_45590);
nand UO_3611 (O_3611,N_45080,N_45486);
or UO_3612 (O_3612,N_46796,N_47678);
and UO_3613 (O_3613,N_49776,N_45845);
xnor UO_3614 (O_3614,N_47212,N_47967);
nor UO_3615 (O_3615,N_45508,N_46695);
xnor UO_3616 (O_3616,N_49144,N_48419);
or UO_3617 (O_3617,N_48529,N_46585);
and UO_3618 (O_3618,N_45882,N_49013);
nor UO_3619 (O_3619,N_48007,N_49819);
nor UO_3620 (O_3620,N_49057,N_48660);
or UO_3621 (O_3621,N_46283,N_49073);
nand UO_3622 (O_3622,N_47926,N_49117);
and UO_3623 (O_3623,N_45790,N_48626);
nand UO_3624 (O_3624,N_49883,N_46538);
or UO_3625 (O_3625,N_46697,N_48298);
xnor UO_3626 (O_3626,N_45615,N_48648);
nor UO_3627 (O_3627,N_49411,N_45048);
or UO_3628 (O_3628,N_47706,N_46196);
nor UO_3629 (O_3629,N_47169,N_45027);
or UO_3630 (O_3630,N_46867,N_45721);
and UO_3631 (O_3631,N_49311,N_46542);
nand UO_3632 (O_3632,N_46655,N_46452);
and UO_3633 (O_3633,N_46513,N_48103);
and UO_3634 (O_3634,N_48290,N_48030);
and UO_3635 (O_3635,N_45039,N_46709);
nor UO_3636 (O_3636,N_48072,N_48838);
or UO_3637 (O_3637,N_46482,N_49857);
xnor UO_3638 (O_3638,N_45503,N_45249);
and UO_3639 (O_3639,N_47836,N_46505);
or UO_3640 (O_3640,N_48127,N_48438);
xnor UO_3641 (O_3641,N_45961,N_46573);
and UO_3642 (O_3642,N_47213,N_49416);
xnor UO_3643 (O_3643,N_45109,N_45986);
xor UO_3644 (O_3644,N_48501,N_49829);
and UO_3645 (O_3645,N_48167,N_45261);
and UO_3646 (O_3646,N_45664,N_49849);
xnor UO_3647 (O_3647,N_46710,N_49193);
nor UO_3648 (O_3648,N_48522,N_45401);
nand UO_3649 (O_3649,N_47811,N_49106);
nor UO_3650 (O_3650,N_48132,N_46780);
xnor UO_3651 (O_3651,N_48823,N_46005);
and UO_3652 (O_3652,N_45940,N_48186);
and UO_3653 (O_3653,N_49277,N_47391);
or UO_3654 (O_3654,N_48462,N_48030);
and UO_3655 (O_3655,N_48381,N_48158);
nand UO_3656 (O_3656,N_45374,N_48155);
and UO_3657 (O_3657,N_45563,N_45307);
nand UO_3658 (O_3658,N_45800,N_48537);
nand UO_3659 (O_3659,N_47750,N_48408);
nand UO_3660 (O_3660,N_49163,N_45070);
nand UO_3661 (O_3661,N_46096,N_46147);
xnor UO_3662 (O_3662,N_49235,N_46262);
xor UO_3663 (O_3663,N_49552,N_48639);
xnor UO_3664 (O_3664,N_49540,N_45304);
nand UO_3665 (O_3665,N_47208,N_45093);
nor UO_3666 (O_3666,N_48585,N_47581);
xnor UO_3667 (O_3667,N_47112,N_49841);
xnor UO_3668 (O_3668,N_47076,N_45586);
and UO_3669 (O_3669,N_45246,N_47817);
nor UO_3670 (O_3670,N_46836,N_46743);
nor UO_3671 (O_3671,N_45762,N_45765);
or UO_3672 (O_3672,N_45240,N_45311);
nor UO_3673 (O_3673,N_45996,N_49665);
or UO_3674 (O_3674,N_45992,N_47676);
nor UO_3675 (O_3675,N_47831,N_46846);
nand UO_3676 (O_3676,N_46927,N_45131);
nor UO_3677 (O_3677,N_46324,N_47606);
nand UO_3678 (O_3678,N_46723,N_48426);
nor UO_3679 (O_3679,N_48372,N_48444);
nor UO_3680 (O_3680,N_45784,N_48189);
nand UO_3681 (O_3681,N_48140,N_46552);
or UO_3682 (O_3682,N_45590,N_48972);
or UO_3683 (O_3683,N_49746,N_45671);
nand UO_3684 (O_3684,N_45691,N_48172);
xor UO_3685 (O_3685,N_49233,N_45846);
and UO_3686 (O_3686,N_47704,N_49954);
nand UO_3687 (O_3687,N_45140,N_47549);
xnor UO_3688 (O_3688,N_45658,N_49359);
and UO_3689 (O_3689,N_49731,N_46769);
and UO_3690 (O_3690,N_46926,N_49553);
xnor UO_3691 (O_3691,N_47887,N_46787);
and UO_3692 (O_3692,N_49150,N_49897);
or UO_3693 (O_3693,N_49026,N_46635);
nor UO_3694 (O_3694,N_49296,N_48341);
and UO_3695 (O_3695,N_46534,N_45421);
xnor UO_3696 (O_3696,N_48276,N_46915);
nor UO_3697 (O_3697,N_46361,N_48666);
nand UO_3698 (O_3698,N_46282,N_46098);
or UO_3699 (O_3699,N_45204,N_46586);
nand UO_3700 (O_3700,N_48640,N_46742);
or UO_3701 (O_3701,N_45049,N_46936);
xor UO_3702 (O_3702,N_49902,N_45116);
or UO_3703 (O_3703,N_48985,N_49460);
and UO_3704 (O_3704,N_48018,N_47595);
and UO_3705 (O_3705,N_48025,N_49373);
or UO_3706 (O_3706,N_47900,N_48986);
xor UO_3707 (O_3707,N_45168,N_48484);
nand UO_3708 (O_3708,N_49273,N_48620);
nand UO_3709 (O_3709,N_49971,N_45484);
and UO_3710 (O_3710,N_49492,N_47684);
xor UO_3711 (O_3711,N_45071,N_49057);
nand UO_3712 (O_3712,N_49539,N_46777);
nand UO_3713 (O_3713,N_46592,N_47188);
xor UO_3714 (O_3714,N_48713,N_45973);
xor UO_3715 (O_3715,N_48651,N_45335);
or UO_3716 (O_3716,N_48288,N_46713);
xnor UO_3717 (O_3717,N_49615,N_49596);
nor UO_3718 (O_3718,N_45089,N_49501);
nor UO_3719 (O_3719,N_48207,N_46202);
nand UO_3720 (O_3720,N_46909,N_47487);
or UO_3721 (O_3721,N_46423,N_47654);
nor UO_3722 (O_3722,N_48588,N_49194);
nor UO_3723 (O_3723,N_45261,N_46536);
xnor UO_3724 (O_3724,N_49916,N_49180);
nand UO_3725 (O_3725,N_49737,N_45273);
nor UO_3726 (O_3726,N_46997,N_47036);
nand UO_3727 (O_3727,N_46456,N_46264);
nor UO_3728 (O_3728,N_46822,N_45654);
or UO_3729 (O_3729,N_49052,N_46018);
nand UO_3730 (O_3730,N_48873,N_48668);
xor UO_3731 (O_3731,N_49674,N_45640);
nor UO_3732 (O_3732,N_45242,N_46440);
or UO_3733 (O_3733,N_46330,N_46250);
or UO_3734 (O_3734,N_46747,N_47019);
and UO_3735 (O_3735,N_45832,N_47880);
xor UO_3736 (O_3736,N_45466,N_45069);
or UO_3737 (O_3737,N_48109,N_47758);
or UO_3738 (O_3738,N_48518,N_45509);
xnor UO_3739 (O_3739,N_48072,N_47728);
nand UO_3740 (O_3740,N_48547,N_49031);
and UO_3741 (O_3741,N_47876,N_49014);
or UO_3742 (O_3742,N_47912,N_49120);
nor UO_3743 (O_3743,N_48538,N_47390);
and UO_3744 (O_3744,N_46334,N_49070);
nand UO_3745 (O_3745,N_46787,N_45106);
or UO_3746 (O_3746,N_45076,N_46864);
nand UO_3747 (O_3747,N_45031,N_48514);
or UO_3748 (O_3748,N_48114,N_48659);
and UO_3749 (O_3749,N_47618,N_48133);
and UO_3750 (O_3750,N_48202,N_48416);
xor UO_3751 (O_3751,N_49668,N_47954);
nand UO_3752 (O_3752,N_46507,N_46988);
xnor UO_3753 (O_3753,N_47961,N_46854);
nand UO_3754 (O_3754,N_48421,N_45909);
nor UO_3755 (O_3755,N_45857,N_45363);
and UO_3756 (O_3756,N_47598,N_46092);
nor UO_3757 (O_3757,N_48760,N_45667);
nand UO_3758 (O_3758,N_45161,N_49685);
nor UO_3759 (O_3759,N_48053,N_47052);
or UO_3760 (O_3760,N_45436,N_47906);
or UO_3761 (O_3761,N_45890,N_49740);
xor UO_3762 (O_3762,N_46499,N_46308);
and UO_3763 (O_3763,N_45192,N_47969);
xnor UO_3764 (O_3764,N_47456,N_47155);
nand UO_3765 (O_3765,N_47949,N_47163);
and UO_3766 (O_3766,N_49190,N_47707);
or UO_3767 (O_3767,N_49723,N_49935);
and UO_3768 (O_3768,N_45281,N_47643);
xnor UO_3769 (O_3769,N_45243,N_48103);
and UO_3770 (O_3770,N_46822,N_48753);
and UO_3771 (O_3771,N_47978,N_45674);
nand UO_3772 (O_3772,N_49073,N_47572);
nor UO_3773 (O_3773,N_47969,N_48452);
or UO_3774 (O_3774,N_49798,N_47317);
nand UO_3775 (O_3775,N_46100,N_45971);
or UO_3776 (O_3776,N_48936,N_47621);
xor UO_3777 (O_3777,N_45092,N_47464);
and UO_3778 (O_3778,N_49404,N_45788);
or UO_3779 (O_3779,N_45760,N_49131);
xor UO_3780 (O_3780,N_48564,N_48580);
nand UO_3781 (O_3781,N_47660,N_45127);
nand UO_3782 (O_3782,N_49395,N_46281);
xnor UO_3783 (O_3783,N_48553,N_49867);
xnor UO_3784 (O_3784,N_46050,N_47163);
and UO_3785 (O_3785,N_46499,N_45192);
and UO_3786 (O_3786,N_46313,N_46526);
or UO_3787 (O_3787,N_48052,N_48195);
nor UO_3788 (O_3788,N_46671,N_49645);
nor UO_3789 (O_3789,N_46420,N_49137);
or UO_3790 (O_3790,N_46156,N_49649);
and UO_3791 (O_3791,N_49345,N_49287);
nand UO_3792 (O_3792,N_45645,N_46204);
xor UO_3793 (O_3793,N_49024,N_46044);
nand UO_3794 (O_3794,N_46639,N_46545);
and UO_3795 (O_3795,N_47420,N_45599);
nand UO_3796 (O_3796,N_49605,N_46035);
xor UO_3797 (O_3797,N_46944,N_45131);
nand UO_3798 (O_3798,N_46357,N_49848);
and UO_3799 (O_3799,N_47488,N_45873);
xnor UO_3800 (O_3800,N_47068,N_48986);
nor UO_3801 (O_3801,N_48387,N_48622);
and UO_3802 (O_3802,N_47390,N_49935);
and UO_3803 (O_3803,N_45026,N_48884);
or UO_3804 (O_3804,N_49609,N_49976);
xor UO_3805 (O_3805,N_47887,N_45349);
xor UO_3806 (O_3806,N_48153,N_46764);
or UO_3807 (O_3807,N_45839,N_45905);
nor UO_3808 (O_3808,N_46723,N_49108);
and UO_3809 (O_3809,N_47954,N_48100);
and UO_3810 (O_3810,N_45297,N_48101);
and UO_3811 (O_3811,N_47671,N_48170);
xor UO_3812 (O_3812,N_47552,N_46443);
or UO_3813 (O_3813,N_45129,N_48591);
xnor UO_3814 (O_3814,N_46013,N_45509);
nor UO_3815 (O_3815,N_46797,N_46319);
nor UO_3816 (O_3816,N_45161,N_46521);
nand UO_3817 (O_3817,N_47726,N_47445);
nor UO_3818 (O_3818,N_47999,N_45425);
or UO_3819 (O_3819,N_49428,N_46160);
nand UO_3820 (O_3820,N_49206,N_49147);
nand UO_3821 (O_3821,N_46541,N_45307);
or UO_3822 (O_3822,N_49706,N_49577);
or UO_3823 (O_3823,N_49459,N_47382);
xnor UO_3824 (O_3824,N_46392,N_46734);
nor UO_3825 (O_3825,N_48577,N_47238);
nand UO_3826 (O_3826,N_47592,N_46427);
or UO_3827 (O_3827,N_48675,N_45299);
and UO_3828 (O_3828,N_45401,N_46764);
nor UO_3829 (O_3829,N_49700,N_45808);
and UO_3830 (O_3830,N_49035,N_49947);
and UO_3831 (O_3831,N_46191,N_46017);
xnor UO_3832 (O_3832,N_47038,N_45777);
or UO_3833 (O_3833,N_46482,N_49964);
or UO_3834 (O_3834,N_47255,N_46081);
nor UO_3835 (O_3835,N_45302,N_48811);
nor UO_3836 (O_3836,N_47608,N_49552);
and UO_3837 (O_3837,N_46182,N_47492);
nor UO_3838 (O_3838,N_46197,N_47354);
or UO_3839 (O_3839,N_47574,N_49202);
nand UO_3840 (O_3840,N_48339,N_46046);
nand UO_3841 (O_3841,N_48200,N_47831);
nor UO_3842 (O_3842,N_47594,N_46449);
nor UO_3843 (O_3843,N_45189,N_45082);
or UO_3844 (O_3844,N_47014,N_48213);
or UO_3845 (O_3845,N_49175,N_46124);
xor UO_3846 (O_3846,N_47665,N_45139);
and UO_3847 (O_3847,N_45130,N_46630);
nand UO_3848 (O_3848,N_47391,N_46294);
or UO_3849 (O_3849,N_47197,N_45969);
xnor UO_3850 (O_3850,N_47960,N_47794);
and UO_3851 (O_3851,N_46715,N_47853);
xor UO_3852 (O_3852,N_49541,N_49943);
or UO_3853 (O_3853,N_47366,N_46824);
and UO_3854 (O_3854,N_47654,N_47165);
nand UO_3855 (O_3855,N_49166,N_45561);
xnor UO_3856 (O_3856,N_47063,N_48183);
xnor UO_3857 (O_3857,N_48887,N_46721);
or UO_3858 (O_3858,N_46029,N_48243);
xor UO_3859 (O_3859,N_49015,N_47157);
and UO_3860 (O_3860,N_46976,N_46705);
nor UO_3861 (O_3861,N_48330,N_48407);
nor UO_3862 (O_3862,N_49222,N_47446);
nor UO_3863 (O_3863,N_45686,N_49463);
or UO_3864 (O_3864,N_45785,N_49750);
xnor UO_3865 (O_3865,N_47374,N_49881);
nand UO_3866 (O_3866,N_47106,N_45989);
or UO_3867 (O_3867,N_45654,N_45232);
or UO_3868 (O_3868,N_47562,N_47643);
nand UO_3869 (O_3869,N_49959,N_49604);
xor UO_3870 (O_3870,N_49137,N_45526);
and UO_3871 (O_3871,N_46691,N_49974);
nand UO_3872 (O_3872,N_45720,N_48765);
nand UO_3873 (O_3873,N_46269,N_48731);
nor UO_3874 (O_3874,N_47879,N_49798);
and UO_3875 (O_3875,N_49968,N_46758);
nand UO_3876 (O_3876,N_46115,N_45500);
xor UO_3877 (O_3877,N_47267,N_49614);
and UO_3878 (O_3878,N_45728,N_49389);
and UO_3879 (O_3879,N_49052,N_46201);
nand UO_3880 (O_3880,N_48201,N_47967);
xnor UO_3881 (O_3881,N_47659,N_49027);
xor UO_3882 (O_3882,N_49286,N_49599);
nor UO_3883 (O_3883,N_47766,N_46894);
xor UO_3884 (O_3884,N_47719,N_47155);
or UO_3885 (O_3885,N_49498,N_49967);
nor UO_3886 (O_3886,N_46325,N_48054);
nor UO_3887 (O_3887,N_48120,N_49098);
nand UO_3888 (O_3888,N_46431,N_48539);
xor UO_3889 (O_3889,N_48662,N_49432);
nor UO_3890 (O_3890,N_45642,N_49715);
or UO_3891 (O_3891,N_49126,N_46079);
and UO_3892 (O_3892,N_45022,N_47989);
xor UO_3893 (O_3893,N_47990,N_47523);
nor UO_3894 (O_3894,N_49893,N_47022);
nor UO_3895 (O_3895,N_46047,N_45621);
nor UO_3896 (O_3896,N_49287,N_48217);
nor UO_3897 (O_3897,N_48989,N_48156);
and UO_3898 (O_3898,N_45806,N_47804);
nor UO_3899 (O_3899,N_47639,N_46973);
nand UO_3900 (O_3900,N_49794,N_45919);
nor UO_3901 (O_3901,N_48700,N_45856);
xor UO_3902 (O_3902,N_46357,N_47613);
xnor UO_3903 (O_3903,N_49942,N_49269);
and UO_3904 (O_3904,N_49234,N_48039);
and UO_3905 (O_3905,N_45332,N_45319);
nand UO_3906 (O_3906,N_49852,N_49446);
and UO_3907 (O_3907,N_46977,N_45191);
or UO_3908 (O_3908,N_47795,N_48833);
or UO_3909 (O_3909,N_48187,N_45597);
xnor UO_3910 (O_3910,N_46697,N_48855);
nor UO_3911 (O_3911,N_46398,N_47186);
and UO_3912 (O_3912,N_46214,N_46929);
xor UO_3913 (O_3913,N_46965,N_47817);
xnor UO_3914 (O_3914,N_45398,N_48094);
and UO_3915 (O_3915,N_49601,N_48970);
nand UO_3916 (O_3916,N_45040,N_45481);
nor UO_3917 (O_3917,N_47424,N_49205);
or UO_3918 (O_3918,N_49787,N_48528);
nor UO_3919 (O_3919,N_46152,N_45335);
and UO_3920 (O_3920,N_48303,N_49495);
nand UO_3921 (O_3921,N_47068,N_49337);
or UO_3922 (O_3922,N_46855,N_49916);
nand UO_3923 (O_3923,N_48077,N_47733);
nand UO_3924 (O_3924,N_46830,N_49050);
or UO_3925 (O_3925,N_47769,N_46236);
nand UO_3926 (O_3926,N_45006,N_49681);
and UO_3927 (O_3927,N_45159,N_46677);
nor UO_3928 (O_3928,N_48771,N_45410);
nand UO_3929 (O_3929,N_49246,N_45831);
xor UO_3930 (O_3930,N_46928,N_49903);
nor UO_3931 (O_3931,N_49430,N_46958);
and UO_3932 (O_3932,N_49351,N_47014);
xnor UO_3933 (O_3933,N_45953,N_48448);
nor UO_3934 (O_3934,N_47796,N_47120);
xnor UO_3935 (O_3935,N_48068,N_45739);
xnor UO_3936 (O_3936,N_48168,N_45453);
nor UO_3937 (O_3937,N_49675,N_45170);
or UO_3938 (O_3938,N_49339,N_48359);
nand UO_3939 (O_3939,N_48466,N_48899);
or UO_3940 (O_3940,N_46568,N_45034);
xnor UO_3941 (O_3941,N_49975,N_47634);
xor UO_3942 (O_3942,N_46140,N_45386);
or UO_3943 (O_3943,N_49932,N_49239);
nor UO_3944 (O_3944,N_49905,N_49239);
nor UO_3945 (O_3945,N_48243,N_47225);
nand UO_3946 (O_3946,N_47862,N_45387);
or UO_3947 (O_3947,N_47511,N_47434);
xor UO_3948 (O_3948,N_47090,N_49218);
and UO_3949 (O_3949,N_47244,N_48897);
nor UO_3950 (O_3950,N_48545,N_48284);
or UO_3951 (O_3951,N_48698,N_48947);
or UO_3952 (O_3952,N_46404,N_48696);
or UO_3953 (O_3953,N_49864,N_46205);
or UO_3954 (O_3954,N_45282,N_46730);
and UO_3955 (O_3955,N_46079,N_45075);
xor UO_3956 (O_3956,N_48512,N_49895);
and UO_3957 (O_3957,N_47946,N_46218);
or UO_3958 (O_3958,N_48158,N_45809);
or UO_3959 (O_3959,N_45352,N_48067);
or UO_3960 (O_3960,N_49692,N_47413);
and UO_3961 (O_3961,N_49233,N_47483);
and UO_3962 (O_3962,N_45637,N_45994);
nor UO_3963 (O_3963,N_45370,N_45236);
nand UO_3964 (O_3964,N_45416,N_49154);
nand UO_3965 (O_3965,N_48105,N_48799);
nor UO_3966 (O_3966,N_49702,N_46274);
or UO_3967 (O_3967,N_47573,N_47748);
nand UO_3968 (O_3968,N_48431,N_47997);
and UO_3969 (O_3969,N_48011,N_49637);
xor UO_3970 (O_3970,N_45190,N_46737);
or UO_3971 (O_3971,N_47606,N_48711);
xor UO_3972 (O_3972,N_45285,N_47722);
nor UO_3973 (O_3973,N_48662,N_48005);
and UO_3974 (O_3974,N_47822,N_45577);
nor UO_3975 (O_3975,N_47077,N_48625);
xor UO_3976 (O_3976,N_46702,N_49083);
and UO_3977 (O_3977,N_48819,N_47189);
or UO_3978 (O_3978,N_47108,N_46771);
nand UO_3979 (O_3979,N_48239,N_48699);
xor UO_3980 (O_3980,N_49190,N_48419);
nor UO_3981 (O_3981,N_49654,N_46432);
or UO_3982 (O_3982,N_49513,N_48685);
xnor UO_3983 (O_3983,N_45983,N_47006);
xnor UO_3984 (O_3984,N_48651,N_49113);
or UO_3985 (O_3985,N_46153,N_49925);
nand UO_3986 (O_3986,N_47266,N_48372);
and UO_3987 (O_3987,N_46885,N_49056);
and UO_3988 (O_3988,N_49201,N_48921);
or UO_3989 (O_3989,N_48551,N_45408);
or UO_3990 (O_3990,N_46799,N_47024);
and UO_3991 (O_3991,N_46987,N_46931);
nor UO_3992 (O_3992,N_46965,N_49275);
nand UO_3993 (O_3993,N_48616,N_48150);
xor UO_3994 (O_3994,N_49026,N_46277);
nand UO_3995 (O_3995,N_45441,N_49438);
nand UO_3996 (O_3996,N_47471,N_48407);
nor UO_3997 (O_3997,N_48106,N_49894);
nand UO_3998 (O_3998,N_45147,N_48573);
or UO_3999 (O_3999,N_46740,N_48542);
xor UO_4000 (O_4000,N_47798,N_49824);
and UO_4001 (O_4001,N_46322,N_47912);
nand UO_4002 (O_4002,N_48908,N_45227);
nand UO_4003 (O_4003,N_48692,N_49032);
nor UO_4004 (O_4004,N_46652,N_46149);
and UO_4005 (O_4005,N_46415,N_47035);
nand UO_4006 (O_4006,N_49533,N_49610);
and UO_4007 (O_4007,N_49064,N_47097);
nor UO_4008 (O_4008,N_46197,N_45354);
nor UO_4009 (O_4009,N_49777,N_45715);
xor UO_4010 (O_4010,N_47824,N_47451);
and UO_4011 (O_4011,N_46693,N_47109);
and UO_4012 (O_4012,N_46685,N_47154);
nor UO_4013 (O_4013,N_45916,N_45934);
or UO_4014 (O_4014,N_45779,N_46740);
and UO_4015 (O_4015,N_47282,N_48102);
or UO_4016 (O_4016,N_45230,N_46845);
nand UO_4017 (O_4017,N_48737,N_46009);
xnor UO_4018 (O_4018,N_47812,N_45325);
and UO_4019 (O_4019,N_49115,N_45786);
nor UO_4020 (O_4020,N_47028,N_48415);
xnor UO_4021 (O_4021,N_46126,N_45552);
xnor UO_4022 (O_4022,N_47479,N_46010);
or UO_4023 (O_4023,N_45662,N_48837);
nor UO_4024 (O_4024,N_49645,N_49881);
nand UO_4025 (O_4025,N_49447,N_45150);
nor UO_4026 (O_4026,N_45775,N_48496);
nand UO_4027 (O_4027,N_47581,N_49956);
nor UO_4028 (O_4028,N_49703,N_47737);
nand UO_4029 (O_4029,N_46580,N_49181);
nand UO_4030 (O_4030,N_48422,N_47998);
and UO_4031 (O_4031,N_48279,N_46625);
and UO_4032 (O_4032,N_46177,N_45200);
and UO_4033 (O_4033,N_45084,N_45242);
xor UO_4034 (O_4034,N_49576,N_47417);
xnor UO_4035 (O_4035,N_48885,N_46481);
nand UO_4036 (O_4036,N_48196,N_49900);
nor UO_4037 (O_4037,N_45201,N_47471);
nor UO_4038 (O_4038,N_49418,N_46256);
nor UO_4039 (O_4039,N_46360,N_49975);
nand UO_4040 (O_4040,N_46843,N_47240);
xnor UO_4041 (O_4041,N_45940,N_48015);
or UO_4042 (O_4042,N_45588,N_45415);
nand UO_4043 (O_4043,N_49377,N_49726);
xor UO_4044 (O_4044,N_49240,N_49870);
nor UO_4045 (O_4045,N_47663,N_48248);
or UO_4046 (O_4046,N_46368,N_49630);
or UO_4047 (O_4047,N_47149,N_49298);
and UO_4048 (O_4048,N_49688,N_46959);
nor UO_4049 (O_4049,N_45269,N_45095);
xnor UO_4050 (O_4050,N_49883,N_48126);
or UO_4051 (O_4051,N_48937,N_48514);
or UO_4052 (O_4052,N_47567,N_48487);
nand UO_4053 (O_4053,N_45005,N_47473);
or UO_4054 (O_4054,N_47956,N_46876);
xor UO_4055 (O_4055,N_48611,N_48599);
nor UO_4056 (O_4056,N_48647,N_46838);
and UO_4057 (O_4057,N_47753,N_47400);
and UO_4058 (O_4058,N_49260,N_49813);
nand UO_4059 (O_4059,N_48306,N_49118);
or UO_4060 (O_4060,N_47588,N_49452);
and UO_4061 (O_4061,N_46781,N_45728);
nor UO_4062 (O_4062,N_48344,N_45934);
nor UO_4063 (O_4063,N_48917,N_48242);
xor UO_4064 (O_4064,N_48510,N_45731);
nor UO_4065 (O_4065,N_49858,N_47953);
nor UO_4066 (O_4066,N_45886,N_47120);
nand UO_4067 (O_4067,N_45042,N_45406);
or UO_4068 (O_4068,N_45481,N_49594);
nand UO_4069 (O_4069,N_45473,N_49132);
xor UO_4070 (O_4070,N_49321,N_46465);
nor UO_4071 (O_4071,N_48540,N_47398);
nand UO_4072 (O_4072,N_48639,N_45198);
xnor UO_4073 (O_4073,N_45546,N_45412);
nor UO_4074 (O_4074,N_46875,N_48286);
and UO_4075 (O_4075,N_48318,N_45732);
nor UO_4076 (O_4076,N_47779,N_46485);
xor UO_4077 (O_4077,N_48611,N_47353);
and UO_4078 (O_4078,N_46492,N_45241);
nor UO_4079 (O_4079,N_48984,N_47962);
nor UO_4080 (O_4080,N_46815,N_46672);
or UO_4081 (O_4081,N_47293,N_47971);
and UO_4082 (O_4082,N_48194,N_46396);
or UO_4083 (O_4083,N_48468,N_45972);
nor UO_4084 (O_4084,N_49763,N_46668);
xor UO_4085 (O_4085,N_49432,N_47910);
or UO_4086 (O_4086,N_46803,N_45066);
nand UO_4087 (O_4087,N_48198,N_46574);
nand UO_4088 (O_4088,N_48497,N_49830);
and UO_4089 (O_4089,N_46857,N_47279);
nand UO_4090 (O_4090,N_49385,N_45237);
and UO_4091 (O_4091,N_48113,N_47375);
or UO_4092 (O_4092,N_46845,N_49492);
nand UO_4093 (O_4093,N_45089,N_45234);
nand UO_4094 (O_4094,N_46842,N_49761);
or UO_4095 (O_4095,N_46101,N_49458);
and UO_4096 (O_4096,N_48117,N_46731);
and UO_4097 (O_4097,N_47366,N_48770);
or UO_4098 (O_4098,N_49226,N_46145);
and UO_4099 (O_4099,N_45575,N_46596);
or UO_4100 (O_4100,N_46754,N_45833);
or UO_4101 (O_4101,N_49127,N_48435);
nor UO_4102 (O_4102,N_48843,N_47006);
and UO_4103 (O_4103,N_48713,N_48275);
nand UO_4104 (O_4104,N_46034,N_47658);
or UO_4105 (O_4105,N_48347,N_45647);
nand UO_4106 (O_4106,N_45702,N_49180);
nand UO_4107 (O_4107,N_48491,N_45466);
nand UO_4108 (O_4108,N_46138,N_45740);
nor UO_4109 (O_4109,N_47437,N_49183);
nor UO_4110 (O_4110,N_46796,N_45815);
and UO_4111 (O_4111,N_48321,N_45996);
and UO_4112 (O_4112,N_47139,N_46315);
nand UO_4113 (O_4113,N_45171,N_48139);
nand UO_4114 (O_4114,N_45942,N_45901);
or UO_4115 (O_4115,N_45139,N_45896);
xor UO_4116 (O_4116,N_49736,N_46555);
or UO_4117 (O_4117,N_48179,N_48650);
or UO_4118 (O_4118,N_45172,N_48963);
or UO_4119 (O_4119,N_49900,N_48878);
and UO_4120 (O_4120,N_49692,N_49541);
nand UO_4121 (O_4121,N_45621,N_45323);
xnor UO_4122 (O_4122,N_48797,N_49956);
or UO_4123 (O_4123,N_45016,N_45067);
or UO_4124 (O_4124,N_46559,N_47991);
or UO_4125 (O_4125,N_46308,N_46893);
xor UO_4126 (O_4126,N_49094,N_47324);
and UO_4127 (O_4127,N_47357,N_45294);
xor UO_4128 (O_4128,N_48027,N_46109);
nand UO_4129 (O_4129,N_48176,N_45725);
xor UO_4130 (O_4130,N_48925,N_49476);
nor UO_4131 (O_4131,N_45065,N_49107);
nor UO_4132 (O_4132,N_46058,N_45091);
or UO_4133 (O_4133,N_46613,N_45519);
xnor UO_4134 (O_4134,N_46460,N_46372);
and UO_4135 (O_4135,N_49948,N_45459);
xor UO_4136 (O_4136,N_49762,N_45411);
nand UO_4137 (O_4137,N_46550,N_47564);
or UO_4138 (O_4138,N_48025,N_48120);
xor UO_4139 (O_4139,N_49755,N_48045);
nor UO_4140 (O_4140,N_48033,N_47219);
nand UO_4141 (O_4141,N_46479,N_48082);
xnor UO_4142 (O_4142,N_46612,N_49370);
and UO_4143 (O_4143,N_47723,N_47747);
or UO_4144 (O_4144,N_46934,N_47908);
xor UO_4145 (O_4145,N_48838,N_48609);
xnor UO_4146 (O_4146,N_45800,N_49332);
nor UO_4147 (O_4147,N_47623,N_47359);
nand UO_4148 (O_4148,N_48661,N_47686);
or UO_4149 (O_4149,N_46521,N_47173);
or UO_4150 (O_4150,N_46888,N_45172);
nand UO_4151 (O_4151,N_45358,N_48932);
and UO_4152 (O_4152,N_45042,N_46645);
xor UO_4153 (O_4153,N_47223,N_46738);
nand UO_4154 (O_4154,N_49816,N_48307);
and UO_4155 (O_4155,N_46245,N_45807);
nor UO_4156 (O_4156,N_45968,N_48564);
nand UO_4157 (O_4157,N_48612,N_49061);
or UO_4158 (O_4158,N_46605,N_48586);
or UO_4159 (O_4159,N_49002,N_48733);
nor UO_4160 (O_4160,N_49495,N_45624);
and UO_4161 (O_4161,N_49637,N_46272);
xnor UO_4162 (O_4162,N_47882,N_46728);
nor UO_4163 (O_4163,N_46474,N_45243);
nand UO_4164 (O_4164,N_48508,N_46192);
xnor UO_4165 (O_4165,N_45386,N_47324);
nand UO_4166 (O_4166,N_49245,N_49269);
and UO_4167 (O_4167,N_49182,N_47168);
or UO_4168 (O_4168,N_45661,N_46996);
nand UO_4169 (O_4169,N_48201,N_46807);
nor UO_4170 (O_4170,N_47246,N_46592);
and UO_4171 (O_4171,N_49545,N_49884);
and UO_4172 (O_4172,N_49181,N_49939);
nand UO_4173 (O_4173,N_48146,N_47893);
and UO_4174 (O_4174,N_45686,N_46833);
nand UO_4175 (O_4175,N_48640,N_46116);
and UO_4176 (O_4176,N_47547,N_48099);
xor UO_4177 (O_4177,N_48498,N_47340);
or UO_4178 (O_4178,N_47298,N_49826);
xnor UO_4179 (O_4179,N_46622,N_47789);
xor UO_4180 (O_4180,N_48078,N_49455);
nand UO_4181 (O_4181,N_45023,N_45413);
nand UO_4182 (O_4182,N_46375,N_49929);
and UO_4183 (O_4183,N_46476,N_49868);
or UO_4184 (O_4184,N_48162,N_49438);
nor UO_4185 (O_4185,N_47099,N_47224);
and UO_4186 (O_4186,N_49550,N_47880);
xor UO_4187 (O_4187,N_48359,N_46674);
xor UO_4188 (O_4188,N_48076,N_48363);
nand UO_4189 (O_4189,N_49072,N_47482);
nor UO_4190 (O_4190,N_47069,N_46689);
xnor UO_4191 (O_4191,N_46134,N_49400);
or UO_4192 (O_4192,N_48374,N_49188);
or UO_4193 (O_4193,N_45812,N_47207);
or UO_4194 (O_4194,N_49688,N_49355);
and UO_4195 (O_4195,N_47162,N_49872);
nor UO_4196 (O_4196,N_46746,N_49364);
and UO_4197 (O_4197,N_48536,N_45706);
nor UO_4198 (O_4198,N_49613,N_45878);
or UO_4199 (O_4199,N_45949,N_48000);
nor UO_4200 (O_4200,N_49460,N_49236);
or UO_4201 (O_4201,N_45241,N_48815);
nor UO_4202 (O_4202,N_45406,N_49732);
or UO_4203 (O_4203,N_49911,N_45727);
nand UO_4204 (O_4204,N_46344,N_45281);
nand UO_4205 (O_4205,N_45544,N_48949);
or UO_4206 (O_4206,N_45188,N_46895);
xor UO_4207 (O_4207,N_47163,N_46134);
xnor UO_4208 (O_4208,N_46283,N_46237);
or UO_4209 (O_4209,N_45632,N_48365);
or UO_4210 (O_4210,N_49736,N_45138);
or UO_4211 (O_4211,N_48510,N_45301);
and UO_4212 (O_4212,N_46191,N_46073);
nor UO_4213 (O_4213,N_45930,N_47347);
nand UO_4214 (O_4214,N_46594,N_46263);
and UO_4215 (O_4215,N_46398,N_47105);
nor UO_4216 (O_4216,N_46276,N_47484);
nor UO_4217 (O_4217,N_48893,N_46389);
xnor UO_4218 (O_4218,N_49843,N_47071);
nor UO_4219 (O_4219,N_48259,N_48573);
nor UO_4220 (O_4220,N_46023,N_47201);
and UO_4221 (O_4221,N_48329,N_48409);
nor UO_4222 (O_4222,N_47757,N_48153);
xor UO_4223 (O_4223,N_46799,N_47944);
and UO_4224 (O_4224,N_48291,N_49582);
nand UO_4225 (O_4225,N_46375,N_46886);
nor UO_4226 (O_4226,N_49356,N_48797);
xnor UO_4227 (O_4227,N_48857,N_45498);
nand UO_4228 (O_4228,N_47267,N_46579);
nor UO_4229 (O_4229,N_46430,N_49616);
xor UO_4230 (O_4230,N_49369,N_45317);
and UO_4231 (O_4231,N_46409,N_49455);
and UO_4232 (O_4232,N_45856,N_49339);
xnor UO_4233 (O_4233,N_47633,N_45838);
or UO_4234 (O_4234,N_49431,N_47386);
nand UO_4235 (O_4235,N_48721,N_46674);
or UO_4236 (O_4236,N_45736,N_47439);
and UO_4237 (O_4237,N_49450,N_47846);
xor UO_4238 (O_4238,N_49350,N_47678);
xor UO_4239 (O_4239,N_49120,N_45036);
nor UO_4240 (O_4240,N_46905,N_46818);
and UO_4241 (O_4241,N_49491,N_46148);
and UO_4242 (O_4242,N_47307,N_46900);
xor UO_4243 (O_4243,N_47752,N_49495);
nand UO_4244 (O_4244,N_45225,N_48029);
or UO_4245 (O_4245,N_45761,N_45599);
nor UO_4246 (O_4246,N_47457,N_46933);
nor UO_4247 (O_4247,N_47941,N_45312);
xor UO_4248 (O_4248,N_48094,N_48692);
or UO_4249 (O_4249,N_48283,N_46560);
and UO_4250 (O_4250,N_47428,N_48231);
and UO_4251 (O_4251,N_49039,N_47754);
nand UO_4252 (O_4252,N_48504,N_45639);
nand UO_4253 (O_4253,N_47142,N_46076);
nand UO_4254 (O_4254,N_46051,N_49699);
nor UO_4255 (O_4255,N_45485,N_49263);
xnor UO_4256 (O_4256,N_48926,N_46884);
or UO_4257 (O_4257,N_45100,N_46658);
nand UO_4258 (O_4258,N_46481,N_49209);
nor UO_4259 (O_4259,N_49617,N_45153);
xnor UO_4260 (O_4260,N_49128,N_48974);
nand UO_4261 (O_4261,N_47052,N_47311);
nor UO_4262 (O_4262,N_47162,N_45362);
xnor UO_4263 (O_4263,N_46901,N_46132);
xnor UO_4264 (O_4264,N_47136,N_45124);
nor UO_4265 (O_4265,N_46056,N_48470);
or UO_4266 (O_4266,N_46923,N_45476);
and UO_4267 (O_4267,N_46831,N_47709);
xor UO_4268 (O_4268,N_47643,N_46116);
and UO_4269 (O_4269,N_46928,N_49522);
and UO_4270 (O_4270,N_46710,N_49926);
and UO_4271 (O_4271,N_45085,N_48445);
xnor UO_4272 (O_4272,N_45678,N_45438);
and UO_4273 (O_4273,N_49001,N_48222);
nand UO_4274 (O_4274,N_46567,N_46919);
and UO_4275 (O_4275,N_49786,N_49292);
nor UO_4276 (O_4276,N_48907,N_48363);
or UO_4277 (O_4277,N_47135,N_47447);
or UO_4278 (O_4278,N_46056,N_49007);
or UO_4279 (O_4279,N_48259,N_45331);
and UO_4280 (O_4280,N_49220,N_48878);
nand UO_4281 (O_4281,N_47837,N_49567);
xnor UO_4282 (O_4282,N_46046,N_47839);
or UO_4283 (O_4283,N_47317,N_46091);
xor UO_4284 (O_4284,N_45015,N_45562);
nand UO_4285 (O_4285,N_48964,N_48473);
xnor UO_4286 (O_4286,N_48849,N_46765);
nor UO_4287 (O_4287,N_47785,N_46513);
or UO_4288 (O_4288,N_45345,N_47363);
or UO_4289 (O_4289,N_49627,N_49488);
and UO_4290 (O_4290,N_46761,N_48201);
xnor UO_4291 (O_4291,N_45410,N_45804);
nor UO_4292 (O_4292,N_48624,N_49853);
xor UO_4293 (O_4293,N_45806,N_48457);
xnor UO_4294 (O_4294,N_47159,N_46471);
nand UO_4295 (O_4295,N_48941,N_48958);
or UO_4296 (O_4296,N_45882,N_46462);
and UO_4297 (O_4297,N_46387,N_47712);
and UO_4298 (O_4298,N_45116,N_49833);
xor UO_4299 (O_4299,N_46880,N_49414);
nor UO_4300 (O_4300,N_48504,N_46709);
or UO_4301 (O_4301,N_46182,N_49200);
or UO_4302 (O_4302,N_45620,N_46823);
or UO_4303 (O_4303,N_47073,N_48151);
nand UO_4304 (O_4304,N_47919,N_46000);
or UO_4305 (O_4305,N_49539,N_49970);
and UO_4306 (O_4306,N_47077,N_48199);
xnor UO_4307 (O_4307,N_46236,N_45425);
nor UO_4308 (O_4308,N_49631,N_49594);
nor UO_4309 (O_4309,N_45188,N_46038);
xnor UO_4310 (O_4310,N_49971,N_47451);
and UO_4311 (O_4311,N_48960,N_49192);
or UO_4312 (O_4312,N_47473,N_46379);
nand UO_4313 (O_4313,N_47414,N_47596);
or UO_4314 (O_4314,N_47965,N_48859);
nor UO_4315 (O_4315,N_48980,N_46186);
nor UO_4316 (O_4316,N_47533,N_48569);
nand UO_4317 (O_4317,N_46332,N_48843);
xor UO_4318 (O_4318,N_47708,N_47630);
nor UO_4319 (O_4319,N_46254,N_45051);
nand UO_4320 (O_4320,N_45007,N_46418);
xor UO_4321 (O_4321,N_45847,N_47344);
nor UO_4322 (O_4322,N_46951,N_48201);
and UO_4323 (O_4323,N_48899,N_47456);
xnor UO_4324 (O_4324,N_49493,N_48319);
nor UO_4325 (O_4325,N_48005,N_46861);
and UO_4326 (O_4326,N_47524,N_47033);
nand UO_4327 (O_4327,N_45272,N_45785);
nor UO_4328 (O_4328,N_46269,N_45001);
nor UO_4329 (O_4329,N_46822,N_46763);
or UO_4330 (O_4330,N_46284,N_47158);
nand UO_4331 (O_4331,N_45906,N_49448);
xor UO_4332 (O_4332,N_45392,N_49203);
xnor UO_4333 (O_4333,N_49688,N_49481);
nand UO_4334 (O_4334,N_47900,N_48588);
xnor UO_4335 (O_4335,N_45338,N_47449);
or UO_4336 (O_4336,N_48288,N_48645);
nor UO_4337 (O_4337,N_49610,N_48413);
or UO_4338 (O_4338,N_48558,N_48625);
nand UO_4339 (O_4339,N_48145,N_47541);
nor UO_4340 (O_4340,N_46110,N_49257);
or UO_4341 (O_4341,N_46750,N_48860);
nand UO_4342 (O_4342,N_45015,N_49679);
nor UO_4343 (O_4343,N_47950,N_49903);
nand UO_4344 (O_4344,N_47066,N_45451);
xnor UO_4345 (O_4345,N_47513,N_46121);
nor UO_4346 (O_4346,N_49605,N_45481);
nand UO_4347 (O_4347,N_46476,N_47896);
nand UO_4348 (O_4348,N_49784,N_46831);
nor UO_4349 (O_4349,N_45993,N_48700);
nor UO_4350 (O_4350,N_48149,N_49407);
and UO_4351 (O_4351,N_45793,N_45596);
xnor UO_4352 (O_4352,N_47147,N_45192);
and UO_4353 (O_4353,N_47581,N_49290);
nor UO_4354 (O_4354,N_48750,N_48099);
xnor UO_4355 (O_4355,N_49087,N_48144);
and UO_4356 (O_4356,N_48960,N_46602);
xnor UO_4357 (O_4357,N_47963,N_45430);
or UO_4358 (O_4358,N_48679,N_46566);
nor UO_4359 (O_4359,N_46945,N_49021);
or UO_4360 (O_4360,N_48957,N_45266);
and UO_4361 (O_4361,N_45718,N_47330);
nor UO_4362 (O_4362,N_48736,N_46042);
xor UO_4363 (O_4363,N_48412,N_49562);
xnor UO_4364 (O_4364,N_48041,N_47510);
or UO_4365 (O_4365,N_45088,N_48552);
or UO_4366 (O_4366,N_45250,N_48455);
or UO_4367 (O_4367,N_45791,N_45654);
nor UO_4368 (O_4368,N_45451,N_48717);
nor UO_4369 (O_4369,N_49989,N_48064);
nand UO_4370 (O_4370,N_49778,N_49127);
nand UO_4371 (O_4371,N_46505,N_46084);
nand UO_4372 (O_4372,N_48745,N_48393);
nor UO_4373 (O_4373,N_45022,N_47323);
xor UO_4374 (O_4374,N_49287,N_46825);
nor UO_4375 (O_4375,N_45149,N_48560);
nand UO_4376 (O_4376,N_47991,N_47695);
xnor UO_4377 (O_4377,N_47431,N_49257);
nand UO_4378 (O_4378,N_48345,N_45668);
xor UO_4379 (O_4379,N_45199,N_46038);
or UO_4380 (O_4380,N_47557,N_46853);
nand UO_4381 (O_4381,N_47467,N_46699);
xor UO_4382 (O_4382,N_48160,N_46527);
or UO_4383 (O_4383,N_49939,N_48393);
nand UO_4384 (O_4384,N_48085,N_48247);
nand UO_4385 (O_4385,N_47814,N_46839);
xnor UO_4386 (O_4386,N_45578,N_45534);
nand UO_4387 (O_4387,N_49630,N_46736);
nor UO_4388 (O_4388,N_46463,N_45021);
or UO_4389 (O_4389,N_45533,N_49160);
and UO_4390 (O_4390,N_47664,N_45807);
nor UO_4391 (O_4391,N_46650,N_49074);
or UO_4392 (O_4392,N_47752,N_49857);
and UO_4393 (O_4393,N_46383,N_47302);
or UO_4394 (O_4394,N_46167,N_49034);
xor UO_4395 (O_4395,N_48158,N_47613);
or UO_4396 (O_4396,N_48606,N_45471);
nor UO_4397 (O_4397,N_47489,N_45470);
and UO_4398 (O_4398,N_48561,N_48839);
nand UO_4399 (O_4399,N_48738,N_46689);
or UO_4400 (O_4400,N_48556,N_47694);
xor UO_4401 (O_4401,N_45722,N_47587);
or UO_4402 (O_4402,N_46684,N_48532);
or UO_4403 (O_4403,N_45471,N_49843);
xnor UO_4404 (O_4404,N_49685,N_49686);
xnor UO_4405 (O_4405,N_46694,N_46734);
nor UO_4406 (O_4406,N_47965,N_48422);
xnor UO_4407 (O_4407,N_48790,N_49357);
nand UO_4408 (O_4408,N_47064,N_47525);
nor UO_4409 (O_4409,N_49939,N_45176);
nor UO_4410 (O_4410,N_49180,N_49247);
nor UO_4411 (O_4411,N_48620,N_48519);
nor UO_4412 (O_4412,N_46813,N_49775);
nand UO_4413 (O_4413,N_48911,N_45843);
xnor UO_4414 (O_4414,N_47919,N_49982);
and UO_4415 (O_4415,N_46011,N_45056);
nand UO_4416 (O_4416,N_45125,N_48669);
nor UO_4417 (O_4417,N_47792,N_48640);
and UO_4418 (O_4418,N_49767,N_49827);
and UO_4419 (O_4419,N_47635,N_47613);
nor UO_4420 (O_4420,N_45916,N_49567);
or UO_4421 (O_4421,N_49453,N_49297);
or UO_4422 (O_4422,N_46925,N_45398);
nor UO_4423 (O_4423,N_46493,N_49124);
nor UO_4424 (O_4424,N_45639,N_48716);
xnor UO_4425 (O_4425,N_48630,N_48983);
xor UO_4426 (O_4426,N_46813,N_45208);
and UO_4427 (O_4427,N_45412,N_49206);
and UO_4428 (O_4428,N_49445,N_47320);
nand UO_4429 (O_4429,N_47818,N_46430);
nor UO_4430 (O_4430,N_45167,N_47212);
or UO_4431 (O_4431,N_48567,N_45384);
and UO_4432 (O_4432,N_49135,N_47417);
nor UO_4433 (O_4433,N_49180,N_46987);
nor UO_4434 (O_4434,N_48788,N_46787);
xor UO_4435 (O_4435,N_49302,N_46074);
or UO_4436 (O_4436,N_45031,N_49008);
nor UO_4437 (O_4437,N_49860,N_48838);
nor UO_4438 (O_4438,N_47558,N_48178);
xnor UO_4439 (O_4439,N_46293,N_46645);
or UO_4440 (O_4440,N_45668,N_45825);
or UO_4441 (O_4441,N_46573,N_46609);
nand UO_4442 (O_4442,N_49368,N_46620);
or UO_4443 (O_4443,N_48677,N_47434);
xnor UO_4444 (O_4444,N_45899,N_48706);
nor UO_4445 (O_4445,N_46990,N_48143);
xnor UO_4446 (O_4446,N_48952,N_48651);
or UO_4447 (O_4447,N_49993,N_48068);
xnor UO_4448 (O_4448,N_46143,N_46509);
or UO_4449 (O_4449,N_47655,N_45124);
xor UO_4450 (O_4450,N_45469,N_46906);
nor UO_4451 (O_4451,N_46844,N_46351);
nand UO_4452 (O_4452,N_48992,N_46401);
or UO_4453 (O_4453,N_47506,N_48167);
and UO_4454 (O_4454,N_46025,N_45882);
nor UO_4455 (O_4455,N_45285,N_49357);
and UO_4456 (O_4456,N_46193,N_46085);
and UO_4457 (O_4457,N_46755,N_49928);
nand UO_4458 (O_4458,N_46096,N_47127);
and UO_4459 (O_4459,N_47985,N_45311);
xnor UO_4460 (O_4460,N_48229,N_49063);
xnor UO_4461 (O_4461,N_46653,N_45735);
xor UO_4462 (O_4462,N_48141,N_47728);
xnor UO_4463 (O_4463,N_48320,N_48512);
nor UO_4464 (O_4464,N_47893,N_46960);
or UO_4465 (O_4465,N_45079,N_48781);
nand UO_4466 (O_4466,N_47875,N_46756);
nor UO_4467 (O_4467,N_48656,N_45525);
nor UO_4468 (O_4468,N_46555,N_46206);
and UO_4469 (O_4469,N_48811,N_48350);
and UO_4470 (O_4470,N_47083,N_46871);
or UO_4471 (O_4471,N_49400,N_47653);
nand UO_4472 (O_4472,N_46812,N_45925);
or UO_4473 (O_4473,N_45641,N_49105);
or UO_4474 (O_4474,N_47688,N_48056);
nor UO_4475 (O_4475,N_48187,N_46516);
or UO_4476 (O_4476,N_49422,N_47276);
or UO_4477 (O_4477,N_46145,N_45907);
nand UO_4478 (O_4478,N_47583,N_45470);
xor UO_4479 (O_4479,N_49139,N_47960);
xnor UO_4480 (O_4480,N_45562,N_48894);
or UO_4481 (O_4481,N_45883,N_48673);
and UO_4482 (O_4482,N_48932,N_46152);
or UO_4483 (O_4483,N_45297,N_48354);
xor UO_4484 (O_4484,N_48717,N_46664);
or UO_4485 (O_4485,N_46461,N_49458);
or UO_4486 (O_4486,N_47955,N_49066);
xor UO_4487 (O_4487,N_46885,N_49482);
nand UO_4488 (O_4488,N_49847,N_49556);
nand UO_4489 (O_4489,N_46420,N_46095);
nor UO_4490 (O_4490,N_46746,N_46419);
and UO_4491 (O_4491,N_46468,N_49610);
and UO_4492 (O_4492,N_47881,N_49483);
xor UO_4493 (O_4493,N_49604,N_48813);
nand UO_4494 (O_4494,N_46927,N_47857);
and UO_4495 (O_4495,N_45337,N_49443);
xor UO_4496 (O_4496,N_47386,N_45233);
xor UO_4497 (O_4497,N_46399,N_47996);
and UO_4498 (O_4498,N_45890,N_45281);
and UO_4499 (O_4499,N_45991,N_47802);
xor UO_4500 (O_4500,N_49431,N_48945);
xor UO_4501 (O_4501,N_47137,N_49728);
or UO_4502 (O_4502,N_48748,N_46187);
and UO_4503 (O_4503,N_49566,N_46529);
or UO_4504 (O_4504,N_49128,N_46976);
or UO_4505 (O_4505,N_45907,N_48084);
or UO_4506 (O_4506,N_48996,N_48816);
nor UO_4507 (O_4507,N_49005,N_47823);
nor UO_4508 (O_4508,N_49088,N_46761);
and UO_4509 (O_4509,N_46920,N_45584);
or UO_4510 (O_4510,N_46023,N_46416);
and UO_4511 (O_4511,N_47038,N_49402);
nand UO_4512 (O_4512,N_48509,N_48926);
nor UO_4513 (O_4513,N_49649,N_47314);
or UO_4514 (O_4514,N_45516,N_46050);
xor UO_4515 (O_4515,N_47776,N_48549);
or UO_4516 (O_4516,N_48599,N_48628);
and UO_4517 (O_4517,N_47182,N_49701);
and UO_4518 (O_4518,N_48669,N_48980);
and UO_4519 (O_4519,N_46465,N_45914);
or UO_4520 (O_4520,N_48446,N_46887);
nor UO_4521 (O_4521,N_46664,N_48534);
nand UO_4522 (O_4522,N_46964,N_47268);
nand UO_4523 (O_4523,N_48832,N_45308);
and UO_4524 (O_4524,N_46317,N_48711);
nor UO_4525 (O_4525,N_48942,N_48796);
or UO_4526 (O_4526,N_46711,N_47633);
nand UO_4527 (O_4527,N_45632,N_46571);
nand UO_4528 (O_4528,N_47695,N_47677);
or UO_4529 (O_4529,N_47279,N_48260);
nand UO_4530 (O_4530,N_45543,N_49383);
nand UO_4531 (O_4531,N_47808,N_47217);
xnor UO_4532 (O_4532,N_48536,N_45439);
nor UO_4533 (O_4533,N_47017,N_49066);
nor UO_4534 (O_4534,N_48231,N_46263);
nor UO_4535 (O_4535,N_48687,N_47116);
xnor UO_4536 (O_4536,N_46970,N_47158);
and UO_4537 (O_4537,N_49051,N_48912);
xor UO_4538 (O_4538,N_48578,N_46080);
and UO_4539 (O_4539,N_47564,N_48844);
nor UO_4540 (O_4540,N_45341,N_45149);
nand UO_4541 (O_4541,N_47895,N_46158);
and UO_4542 (O_4542,N_45514,N_46886);
nand UO_4543 (O_4543,N_46439,N_49322);
or UO_4544 (O_4544,N_45593,N_45367);
and UO_4545 (O_4545,N_49332,N_46949);
and UO_4546 (O_4546,N_46911,N_48517);
and UO_4547 (O_4547,N_47441,N_46612);
nor UO_4548 (O_4548,N_47992,N_45400);
xnor UO_4549 (O_4549,N_48753,N_46594);
nand UO_4550 (O_4550,N_48053,N_48169);
and UO_4551 (O_4551,N_48853,N_47327);
or UO_4552 (O_4552,N_48297,N_49374);
nand UO_4553 (O_4553,N_48838,N_46468);
nand UO_4554 (O_4554,N_49608,N_48146);
and UO_4555 (O_4555,N_45675,N_47805);
xor UO_4556 (O_4556,N_46596,N_45700);
or UO_4557 (O_4557,N_47088,N_47738);
xor UO_4558 (O_4558,N_49034,N_46430);
nand UO_4559 (O_4559,N_45188,N_45339);
or UO_4560 (O_4560,N_47740,N_46480);
nor UO_4561 (O_4561,N_47301,N_45255);
and UO_4562 (O_4562,N_48329,N_48151);
nand UO_4563 (O_4563,N_48196,N_45255);
nor UO_4564 (O_4564,N_45822,N_47148);
nand UO_4565 (O_4565,N_48595,N_45676);
nor UO_4566 (O_4566,N_47253,N_46040);
and UO_4567 (O_4567,N_45996,N_45718);
nor UO_4568 (O_4568,N_45306,N_45018);
xor UO_4569 (O_4569,N_47629,N_47787);
nand UO_4570 (O_4570,N_49976,N_49890);
nand UO_4571 (O_4571,N_47074,N_49060);
or UO_4572 (O_4572,N_45683,N_49488);
nand UO_4573 (O_4573,N_45261,N_45444);
and UO_4574 (O_4574,N_48797,N_48413);
nand UO_4575 (O_4575,N_49745,N_45039);
and UO_4576 (O_4576,N_46984,N_45913);
nand UO_4577 (O_4577,N_48952,N_49927);
xnor UO_4578 (O_4578,N_45384,N_46057);
nor UO_4579 (O_4579,N_48919,N_47463);
xor UO_4580 (O_4580,N_48419,N_47265);
xnor UO_4581 (O_4581,N_46318,N_49283);
and UO_4582 (O_4582,N_49924,N_45873);
or UO_4583 (O_4583,N_47268,N_48504);
xnor UO_4584 (O_4584,N_47543,N_46955);
xor UO_4585 (O_4585,N_48172,N_47552);
nand UO_4586 (O_4586,N_47390,N_46476);
or UO_4587 (O_4587,N_45306,N_48214);
xnor UO_4588 (O_4588,N_48465,N_48846);
nor UO_4589 (O_4589,N_49547,N_47966);
or UO_4590 (O_4590,N_45585,N_49882);
xnor UO_4591 (O_4591,N_49887,N_46609);
and UO_4592 (O_4592,N_48615,N_47826);
nor UO_4593 (O_4593,N_48067,N_46828);
nor UO_4594 (O_4594,N_45108,N_46558);
or UO_4595 (O_4595,N_46248,N_47980);
or UO_4596 (O_4596,N_49161,N_49389);
nor UO_4597 (O_4597,N_47752,N_49986);
or UO_4598 (O_4598,N_49132,N_48356);
xnor UO_4599 (O_4599,N_45330,N_49971);
or UO_4600 (O_4600,N_47588,N_48539);
or UO_4601 (O_4601,N_46195,N_49569);
nor UO_4602 (O_4602,N_47082,N_48105);
nor UO_4603 (O_4603,N_49995,N_48116);
or UO_4604 (O_4604,N_48849,N_48896);
and UO_4605 (O_4605,N_49994,N_48389);
nand UO_4606 (O_4606,N_46852,N_48517);
and UO_4607 (O_4607,N_46856,N_46413);
and UO_4608 (O_4608,N_45548,N_48130);
and UO_4609 (O_4609,N_45052,N_47963);
and UO_4610 (O_4610,N_48224,N_46484);
nand UO_4611 (O_4611,N_46592,N_46972);
nor UO_4612 (O_4612,N_48444,N_47545);
or UO_4613 (O_4613,N_47132,N_48586);
or UO_4614 (O_4614,N_47248,N_49481);
nor UO_4615 (O_4615,N_49965,N_48906);
xor UO_4616 (O_4616,N_46656,N_49608);
or UO_4617 (O_4617,N_46244,N_47758);
nor UO_4618 (O_4618,N_47922,N_48977);
and UO_4619 (O_4619,N_46740,N_49095);
nor UO_4620 (O_4620,N_49798,N_45466);
xor UO_4621 (O_4621,N_46449,N_47569);
and UO_4622 (O_4622,N_48548,N_46763);
and UO_4623 (O_4623,N_47928,N_47361);
or UO_4624 (O_4624,N_47281,N_45542);
and UO_4625 (O_4625,N_47690,N_48391);
xnor UO_4626 (O_4626,N_47541,N_48376);
or UO_4627 (O_4627,N_46852,N_47517);
nor UO_4628 (O_4628,N_45409,N_46140);
nand UO_4629 (O_4629,N_49996,N_48487);
nand UO_4630 (O_4630,N_48582,N_45121);
and UO_4631 (O_4631,N_49477,N_47041);
xnor UO_4632 (O_4632,N_48488,N_48915);
and UO_4633 (O_4633,N_45185,N_47169);
nand UO_4634 (O_4634,N_48364,N_47301);
and UO_4635 (O_4635,N_46200,N_46793);
and UO_4636 (O_4636,N_49720,N_46027);
xnor UO_4637 (O_4637,N_49612,N_47417);
xor UO_4638 (O_4638,N_47319,N_49709);
nor UO_4639 (O_4639,N_47746,N_45592);
nand UO_4640 (O_4640,N_48752,N_48036);
or UO_4641 (O_4641,N_45178,N_49796);
xnor UO_4642 (O_4642,N_49043,N_49503);
nor UO_4643 (O_4643,N_45367,N_45555);
nand UO_4644 (O_4644,N_45753,N_48326);
nand UO_4645 (O_4645,N_48256,N_49558);
nand UO_4646 (O_4646,N_48248,N_48898);
nand UO_4647 (O_4647,N_48978,N_47792);
and UO_4648 (O_4648,N_46254,N_45934);
nor UO_4649 (O_4649,N_47356,N_49911);
or UO_4650 (O_4650,N_48731,N_47014);
xor UO_4651 (O_4651,N_49435,N_47705);
nand UO_4652 (O_4652,N_45680,N_46688);
xor UO_4653 (O_4653,N_48819,N_48939);
nand UO_4654 (O_4654,N_46581,N_46130);
and UO_4655 (O_4655,N_49085,N_47436);
xor UO_4656 (O_4656,N_46846,N_47832);
xnor UO_4657 (O_4657,N_46132,N_46731);
or UO_4658 (O_4658,N_47382,N_45515);
or UO_4659 (O_4659,N_48526,N_46518);
xor UO_4660 (O_4660,N_45018,N_48306);
or UO_4661 (O_4661,N_46324,N_48849);
nand UO_4662 (O_4662,N_48604,N_45434);
and UO_4663 (O_4663,N_47641,N_49625);
or UO_4664 (O_4664,N_47088,N_49020);
xor UO_4665 (O_4665,N_45516,N_45172);
or UO_4666 (O_4666,N_48731,N_45489);
nand UO_4667 (O_4667,N_49531,N_48624);
nor UO_4668 (O_4668,N_48556,N_49808);
and UO_4669 (O_4669,N_47798,N_45199);
and UO_4670 (O_4670,N_46399,N_47123);
nand UO_4671 (O_4671,N_49126,N_49124);
xnor UO_4672 (O_4672,N_49507,N_45471);
and UO_4673 (O_4673,N_47367,N_48223);
and UO_4674 (O_4674,N_47525,N_49581);
xor UO_4675 (O_4675,N_46526,N_47515);
and UO_4676 (O_4676,N_45773,N_47663);
or UO_4677 (O_4677,N_47933,N_46511);
and UO_4678 (O_4678,N_46122,N_46753);
nand UO_4679 (O_4679,N_48864,N_49668);
xnor UO_4680 (O_4680,N_48233,N_46884);
xnor UO_4681 (O_4681,N_46317,N_47361);
nor UO_4682 (O_4682,N_47150,N_48947);
and UO_4683 (O_4683,N_48461,N_49862);
or UO_4684 (O_4684,N_48870,N_46864);
and UO_4685 (O_4685,N_46934,N_48759);
xor UO_4686 (O_4686,N_47277,N_45116);
xnor UO_4687 (O_4687,N_45106,N_48586);
nor UO_4688 (O_4688,N_47953,N_45466);
nand UO_4689 (O_4689,N_49874,N_45599);
nand UO_4690 (O_4690,N_47237,N_45964);
nand UO_4691 (O_4691,N_46522,N_49301);
nand UO_4692 (O_4692,N_47827,N_45035);
or UO_4693 (O_4693,N_45793,N_49255);
nor UO_4694 (O_4694,N_48393,N_49488);
xor UO_4695 (O_4695,N_48659,N_45122);
xor UO_4696 (O_4696,N_47778,N_46761);
xor UO_4697 (O_4697,N_45594,N_49673);
and UO_4698 (O_4698,N_47956,N_46871);
nor UO_4699 (O_4699,N_46687,N_46292);
or UO_4700 (O_4700,N_47451,N_46441);
or UO_4701 (O_4701,N_49985,N_46999);
nand UO_4702 (O_4702,N_48333,N_48924);
xnor UO_4703 (O_4703,N_46035,N_49131);
nor UO_4704 (O_4704,N_48182,N_48681);
nor UO_4705 (O_4705,N_46251,N_45629);
and UO_4706 (O_4706,N_47454,N_45686);
and UO_4707 (O_4707,N_46048,N_45588);
xor UO_4708 (O_4708,N_49969,N_48863);
and UO_4709 (O_4709,N_46627,N_49534);
or UO_4710 (O_4710,N_46279,N_48838);
nor UO_4711 (O_4711,N_46675,N_48758);
or UO_4712 (O_4712,N_47342,N_48783);
nor UO_4713 (O_4713,N_46657,N_48762);
nor UO_4714 (O_4714,N_45007,N_46707);
or UO_4715 (O_4715,N_46935,N_46204);
or UO_4716 (O_4716,N_46688,N_47056);
xnor UO_4717 (O_4717,N_47652,N_48619);
and UO_4718 (O_4718,N_45914,N_49296);
xnor UO_4719 (O_4719,N_48752,N_48551);
xor UO_4720 (O_4720,N_48957,N_45041);
and UO_4721 (O_4721,N_48207,N_46597);
xnor UO_4722 (O_4722,N_46328,N_48635);
or UO_4723 (O_4723,N_48137,N_48769);
nand UO_4724 (O_4724,N_47603,N_45694);
nor UO_4725 (O_4725,N_48450,N_48996);
or UO_4726 (O_4726,N_46728,N_48846);
nor UO_4727 (O_4727,N_49466,N_48403);
or UO_4728 (O_4728,N_47234,N_46832);
nand UO_4729 (O_4729,N_48037,N_49074);
or UO_4730 (O_4730,N_47700,N_45117);
nor UO_4731 (O_4731,N_46118,N_47915);
nor UO_4732 (O_4732,N_46144,N_48137);
nand UO_4733 (O_4733,N_49607,N_47421);
nor UO_4734 (O_4734,N_46818,N_49943);
or UO_4735 (O_4735,N_46156,N_49999);
nor UO_4736 (O_4736,N_49923,N_46951);
nand UO_4737 (O_4737,N_45997,N_49396);
nor UO_4738 (O_4738,N_49263,N_48746);
or UO_4739 (O_4739,N_49116,N_46225);
xnor UO_4740 (O_4740,N_49096,N_48864);
nor UO_4741 (O_4741,N_46680,N_48335);
or UO_4742 (O_4742,N_45585,N_49751);
or UO_4743 (O_4743,N_46353,N_49917);
nand UO_4744 (O_4744,N_47486,N_49453);
xor UO_4745 (O_4745,N_48147,N_47946);
nand UO_4746 (O_4746,N_48140,N_46810);
xnor UO_4747 (O_4747,N_46917,N_46733);
nand UO_4748 (O_4748,N_49612,N_48018);
and UO_4749 (O_4749,N_48489,N_48505);
nor UO_4750 (O_4750,N_48125,N_48834);
nor UO_4751 (O_4751,N_46000,N_49757);
or UO_4752 (O_4752,N_46310,N_48987);
nand UO_4753 (O_4753,N_47457,N_45503);
and UO_4754 (O_4754,N_46813,N_48764);
and UO_4755 (O_4755,N_45774,N_47350);
xnor UO_4756 (O_4756,N_45662,N_45834);
and UO_4757 (O_4757,N_45567,N_45987);
and UO_4758 (O_4758,N_48519,N_46803);
or UO_4759 (O_4759,N_48286,N_46358);
nor UO_4760 (O_4760,N_47562,N_45893);
and UO_4761 (O_4761,N_47590,N_46047);
or UO_4762 (O_4762,N_45498,N_48273);
nand UO_4763 (O_4763,N_48635,N_45230);
and UO_4764 (O_4764,N_45149,N_49966);
nand UO_4765 (O_4765,N_46017,N_47959);
nand UO_4766 (O_4766,N_48918,N_49876);
and UO_4767 (O_4767,N_48998,N_45115);
xnor UO_4768 (O_4768,N_47646,N_49687);
nor UO_4769 (O_4769,N_45464,N_48802);
nor UO_4770 (O_4770,N_48713,N_46274);
nor UO_4771 (O_4771,N_48113,N_45951);
or UO_4772 (O_4772,N_48387,N_47549);
nor UO_4773 (O_4773,N_45957,N_46444);
nand UO_4774 (O_4774,N_47705,N_45679);
nor UO_4775 (O_4775,N_49797,N_49947);
xnor UO_4776 (O_4776,N_47347,N_47843);
or UO_4777 (O_4777,N_48069,N_46830);
nor UO_4778 (O_4778,N_49596,N_46763);
and UO_4779 (O_4779,N_48600,N_47925);
xor UO_4780 (O_4780,N_48931,N_45344);
nand UO_4781 (O_4781,N_47710,N_49476);
xnor UO_4782 (O_4782,N_47803,N_45174);
or UO_4783 (O_4783,N_48545,N_46057);
nand UO_4784 (O_4784,N_47410,N_47667);
and UO_4785 (O_4785,N_48081,N_48930);
or UO_4786 (O_4786,N_46402,N_45474);
nor UO_4787 (O_4787,N_45762,N_49166);
xor UO_4788 (O_4788,N_46877,N_47500);
or UO_4789 (O_4789,N_46884,N_46647);
and UO_4790 (O_4790,N_46812,N_45414);
xor UO_4791 (O_4791,N_48826,N_48119);
or UO_4792 (O_4792,N_49551,N_48412);
nor UO_4793 (O_4793,N_49947,N_49786);
xnor UO_4794 (O_4794,N_48936,N_47878);
or UO_4795 (O_4795,N_47012,N_49159);
xnor UO_4796 (O_4796,N_46084,N_47353);
or UO_4797 (O_4797,N_47316,N_47331);
or UO_4798 (O_4798,N_47718,N_47548);
nand UO_4799 (O_4799,N_47542,N_47116);
or UO_4800 (O_4800,N_48828,N_48631);
nand UO_4801 (O_4801,N_48372,N_48921);
nand UO_4802 (O_4802,N_46048,N_48737);
xor UO_4803 (O_4803,N_48012,N_48904);
or UO_4804 (O_4804,N_45534,N_45511);
or UO_4805 (O_4805,N_47120,N_49280);
xnor UO_4806 (O_4806,N_45709,N_45771);
nor UO_4807 (O_4807,N_48270,N_47345);
nand UO_4808 (O_4808,N_49043,N_47677);
or UO_4809 (O_4809,N_46653,N_45730);
nor UO_4810 (O_4810,N_47499,N_46514);
and UO_4811 (O_4811,N_49804,N_49209);
or UO_4812 (O_4812,N_46436,N_46593);
nor UO_4813 (O_4813,N_48716,N_46731);
or UO_4814 (O_4814,N_49639,N_45803);
nor UO_4815 (O_4815,N_49907,N_49157);
nand UO_4816 (O_4816,N_49639,N_47501);
nand UO_4817 (O_4817,N_46582,N_45329);
nor UO_4818 (O_4818,N_45478,N_48481);
nor UO_4819 (O_4819,N_45816,N_46935);
or UO_4820 (O_4820,N_45558,N_49521);
xor UO_4821 (O_4821,N_47134,N_47421);
or UO_4822 (O_4822,N_49042,N_49728);
or UO_4823 (O_4823,N_48708,N_49784);
or UO_4824 (O_4824,N_49941,N_45561);
and UO_4825 (O_4825,N_48195,N_49478);
nand UO_4826 (O_4826,N_47691,N_48713);
nand UO_4827 (O_4827,N_46698,N_49231);
nand UO_4828 (O_4828,N_45675,N_46491);
xor UO_4829 (O_4829,N_49015,N_47115);
and UO_4830 (O_4830,N_48433,N_46415);
xor UO_4831 (O_4831,N_46215,N_48893);
nor UO_4832 (O_4832,N_45926,N_45830);
nand UO_4833 (O_4833,N_45135,N_48919);
or UO_4834 (O_4834,N_46807,N_49835);
xnor UO_4835 (O_4835,N_48368,N_46801);
xor UO_4836 (O_4836,N_47546,N_48415);
nor UO_4837 (O_4837,N_49634,N_47891);
nand UO_4838 (O_4838,N_47758,N_45038);
or UO_4839 (O_4839,N_45028,N_45229);
or UO_4840 (O_4840,N_46606,N_46688);
nor UO_4841 (O_4841,N_49322,N_47384);
or UO_4842 (O_4842,N_48446,N_47353);
nand UO_4843 (O_4843,N_46755,N_48516);
nor UO_4844 (O_4844,N_45944,N_46694);
and UO_4845 (O_4845,N_49987,N_47245);
xnor UO_4846 (O_4846,N_46575,N_48004);
xor UO_4847 (O_4847,N_47082,N_45101);
xnor UO_4848 (O_4848,N_47178,N_46217);
and UO_4849 (O_4849,N_49463,N_49140);
nor UO_4850 (O_4850,N_46163,N_46014);
xnor UO_4851 (O_4851,N_49600,N_46419);
or UO_4852 (O_4852,N_45439,N_46133);
and UO_4853 (O_4853,N_48548,N_48834);
and UO_4854 (O_4854,N_49600,N_46838);
or UO_4855 (O_4855,N_49769,N_48407);
nor UO_4856 (O_4856,N_45269,N_49423);
nor UO_4857 (O_4857,N_45991,N_48146);
xor UO_4858 (O_4858,N_48945,N_47546);
xor UO_4859 (O_4859,N_48234,N_46176);
nand UO_4860 (O_4860,N_47957,N_48263);
nand UO_4861 (O_4861,N_46209,N_48198);
or UO_4862 (O_4862,N_46915,N_49027);
nor UO_4863 (O_4863,N_46338,N_47786);
xor UO_4864 (O_4864,N_49590,N_49393);
nor UO_4865 (O_4865,N_46192,N_47198);
nor UO_4866 (O_4866,N_46759,N_46068);
xnor UO_4867 (O_4867,N_45622,N_49345);
nor UO_4868 (O_4868,N_49064,N_45552);
or UO_4869 (O_4869,N_45149,N_48247);
nand UO_4870 (O_4870,N_48282,N_45931);
xor UO_4871 (O_4871,N_48180,N_49789);
and UO_4872 (O_4872,N_47424,N_45112);
xnor UO_4873 (O_4873,N_47982,N_45273);
or UO_4874 (O_4874,N_49011,N_48945);
nor UO_4875 (O_4875,N_45306,N_45044);
nor UO_4876 (O_4876,N_47617,N_48659);
or UO_4877 (O_4877,N_47685,N_45827);
and UO_4878 (O_4878,N_46604,N_49783);
or UO_4879 (O_4879,N_48413,N_49941);
or UO_4880 (O_4880,N_46642,N_48117);
nor UO_4881 (O_4881,N_49010,N_49922);
nor UO_4882 (O_4882,N_48693,N_45326);
and UO_4883 (O_4883,N_49422,N_49187);
xnor UO_4884 (O_4884,N_49644,N_49779);
nor UO_4885 (O_4885,N_45395,N_48326);
or UO_4886 (O_4886,N_49195,N_49701);
nand UO_4887 (O_4887,N_45735,N_46076);
nor UO_4888 (O_4888,N_46959,N_48890);
nand UO_4889 (O_4889,N_46524,N_47015);
nor UO_4890 (O_4890,N_49630,N_46657);
nor UO_4891 (O_4891,N_47941,N_46413);
and UO_4892 (O_4892,N_48448,N_45600);
nand UO_4893 (O_4893,N_48420,N_49714);
or UO_4894 (O_4894,N_48440,N_48696);
and UO_4895 (O_4895,N_46489,N_47030);
and UO_4896 (O_4896,N_49699,N_48401);
nand UO_4897 (O_4897,N_49405,N_46008);
and UO_4898 (O_4898,N_46511,N_45592);
nand UO_4899 (O_4899,N_45794,N_47745);
and UO_4900 (O_4900,N_48505,N_46611);
nand UO_4901 (O_4901,N_47305,N_46378);
and UO_4902 (O_4902,N_49091,N_45495);
xor UO_4903 (O_4903,N_48249,N_46997);
nor UO_4904 (O_4904,N_49229,N_45664);
and UO_4905 (O_4905,N_47635,N_49669);
or UO_4906 (O_4906,N_46909,N_48278);
nand UO_4907 (O_4907,N_46663,N_45686);
or UO_4908 (O_4908,N_45701,N_49820);
xor UO_4909 (O_4909,N_46545,N_45829);
xor UO_4910 (O_4910,N_45907,N_46406);
or UO_4911 (O_4911,N_48155,N_49412);
or UO_4912 (O_4912,N_46616,N_47752);
nor UO_4913 (O_4913,N_48999,N_47071);
or UO_4914 (O_4914,N_49718,N_48540);
nor UO_4915 (O_4915,N_47131,N_48617);
and UO_4916 (O_4916,N_48543,N_45107);
xnor UO_4917 (O_4917,N_48226,N_46034);
nand UO_4918 (O_4918,N_46439,N_48853);
nand UO_4919 (O_4919,N_46893,N_49810);
nand UO_4920 (O_4920,N_47212,N_48308);
nand UO_4921 (O_4921,N_49780,N_46277);
nand UO_4922 (O_4922,N_45196,N_48117);
nand UO_4923 (O_4923,N_45310,N_48658);
or UO_4924 (O_4924,N_46414,N_47571);
and UO_4925 (O_4925,N_48214,N_49120);
nor UO_4926 (O_4926,N_45887,N_45333);
or UO_4927 (O_4927,N_49142,N_47107);
xor UO_4928 (O_4928,N_46556,N_47534);
xnor UO_4929 (O_4929,N_46429,N_45490);
or UO_4930 (O_4930,N_46761,N_47854);
and UO_4931 (O_4931,N_45305,N_46297);
nand UO_4932 (O_4932,N_49629,N_49878);
and UO_4933 (O_4933,N_45941,N_45373);
xnor UO_4934 (O_4934,N_47663,N_46337);
nor UO_4935 (O_4935,N_47673,N_45489);
nor UO_4936 (O_4936,N_49253,N_47163);
or UO_4937 (O_4937,N_49438,N_48295);
nor UO_4938 (O_4938,N_48910,N_49612);
or UO_4939 (O_4939,N_49087,N_46857);
nor UO_4940 (O_4940,N_45868,N_49165);
nor UO_4941 (O_4941,N_45583,N_49562);
and UO_4942 (O_4942,N_49742,N_45245);
xor UO_4943 (O_4943,N_45326,N_48009);
xor UO_4944 (O_4944,N_48801,N_46006);
nand UO_4945 (O_4945,N_45984,N_49623);
and UO_4946 (O_4946,N_48548,N_48549);
or UO_4947 (O_4947,N_48647,N_46461);
nor UO_4948 (O_4948,N_46311,N_47149);
nand UO_4949 (O_4949,N_49090,N_46133);
and UO_4950 (O_4950,N_45450,N_47080);
xor UO_4951 (O_4951,N_47627,N_47925);
and UO_4952 (O_4952,N_48298,N_48074);
and UO_4953 (O_4953,N_47414,N_48568);
xor UO_4954 (O_4954,N_46673,N_47168);
nor UO_4955 (O_4955,N_49825,N_47637);
xor UO_4956 (O_4956,N_49767,N_47033);
xor UO_4957 (O_4957,N_46870,N_46719);
and UO_4958 (O_4958,N_45307,N_46988);
nor UO_4959 (O_4959,N_48769,N_49738);
or UO_4960 (O_4960,N_48808,N_46018);
nand UO_4961 (O_4961,N_48016,N_49996);
nand UO_4962 (O_4962,N_45247,N_46860);
and UO_4963 (O_4963,N_49553,N_49866);
or UO_4964 (O_4964,N_45251,N_46620);
xor UO_4965 (O_4965,N_46201,N_48642);
nor UO_4966 (O_4966,N_49587,N_46495);
or UO_4967 (O_4967,N_46683,N_47119);
or UO_4968 (O_4968,N_45700,N_47465);
nand UO_4969 (O_4969,N_48661,N_47613);
or UO_4970 (O_4970,N_45433,N_47521);
or UO_4971 (O_4971,N_46391,N_47608);
nand UO_4972 (O_4972,N_47372,N_47301);
nor UO_4973 (O_4973,N_45127,N_46590);
and UO_4974 (O_4974,N_47147,N_47952);
or UO_4975 (O_4975,N_46570,N_45229);
nand UO_4976 (O_4976,N_45172,N_46674);
and UO_4977 (O_4977,N_49749,N_47009);
xnor UO_4978 (O_4978,N_45768,N_45478);
nand UO_4979 (O_4979,N_48677,N_49670);
xor UO_4980 (O_4980,N_47829,N_49614);
and UO_4981 (O_4981,N_49148,N_46388);
nor UO_4982 (O_4982,N_45787,N_45902);
or UO_4983 (O_4983,N_47767,N_45626);
nor UO_4984 (O_4984,N_48082,N_49746);
nor UO_4985 (O_4985,N_45974,N_45577);
nor UO_4986 (O_4986,N_46263,N_45917);
or UO_4987 (O_4987,N_46484,N_45706);
nand UO_4988 (O_4988,N_46676,N_47977);
or UO_4989 (O_4989,N_47835,N_48509);
or UO_4990 (O_4990,N_47938,N_46633);
xor UO_4991 (O_4991,N_49611,N_46402);
and UO_4992 (O_4992,N_48478,N_46600);
nand UO_4993 (O_4993,N_49763,N_48024);
nor UO_4994 (O_4994,N_49931,N_46855);
nor UO_4995 (O_4995,N_48850,N_47483);
nand UO_4996 (O_4996,N_47363,N_49439);
or UO_4997 (O_4997,N_49441,N_45303);
and UO_4998 (O_4998,N_45214,N_48289);
nor UO_4999 (O_4999,N_46285,N_49689);
endmodule