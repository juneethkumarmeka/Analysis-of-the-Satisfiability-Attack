module basic_500_3000_500_50_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_420,In_448);
and U1 (N_1,In_125,In_313);
and U2 (N_2,In_370,In_88);
nand U3 (N_3,In_426,In_309);
nor U4 (N_4,In_481,In_16);
or U5 (N_5,In_432,In_207);
nor U6 (N_6,In_133,In_337);
and U7 (N_7,In_410,In_32);
nor U8 (N_8,In_163,In_222);
nor U9 (N_9,In_324,In_76);
and U10 (N_10,In_327,In_78);
nor U11 (N_11,In_155,In_300);
nand U12 (N_12,In_77,In_454);
xor U13 (N_13,In_306,In_232);
and U14 (N_14,In_376,In_67);
and U15 (N_15,In_457,In_434);
nor U16 (N_16,In_68,In_120);
or U17 (N_17,In_165,In_196);
and U18 (N_18,In_170,In_275);
or U19 (N_19,In_246,In_399);
nand U20 (N_20,In_267,In_50);
nand U21 (N_21,In_189,In_494);
nand U22 (N_22,In_462,In_418);
xnor U23 (N_23,In_31,In_72);
xnor U24 (N_24,In_202,In_444);
and U25 (N_25,In_354,In_447);
nand U26 (N_26,In_11,In_223);
and U27 (N_27,In_391,In_497);
nand U28 (N_28,In_18,In_393);
xor U29 (N_29,In_6,In_171);
nand U30 (N_30,In_211,In_105);
nor U31 (N_31,In_152,In_241);
xor U32 (N_32,In_35,In_179);
or U33 (N_33,In_84,In_27);
nor U34 (N_34,In_363,In_26);
nand U35 (N_35,In_452,In_279);
and U36 (N_36,In_383,In_262);
nor U37 (N_37,In_66,In_28);
nand U38 (N_38,In_90,In_479);
and U39 (N_39,In_29,In_71);
and U40 (N_40,In_178,In_149);
xnor U41 (N_41,In_417,In_231);
nand U42 (N_42,In_386,In_419);
nand U43 (N_43,In_406,In_69);
nor U44 (N_44,In_480,In_312);
and U45 (N_45,In_98,In_377);
or U46 (N_46,In_25,In_79);
nor U47 (N_47,In_161,In_297);
nand U48 (N_48,In_103,In_298);
or U49 (N_49,In_290,In_226);
nand U50 (N_50,In_319,In_325);
xor U51 (N_51,In_473,In_151);
nand U52 (N_52,In_214,In_58);
xnor U53 (N_53,In_199,In_48);
nor U54 (N_54,In_437,In_174);
nand U55 (N_55,In_43,In_445);
nand U56 (N_56,In_466,In_156);
and U57 (N_57,In_200,In_299);
and U58 (N_58,In_331,In_157);
or U59 (N_59,In_233,In_381);
nor U60 (N_60,In_358,In_276);
or U61 (N_61,In_465,N_15);
or U62 (N_62,In_96,In_115);
nand U63 (N_63,In_459,In_51);
nand U64 (N_64,In_345,N_52);
or U65 (N_65,In_340,In_476);
nor U66 (N_66,In_140,In_209);
or U67 (N_67,In_326,In_158);
xnor U68 (N_68,In_339,In_487);
or U69 (N_69,In_414,In_413);
xor U70 (N_70,N_2,In_273);
nand U71 (N_71,In_0,In_239);
nor U72 (N_72,In_236,In_373);
and U73 (N_73,N_30,In_488);
or U74 (N_74,In_284,In_94);
nand U75 (N_75,In_34,N_6);
nor U76 (N_76,In_364,In_63);
or U77 (N_77,N_12,In_95);
and U78 (N_78,In_320,In_382);
nand U79 (N_79,In_142,In_441);
and U80 (N_80,In_243,In_408);
nand U81 (N_81,N_57,In_294);
or U82 (N_82,N_13,In_99);
nand U83 (N_83,In_45,In_416);
xor U84 (N_84,In_153,In_40);
nand U85 (N_85,In_485,In_277);
nand U86 (N_86,In_201,In_291);
nand U87 (N_87,N_19,In_283);
nand U88 (N_88,In_74,In_102);
nor U89 (N_89,In_59,N_3);
or U90 (N_90,In_5,In_435);
nor U91 (N_91,In_144,In_440);
nor U92 (N_92,In_57,In_311);
xor U93 (N_93,In_65,In_55);
or U94 (N_94,In_124,In_130);
xnor U95 (N_95,In_169,In_463);
and U96 (N_96,In_367,In_475);
and U97 (N_97,In_372,In_258);
nor U98 (N_98,In_310,In_353);
or U99 (N_99,In_173,In_177);
nor U100 (N_100,In_371,N_21);
nor U101 (N_101,In_346,N_53);
xor U102 (N_102,In_350,In_37);
nor U103 (N_103,N_0,In_316);
nor U104 (N_104,In_164,In_315);
and U105 (N_105,In_126,N_47);
or U106 (N_106,In_47,In_46);
xnor U107 (N_107,In_288,In_464);
nor U108 (N_108,In_398,N_44);
nand U109 (N_109,In_104,In_280);
and U110 (N_110,In_317,In_217);
xnor U111 (N_111,In_123,In_42);
or U112 (N_112,In_355,In_287);
and U113 (N_113,In_184,In_368);
nor U114 (N_114,In_251,In_139);
nor U115 (N_115,In_458,In_237);
or U116 (N_116,In_396,In_54);
nor U117 (N_117,In_235,In_166);
xor U118 (N_118,In_147,N_34);
nand U119 (N_119,N_59,In_110);
nor U120 (N_120,N_8,In_425);
nand U121 (N_121,In_266,In_121);
and U122 (N_122,In_255,In_292);
nand U123 (N_123,In_119,N_72);
xor U124 (N_124,N_77,In_19);
nand U125 (N_125,N_113,N_54);
and U126 (N_126,In_187,In_343);
or U127 (N_127,In_181,N_86);
nor U128 (N_128,In_248,In_449);
nand U129 (N_129,In_415,In_256);
nand U130 (N_130,In_385,In_438);
or U131 (N_131,In_114,N_46);
nand U132 (N_132,N_85,In_225);
and U133 (N_133,In_210,N_18);
nand U134 (N_134,In_433,In_221);
or U135 (N_135,In_384,N_78);
and U136 (N_136,In_271,In_428);
or U137 (N_137,In_356,In_351);
or U138 (N_138,In_112,N_24);
nand U139 (N_139,In_213,In_427);
nor U140 (N_140,In_92,In_492);
nor U141 (N_141,In_93,In_182);
nor U142 (N_142,N_32,N_80);
and U143 (N_143,In_249,In_3);
nor U144 (N_144,In_36,In_108);
and U145 (N_145,In_264,In_146);
and U146 (N_146,In_135,N_70);
nand U147 (N_147,In_302,In_349);
nor U148 (N_148,N_56,N_49);
nor U149 (N_149,In_205,In_424);
or U150 (N_150,In_453,In_228);
nand U151 (N_151,N_45,N_92);
nor U152 (N_152,In_357,N_50);
nand U153 (N_153,In_293,In_131);
or U154 (N_154,In_304,In_482);
nor U155 (N_155,In_446,In_484);
and U156 (N_156,In_73,In_215);
nor U157 (N_157,N_41,In_474);
xnor U158 (N_158,In_362,In_122);
and U159 (N_159,In_62,In_483);
nor U160 (N_160,In_378,N_95);
nand U161 (N_161,In_344,In_183);
nor U162 (N_162,In_100,N_69);
xnor U163 (N_163,In_188,In_336);
nand U164 (N_164,In_176,In_301);
and U165 (N_165,In_456,In_366);
and U166 (N_166,N_90,N_83);
nor U167 (N_167,In_13,In_22);
xor U168 (N_168,In_407,In_137);
nor U169 (N_169,In_422,N_76);
and U170 (N_170,In_83,In_186);
nand U171 (N_171,N_25,In_192);
nor U172 (N_172,In_278,In_1);
nor U173 (N_173,N_101,In_87);
xor U174 (N_174,In_134,N_79);
and U175 (N_175,In_250,N_42);
nor U176 (N_176,In_49,In_431);
or U177 (N_177,In_91,N_60);
or U178 (N_178,N_105,In_314);
and U179 (N_179,In_116,In_64);
nand U180 (N_180,N_130,N_63);
or U181 (N_181,In_308,In_259);
nand U182 (N_182,N_87,N_96);
or U183 (N_183,In_9,N_135);
or U184 (N_184,In_252,In_208);
xnor U185 (N_185,N_51,In_80);
nand U186 (N_186,In_60,In_175);
nor U187 (N_187,N_89,N_117);
nand U188 (N_188,In_20,In_109);
or U189 (N_189,N_128,In_61);
and U190 (N_190,In_374,N_163);
or U191 (N_191,In_86,In_220);
and U192 (N_192,N_168,In_334);
or U193 (N_193,N_33,In_127);
and U194 (N_194,N_166,N_74);
and U195 (N_195,N_178,In_421);
nor U196 (N_196,In_148,In_97);
and U197 (N_197,In_491,In_14);
nand U198 (N_198,In_490,N_124);
or U199 (N_199,In_234,In_162);
and U200 (N_200,N_103,N_29);
nand U201 (N_201,In_160,In_113);
and U202 (N_202,N_7,In_429);
or U203 (N_203,In_85,N_37);
and U204 (N_204,In_75,In_359);
or U205 (N_205,In_154,N_141);
nand U206 (N_206,In_450,N_114);
nand U207 (N_207,In_106,In_24);
or U208 (N_208,In_8,N_1);
and U209 (N_209,In_471,In_361);
nand U210 (N_210,N_164,In_159);
xor U211 (N_211,In_30,In_305);
nand U212 (N_212,N_104,In_388);
or U213 (N_213,N_26,In_338);
nor U214 (N_214,N_116,N_48);
nor U215 (N_215,N_82,N_115);
nand U216 (N_216,N_153,N_17);
nor U217 (N_217,N_23,In_7);
or U218 (N_218,In_39,N_161);
nand U219 (N_219,In_442,In_289);
nand U220 (N_220,N_100,In_468);
nand U221 (N_221,In_321,In_81);
nand U222 (N_222,In_107,In_369);
or U223 (N_223,In_496,In_461);
nor U224 (N_224,In_129,In_38);
nand U225 (N_225,In_470,In_82);
nand U226 (N_226,N_71,In_455);
nand U227 (N_227,N_110,In_227);
and U228 (N_228,N_132,In_402);
or U229 (N_229,In_128,N_91);
nand U230 (N_230,N_39,In_477);
or U231 (N_231,In_307,In_229);
or U232 (N_232,N_66,N_5);
nor U233 (N_233,N_11,N_108);
and U234 (N_234,N_22,In_333);
nand U235 (N_235,In_436,N_120);
nand U236 (N_236,N_84,N_88);
nor U237 (N_237,In_411,In_412);
nor U238 (N_238,In_286,In_197);
xnor U239 (N_239,N_129,N_139);
nor U240 (N_240,N_195,In_423);
xnor U241 (N_241,In_323,In_41);
and U242 (N_242,In_193,N_68);
or U243 (N_243,N_16,In_2);
and U244 (N_244,N_222,N_191);
nor U245 (N_245,N_155,In_141);
nand U246 (N_246,In_499,In_272);
nand U247 (N_247,In_167,N_189);
nand U248 (N_248,In_430,N_165);
or U249 (N_249,In_136,In_270);
or U250 (N_250,N_215,N_109);
and U251 (N_251,N_150,N_190);
or U252 (N_252,In_469,N_145);
nor U253 (N_253,N_185,In_260);
xnor U254 (N_254,N_20,N_202);
nand U255 (N_255,In_242,In_281);
nor U256 (N_256,In_203,In_269);
and U257 (N_257,N_234,N_206);
nor U258 (N_258,N_118,N_111);
and U259 (N_259,N_61,N_158);
nor U260 (N_260,N_193,N_169);
or U261 (N_261,In_392,In_387);
and U262 (N_262,In_143,N_123);
and U263 (N_263,N_94,N_156);
nand U264 (N_264,In_212,N_73);
nor U265 (N_265,In_352,N_93);
or U266 (N_266,In_467,N_233);
nand U267 (N_267,N_147,In_70);
or U268 (N_268,N_170,N_154);
or U269 (N_269,In_89,In_395);
or U270 (N_270,N_229,In_132);
or U271 (N_271,N_194,N_102);
or U272 (N_272,N_220,N_131);
or U273 (N_273,N_188,In_194);
nand U274 (N_274,In_44,In_253);
and U275 (N_275,N_237,In_365);
nand U276 (N_276,In_403,In_268);
nor U277 (N_277,In_191,In_360);
xnor U278 (N_278,N_196,N_173);
and U279 (N_279,N_227,N_213);
and U280 (N_280,In_261,In_172);
and U281 (N_281,N_159,N_223);
or U282 (N_282,In_21,In_10);
or U283 (N_283,N_99,In_218);
or U284 (N_284,In_443,In_195);
nand U285 (N_285,In_238,N_162);
xnor U286 (N_286,N_209,N_127);
xor U287 (N_287,In_263,In_451);
or U288 (N_288,In_390,In_240);
or U289 (N_289,In_282,N_62);
nor U290 (N_290,N_219,N_126);
and U291 (N_291,N_143,N_67);
nand U292 (N_292,In_285,In_303);
and U293 (N_293,In_472,In_168);
xnor U294 (N_294,In_332,N_187);
or U295 (N_295,N_112,In_254);
and U296 (N_296,N_212,N_204);
nand U297 (N_297,In_498,In_329);
and U298 (N_298,N_199,In_295);
and U299 (N_299,N_14,N_119);
nand U300 (N_300,N_291,N_250);
and U301 (N_301,In_247,In_198);
or U302 (N_302,N_217,N_172);
xnor U303 (N_303,N_121,N_261);
xor U304 (N_304,N_293,In_244);
and U305 (N_305,N_275,N_133);
xor U306 (N_306,N_97,In_230);
nor U307 (N_307,N_174,In_348);
and U308 (N_308,N_176,In_439);
nand U309 (N_309,N_268,N_122);
or U310 (N_310,In_245,N_65);
nand U311 (N_311,N_267,N_228);
and U312 (N_312,N_273,N_277);
nand U313 (N_313,In_322,N_207);
nand U314 (N_314,N_260,N_266);
or U315 (N_315,N_245,N_257);
nor U316 (N_316,In_4,In_274);
nor U317 (N_317,N_278,In_389);
or U318 (N_318,N_272,In_341);
or U319 (N_319,N_242,In_204);
and U320 (N_320,N_270,N_10);
or U321 (N_321,N_274,N_40);
or U322 (N_322,In_400,N_232);
nor U323 (N_323,N_146,N_179);
nor U324 (N_324,In_493,In_145);
nand U325 (N_325,N_286,N_231);
xnor U326 (N_326,N_31,N_98);
xor U327 (N_327,N_151,N_148);
and U328 (N_328,N_253,N_249);
nand U329 (N_329,N_180,N_281);
nor U330 (N_330,N_27,N_280);
and U331 (N_331,N_64,In_101);
and U332 (N_332,N_283,N_299);
nor U333 (N_333,N_216,N_271);
nand U334 (N_334,In_478,In_15);
and U335 (N_335,N_251,N_138);
nand U336 (N_336,N_201,N_203);
xnor U337 (N_337,N_269,N_43);
or U338 (N_338,In_111,N_197);
or U339 (N_339,N_28,N_235);
or U340 (N_340,In_190,In_401);
nor U341 (N_341,N_149,In_53);
or U342 (N_342,N_171,N_4);
or U343 (N_343,N_183,N_142);
and U344 (N_344,N_160,N_137);
nand U345 (N_345,N_288,In_404);
nand U346 (N_346,In_118,N_247);
nand U347 (N_347,N_282,In_56);
or U348 (N_348,N_264,N_290);
nor U349 (N_349,In_397,N_186);
nor U350 (N_350,N_297,N_254);
or U351 (N_351,N_144,N_218);
and U352 (N_352,N_36,In_335);
xor U353 (N_353,N_198,N_248);
and U354 (N_354,N_9,N_262);
nand U355 (N_355,N_292,N_157);
and U356 (N_356,N_298,N_182);
nor U357 (N_357,N_210,N_107);
nor U358 (N_358,In_405,N_224);
or U359 (N_359,N_276,N_208);
or U360 (N_360,N_329,N_308);
xor U361 (N_361,N_334,In_296);
and U362 (N_362,N_342,N_318);
nand U363 (N_363,N_284,N_306);
xor U364 (N_364,N_184,In_265);
nand U365 (N_365,N_301,In_495);
and U366 (N_366,In_33,N_305);
nand U367 (N_367,N_357,N_226);
nor U368 (N_368,N_300,N_352);
and U369 (N_369,N_75,N_279);
nand U370 (N_370,N_309,N_175);
or U371 (N_371,N_327,N_255);
or U372 (N_372,In_219,In_185);
or U373 (N_373,In_257,In_180);
or U374 (N_374,In_150,N_287);
and U375 (N_375,N_343,N_259);
nor U376 (N_376,N_35,N_238);
and U377 (N_377,N_295,N_346);
and U378 (N_378,N_256,N_140);
nand U379 (N_379,In_117,N_349);
nor U380 (N_380,N_134,N_152);
or U381 (N_381,N_244,N_200);
nor U382 (N_382,N_177,N_335);
nand U383 (N_383,N_347,N_230);
nor U384 (N_384,In_394,N_265);
nor U385 (N_385,N_302,N_311);
or U386 (N_386,N_354,N_225);
and U387 (N_387,N_323,N_341);
and U388 (N_388,N_317,N_38);
nor U389 (N_389,N_221,N_350);
nor U390 (N_390,N_313,N_181);
nor U391 (N_391,N_322,N_340);
or U392 (N_392,N_211,N_55);
xnor U393 (N_393,N_351,N_315);
nand U394 (N_394,N_214,In_409);
or U395 (N_395,N_304,N_258);
nor U396 (N_396,In_460,In_23);
xor U397 (N_397,N_333,N_58);
nor U398 (N_398,N_359,In_379);
xnor U399 (N_399,In_375,In_380);
or U400 (N_400,N_136,N_240);
nand U401 (N_401,N_263,In_12);
nand U402 (N_402,N_285,N_303);
and U403 (N_403,N_252,N_192);
nor U404 (N_404,N_326,N_243);
and U405 (N_405,N_336,N_321);
and U406 (N_406,In_224,In_138);
xor U407 (N_407,In_52,N_356);
nand U408 (N_408,N_307,N_325);
or U409 (N_409,N_337,N_239);
nor U410 (N_410,N_358,N_167);
nand U411 (N_411,In_347,N_353);
and U412 (N_412,N_330,In_206);
nand U413 (N_413,N_344,N_246);
or U414 (N_414,N_236,N_289);
and U415 (N_415,N_348,In_17);
nand U416 (N_416,N_81,N_205);
nor U417 (N_417,In_489,In_342);
or U418 (N_418,N_320,In_330);
nand U419 (N_419,N_241,N_345);
nor U420 (N_420,N_296,N_406);
nor U421 (N_421,N_414,N_360);
nor U422 (N_422,N_398,N_416);
nor U423 (N_423,N_370,N_364);
and U424 (N_424,N_418,N_413);
nand U425 (N_425,N_384,N_381);
nor U426 (N_426,N_368,N_404);
or U427 (N_427,N_377,In_318);
and U428 (N_428,N_362,N_312);
nor U429 (N_429,N_393,N_379);
and U430 (N_430,N_412,N_372);
xnor U431 (N_431,N_324,N_310);
nand U432 (N_432,N_401,N_399);
nor U433 (N_433,N_397,N_392);
or U434 (N_434,N_316,N_374);
and U435 (N_435,N_396,In_328);
nand U436 (N_436,N_408,N_386);
xnor U437 (N_437,N_383,N_387);
and U438 (N_438,N_376,N_371);
nand U439 (N_439,N_125,N_339);
nand U440 (N_440,N_411,N_403);
nand U441 (N_441,N_400,N_391);
and U442 (N_442,N_419,N_328);
nand U443 (N_443,N_314,N_389);
nor U444 (N_444,N_331,N_378);
nand U445 (N_445,N_367,N_407);
nand U446 (N_446,N_366,N_390);
and U447 (N_447,In_486,In_216);
or U448 (N_448,N_417,N_106);
nor U449 (N_449,N_380,N_369);
and U450 (N_450,N_319,N_361);
nand U451 (N_451,N_388,N_294);
nor U452 (N_452,N_363,N_395);
and U453 (N_453,N_332,N_409);
xnor U454 (N_454,N_394,N_373);
and U455 (N_455,N_365,N_338);
or U456 (N_456,N_385,N_415);
or U457 (N_457,N_402,N_405);
xor U458 (N_458,N_382,N_375);
nor U459 (N_459,N_355,N_410);
nand U460 (N_460,N_370,N_375);
and U461 (N_461,N_364,N_399);
nand U462 (N_462,N_396,N_387);
or U463 (N_463,N_386,N_366);
nor U464 (N_464,N_365,N_413);
or U465 (N_465,N_369,N_338);
or U466 (N_466,N_395,N_375);
and U467 (N_467,N_376,N_372);
nand U468 (N_468,N_405,In_318);
and U469 (N_469,N_387,N_411);
nand U470 (N_470,N_390,N_339);
or U471 (N_471,N_316,N_396);
nor U472 (N_472,N_405,N_400);
nand U473 (N_473,N_406,N_389);
and U474 (N_474,N_393,N_404);
nand U475 (N_475,In_328,N_394);
nor U476 (N_476,N_392,N_319);
or U477 (N_477,N_385,N_331);
or U478 (N_478,N_381,N_372);
and U479 (N_479,N_324,N_360);
xor U480 (N_480,N_458,N_465);
nand U481 (N_481,N_436,N_455);
nor U482 (N_482,N_440,N_459);
nand U483 (N_483,N_477,N_431);
nand U484 (N_484,N_442,N_470);
and U485 (N_485,N_427,N_438);
and U486 (N_486,N_426,N_448);
or U487 (N_487,N_453,N_443);
nand U488 (N_488,N_422,N_446);
or U489 (N_489,N_423,N_454);
nand U490 (N_490,N_437,N_474);
xor U491 (N_491,N_441,N_420);
and U492 (N_492,N_435,N_449);
xor U493 (N_493,N_462,N_456);
nor U494 (N_494,N_428,N_468);
or U495 (N_495,N_445,N_472);
and U496 (N_496,N_463,N_447);
and U497 (N_497,N_479,N_476);
xor U498 (N_498,N_473,N_471);
and U499 (N_499,N_460,N_464);
nand U500 (N_500,N_452,N_478);
nor U501 (N_501,N_430,N_432);
or U502 (N_502,N_461,N_469);
or U503 (N_503,N_466,N_421);
nor U504 (N_504,N_429,N_450);
nor U505 (N_505,N_475,N_434);
nor U506 (N_506,N_439,N_425);
and U507 (N_507,N_424,N_467);
nand U508 (N_508,N_433,N_457);
or U509 (N_509,N_444,N_451);
xnor U510 (N_510,N_459,N_428);
nor U511 (N_511,N_435,N_478);
and U512 (N_512,N_423,N_447);
nor U513 (N_513,N_452,N_462);
nor U514 (N_514,N_451,N_454);
and U515 (N_515,N_424,N_470);
nand U516 (N_516,N_442,N_453);
or U517 (N_517,N_463,N_454);
and U518 (N_518,N_445,N_447);
xnor U519 (N_519,N_446,N_449);
or U520 (N_520,N_478,N_429);
xor U521 (N_521,N_450,N_421);
nor U522 (N_522,N_458,N_445);
nand U523 (N_523,N_442,N_451);
nand U524 (N_524,N_471,N_470);
or U525 (N_525,N_473,N_432);
nor U526 (N_526,N_453,N_456);
nor U527 (N_527,N_467,N_435);
xor U528 (N_528,N_471,N_441);
nand U529 (N_529,N_479,N_436);
and U530 (N_530,N_445,N_462);
nand U531 (N_531,N_477,N_465);
xnor U532 (N_532,N_449,N_438);
or U533 (N_533,N_438,N_423);
nor U534 (N_534,N_466,N_427);
and U535 (N_535,N_426,N_421);
nor U536 (N_536,N_449,N_443);
nor U537 (N_537,N_444,N_450);
or U538 (N_538,N_423,N_449);
and U539 (N_539,N_420,N_460);
nor U540 (N_540,N_493,N_539);
nor U541 (N_541,N_498,N_521);
and U542 (N_542,N_513,N_523);
and U543 (N_543,N_519,N_481);
xor U544 (N_544,N_518,N_510);
nor U545 (N_545,N_487,N_530);
and U546 (N_546,N_503,N_489);
nand U547 (N_547,N_497,N_531);
nor U548 (N_548,N_505,N_506);
and U549 (N_549,N_526,N_496);
or U550 (N_550,N_480,N_534);
nor U551 (N_551,N_528,N_501);
and U552 (N_552,N_514,N_516);
nand U553 (N_553,N_484,N_525);
nor U554 (N_554,N_520,N_486);
nand U555 (N_555,N_509,N_500);
or U556 (N_556,N_512,N_504);
or U557 (N_557,N_511,N_522);
xnor U558 (N_558,N_502,N_490);
and U559 (N_559,N_499,N_529);
and U560 (N_560,N_515,N_491);
or U561 (N_561,N_538,N_536);
nor U562 (N_562,N_533,N_488);
nand U563 (N_563,N_485,N_508);
nand U564 (N_564,N_537,N_532);
xor U565 (N_565,N_517,N_535);
nor U566 (N_566,N_507,N_482);
nor U567 (N_567,N_495,N_524);
nor U568 (N_568,N_494,N_492);
xnor U569 (N_569,N_527,N_483);
nand U570 (N_570,N_535,N_518);
nor U571 (N_571,N_481,N_527);
and U572 (N_572,N_521,N_538);
and U573 (N_573,N_512,N_509);
nand U574 (N_574,N_531,N_510);
xor U575 (N_575,N_487,N_512);
nand U576 (N_576,N_526,N_538);
and U577 (N_577,N_484,N_480);
or U578 (N_578,N_508,N_538);
and U579 (N_579,N_486,N_537);
and U580 (N_580,N_495,N_522);
nand U581 (N_581,N_515,N_481);
nor U582 (N_582,N_485,N_539);
xor U583 (N_583,N_487,N_529);
and U584 (N_584,N_529,N_503);
xor U585 (N_585,N_504,N_534);
nand U586 (N_586,N_534,N_517);
and U587 (N_587,N_532,N_530);
nand U588 (N_588,N_518,N_480);
nand U589 (N_589,N_538,N_511);
nand U590 (N_590,N_505,N_496);
and U591 (N_591,N_516,N_519);
nor U592 (N_592,N_532,N_522);
xnor U593 (N_593,N_508,N_528);
nand U594 (N_594,N_524,N_522);
and U595 (N_595,N_492,N_482);
nor U596 (N_596,N_491,N_486);
or U597 (N_597,N_520,N_511);
nor U598 (N_598,N_524,N_513);
nor U599 (N_599,N_529,N_496);
nor U600 (N_600,N_547,N_548);
or U601 (N_601,N_552,N_558);
nor U602 (N_602,N_550,N_559);
nand U603 (N_603,N_541,N_567);
or U604 (N_604,N_580,N_557);
nor U605 (N_605,N_562,N_561);
or U606 (N_606,N_588,N_577);
and U607 (N_607,N_573,N_576);
or U608 (N_608,N_597,N_575);
nand U609 (N_609,N_551,N_595);
nand U610 (N_610,N_590,N_564);
nand U611 (N_611,N_589,N_572);
nand U612 (N_612,N_545,N_598);
or U613 (N_613,N_581,N_543);
nand U614 (N_614,N_586,N_583);
or U615 (N_615,N_579,N_570);
or U616 (N_616,N_594,N_596);
nor U617 (N_617,N_540,N_571);
xor U618 (N_618,N_568,N_563);
or U619 (N_619,N_554,N_591);
xor U620 (N_620,N_578,N_546);
nand U621 (N_621,N_549,N_587);
nand U622 (N_622,N_585,N_566);
nor U623 (N_623,N_599,N_565);
or U624 (N_624,N_593,N_560);
nand U625 (N_625,N_553,N_582);
and U626 (N_626,N_556,N_584);
nand U627 (N_627,N_542,N_555);
or U628 (N_628,N_574,N_544);
or U629 (N_629,N_592,N_569);
or U630 (N_630,N_584,N_581);
and U631 (N_631,N_569,N_566);
and U632 (N_632,N_572,N_585);
nand U633 (N_633,N_595,N_572);
and U634 (N_634,N_544,N_573);
and U635 (N_635,N_598,N_597);
and U636 (N_636,N_552,N_563);
nand U637 (N_637,N_589,N_582);
nand U638 (N_638,N_582,N_576);
xnor U639 (N_639,N_582,N_543);
or U640 (N_640,N_563,N_555);
or U641 (N_641,N_575,N_572);
and U642 (N_642,N_586,N_575);
or U643 (N_643,N_564,N_592);
nor U644 (N_644,N_548,N_572);
xnor U645 (N_645,N_573,N_584);
nand U646 (N_646,N_587,N_578);
or U647 (N_647,N_573,N_563);
or U648 (N_648,N_547,N_569);
nor U649 (N_649,N_583,N_574);
and U650 (N_650,N_588,N_575);
nor U651 (N_651,N_581,N_549);
and U652 (N_652,N_595,N_583);
nor U653 (N_653,N_599,N_552);
or U654 (N_654,N_594,N_576);
nand U655 (N_655,N_552,N_575);
or U656 (N_656,N_592,N_597);
and U657 (N_657,N_585,N_560);
or U658 (N_658,N_540,N_568);
and U659 (N_659,N_549,N_583);
xor U660 (N_660,N_604,N_600);
nor U661 (N_661,N_613,N_608);
and U662 (N_662,N_646,N_633);
and U663 (N_663,N_622,N_615);
and U664 (N_664,N_639,N_624);
nor U665 (N_665,N_630,N_601);
nor U666 (N_666,N_644,N_652);
and U667 (N_667,N_642,N_602);
nand U668 (N_668,N_620,N_626);
nor U669 (N_669,N_659,N_610);
or U670 (N_670,N_636,N_623);
nor U671 (N_671,N_629,N_654);
xor U672 (N_672,N_632,N_638);
or U673 (N_673,N_647,N_617);
and U674 (N_674,N_637,N_627);
or U675 (N_675,N_603,N_614);
xor U676 (N_676,N_653,N_640);
or U677 (N_677,N_635,N_643);
nor U678 (N_678,N_649,N_628);
nor U679 (N_679,N_606,N_609);
or U680 (N_680,N_621,N_619);
and U681 (N_681,N_648,N_650);
and U682 (N_682,N_605,N_655);
nand U683 (N_683,N_645,N_658);
and U684 (N_684,N_607,N_618);
nand U685 (N_685,N_631,N_641);
nand U686 (N_686,N_656,N_657);
and U687 (N_687,N_625,N_634);
xor U688 (N_688,N_612,N_616);
xnor U689 (N_689,N_611,N_651);
nand U690 (N_690,N_606,N_648);
nand U691 (N_691,N_657,N_616);
and U692 (N_692,N_645,N_606);
and U693 (N_693,N_600,N_618);
or U694 (N_694,N_622,N_618);
nor U695 (N_695,N_624,N_604);
or U696 (N_696,N_601,N_658);
nor U697 (N_697,N_627,N_623);
xor U698 (N_698,N_604,N_601);
and U699 (N_699,N_622,N_651);
and U700 (N_700,N_645,N_641);
xnor U701 (N_701,N_633,N_619);
nand U702 (N_702,N_654,N_648);
xor U703 (N_703,N_653,N_620);
and U704 (N_704,N_639,N_610);
or U705 (N_705,N_640,N_601);
nand U706 (N_706,N_619,N_646);
nor U707 (N_707,N_653,N_610);
or U708 (N_708,N_640,N_636);
or U709 (N_709,N_620,N_652);
or U710 (N_710,N_653,N_651);
nor U711 (N_711,N_608,N_642);
nand U712 (N_712,N_649,N_629);
nor U713 (N_713,N_614,N_630);
xor U714 (N_714,N_657,N_650);
or U715 (N_715,N_635,N_653);
and U716 (N_716,N_636,N_602);
or U717 (N_717,N_609,N_637);
nand U718 (N_718,N_651,N_603);
nand U719 (N_719,N_628,N_634);
xor U720 (N_720,N_701,N_663);
and U721 (N_721,N_662,N_714);
and U722 (N_722,N_692,N_677);
nor U723 (N_723,N_667,N_689);
and U724 (N_724,N_703,N_676);
nor U725 (N_725,N_660,N_695);
nor U726 (N_726,N_688,N_718);
nor U727 (N_727,N_671,N_697);
and U728 (N_728,N_680,N_672);
nor U729 (N_729,N_690,N_670);
nor U730 (N_730,N_717,N_674);
and U731 (N_731,N_700,N_693);
nor U732 (N_732,N_687,N_707);
nand U733 (N_733,N_709,N_708);
and U734 (N_734,N_686,N_694);
and U735 (N_735,N_668,N_716);
nor U736 (N_736,N_696,N_705);
nand U737 (N_737,N_685,N_699);
and U738 (N_738,N_711,N_710);
and U739 (N_739,N_683,N_715);
xor U740 (N_740,N_679,N_691);
and U741 (N_741,N_665,N_719);
xnor U742 (N_742,N_713,N_664);
nor U743 (N_743,N_706,N_682);
xor U744 (N_744,N_661,N_712);
and U745 (N_745,N_666,N_673);
and U746 (N_746,N_704,N_675);
nor U747 (N_747,N_669,N_702);
or U748 (N_748,N_681,N_684);
nand U749 (N_749,N_678,N_698);
and U750 (N_750,N_686,N_662);
or U751 (N_751,N_670,N_671);
nand U752 (N_752,N_696,N_679);
and U753 (N_753,N_660,N_694);
nor U754 (N_754,N_685,N_681);
nor U755 (N_755,N_714,N_684);
or U756 (N_756,N_699,N_663);
and U757 (N_757,N_707,N_669);
or U758 (N_758,N_663,N_685);
nand U759 (N_759,N_674,N_706);
and U760 (N_760,N_715,N_679);
nand U761 (N_761,N_703,N_694);
or U762 (N_762,N_680,N_660);
nor U763 (N_763,N_691,N_716);
xnor U764 (N_764,N_714,N_700);
or U765 (N_765,N_678,N_708);
nand U766 (N_766,N_711,N_673);
nand U767 (N_767,N_706,N_704);
nand U768 (N_768,N_676,N_664);
xnor U769 (N_769,N_699,N_669);
or U770 (N_770,N_666,N_670);
xor U771 (N_771,N_670,N_677);
xnor U772 (N_772,N_699,N_705);
nor U773 (N_773,N_710,N_709);
and U774 (N_774,N_692,N_674);
and U775 (N_775,N_673,N_693);
nand U776 (N_776,N_712,N_701);
and U777 (N_777,N_682,N_689);
and U778 (N_778,N_674,N_681);
and U779 (N_779,N_683,N_680);
and U780 (N_780,N_743,N_744);
xor U781 (N_781,N_735,N_745);
and U782 (N_782,N_754,N_779);
and U783 (N_783,N_727,N_750);
and U784 (N_784,N_740,N_766);
or U785 (N_785,N_767,N_731);
and U786 (N_786,N_776,N_763);
xor U787 (N_787,N_771,N_778);
xnor U788 (N_788,N_733,N_737);
or U789 (N_789,N_747,N_724);
or U790 (N_790,N_755,N_736);
and U791 (N_791,N_738,N_762);
or U792 (N_792,N_764,N_726);
nand U793 (N_793,N_732,N_772);
nor U794 (N_794,N_720,N_752);
nor U795 (N_795,N_760,N_770);
or U796 (N_796,N_769,N_742);
nand U797 (N_797,N_739,N_723);
and U798 (N_798,N_721,N_758);
and U799 (N_799,N_768,N_728);
nor U800 (N_800,N_765,N_730);
xnor U801 (N_801,N_756,N_757);
nor U802 (N_802,N_748,N_759);
nor U803 (N_803,N_761,N_753);
nor U804 (N_804,N_741,N_751);
nand U805 (N_805,N_729,N_774);
and U806 (N_806,N_734,N_777);
and U807 (N_807,N_746,N_722);
nand U808 (N_808,N_725,N_773);
nor U809 (N_809,N_775,N_749);
nor U810 (N_810,N_776,N_723);
nand U811 (N_811,N_738,N_772);
and U812 (N_812,N_728,N_738);
or U813 (N_813,N_732,N_744);
or U814 (N_814,N_777,N_725);
or U815 (N_815,N_739,N_741);
or U816 (N_816,N_772,N_752);
nand U817 (N_817,N_762,N_760);
nand U818 (N_818,N_729,N_724);
or U819 (N_819,N_726,N_742);
or U820 (N_820,N_776,N_779);
xor U821 (N_821,N_772,N_764);
or U822 (N_822,N_752,N_728);
nor U823 (N_823,N_770,N_759);
nand U824 (N_824,N_742,N_725);
and U825 (N_825,N_738,N_775);
nand U826 (N_826,N_743,N_771);
and U827 (N_827,N_759,N_738);
or U828 (N_828,N_759,N_741);
nand U829 (N_829,N_758,N_755);
xnor U830 (N_830,N_748,N_732);
or U831 (N_831,N_764,N_724);
nor U832 (N_832,N_721,N_734);
or U833 (N_833,N_737,N_754);
nand U834 (N_834,N_730,N_778);
nand U835 (N_835,N_731,N_770);
and U836 (N_836,N_756,N_754);
or U837 (N_837,N_735,N_723);
nor U838 (N_838,N_776,N_735);
nand U839 (N_839,N_737,N_740);
nand U840 (N_840,N_824,N_815);
and U841 (N_841,N_796,N_838);
and U842 (N_842,N_803,N_825);
or U843 (N_843,N_822,N_823);
nand U844 (N_844,N_814,N_811);
or U845 (N_845,N_787,N_812);
nor U846 (N_846,N_816,N_802);
and U847 (N_847,N_783,N_817);
nand U848 (N_848,N_791,N_788);
or U849 (N_849,N_789,N_820);
and U850 (N_850,N_781,N_828);
nor U851 (N_851,N_813,N_806);
and U852 (N_852,N_829,N_826);
or U853 (N_853,N_784,N_794);
and U854 (N_854,N_834,N_836);
nand U855 (N_855,N_833,N_830);
nor U856 (N_856,N_798,N_818);
or U857 (N_857,N_795,N_821);
nand U858 (N_858,N_800,N_797);
nor U859 (N_859,N_807,N_837);
or U860 (N_860,N_832,N_792);
nor U861 (N_861,N_804,N_805);
nand U862 (N_862,N_808,N_831);
nand U863 (N_863,N_827,N_786);
nor U864 (N_864,N_839,N_809);
or U865 (N_865,N_835,N_819);
nand U866 (N_866,N_801,N_799);
nand U867 (N_867,N_785,N_780);
and U868 (N_868,N_790,N_782);
and U869 (N_869,N_810,N_793);
or U870 (N_870,N_789,N_785);
or U871 (N_871,N_790,N_797);
nor U872 (N_872,N_806,N_812);
nand U873 (N_873,N_788,N_839);
xnor U874 (N_874,N_817,N_793);
and U875 (N_875,N_801,N_812);
nand U876 (N_876,N_794,N_811);
xnor U877 (N_877,N_789,N_835);
and U878 (N_878,N_832,N_805);
nor U879 (N_879,N_804,N_806);
or U880 (N_880,N_787,N_813);
or U881 (N_881,N_830,N_820);
xnor U882 (N_882,N_794,N_806);
nand U883 (N_883,N_787,N_801);
and U884 (N_884,N_838,N_799);
and U885 (N_885,N_809,N_789);
nor U886 (N_886,N_806,N_815);
nor U887 (N_887,N_839,N_787);
nand U888 (N_888,N_828,N_795);
xnor U889 (N_889,N_797,N_799);
nor U890 (N_890,N_789,N_830);
nand U891 (N_891,N_796,N_836);
or U892 (N_892,N_825,N_808);
and U893 (N_893,N_822,N_795);
nor U894 (N_894,N_803,N_807);
nor U895 (N_895,N_780,N_830);
nand U896 (N_896,N_831,N_830);
or U897 (N_897,N_780,N_823);
nand U898 (N_898,N_793,N_826);
and U899 (N_899,N_829,N_832);
and U900 (N_900,N_894,N_844);
xor U901 (N_901,N_878,N_874);
xor U902 (N_902,N_893,N_852);
or U903 (N_903,N_889,N_876);
or U904 (N_904,N_866,N_880);
nand U905 (N_905,N_873,N_860);
or U906 (N_906,N_885,N_892);
nor U907 (N_907,N_845,N_898);
and U908 (N_908,N_862,N_842);
and U909 (N_909,N_850,N_888);
nor U910 (N_910,N_869,N_847);
nand U911 (N_911,N_849,N_890);
nor U912 (N_912,N_858,N_879);
nor U913 (N_913,N_895,N_896);
nor U914 (N_914,N_863,N_841);
and U915 (N_915,N_843,N_897);
nand U916 (N_916,N_848,N_857);
and U917 (N_917,N_899,N_871);
nand U918 (N_918,N_881,N_861);
or U919 (N_919,N_846,N_872);
and U920 (N_920,N_851,N_884);
xor U921 (N_921,N_864,N_865);
or U922 (N_922,N_859,N_854);
nor U923 (N_923,N_882,N_867);
and U924 (N_924,N_840,N_883);
nor U925 (N_925,N_855,N_868);
nor U926 (N_926,N_886,N_887);
or U927 (N_927,N_856,N_877);
or U928 (N_928,N_870,N_875);
nand U929 (N_929,N_853,N_891);
or U930 (N_930,N_892,N_865);
and U931 (N_931,N_885,N_882);
or U932 (N_932,N_881,N_853);
or U933 (N_933,N_866,N_890);
and U934 (N_934,N_891,N_840);
nor U935 (N_935,N_854,N_881);
or U936 (N_936,N_898,N_858);
nor U937 (N_937,N_879,N_891);
or U938 (N_938,N_883,N_856);
nor U939 (N_939,N_869,N_858);
nand U940 (N_940,N_875,N_858);
or U941 (N_941,N_899,N_853);
xnor U942 (N_942,N_887,N_840);
nor U943 (N_943,N_859,N_897);
nand U944 (N_944,N_879,N_865);
nor U945 (N_945,N_871,N_869);
and U946 (N_946,N_850,N_899);
nor U947 (N_947,N_866,N_869);
or U948 (N_948,N_870,N_888);
or U949 (N_949,N_849,N_850);
and U950 (N_950,N_873,N_866);
nand U951 (N_951,N_860,N_895);
nor U952 (N_952,N_868,N_865);
nand U953 (N_953,N_859,N_856);
nor U954 (N_954,N_861,N_849);
or U955 (N_955,N_880,N_864);
nor U956 (N_956,N_877,N_850);
nand U957 (N_957,N_884,N_891);
and U958 (N_958,N_855,N_885);
nor U959 (N_959,N_857,N_894);
and U960 (N_960,N_940,N_908);
nand U961 (N_961,N_952,N_949);
nor U962 (N_962,N_910,N_913);
or U963 (N_963,N_958,N_911);
or U964 (N_964,N_917,N_923);
or U965 (N_965,N_934,N_932);
or U966 (N_966,N_936,N_921);
or U967 (N_967,N_955,N_926);
nor U968 (N_968,N_914,N_950);
nand U969 (N_969,N_945,N_944);
nand U970 (N_970,N_937,N_951);
nor U971 (N_971,N_942,N_941);
xor U972 (N_972,N_918,N_954);
nand U973 (N_973,N_931,N_901);
nand U974 (N_974,N_922,N_930);
xnor U975 (N_975,N_948,N_956);
and U976 (N_976,N_957,N_959);
nand U977 (N_977,N_929,N_935);
and U978 (N_978,N_920,N_900);
xnor U979 (N_979,N_928,N_912);
and U980 (N_980,N_947,N_905);
nor U981 (N_981,N_953,N_919);
or U982 (N_982,N_925,N_927);
nor U983 (N_983,N_924,N_903);
nand U984 (N_984,N_916,N_909);
nor U985 (N_985,N_907,N_915);
xnor U986 (N_986,N_933,N_902);
and U987 (N_987,N_939,N_904);
xnor U988 (N_988,N_943,N_938);
xor U989 (N_989,N_946,N_906);
nand U990 (N_990,N_918,N_912);
xnor U991 (N_991,N_952,N_957);
or U992 (N_992,N_912,N_930);
or U993 (N_993,N_910,N_947);
or U994 (N_994,N_957,N_923);
or U995 (N_995,N_918,N_915);
and U996 (N_996,N_922,N_949);
nor U997 (N_997,N_924,N_923);
or U998 (N_998,N_937,N_911);
or U999 (N_999,N_923,N_914);
and U1000 (N_1000,N_958,N_954);
nor U1001 (N_1001,N_926,N_941);
nor U1002 (N_1002,N_946,N_924);
and U1003 (N_1003,N_946,N_959);
or U1004 (N_1004,N_933,N_946);
or U1005 (N_1005,N_934,N_936);
or U1006 (N_1006,N_957,N_920);
or U1007 (N_1007,N_906,N_915);
nand U1008 (N_1008,N_944,N_907);
and U1009 (N_1009,N_923,N_938);
or U1010 (N_1010,N_951,N_952);
and U1011 (N_1011,N_909,N_948);
nor U1012 (N_1012,N_926,N_952);
nor U1013 (N_1013,N_905,N_938);
and U1014 (N_1014,N_958,N_925);
or U1015 (N_1015,N_902,N_956);
and U1016 (N_1016,N_914,N_943);
and U1017 (N_1017,N_941,N_922);
or U1018 (N_1018,N_901,N_954);
nand U1019 (N_1019,N_927,N_949);
xor U1020 (N_1020,N_960,N_987);
nor U1021 (N_1021,N_992,N_1010);
nor U1022 (N_1022,N_966,N_1008);
nor U1023 (N_1023,N_970,N_1006);
nand U1024 (N_1024,N_974,N_986);
nor U1025 (N_1025,N_962,N_973);
and U1026 (N_1026,N_975,N_990);
nor U1027 (N_1027,N_1018,N_1012);
xor U1028 (N_1028,N_983,N_988);
xnor U1029 (N_1029,N_1016,N_1009);
nand U1030 (N_1030,N_991,N_976);
and U1031 (N_1031,N_961,N_985);
nor U1032 (N_1032,N_971,N_996);
and U1033 (N_1033,N_1003,N_1019);
nand U1034 (N_1034,N_1004,N_978);
nor U1035 (N_1035,N_1015,N_980);
or U1036 (N_1036,N_963,N_979);
and U1037 (N_1037,N_1007,N_984);
nand U1038 (N_1038,N_993,N_1011);
or U1039 (N_1039,N_998,N_1001);
nand U1040 (N_1040,N_977,N_967);
nor U1041 (N_1041,N_968,N_989);
or U1042 (N_1042,N_969,N_994);
or U1043 (N_1043,N_1000,N_972);
or U1044 (N_1044,N_965,N_1014);
or U1045 (N_1045,N_995,N_1005);
or U1046 (N_1046,N_1002,N_982);
nor U1047 (N_1047,N_981,N_964);
nor U1048 (N_1048,N_997,N_1017);
nand U1049 (N_1049,N_1013,N_999);
or U1050 (N_1050,N_989,N_996);
xor U1051 (N_1051,N_961,N_1005);
nand U1052 (N_1052,N_994,N_971);
nor U1053 (N_1053,N_1012,N_1015);
or U1054 (N_1054,N_976,N_1017);
nand U1055 (N_1055,N_996,N_965);
and U1056 (N_1056,N_980,N_1017);
nand U1057 (N_1057,N_974,N_981);
and U1058 (N_1058,N_967,N_1013);
or U1059 (N_1059,N_1012,N_1008);
nor U1060 (N_1060,N_1013,N_980);
nand U1061 (N_1061,N_1011,N_961);
xor U1062 (N_1062,N_1011,N_985);
nand U1063 (N_1063,N_1011,N_1015);
xnor U1064 (N_1064,N_990,N_989);
or U1065 (N_1065,N_974,N_1003);
nand U1066 (N_1066,N_993,N_964);
and U1067 (N_1067,N_961,N_966);
nand U1068 (N_1068,N_999,N_1001);
xnor U1069 (N_1069,N_1016,N_980);
nor U1070 (N_1070,N_993,N_971);
and U1071 (N_1071,N_1016,N_997);
xnor U1072 (N_1072,N_978,N_991);
nor U1073 (N_1073,N_1002,N_1001);
nor U1074 (N_1074,N_1017,N_982);
nand U1075 (N_1075,N_979,N_965);
or U1076 (N_1076,N_1001,N_982);
or U1077 (N_1077,N_985,N_966);
and U1078 (N_1078,N_1012,N_984);
nand U1079 (N_1079,N_1013,N_982);
or U1080 (N_1080,N_1052,N_1048);
or U1081 (N_1081,N_1063,N_1030);
nand U1082 (N_1082,N_1042,N_1074);
or U1083 (N_1083,N_1031,N_1065);
nor U1084 (N_1084,N_1047,N_1045);
nand U1085 (N_1085,N_1072,N_1036);
nor U1086 (N_1086,N_1073,N_1025);
and U1087 (N_1087,N_1044,N_1024);
or U1088 (N_1088,N_1054,N_1027);
nor U1089 (N_1089,N_1071,N_1061);
nand U1090 (N_1090,N_1037,N_1053);
and U1091 (N_1091,N_1079,N_1041);
xnor U1092 (N_1092,N_1051,N_1066);
nand U1093 (N_1093,N_1028,N_1075);
nand U1094 (N_1094,N_1035,N_1020);
nor U1095 (N_1095,N_1068,N_1039);
xor U1096 (N_1096,N_1050,N_1077);
nor U1097 (N_1097,N_1067,N_1078);
nand U1098 (N_1098,N_1043,N_1056);
and U1099 (N_1099,N_1026,N_1060);
nor U1100 (N_1100,N_1033,N_1057);
and U1101 (N_1101,N_1055,N_1064);
or U1102 (N_1102,N_1046,N_1023);
and U1103 (N_1103,N_1049,N_1058);
and U1104 (N_1104,N_1032,N_1029);
xor U1105 (N_1105,N_1040,N_1034);
xnor U1106 (N_1106,N_1022,N_1062);
nor U1107 (N_1107,N_1059,N_1070);
nor U1108 (N_1108,N_1021,N_1038);
nand U1109 (N_1109,N_1069,N_1076);
and U1110 (N_1110,N_1036,N_1063);
nand U1111 (N_1111,N_1065,N_1050);
or U1112 (N_1112,N_1040,N_1035);
nand U1113 (N_1113,N_1045,N_1037);
nor U1114 (N_1114,N_1054,N_1064);
and U1115 (N_1115,N_1034,N_1059);
and U1116 (N_1116,N_1050,N_1074);
nor U1117 (N_1117,N_1073,N_1048);
and U1118 (N_1118,N_1055,N_1022);
nor U1119 (N_1119,N_1054,N_1052);
nand U1120 (N_1120,N_1026,N_1020);
or U1121 (N_1121,N_1062,N_1040);
nand U1122 (N_1122,N_1061,N_1045);
and U1123 (N_1123,N_1058,N_1034);
nand U1124 (N_1124,N_1069,N_1032);
nor U1125 (N_1125,N_1046,N_1058);
xor U1126 (N_1126,N_1073,N_1031);
nor U1127 (N_1127,N_1044,N_1045);
xnor U1128 (N_1128,N_1047,N_1072);
nand U1129 (N_1129,N_1028,N_1022);
and U1130 (N_1130,N_1034,N_1075);
xor U1131 (N_1131,N_1049,N_1023);
nor U1132 (N_1132,N_1022,N_1051);
and U1133 (N_1133,N_1022,N_1073);
nand U1134 (N_1134,N_1064,N_1027);
nor U1135 (N_1135,N_1053,N_1061);
nand U1136 (N_1136,N_1057,N_1051);
and U1137 (N_1137,N_1079,N_1048);
nor U1138 (N_1138,N_1073,N_1052);
xor U1139 (N_1139,N_1061,N_1078);
nand U1140 (N_1140,N_1130,N_1133);
nand U1141 (N_1141,N_1122,N_1115);
or U1142 (N_1142,N_1086,N_1134);
nand U1143 (N_1143,N_1128,N_1091);
xnor U1144 (N_1144,N_1129,N_1104);
nand U1145 (N_1145,N_1111,N_1095);
xnor U1146 (N_1146,N_1102,N_1120);
or U1147 (N_1147,N_1125,N_1110);
and U1148 (N_1148,N_1084,N_1121);
or U1149 (N_1149,N_1096,N_1097);
nor U1150 (N_1150,N_1119,N_1105);
xor U1151 (N_1151,N_1092,N_1116);
nor U1152 (N_1152,N_1139,N_1107);
and U1153 (N_1153,N_1085,N_1117);
nor U1154 (N_1154,N_1082,N_1098);
nand U1155 (N_1155,N_1131,N_1124);
and U1156 (N_1156,N_1112,N_1132);
and U1157 (N_1157,N_1100,N_1108);
or U1158 (N_1158,N_1081,N_1113);
xnor U1159 (N_1159,N_1103,N_1137);
nand U1160 (N_1160,N_1094,N_1118);
nor U1161 (N_1161,N_1126,N_1123);
and U1162 (N_1162,N_1090,N_1106);
or U1163 (N_1163,N_1087,N_1135);
and U1164 (N_1164,N_1138,N_1109);
and U1165 (N_1165,N_1099,N_1136);
nor U1166 (N_1166,N_1101,N_1083);
and U1167 (N_1167,N_1127,N_1088);
or U1168 (N_1168,N_1080,N_1089);
or U1169 (N_1169,N_1114,N_1093);
xor U1170 (N_1170,N_1112,N_1111);
and U1171 (N_1171,N_1131,N_1116);
or U1172 (N_1172,N_1097,N_1108);
nor U1173 (N_1173,N_1092,N_1133);
nand U1174 (N_1174,N_1123,N_1102);
or U1175 (N_1175,N_1119,N_1133);
nand U1176 (N_1176,N_1122,N_1080);
nand U1177 (N_1177,N_1132,N_1090);
nor U1178 (N_1178,N_1093,N_1118);
or U1179 (N_1179,N_1099,N_1087);
nor U1180 (N_1180,N_1108,N_1128);
nor U1181 (N_1181,N_1104,N_1106);
nand U1182 (N_1182,N_1119,N_1115);
or U1183 (N_1183,N_1104,N_1130);
nor U1184 (N_1184,N_1086,N_1108);
and U1185 (N_1185,N_1098,N_1108);
and U1186 (N_1186,N_1108,N_1091);
and U1187 (N_1187,N_1114,N_1088);
nor U1188 (N_1188,N_1114,N_1119);
nor U1189 (N_1189,N_1089,N_1118);
nor U1190 (N_1190,N_1086,N_1126);
nand U1191 (N_1191,N_1101,N_1112);
nor U1192 (N_1192,N_1088,N_1111);
and U1193 (N_1193,N_1130,N_1084);
nand U1194 (N_1194,N_1133,N_1088);
nand U1195 (N_1195,N_1102,N_1082);
and U1196 (N_1196,N_1082,N_1088);
xor U1197 (N_1197,N_1104,N_1123);
and U1198 (N_1198,N_1097,N_1128);
xor U1199 (N_1199,N_1121,N_1091);
and U1200 (N_1200,N_1164,N_1188);
nand U1201 (N_1201,N_1163,N_1186);
nand U1202 (N_1202,N_1157,N_1192);
nor U1203 (N_1203,N_1170,N_1160);
and U1204 (N_1204,N_1151,N_1142);
or U1205 (N_1205,N_1149,N_1177);
nor U1206 (N_1206,N_1171,N_1155);
nor U1207 (N_1207,N_1181,N_1145);
or U1208 (N_1208,N_1175,N_1174);
nand U1209 (N_1209,N_1180,N_1189);
and U1210 (N_1210,N_1150,N_1185);
nor U1211 (N_1211,N_1153,N_1154);
and U1212 (N_1212,N_1197,N_1162);
nor U1213 (N_1213,N_1173,N_1141);
nand U1214 (N_1214,N_1159,N_1167);
and U1215 (N_1215,N_1191,N_1156);
xor U1216 (N_1216,N_1187,N_1194);
xnor U1217 (N_1217,N_1172,N_1182);
nand U1218 (N_1218,N_1148,N_1190);
and U1219 (N_1219,N_1152,N_1179);
nand U1220 (N_1220,N_1158,N_1199);
and U1221 (N_1221,N_1144,N_1178);
or U1222 (N_1222,N_1143,N_1146);
and U1223 (N_1223,N_1183,N_1184);
or U1224 (N_1224,N_1198,N_1168);
nand U1225 (N_1225,N_1165,N_1161);
nor U1226 (N_1226,N_1195,N_1147);
and U1227 (N_1227,N_1193,N_1196);
and U1228 (N_1228,N_1140,N_1176);
and U1229 (N_1229,N_1169,N_1166);
or U1230 (N_1230,N_1169,N_1145);
and U1231 (N_1231,N_1153,N_1162);
and U1232 (N_1232,N_1191,N_1194);
or U1233 (N_1233,N_1159,N_1149);
or U1234 (N_1234,N_1186,N_1169);
or U1235 (N_1235,N_1171,N_1185);
nor U1236 (N_1236,N_1144,N_1185);
nand U1237 (N_1237,N_1167,N_1181);
nand U1238 (N_1238,N_1177,N_1195);
or U1239 (N_1239,N_1175,N_1141);
nor U1240 (N_1240,N_1141,N_1181);
and U1241 (N_1241,N_1145,N_1191);
nand U1242 (N_1242,N_1174,N_1151);
and U1243 (N_1243,N_1147,N_1180);
or U1244 (N_1244,N_1179,N_1181);
nand U1245 (N_1245,N_1148,N_1187);
or U1246 (N_1246,N_1157,N_1195);
xnor U1247 (N_1247,N_1159,N_1180);
nand U1248 (N_1248,N_1164,N_1183);
xnor U1249 (N_1249,N_1143,N_1183);
and U1250 (N_1250,N_1173,N_1199);
and U1251 (N_1251,N_1171,N_1153);
and U1252 (N_1252,N_1178,N_1184);
or U1253 (N_1253,N_1184,N_1177);
nand U1254 (N_1254,N_1187,N_1186);
or U1255 (N_1255,N_1154,N_1183);
nor U1256 (N_1256,N_1184,N_1168);
xnor U1257 (N_1257,N_1198,N_1199);
nor U1258 (N_1258,N_1176,N_1167);
nand U1259 (N_1259,N_1167,N_1160);
or U1260 (N_1260,N_1210,N_1215);
and U1261 (N_1261,N_1219,N_1201);
and U1262 (N_1262,N_1250,N_1239);
nor U1263 (N_1263,N_1223,N_1206);
and U1264 (N_1264,N_1212,N_1238);
and U1265 (N_1265,N_1229,N_1205);
nand U1266 (N_1266,N_1257,N_1222);
nand U1267 (N_1267,N_1243,N_1211);
or U1268 (N_1268,N_1214,N_1259);
nand U1269 (N_1269,N_1233,N_1253);
nand U1270 (N_1270,N_1240,N_1220);
nor U1271 (N_1271,N_1207,N_1232);
nand U1272 (N_1272,N_1230,N_1221);
nor U1273 (N_1273,N_1209,N_1216);
nand U1274 (N_1274,N_1245,N_1225);
or U1275 (N_1275,N_1246,N_1256);
nor U1276 (N_1276,N_1217,N_1248);
nor U1277 (N_1277,N_1227,N_1247);
and U1278 (N_1278,N_1244,N_1249);
or U1279 (N_1279,N_1236,N_1213);
nor U1280 (N_1280,N_1202,N_1235);
nand U1281 (N_1281,N_1241,N_1218);
nand U1282 (N_1282,N_1258,N_1204);
and U1283 (N_1283,N_1252,N_1251);
and U1284 (N_1284,N_1242,N_1255);
nor U1285 (N_1285,N_1208,N_1231);
and U1286 (N_1286,N_1200,N_1254);
nor U1287 (N_1287,N_1224,N_1234);
and U1288 (N_1288,N_1237,N_1203);
nand U1289 (N_1289,N_1226,N_1228);
or U1290 (N_1290,N_1212,N_1218);
nand U1291 (N_1291,N_1258,N_1252);
xnor U1292 (N_1292,N_1231,N_1247);
and U1293 (N_1293,N_1227,N_1244);
nand U1294 (N_1294,N_1220,N_1219);
nor U1295 (N_1295,N_1218,N_1221);
nor U1296 (N_1296,N_1252,N_1243);
nor U1297 (N_1297,N_1235,N_1228);
and U1298 (N_1298,N_1228,N_1211);
and U1299 (N_1299,N_1250,N_1234);
or U1300 (N_1300,N_1204,N_1233);
or U1301 (N_1301,N_1233,N_1208);
nor U1302 (N_1302,N_1247,N_1241);
or U1303 (N_1303,N_1218,N_1244);
nand U1304 (N_1304,N_1206,N_1209);
or U1305 (N_1305,N_1213,N_1201);
and U1306 (N_1306,N_1254,N_1232);
or U1307 (N_1307,N_1236,N_1217);
nor U1308 (N_1308,N_1258,N_1234);
and U1309 (N_1309,N_1245,N_1217);
or U1310 (N_1310,N_1227,N_1256);
or U1311 (N_1311,N_1239,N_1224);
nand U1312 (N_1312,N_1229,N_1210);
nand U1313 (N_1313,N_1242,N_1238);
or U1314 (N_1314,N_1233,N_1225);
nand U1315 (N_1315,N_1212,N_1254);
nor U1316 (N_1316,N_1200,N_1221);
nor U1317 (N_1317,N_1213,N_1251);
or U1318 (N_1318,N_1220,N_1233);
nand U1319 (N_1319,N_1226,N_1239);
nand U1320 (N_1320,N_1263,N_1288);
nand U1321 (N_1321,N_1298,N_1317);
nor U1322 (N_1322,N_1264,N_1292);
xor U1323 (N_1323,N_1268,N_1294);
and U1324 (N_1324,N_1319,N_1303);
nor U1325 (N_1325,N_1287,N_1316);
or U1326 (N_1326,N_1290,N_1265);
nand U1327 (N_1327,N_1299,N_1286);
nand U1328 (N_1328,N_1289,N_1270);
nor U1329 (N_1329,N_1310,N_1275);
or U1330 (N_1330,N_1295,N_1279);
or U1331 (N_1331,N_1273,N_1269);
xnor U1332 (N_1332,N_1282,N_1284);
or U1333 (N_1333,N_1283,N_1309);
nor U1334 (N_1334,N_1278,N_1306);
and U1335 (N_1335,N_1267,N_1296);
or U1336 (N_1336,N_1272,N_1312);
or U1337 (N_1337,N_1314,N_1271);
nor U1338 (N_1338,N_1281,N_1280);
or U1339 (N_1339,N_1293,N_1305);
nor U1340 (N_1340,N_1262,N_1291);
nand U1341 (N_1341,N_1313,N_1311);
and U1342 (N_1342,N_1276,N_1302);
or U1343 (N_1343,N_1297,N_1285);
or U1344 (N_1344,N_1304,N_1300);
and U1345 (N_1345,N_1315,N_1274);
and U1346 (N_1346,N_1260,N_1318);
nor U1347 (N_1347,N_1277,N_1307);
and U1348 (N_1348,N_1301,N_1261);
and U1349 (N_1349,N_1308,N_1266);
nand U1350 (N_1350,N_1311,N_1310);
or U1351 (N_1351,N_1318,N_1270);
and U1352 (N_1352,N_1281,N_1295);
nand U1353 (N_1353,N_1308,N_1317);
nor U1354 (N_1354,N_1286,N_1279);
nor U1355 (N_1355,N_1303,N_1264);
and U1356 (N_1356,N_1276,N_1301);
nand U1357 (N_1357,N_1273,N_1278);
nor U1358 (N_1358,N_1315,N_1271);
or U1359 (N_1359,N_1262,N_1265);
or U1360 (N_1360,N_1302,N_1281);
nand U1361 (N_1361,N_1267,N_1314);
or U1362 (N_1362,N_1279,N_1267);
or U1363 (N_1363,N_1269,N_1316);
nand U1364 (N_1364,N_1281,N_1273);
and U1365 (N_1365,N_1319,N_1283);
or U1366 (N_1366,N_1263,N_1302);
nand U1367 (N_1367,N_1285,N_1289);
nand U1368 (N_1368,N_1319,N_1314);
or U1369 (N_1369,N_1297,N_1316);
and U1370 (N_1370,N_1275,N_1293);
xor U1371 (N_1371,N_1297,N_1313);
and U1372 (N_1372,N_1272,N_1268);
nor U1373 (N_1373,N_1318,N_1266);
and U1374 (N_1374,N_1302,N_1269);
and U1375 (N_1375,N_1290,N_1261);
nor U1376 (N_1376,N_1273,N_1314);
and U1377 (N_1377,N_1304,N_1275);
nand U1378 (N_1378,N_1265,N_1293);
nand U1379 (N_1379,N_1302,N_1310);
nand U1380 (N_1380,N_1371,N_1340);
xnor U1381 (N_1381,N_1344,N_1338);
nor U1382 (N_1382,N_1347,N_1360);
nand U1383 (N_1383,N_1362,N_1370);
nand U1384 (N_1384,N_1349,N_1379);
nor U1385 (N_1385,N_1335,N_1374);
nor U1386 (N_1386,N_1327,N_1350);
xor U1387 (N_1387,N_1341,N_1378);
nor U1388 (N_1388,N_1323,N_1328);
nand U1389 (N_1389,N_1357,N_1348);
and U1390 (N_1390,N_1377,N_1330);
nand U1391 (N_1391,N_1332,N_1333);
or U1392 (N_1392,N_1342,N_1354);
nor U1393 (N_1393,N_1345,N_1337);
nor U1394 (N_1394,N_1356,N_1366);
and U1395 (N_1395,N_1339,N_1369);
nand U1396 (N_1396,N_1355,N_1352);
and U1397 (N_1397,N_1363,N_1320);
nor U1398 (N_1398,N_1367,N_1334);
nor U1399 (N_1399,N_1358,N_1364);
or U1400 (N_1400,N_1372,N_1361);
or U1401 (N_1401,N_1326,N_1325);
or U1402 (N_1402,N_1321,N_1353);
nor U1403 (N_1403,N_1375,N_1346);
nor U1404 (N_1404,N_1324,N_1343);
and U1405 (N_1405,N_1322,N_1365);
xor U1406 (N_1406,N_1331,N_1359);
or U1407 (N_1407,N_1336,N_1368);
and U1408 (N_1408,N_1329,N_1373);
nand U1409 (N_1409,N_1376,N_1351);
or U1410 (N_1410,N_1358,N_1329);
or U1411 (N_1411,N_1320,N_1337);
nor U1412 (N_1412,N_1344,N_1334);
and U1413 (N_1413,N_1332,N_1352);
and U1414 (N_1414,N_1323,N_1342);
and U1415 (N_1415,N_1327,N_1329);
xnor U1416 (N_1416,N_1333,N_1322);
and U1417 (N_1417,N_1379,N_1370);
nand U1418 (N_1418,N_1352,N_1328);
xnor U1419 (N_1419,N_1356,N_1371);
nand U1420 (N_1420,N_1344,N_1337);
xor U1421 (N_1421,N_1342,N_1364);
nor U1422 (N_1422,N_1340,N_1342);
and U1423 (N_1423,N_1324,N_1367);
nand U1424 (N_1424,N_1343,N_1374);
nor U1425 (N_1425,N_1363,N_1366);
nor U1426 (N_1426,N_1366,N_1370);
nor U1427 (N_1427,N_1341,N_1351);
nor U1428 (N_1428,N_1378,N_1365);
nor U1429 (N_1429,N_1361,N_1359);
or U1430 (N_1430,N_1325,N_1351);
or U1431 (N_1431,N_1320,N_1375);
nand U1432 (N_1432,N_1376,N_1354);
and U1433 (N_1433,N_1328,N_1371);
and U1434 (N_1434,N_1329,N_1359);
and U1435 (N_1435,N_1329,N_1361);
and U1436 (N_1436,N_1340,N_1330);
nand U1437 (N_1437,N_1371,N_1368);
or U1438 (N_1438,N_1377,N_1320);
or U1439 (N_1439,N_1374,N_1333);
or U1440 (N_1440,N_1407,N_1409);
or U1441 (N_1441,N_1384,N_1391);
and U1442 (N_1442,N_1426,N_1393);
xnor U1443 (N_1443,N_1429,N_1405);
nand U1444 (N_1444,N_1427,N_1400);
nand U1445 (N_1445,N_1439,N_1401);
or U1446 (N_1446,N_1399,N_1403);
and U1447 (N_1447,N_1423,N_1398);
and U1448 (N_1448,N_1412,N_1385);
and U1449 (N_1449,N_1438,N_1434);
nand U1450 (N_1450,N_1411,N_1437);
or U1451 (N_1451,N_1432,N_1414);
or U1452 (N_1452,N_1431,N_1421);
or U1453 (N_1453,N_1386,N_1420);
xnor U1454 (N_1454,N_1382,N_1389);
nand U1455 (N_1455,N_1404,N_1410);
and U1456 (N_1456,N_1435,N_1380);
nand U1457 (N_1457,N_1418,N_1394);
and U1458 (N_1458,N_1402,N_1397);
and U1459 (N_1459,N_1428,N_1415);
nand U1460 (N_1460,N_1388,N_1419);
nand U1461 (N_1461,N_1422,N_1413);
nor U1462 (N_1462,N_1390,N_1408);
nand U1463 (N_1463,N_1406,N_1416);
nor U1464 (N_1464,N_1387,N_1396);
or U1465 (N_1465,N_1430,N_1424);
and U1466 (N_1466,N_1436,N_1381);
nand U1467 (N_1467,N_1433,N_1395);
or U1468 (N_1468,N_1392,N_1425);
and U1469 (N_1469,N_1383,N_1417);
nand U1470 (N_1470,N_1414,N_1391);
nand U1471 (N_1471,N_1412,N_1408);
nand U1472 (N_1472,N_1404,N_1382);
and U1473 (N_1473,N_1408,N_1405);
nand U1474 (N_1474,N_1431,N_1400);
or U1475 (N_1475,N_1407,N_1408);
and U1476 (N_1476,N_1411,N_1383);
or U1477 (N_1477,N_1434,N_1410);
and U1478 (N_1478,N_1419,N_1416);
and U1479 (N_1479,N_1397,N_1382);
nor U1480 (N_1480,N_1386,N_1394);
and U1481 (N_1481,N_1423,N_1424);
and U1482 (N_1482,N_1384,N_1426);
and U1483 (N_1483,N_1380,N_1416);
and U1484 (N_1484,N_1396,N_1385);
nor U1485 (N_1485,N_1394,N_1388);
xnor U1486 (N_1486,N_1421,N_1386);
nand U1487 (N_1487,N_1384,N_1381);
xnor U1488 (N_1488,N_1406,N_1399);
or U1489 (N_1489,N_1397,N_1434);
and U1490 (N_1490,N_1423,N_1409);
nand U1491 (N_1491,N_1380,N_1401);
and U1492 (N_1492,N_1417,N_1427);
xor U1493 (N_1493,N_1387,N_1397);
nor U1494 (N_1494,N_1389,N_1405);
or U1495 (N_1495,N_1403,N_1408);
nand U1496 (N_1496,N_1412,N_1438);
or U1497 (N_1497,N_1420,N_1411);
and U1498 (N_1498,N_1382,N_1434);
and U1499 (N_1499,N_1392,N_1390);
and U1500 (N_1500,N_1449,N_1442);
and U1501 (N_1501,N_1477,N_1487);
nand U1502 (N_1502,N_1467,N_1447);
nor U1503 (N_1503,N_1455,N_1476);
or U1504 (N_1504,N_1471,N_1499);
and U1505 (N_1505,N_1481,N_1458);
and U1506 (N_1506,N_1492,N_1496);
nor U1507 (N_1507,N_1479,N_1463);
or U1508 (N_1508,N_1443,N_1444);
nor U1509 (N_1509,N_1472,N_1491);
and U1510 (N_1510,N_1450,N_1453);
or U1511 (N_1511,N_1441,N_1493);
nand U1512 (N_1512,N_1462,N_1484);
nand U1513 (N_1513,N_1488,N_1475);
and U1514 (N_1514,N_1497,N_1469);
nor U1515 (N_1515,N_1489,N_1459);
nand U1516 (N_1516,N_1468,N_1483);
or U1517 (N_1517,N_1445,N_1495);
nand U1518 (N_1518,N_1490,N_1486);
xor U1519 (N_1519,N_1474,N_1473);
nand U1520 (N_1520,N_1465,N_1456);
nand U1521 (N_1521,N_1466,N_1494);
and U1522 (N_1522,N_1498,N_1480);
nor U1523 (N_1523,N_1451,N_1461);
or U1524 (N_1524,N_1457,N_1482);
nand U1525 (N_1525,N_1448,N_1452);
xnor U1526 (N_1526,N_1478,N_1446);
nand U1527 (N_1527,N_1485,N_1470);
and U1528 (N_1528,N_1454,N_1464);
and U1529 (N_1529,N_1460,N_1440);
nand U1530 (N_1530,N_1458,N_1478);
and U1531 (N_1531,N_1485,N_1491);
and U1532 (N_1532,N_1451,N_1450);
nor U1533 (N_1533,N_1498,N_1453);
nand U1534 (N_1534,N_1463,N_1498);
and U1535 (N_1535,N_1476,N_1483);
nor U1536 (N_1536,N_1468,N_1488);
and U1537 (N_1537,N_1473,N_1468);
or U1538 (N_1538,N_1477,N_1469);
nor U1539 (N_1539,N_1479,N_1488);
or U1540 (N_1540,N_1456,N_1485);
nand U1541 (N_1541,N_1453,N_1462);
nor U1542 (N_1542,N_1452,N_1494);
nand U1543 (N_1543,N_1446,N_1484);
xor U1544 (N_1544,N_1486,N_1499);
and U1545 (N_1545,N_1454,N_1471);
xnor U1546 (N_1546,N_1494,N_1444);
xnor U1547 (N_1547,N_1442,N_1455);
and U1548 (N_1548,N_1443,N_1450);
nand U1549 (N_1549,N_1478,N_1465);
or U1550 (N_1550,N_1482,N_1471);
nor U1551 (N_1551,N_1455,N_1478);
or U1552 (N_1552,N_1449,N_1447);
and U1553 (N_1553,N_1456,N_1493);
or U1554 (N_1554,N_1487,N_1452);
nor U1555 (N_1555,N_1479,N_1459);
nand U1556 (N_1556,N_1460,N_1464);
xor U1557 (N_1557,N_1460,N_1472);
or U1558 (N_1558,N_1492,N_1443);
or U1559 (N_1559,N_1495,N_1447);
xnor U1560 (N_1560,N_1511,N_1503);
and U1561 (N_1561,N_1536,N_1501);
or U1562 (N_1562,N_1557,N_1547);
and U1563 (N_1563,N_1517,N_1526);
nand U1564 (N_1564,N_1516,N_1520);
or U1565 (N_1565,N_1538,N_1504);
nand U1566 (N_1566,N_1523,N_1543);
and U1567 (N_1567,N_1540,N_1550);
nor U1568 (N_1568,N_1525,N_1558);
nor U1569 (N_1569,N_1500,N_1531);
or U1570 (N_1570,N_1551,N_1522);
and U1571 (N_1571,N_1502,N_1506);
nand U1572 (N_1572,N_1546,N_1544);
and U1573 (N_1573,N_1553,N_1535);
xor U1574 (N_1574,N_1510,N_1527);
or U1575 (N_1575,N_1534,N_1521);
or U1576 (N_1576,N_1513,N_1533);
nand U1577 (N_1577,N_1549,N_1518);
nor U1578 (N_1578,N_1554,N_1528);
and U1579 (N_1579,N_1539,N_1542);
and U1580 (N_1580,N_1537,N_1509);
or U1581 (N_1581,N_1541,N_1552);
and U1582 (N_1582,N_1548,N_1515);
nor U1583 (N_1583,N_1508,N_1529);
nand U1584 (N_1584,N_1514,N_1545);
nand U1585 (N_1585,N_1524,N_1532);
and U1586 (N_1586,N_1556,N_1512);
nor U1587 (N_1587,N_1530,N_1559);
nor U1588 (N_1588,N_1555,N_1519);
or U1589 (N_1589,N_1507,N_1505);
xor U1590 (N_1590,N_1521,N_1523);
nor U1591 (N_1591,N_1548,N_1518);
or U1592 (N_1592,N_1538,N_1505);
and U1593 (N_1593,N_1553,N_1529);
and U1594 (N_1594,N_1559,N_1542);
and U1595 (N_1595,N_1539,N_1509);
and U1596 (N_1596,N_1549,N_1511);
nand U1597 (N_1597,N_1546,N_1530);
or U1598 (N_1598,N_1521,N_1558);
and U1599 (N_1599,N_1558,N_1537);
nor U1600 (N_1600,N_1504,N_1510);
or U1601 (N_1601,N_1542,N_1557);
nand U1602 (N_1602,N_1538,N_1553);
or U1603 (N_1603,N_1552,N_1500);
xnor U1604 (N_1604,N_1558,N_1519);
and U1605 (N_1605,N_1517,N_1553);
or U1606 (N_1606,N_1511,N_1537);
nor U1607 (N_1607,N_1538,N_1502);
or U1608 (N_1608,N_1503,N_1522);
nand U1609 (N_1609,N_1552,N_1531);
nand U1610 (N_1610,N_1538,N_1506);
or U1611 (N_1611,N_1551,N_1526);
nor U1612 (N_1612,N_1515,N_1551);
and U1613 (N_1613,N_1546,N_1503);
xor U1614 (N_1614,N_1527,N_1519);
nand U1615 (N_1615,N_1537,N_1505);
xnor U1616 (N_1616,N_1505,N_1554);
nor U1617 (N_1617,N_1528,N_1521);
nand U1618 (N_1618,N_1518,N_1529);
and U1619 (N_1619,N_1553,N_1555);
and U1620 (N_1620,N_1603,N_1617);
or U1621 (N_1621,N_1575,N_1563);
nor U1622 (N_1622,N_1594,N_1611);
or U1623 (N_1623,N_1583,N_1596);
or U1624 (N_1624,N_1604,N_1577);
nand U1625 (N_1625,N_1586,N_1592);
and U1626 (N_1626,N_1610,N_1560);
or U1627 (N_1627,N_1564,N_1590);
and U1628 (N_1628,N_1567,N_1566);
or U1629 (N_1629,N_1576,N_1599);
nand U1630 (N_1630,N_1578,N_1589);
and U1631 (N_1631,N_1614,N_1595);
nor U1632 (N_1632,N_1608,N_1619);
nand U1633 (N_1633,N_1618,N_1601);
nand U1634 (N_1634,N_1609,N_1591);
nor U1635 (N_1635,N_1572,N_1612);
xnor U1636 (N_1636,N_1561,N_1569);
and U1637 (N_1637,N_1616,N_1579);
nor U1638 (N_1638,N_1580,N_1573);
nor U1639 (N_1639,N_1598,N_1574);
or U1640 (N_1640,N_1605,N_1585);
nand U1641 (N_1641,N_1582,N_1593);
and U1642 (N_1642,N_1581,N_1607);
or U1643 (N_1643,N_1565,N_1602);
nor U1644 (N_1644,N_1568,N_1562);
or U1645 (N_1645,N_1588,N_1584);
nand U1646 (N_1646,N_1600,N_1587);
xnor U1647 (N_1647,N_1615,N_1570);
or U1648 (N_1648,N_1597,N_1613);
and U1649 (N_1649,N_1606,N_1571);
and U1650 (N_1650,N_1576,N_1583);
nor U1651 (N_1651,N_1566,N_1590);
nand U1652 (N_1652,N_1582,N_1597);
nor U1653 (N_1653,N_1603,N_1586);
nand U1654 (N_1654,N_1608,N_1598);
nand U1655 (N_1655,N_1566,N_1618);
and U1656 (N_1656,N_1586,N_1562);
nor U1657 (N_1657,N_1574,N_1612);
and U1658 (N_1658,N_1603,N_1604);
and U1659 (N_1659,N_1569,N_1618);
and U1660 (N_1660,N_1606,N_1589);
nor U1661 (N_1661,N_1612,N_1591);
and U1662 (N_1662,N_1605,N_1577);
nor U1663 (N_1663,N_1575,N_1614);
nor U1664 (N_1664,N_1594,N_1561);
or U1665 (N_1665,N_1567,N_1596);
or U1666 (N_1666,N_1568,N_1610);
or U1667 (N_1667,N_1580,N_1586);
xor U1668 (N_1668,N_1579,N_1581);
nor U1669 (N_1669,N_1568,N_1576);
nor U1670 (N_1670,N_1580,N_1615);
or U1671 (N_1671,N_1601,N_1562);
or U1672 (N_1672,N_1600,N_1570);
or U1673 (N_1673,N_1598,N_1576);
and U1674 (N_1674,N_1590,N_1565);
or U1675 (N_1675,N_1591,N_1560);
nand U1676 (N_1676,N_1616,N_1605);
or U1677 (N_1677,N_1585,N_1580);
nand U1678 (N_1678,N_1615,N_1590);
and U1679 (N_1679,N_1604,N_1578);
nand U1680 (N_1680,N_1632,N_1660);
or U1681 (N_1681,N_1642,N_1637);
xor U1682 (N_1682,N_1638,N_1627);
or U1683 (N_1683,N_1652,N_1670);
or U1684 (N_1684,N_1658,N_1633);
and U1685 (N_1685,N_1657,N_1664);
nor U1686 (N_1686,N_1661,N_1651);
or U1687 (N_1687,N_1675,N_1629);
or U1688 (N_1688,N_1626,N_1656);
or U1689 (N_1689,N_1665,N_1648);
nor U1690 (N_1690,N_1640,N_1659);
or U1691 (N_1691,N_1667,N_1644);
nand U1692 (N_1692,N_1635,N_1639);
or U1693 (N_1693,N_1679,N_1636);
or U1694 (N_1694,N_1643,N_1676);
xnor U1695 (N_1695,N_1671,N_1674);
or U1696 (N_1696,N_1641,N_1677);
nor U1697 (N_1697,N_1622,N_1650);
and U1698 (N_1698,N_1673,N_1631);
or U1699 (N_1699,N_1663,N_1623);
and U1700 (N_1700,N_1653,N_1620);
nor U1701 (N_1701,N_1630,N_1678);
or U1702 (N_1702,N_1624,N_1649);
nor U1703 (N_1703,N_1669,N_1646);
nor U1704 (N_1704,N_1621,N_1668);
nand U1705 (N_1705,N_1647,N_1666);
or U1706 (N_1706,N_1672,N_1655);
or U1707 (N_1707,N_1634,N_1662);
and U1708 (N_1708,N_1654,N_1628);
xor U1709 (N_1709,N_1625,N_1645);
nor U1710 (N_1710,N_1647,N_1624);
or U1711 (N_1711,N_1673,N_1645);
and U1712 (N_1712,N_1656,N_1661);
and U1713 (N_1713,N_1659,N_1633);
nor U1714 (N_1714,N_1665,N_1658);
nand U1715 (N_1715,N_1674,N_1667);
or U1716 (N_1716,N_1626,N_1641);
and U1717 (N_1717,N_1632,N_1662);
nand U1718 (N_1718,N_1640,N_1637);
nand U1719 (N_1719,N_1670,N_1627);
or U1720 (N_1720,N_1679,N_1670);
nand U1721 (N_1721,N_1660,N_1653);
and U1722 (N_1722,N_1641,N_1669);
nand U1723 (N_1723,N_1641,N_1638);
nor U1724 (N_1724,N_1645,N_1634);
nand U1725 (N_1725,N_1667,N_1656);
nand U1726 (N_1726,N_1648,N_1625);
nor U1727 (N_1727,N_1666,N_1672);
and U1728 (N_1728,N_1658,N_1660);
and U1729 (N_1729,N_1634,N_1621);
nor U1730 (N_1730,N_1663,N_1636);
or U1731 (N_1731,N_1662,N_1642);
nor U1732 (N_1732,N_1646,N_1620);
xnor U1733 (N_1733,N_1632,N_1659);
and U1734 (N_1734,N_1632,N_1634);
or U1735 (N_1735,N_1660,N_1622);
and U1736 (N_1736,N_1651,N_1679);
nor U1737 (N_1737,N_1657,N_1641);
or U1738 (N_1738,N_1668,N_1669);
nor U1739 (N_1739,N_1640,N_1652);
xnor U1740 (N_1740,N_1738,N_1736);
nand U1741 (N_1741,N_1739,N_1734);
nand U1742 (N_1742,N_1731,N_1708);
nor U1743 (N_1743,N_1711,N_1727);
or U1744 (N_1744,N_1712,N_1720);
xnor U1745 (N_1745,N_1682,N_1699);
nand U1746 (N_1746,N_1713,N_1721);
nor U1747 (N_1747,N_1722,N_1701);
and U1748 (N_1748,N_1687,N_1715);
and U1749 (N_1749,N_1709,N_1717);
nand U1750 (N_1750,N_1680,N_1697);
and U1751 (N_1751,N_1698,N_1690);
nand U1752 (N_1752,N_1696,N_1732);
nand U1753 (N_1753,N_1694,N_1707);
and U1754 (N_1754,N_1688,N_1704);
and U1755 (N_1755,N_1706,N_1729);
xor U1756 (N_1756,N_1725,N_1689);
nand U1757 (N_1757,N_1705,N_1726);
nor U1758 (N_1758,N_1695,N_1691);
nand U1759 (N_1759,N_1728,N_1685);
nand U1760 (N_1760,N_1714,N_1710);
nand U1761 (N_1761,N_1730,N_1681);
and U1762 (N_1762,N_1684,N_1703);
and U1763 (N_1763,N_1735,N_1686);
nand U1764 (N_1764,N_1700,N_1724);
xor U1765 (N_1765,N_1692,N_1716);
nand U1766 (N_1766,N_1683,N_1702);
or U1767 (N_1767,N_1693,N_1723);
or U1768 (N_1768,N_1733,N_1719);
nor U1769 (N_1769,N_1737,N_1718);
or U1770 (N_1770,N_1715,N_1683);
or U1771 (N_1771,N_1735,N_1721);
and U1772 (N_1772,N_1684,N_1683);
or U1773 (N_1773,N_1739,N_1693);
or U1774 (N_1774,N_1708,N_1736);
xor U1775 (N_1775,N_1733,N_1711);
or U1776 (N_1776,N_1688,N_1712);
xor U1777 (N_1777,N_1733,N_1685);
and U1778 (N_1778,N_1737,N_1728);
nor U1779 (N_1779,N_1734,N_1735);
nand U1780 (N_1780,N_1725,N_1714);
nor U1781 (N_1781,N_1713,N_1709);
xnor U1782 (N_1782,N_1691,N_1728);
and U1783 (N_1783,N_1738,N_1721);
nand U1784 (N_1784,N_1693,N_1733);
and U1785 (N_1785,N_1727,N_1693);
or U1786 (N_1786,N_1695,N_1719);
nor U1787 (N_1787,N_1707,N_1728);
or U1788 (N_1788,N_1731,N_1714);
and U1789 (N_1789,N_1716,N_1727);
nor U1790 (N_1790,N_1710,N_1682);
nand U1791 (N_1791,N_1700,N_1689);
nand U1792 (N_1792,N_1738,N_1688);
nor U1793 (N_1793,N_1702,N_1690);
nor U1794 (N_1794,N_1706,N_1683);
xor U1795 (N_1795,N_1717,N_1726);
nand U1796 (N_1796,N_1717,N_1712);
and U1797 (N_1797,N_1718,N_1725);
nor U1798 (N_1798,N_1717,N_1711);
or U1799 (N_1799,N_1732,N_1695);
nor U1800 (N_1800,N_1784,N_1749);
or U1801 (N_1801,N_1768,N_1789);
xor U1802 (N_1802,N_1793,N_1758);
nand U1803 (N_1803,N_1770,N_1743);
nand U1804 (N_1804,N_1771,N_1776);
or U1805 (N_1805,N_1753,N_1746);
nor U1806 (N_1806,N_1742,N_1775);
nand U1807 (N_1807,N_1765,N_1796);
nor U1808 (N_1808,N_1782,N_1760);
nand U1809 (N_1809,N_1763,N_1747);
nand U1810 (N_1810,N_1798,N_1754);
nand U1811 (N_1811,N_1788,N_1767);
and U1812 (N_1812,N_1792,N_1779);
nor U1813 (N_1813,N_1756,N_1751);
and U1814 (N_1814,N_1791,N_1787);
nand U1815 (N_1815,N_1794,N_1786);
or U1816 (N_1816,N_1781,N_1799);
nand U1817 (N_1817,N_1795,N_1741);
or U1818 (N_1818,N_1750,N_1774);
nand U1819 (N_1819,N_1762,N_1757);
and U1820 (N_1820,N_1772,N_1778);
nor U1821 (N_1821,N_1766,N_1761);
or U1822 (N_1822,N_1790,N_1769);
and U1823 (N_1823,N_1780,N_1752);
nand U1824 (N_1824,N_1759,N_1748);
nand U1825 (N_1825,N_1777,N_1773);
and U1826 (N_1826,N_1740,N_1764);
or U1827 (N_1827,N_1744,N_1785);
and U1828 (N_1828,N_1783,N_1745);
and U1829 (N_1829,N_1755,N_1797);
nand U1830 (N_1830,N_1763,N_1796);
nor U1831 (N_1831,N_1768,N_1754);
or U1832 (N_1832,N_1794,N_1789);
nor U1833 (N_1833,N_1787,N_1755);
or U1834 (N_1834,N_1750,N_1753);
xor U1835 (N_1835,N_1769,N_1744);
and U1836 (N_1836,N_1763,N_1769);
nor U1837 (N_1837,N_1750,N_1772);
nand U1838 (N_1838,N_1776,N_1766);
nor U1839 (N_1839,N_1757,N_1775);
xnor U1840 (N_1840,N_1784,N_1794);
or U1841 (N_1841,N_1788,N_1779);
and U1842 (N_1842,N_1799,N_1786);
or U1843 (N_1843,N_1760,N_1761);
or U1844 (N_1844,N_1741,N_1772);
nand U1845 (N_1845,N_1786,N_1755);
and U1846 (N_1846,N_1778,N_1756);
and U1847 (N_1847,N_1796,N_1742);
xnor U1848 (N_1848,N_1782,N_1748);
or U1849 (N_1849,N_1781,N_1790);
nand U1850 (N_1850,N_1740,N_1772);
and U1851 (N_1851,N_1769,N_1760);
xnor U1852 (N_1852,N_1774,N_1759);
nor U1853 (N_1853,N_1791,N_1743);
or U1854 (N_1854,N_1786,N_1782);
xor U1855 (N_1855,N_1764,N_1797);
xor U1856 (N_1856,N_1775,N_1747);
or U1857 (N_1857,N_1790,N_1740);
and U1858 (N_1858,N_1763,N_1799);
and U1859 (N_1859,N_1792,N_1751);
or U1860 (N_1860,N_1832,N_1836);
nor U1861 (N_1861,N_1853,N_1841);
xnor U1862 (N_1862,N_1835,N_1844);
and U1863 (N_1863,N_1845,N_1803);
or U1864 (N_1864,N_1848,N_1817);
nor U1865 (N_1865,N_1805,N_1849);
nor U1866 (N_1866,N_1851,N_1802);
nand U1867 (N_1867,N_1843,N_1822);
or U1868 (N_1868,N_1810,N_1837);
and U1869 (N_1869,N_1816,N_1856);
nand U1870 (N_1870,N_1808,N_1852);
and U1871 (N_1871,N_1809,N_1850);
and U1872 (N_1872,N_1814,N_1827);
nor U1873 (N_1873,N_1857,N_1819);
or U1874 (N_1874,N_1823,N_1820);
and U1875 (N_1875,N_1824,N_1854);
nand U1876 (N_1876,N_1858,N_1811);
nand U1877 (N_1877,N_1840,N_1855);
nand U1878 (N_1878,N_1812,N_1806);
nand U1879 (N_1879,N_1834,N_1821);
or U1880 (N_1880,N_1818,N_1800);
or U1881 (N_1881,N_1815,N_1833);
nand U1882 (N_1882,N_1826,N_1801);
or U1883 (N_1883,N_1825,N_1828);
nor U1884 (N_1884,N_1831,N_1859);
xnor U1885 (N_1885,N_1838,N_1813);
xor U1886 (N_1886,N_1846,N_1830);
and U1887 (N_1887,N_1804,N_1839);
and U1888 (N_1888,N_1807,N_1847);
nor U1889 (N_1889,N_1842,N_1829);
or U1890 (N_1890,N_1833,N_1839);
or U1891 (N_1891,N_1836,N_1813);
nor U1892 (N_1892,N_1831,N_1837);
and U1893 (N_1893,N_1826,N_1802);
or U1894 (N_1894,N_1844,N_1823);
nand U1895 (N_1895,N_1810,N_1825);
nand U1896 (N_1896,N_1841,N_1848);
or U1897 (N_1897,N_1853,N_1821);
or U1898 (N_1898,N_1807,N_1819);
nor U1899 (N_1899,N_1843,N_1810);
nand U1900 (N_1900,N_1825,N_1822);
nor U1901 (N_1901,N_1805,N_1828);
or U1902 (N_1902,N_1840,N_1831);
nand U1903 (N_1903,N_1832,N_1822);
and U1904 (N_1904,N_1843,N_1815);
xor U1905 (N_1905,N_1823,N_1850);
nand U1906 (N_1906,N_1803,N_1833);
nand U1907 (N_1907,N_1841,N_1832);
xor U1908 (N_1908,N_1839,N_1850);
and U1909 (N_1909,N_1830,N_1825);
xor U1910 (N_1910,N_1802,N_1857);
nand U1911 (N_1911,N_1857,N_1811);
or U1912 (N_1912,N_1825,N_1853);
nand U1913 (N_1913,N_1827,N_1821);
nor U1914 (N_1914,N_1838,N_1839);
nand U1915 (N_1915,N_1814,N_1812);
nor U1916 (N_1916,N_1807,N_1800);
nand U1917 (N_1917,N_1809,N_1857);
or U1918 (N_1918,N_1814,N_1831);
nand U1919 (N_1919,N_1826,N_1840);
and U1920 (N_1920,N_1886,N_1881);
and U1921 (N_1921,N_1883,N_1901);
and U1922 (N_1922,N_1910,N_1868);
and U1923 (N_1923,N_1861,N_1860);
or U1924 (N_1924,N_1911,N_1891);
nand U1925 (N_1925,N_1913,N_1876);
nor U1926 (N_1926,N_1870,N_1897);
or U1927 (N_1927,N_1878,N_1882);
nor U1928 (N_1928,N_1916,N_1917);
nor U1929 (N_1929,N_1915,N_1907);
or U1930 (N_1930,N_1888,N_1874);
and U1931 (N_1931,N_1905,N_1893);
nor U1932 (N_1932,N_1890,N_1877);
and U1933 (N_1933,N_1866,N_1908);
xor U1934 (N_1934,N_1895,N_1912);
and U1935 (N_1935,N_1894,N_1867);
or U1936 (N_1936,N_1871,N_1880);
nand U1937 (N_1937,N_1872,N_1884);
and U1938 (N_1938,N_1869,N_1892);
nor U1939 (N_1939,N_1904,N_1909);
xnor U1940 (N_1940,N_1918,N_1900);
or U1941 (N_1941,N_1887,N_1889);
or U1942 (N_1942,N_1906,N_1862);
nor U1943 (N_1943,N_1914,N_1919);
xor U1944 (N_1944,N_1864,N_1902);
nand U1945 (N_1945,N_1863,N_1899);
nand U1946 (N_1946,N_1873,N_1896);
nand U1947 (N_1947,N_1898,N_1903);
nor U1948 (N_1948,N_1879,N_1875);
or U1949 (N_1949,N_1865,N_1885);
or U1950 (N_1950,N_1863,N_1864);
xnor U1951 (N_1951,N_1913,N_1873);
and U1952 (N_1952,N_1905,N_1901);
nand U1953 (N_1953,N_1860,N_1896);
nand U1954 (N_1954,N_1882,N_1910);
nor U1955 (N_1955,N_1912,N_1863);
and U1956 (N_1956,N_1917,N_1876);
nand U1957 (N_1957,N_1893,N_1886);
or U1958 (N_1958,N_1874,N_1898);
or U1959 (N_1959,N_1866,N_1876);
or U1960 (N_1960,N_1871,N_1888);
and U1961 (N_1961,N_1870,N_1882);
and U1962 (N_1962,N_1903,N_1869);
or U1963 (N_1963,N_1869,N_1906);
or U1964 (N_1964,N_1864,N_1895);
or U1965 (N_1965,N_1885,N_1864);
nand U1966 (N_1966,N_1914,N_1898);
and U1967 (N_1967,N_1916,N_1871);
and U1968 (N_1968,N_1862,N_1919);
or U1969 (N_1969,N_1904,N_1893);
nor U1970 (N_1970,N_1864,N_1913);
nand U1971 (N_1971,N_1885,N_1863);
nand U1972 (N_1972,N_1914,N_1867);
nand U1973 (N_1973,N_1904,N_1911);
xor U1974 (N_1974,N_1914,N_1888);
or U1975 (N_1975,N_1864,N_1875);
nor U1976 (N_1976,N_1876,N_1870);
and U1977 (N_1977,N_1918,N_1916);
nor U1978 (N_1978,N_1871,N_1894);
nand U1979 (N_1979,N_1901,N_1906);
nand U1980 (N_1980,N_1925,N_1941);
and U1981 (N_1981,N_1938,N_1945);
and U1982 (N_1982,N_1940,N_1922);
nor U1983 (N_1983,N_1949,N_1955);
or U1984 (N_1984,N_1964,N_1978);
nor U1985 (N_1985,N_1953,N_1954);
nor U1986 (N_1986,N_1947,N_1957);
nor U1987 (N_1987,N_1951,N_1966);
nand U1988 (N_1988,N_1928,N_1946);
xor U1989 (N_1989,N_1958,N_1932);
and U1990 (N_1990,N_1967,N_1924);
and U1991 (N_1991,N_1969,N_1979);
nor U1992 (N_1992,N_1963,N_1952);
nor U1993 (N_1993,N_1935,N_1972);
nand U1994 (N_1994,N_1936,N_1943);
nand U1995 (N_1995,N_1931,N_1974);
xor U1996 (N_1996,N_1926,N_1973);
or U1997 (N_1997,N_1968,N_1937);
xnor U1998 (N_1998,N_1971,N_1959);
and U1999 (N_1999,N_1956,N_1921);
nand U2000 (N_2000,N_1942,N_1927);
nand U2001 (N_2001,N_1920,N_1948);
and U2002 (N_2002,N_1975,N_1970);
nand U2003 (N_2003,N_1965,N_1976);
xor U2004 (N_2004,N_1930,N_1929);
xnor U2005 (N_2005,N_1944,N_1961);
and U2006 (N_2006,N_1960,N_1950);
and U2007 (N_2007,N_1934,N_1962);
or U2008 (N_2008,N_1939,N_1923);
nand U2009 (N_2009,N_1977,N_1933);
nor U2010 (N_2010,N_1947,N_1948);
xor U2011 (N_2011,N_1931,N_1956);
and U2012 (N_2012,N_1948,N_1938);
nand U2013 (N_2013,N_1951,N_1973);
and U2014 (N_2014,N_1944,N_1921);
nor U2015 (N_2015,N_1931,N_1967);
and U2016 (N_2016,N_1945,N_1929);
nor U2017 (N_2017,N_1962,N_1944);
nand U2018 (N_2018,N_1961,N_1966);
and U2019 (N_2019,N_1971,N_1949);
nand U2020 (N_2020,N_1947,N_1943);
nor U2021 (N_2021,N_1979,N_1978);
nand U2022 (N_2022,N_1976,N_1953);
and U2023 (N_2023,N_1921,N_1979);
nor U2024 (N_2024,N_1940,N_1937);
and U2025 (N_2025,N_1948,N_1940);
nand U2026 (N_2026,N_1970,N_1926);
and U2027 (N_2027,N_1935,N_1957);
nand U2028 (N_2028,N_1941,N_1928);
and U2029 (N_2029,N_1966,N_1944);
nor U2030 (N_2030,N_1926,N_1937);
or U2031 (N_2031,N_1938,N_1921);
nand U2032 (N_2032,N_1959,N_1963);
nor U2033 (N_2033,N_1931,N_1930);
nor U2034 (N_2034,N_1967,N_1944);
nand U2035 (N_2035,N_1941,N_1921);
or U2036 (N_2036,N_1958,N_1962);
nor U2037 (N_2037,N_1921,N_1942);
nand U2038 (N_2038,N_1949,N_1975);
nand U2039 (N_2039,N_1940,N_1975);
nor U2040 (N_2040,N_2002,N_1995);
nor U2041 (N_2041,N_2000,N_2011);
nor U2042 (N_2042,N_2038,N_1984);
and U2043 (N_2043,N_1998,N_1981);
or U2044 (N_2044,N_2016,N_2008);
nor U2045 (N_2045,N_2020,N_2023);
nor U2046 (N_2046,N_2015,N_2012);
or U2047 (N_2047,N_2006,N_2019);
or U2048 (N_2048,N_1993,N_2026);
or U2049 (N_2049,N_2024,N_1988);
or U2050 (N_2050,N_2021,N_2017);
nor U2051 (N_2051,N_2027,N_2030);
and U2052 (N_2052,N_2037,N_1996);
nand U2053 (N_2053,N_2029,N_1982);
and U2054 (N_2054,N_1991,N_1999);
nor U2055 (N_2055,N_1990,N_1985);
nor U2056 (N_2056,N_2004,N_2035);
and U2057 (N_2057,N_2032,N_2003);
nor U2058 (N_2058,N_1997,N_1987);
or U2059 (N_2059,N_2033,N_2007);
and U2060 (N_2060,N_1994,N_2031);
or U2061 (N_2061,N_2018,N_1983);
and U2062 (N_2062,N_2039,N_2022);
or U2063 (N_2063,N_1980,N_2001);
nor U2064 (N_2064,N_1989,N_1992);
xnor U2065 (N_2065,N_2028,N_2036);
nand U2066 (N_2066,N_2005,N_2010);
or U2067 (N_2067,N_2013,N_1986);
nand U2068 (N_2068,N_2014,N_2025);
nor U2069 (N_2069,N_2034,N_2009);
nand U2070 (N_2070,N_2020,N_2029);
and U2071 (N_2071,N_2012,N_1988);
or U2072 (N_2072,N_2007,N_1988);
xor U2073 (N_2073,N_1997,N_1992);
nor U2074 (N_2074,N_1999,N_2028);
xor U2075 (N_2075,N_2003,N_2029);
or U2076 (N_2076,N_1995,N_2014);
or U2077 (N_2077,N_2034,N_2028);
nand U2078 (N_2078,N_2008,N_1995);
and U2079 (N_2079,N_1999,N_1996);
or U2080 (N_2080,N_2038,N_2018);
xor U2081 (N_2081,N_2024,N_2009);
nand U2082 (N_2082,N_2015,N_2033);
xor U2083 (N_2083,N_2022,N_1991);
or U2084 (N_2084,N_2038,N_1999);
xor U2085 (N_2085,N_2028,N_2009);
or U2086 (N_2086,N_2000,N_2028);
nor U2087 (N_2087,N_1987,N_2021);
or U2088 (N_2088,N_1998,N_2019);
nor U2089 (N_2089,N_2013,N_1997);
nand U2090 (N_2090,N_2036,N_2004);
xnor U2091 (N_2091,N_2000,N_2037);
and U2092 (N_2092,N_2033,N_2022);
nor U2093 (N_2093,N_2032,N_2030);
and U2094 (N_2094,N_2017,N_1980);
and U2095 (N_2095,N_2010,N_2009);
or U2096 (N_2096,N_2037,N_2024);
nand U2097 (N_2097,N_1983,N_2020);
nor U2098 (N_2098,N_2039,N_2023);
or U2099 (N_2099,N_2021,N_2030);
xor U2100 (N_2100,N_2090,N_2057);
nand U2101 (N_2101,N_2091,N_2075);
nor U2102 (N_2102,N_2064,N_2060);
nand U2103 (N_2103,N_2063,N_2050);
or U2104 (N_2104,N_2086,N_2099);
and U2105 (N_2105,N_2084,N_2072);
or U2106 (N_2106,N_2073,N_2062);
or U2107 (N_2107,N_2040,N_2041);
or U2108 (N_2108,N_2046,N_2081);
or U2109 (N_2109,N_2045,N_2067);
nand U2110 (N_2110,N_2066,N_2093);
nand U2111 (N_2111,N_2077,N_2055);
or U2112 (N_2112,N_2098,N_2069);
xor U2113 (N_2113,N_2052,N_2083);
or U2114 (N_2114,N_2088,N_2078);
xor U2115 (N_2115,N_2095,N_2048);
and U2116 (N_2116,N_2087,N_2080);
xnor U2117 (N_2117,N_2074,N_2082);
nor U2118 (N_2118,N_2047,N_2070);
nand U2119 (N_2119,N_2092,N_2054);
or U2120 (N_2120,N_2097,N_2065);
or U2121 (N_2121,N_2068,N_2071);
or U2122 (N_2122,N_2043,N_2076);
or U2123 (N_2123,N_2096,N_2085);
nor U2124 (N_2124,N_2044,N_2079);
nand U2125 (N_2125,N_2056,N_2042);
nor U2126 (N_2126,N_2053,N_2094);
nand U2127 (N_2127,N_2061,N_2059);
or U2128 (N_2128,N_2051,N_2089);
or U2129 (N_2129,N_2058,N_2049);
xnor U2130 (N_2130,N_2088,N_2053);
and U2131 (N_2131,N_2074,N_2078);
nand U2132 (N_2132,N_2097,N_2073);
or U2133 (N_2133,N_2066,N_2091);
nand U2134 (N_2134,N_2071,N_2082);
nor U2135 (N_2135,N_2043,N_2082);
or U2136 (N_2136,N_2062,N_2052);
or U2137 (N_2137,N_2061,N_2077);
and U2138 (N_2138,N_2048,N_2071);
or U2139 (N_2139,N_2058,N_2089);
nor U2140 (N_2140,N_2061,N_2071);
and U2141 (N_2141,N_2085,N_2040);
and U2142 (N_2142,N_2092,N_2062);
or U2143 (N_2143,N_2087,N_2049);
and U2144 (N_2144,N_2064,N_2063);
nor U2145 (N_2145,N_2045,N_2071);
and U2146 (N_2146,N_2042,N_2076);
and U2147 (N_2147,N_2096,N_2049);
nor U2148 (N_2148,N_2066,N_2083);
nor U2149 (N_2149,N_2095,N_2094);
and U2150 (N_2150,N_2050,N_2060);
and U2151 (N_2151,N_2051,N_2076);
xnor U2152 (N_2152,N_2050,N_2056);
or U2153 (N_2153,N_2097,N_2082);
nand U2154 (N_2154,N_2075,N_2086);
xnor U2155 (N_2155,N_2098,N_2070);
nor U2156 (N_2156,N_2050,N_2092);
nand U2157 (N_2157,N_2078,N_2063);
and U2158 (N_2158,N_2056,N_2076);
nor U2159 (N_2159,N_2075,N_2061);
nand U2160 (N_2160,N_2100,N_2154);
nand U2161 (N_2161,N_2129,N_2107);
nand U2162 (N_2162,N_2112,N_2102);
nand U2163 (N_2163,N_2106,N_2104);
and U2164 (N_2164,N_2147,N_2155);
or U2165 (N_2165,N_2113,N_2115);
or U2166 (N_2166,N_2145,N_2151);
or U2167 (N_2167,N_2119,N_2121);
nor U2168 (N_2168,N_2123,N_2117);
or U2169 (N_2169,N_2101,N_2120);
and U2170 (N_2170,N_2144,N_2136);
nand U2171 (N_2171,N_2108,N_2139);
or U2172 (N_2172,N_2131,N_2128);
and U2173 (N_2173,N_2124,N_2157);
xnor U2174 (N_2174,N_2148,N_2149);
nor U2175 (N_2175,N_2159,N_2142);
nand U2176 (N_2176,N_2152,N_2118);
nand U2177 (N_2177,N_2122,N_2125);
and U2178 (N_2178,N_2103,N_2110);
nand U2179 (N_2179,N_2146,N_2130);
or U2180 (N_2180,N_2156,N_2109);
nand U2181 (N_2181,N_2134,N_2143);
or U2182 (N_2182,N_2150,N_2111);
nand U2183 (N_2183,N_2137,N_2126);
and U2184 (N_2184,N_2158,N_2138);
and U2185 (N_2185,N_2114,N_2132);
nor U2186 (N_2186,N_2153,N_2105);
nand U2187 (N_2187,N_2140,N_2135);
nor U2188 (N_2188,N_2116,N_2133);
nor U2189 (N_2189,N_2127,N_2141);
and U2190 (N_2190,N_2117,N_2157);
nand U2191 (N_2191,N_2119,N_2102);
nor U2192 (N_2192,N_2125,N_2116);
and U2193 (N_2193,N_2128,N_2118);
nor U2194 (N_2194,N_2119,N_2142);
or U2195 (N_2195,N_2129,N_2153);
nor U2196 (N_2196,N_2156,N_2119);
or U2197 (N_2197,N_2148,N_2100);
nand U2198 (N_2198,N_2115,N_2117);
and U2199 (N_2199,N_2153,N_2143);
or U2200 (N_2200,N_2116,N_2137);
nor U2201 (N_2201,N_2144,N_2108);
nor U2202 (N_2202,N_2132,N_2153);
nand U2203 (N_2203,N_2103,N_2155);
nand U2204 (N_2204,N_2106,N_2122);
xor U2205 (N_2205,N_2144,N_2130);
and U2206 (N_2206,N_2127,N_2101);
nor U2207 (N_2207,N_2149,N_2104);
nor U2208 (N_2208,N_2133,N_2103);
and U2209 (N_2209,N_2140,N_2111);
nand U2210 (N_2210,N_2133,N_2159);
and U2211 (N_2211,N_2105,N_2136);
and U2212 (N_2212,N_2155,N_2150);
xnor U2213 (N_2213,N_2134,N_2147);
nand U2214 (N_2214,N_2113,N_2120);
nor U2215 (N_2215,N_2135,N_2129);
nand U2216 (N_2216,N_2135,N_2148);
and U2217 (N_2217,N_2144,N_2131);
nor U2218 (N_2218,N_2101,N_2111);
nand U2219 (N_2219,N_2111,N_2133);
nand U2220 (N_2220,N_2179,N_2167);
nand U2221 (N_2221,N_2181,N_2205);
or U2222 (N_2222,N_2162,N_2204);
or U2223 (N_2223,N_2194,N_2213);
or U2224 (N_2224,N_2166,N_2180);
nand U2225 (N_2225,N_2212,N_2164);
and U2226 (N_2226,N_2186,N_2219);
or U2227 (N_2227,N_2206,N_2195);
and U2228 (N_2228,N_2176,N_2197);
and U2229 (N_2229,N_2160,N_2173);
nor U2230 (N_2230,N_2211,N_2218);
xor U2231 (N_2231,N_2191,N_2198);
and U2232 (N_2232,N_2193,N_2203);
or U2233 (N_2233,N_2208,N_2183);
and U2234 (N_2234,N_2182,N_2196);
and U2235 (N_2235,N_2214,N_2175);
or U2236 (N_2236,N_2192,N_2190);
nand U2237 (N_2237,N_2168,N_2161);
and U2238 (N_2238,N_2200,N_2163);
or U2239 (N_2239,N_2202,N_2207);
nand U2240 (N_2240,N_2185,N_2184);
and U2241 (N_2241,N_2215,N_2201);
and U2242 (N_2242,N_2174,N_2165);
and U2243 (N_2243,N_2189,N_2172);
nor U2244 (N_2244,N_2209,N_2178);
or U2245 (N_2245,N_2216,N_2188);
and U2246 (N_2246,N_2170,N_2177);
nor U2247 (N_2247,N_2169,N_2187);
nand U2248 (N_2248,N_2171,N_2199);
or U2249 (N_2249,N_2210,N_2217);
nor U2250 (N_2250,N_2197,N_2217);
nor U2251 (N_2251,N_2170,N_2215);
and U2252 (N_2252,N_2213,N_2205);
nor U2253 (N_2253,N_2210,N_2181);
nand U2254 (N_2254,N_2210,N_2203);
or U2255 (N_2255,N_2174,N_2191);
nor U2256 (N_2256,N_2192,N_2208);
nor U2257 (N_2257,N_2196,N_2200);
nand U2258 (N_2258,N_2202,N_2164);
nor U2259 (N_2259,N_2177,N_2200);
nand U2260 (N_2260,N_2166,N_2184);
nor U2261 (N_2261,N_2197,N_2174);
or U2262 (N_2262,N_2180,N_2163);
nor U2263 (N_2263,N_2171,N_2202);
or U2264 (N_2264,N_2170,N_2187);
or U2265 (N_2265,N_2216,N_2170);
and U2266 (N_2266,N_2218,N_2212);
nand U2267 (N_2267,N_2166,N_2203);
nand U2268 (N_2268,N_2183,N_2207);
nand U2269 (N_2269,N_2173,N_2179);
nor U2270 (N_2270,N_2212,N_2179);
nand U2271 (N_2271,N_2217,N_2179);
nor U2272 (N_2272,N_2214,N_2205);
nand U2273 (N_2273,N_2167,N_2212);
and U2274 (N_2274,N_2207,N_2195);
and U2275 (N_2275,N_2189,N_2162);
xnor U2276 (N_2276,N_2162,N_2188);
nor U2277 (N_2277,N_2219,N_2192);
nor U2278 (N_2278,N_2183,N_2195);
nand U2279 (N_2279,N_2218,N_2175);
nand U2280 (N_2280,N_2276,N_2224);
xor U2281 (N_2281,N_2230,N_2257);
and U2282 (N_2282,N_2241,N_2277);
nor U2283 (N_2283,N_2254,N_2266);
nor U2284 (N_2284,N_2221,N_2248);
xor U2285 (N_2285,N_2268,N_2244);
nor U2286 (N_2286,N_2269,N_2223);
or U2287 (N_2287,N_2274,N_2278);
xnor U2288 (N_2288,N_2240,N_2265);
or U2289 (N_2289,N_2238,N_2225);
nand U2290 (N_2290,N_2245,N_2235);
nor U2291 (N_2291,N_2227,N_2271);
nor U2292 (N_2292,N_2263,N_2231);
nand U2293 (N_2293,N_2255,N_2267);
xor U2294 (N_2294,N_2279,N_2220);
or U2295 (N_2295,N_2252,N_2222);
and U2296 (N_2296,N_2234,N_2258);
and U2297 (N_2297,N_2270,N_2273);
nand U2298 (N_2298,N_2260,N_2262);
or U2299 (N_2299,N_2259,N_2247);
nor U2300 (N_2300,N_2242,N_2272);
nor U2301 (N_2301,N_2226,N_2239);
nand U2302 (N_2302,N_2264,N_2251);
nor U2303 (N_2303,N_2236,N_2243);
nor U2304 (N_2304,N_2228,N_2229);
and U2305 (N_2305,N_2237,N_2253);
nor U2306 (N_2306,N_2275,N_2249);
xor U2307 (N_2307,N_2246,N_2233);
or U2308 (N_2308,N_2232,N_2256);
and U2309 (N_2309,N_2250,N_2261);
xnor U2310 (N_2310,N_2237,N_2233);
nand U2311 (N_2311,N_2231,N_2236);
nand U2312 (N_2312,N_2261,N_2254);
or U2313 (N_2313,N_2250,N_2226);
and U2314 (N_2314,N_2221,N_2246);
xnor U2315 (N_2315,N_2247,N_2239);
or U2316 (N_2316,N_2277,N_2221);
and U2317 (N_2317,N_2234,N_2248);
nor U2318 (N_2318,N_2244,N_2228);
and U2319 (N_2319,N_2222,N_2232);
and U2320 (N_2320,N_2263,N_2227);
or U2321 (N_2321,N_2222,N_2261);
and U2322 (N_2322,N_2227,N_2241);
or U2323 (N_2323,N_2226,N_2224);
nor U2324 (N_2324,N_2228,N_2232);
nand U2325 (N_2325,N_2276,N_2275);
nor U2326 (N_2326,N_2244,N_2264);
or U2327 (N_2327,N_2236,N_2227);
or U2328 (N_2328,N_2227,N_2279);
nor U2329 (N_2329,N_2269,N_2236);
and U2330 (N_2330,N_2229,N_2273);
and U2331 (N_2331,N_2264,N_2231);
and U2332 (N_2332,N_2222,N_2244);
and U2333 (N_2333,N_2247,N_2224);
nand U2334 (N_2334,N_2256,N_2279);
nand U2335 (N_2335,N_2252,N_2223);
or U2336 (N_2336,N_2228,N_2243);
or U2337 (N_2337,N_2239,N_2238);
and U2338 (N_2338,N_2230,N_2232);
and U2339 (N_2339,N_2279,N_2223);
or U2340 (N_2340,N_2317,N_2291);
or U2341 (N_2341,N_2337,N_2309);
xnor U2342 (N_2342,N_2332,N_2311);
nand U2343 (N_2343,N_2301,N_2304);
nand U2344 (N_2344,N_2331,N_2329);
and U2345 (N_2345,N_2307,N_2299);
nor U2346 (N_2346,N_2336,N_2308);
xnor U2347 (N_2347,N_2322,N_2316);
nand U2348 (N_2348,N_2286,N_2330);
nor U2349 (N_2349,N_2335,N_2302);
nor U2350 (N_2350,N_2321,N_2282);
or U2351 (N_2351,N_2333,N_2310);
nor U2352 (N_2352,N_2292,N_2328);
nand U2353 (N_2353,N_2320,N_2283);
or U2354 (N_2354,N_2303,N_2289);
and U2355 (N_2355,N_2280,N_2296);
nand U2356 (N_2356,N_2325,N_2295);
and U2357 (N_2357,N_2313,N_2314);
nand U2358 (N_2358,N_2306,N_2281);
or U2359 (N_2359,N_2293,N_2305);
or U2360 (N_2360,N_2319,N_2315);
xor U2361 (N_2361,N_2287,N_2285);
nand U2362 (N_2362,N_2338,N_2298);
nor U2363 (N_2363,N_2318,N_2327);
or U2364 (N_2364,N_2284,N_2326);
or U2365 (N_2365,N_2324,N_2300);
or U2366 (N_2366,N_2312,N_2297);
nor U2367 (N_2367,N_2288,N_2334);
nor U2368 (N_2368,N_2323,N_2339);
and U2369 (N_2369,N_2290,N_2294);
nor U2370 (N_2370,N_2325,N_2288);
and U2371 (N_2371,N_2335,N_2331);
and U2372 (N_2372,N_2336,N_2286);
nand U2373 (N_2373,N_2319,N_2320);
and U2374 (N_2374,N_2297,N_2287);
or U2375 (N_2375,N_2289,N_2284);
or U2376 (N_2376,N_2327,N_2320);
or U2377 (N_2377,N_2292,N_2312);
nand U2378 (N_2378,N_2305,N_2338);
nand U2379 (N_2379,N_2334,N_2329);
nand U2380 (N_2380,N_2338,N_2294);
and U2381 (N_2381,N_2310,N_2299);
or U2382 (N_2382,N_2297,N_2329);
xnor U2383 (N_2383,N_2316,N_2286);
and U2384 (N_2384,N_2306,N_2301);
nand U2385 (N_2385,N_2303,N_2281);
xor U2386 (N_2386,N_2320,N_2321);
and U2387 (N_2387,N_2291,N_2331);
xor U2388 (N_2388,N_2337,N_2328);
nor U2389 (N_2389,N_2290,N_2335);
and U2390 (N_2390,N_2302,N_2336);
and U2391 (N_2391,N_2325,N_2338);
or U2392 (N_2392,N_2316,N_2325);
nand U2393 (N_2393,N_2299,N_2309);
or U2394 (N_2394,N_2295,N_2294);
xor U2395 (N_2395,N_2326,N_2327);
or U2396 (N_2396,N_2321,N_2289);
and U2397 (N_2397,N_2288,N_2331);
xor U2398 (N_2398,N_2291,N_2296);
nor U2399 (N_2399,N_2327,N_2321);
xnor U2400 (N_2400,N_2385,N_2397);
or U2401 (N_2401,N_2393,N_2373);
nand U2402 (N_2402,N_2377,N_2352);
or U2403 (N_2403,N_2361,N_2384);
and U2404 (N_2404,N_2386,N_2376);
nand U2405 (N_2405,N_2398,N_2370);
nor U2406 (N_2406,N_2387,N_2355);
nor U2407 (N_2407,N_2348,N_2342);
and U2408 (N_2408,N_2383,N_2364);
nor U2409 (N_2409,N_2380,N_2375);
or U2410 (N_2410,N_2396,N_2381);
xnor U2411 (N_2411,N_2382,N_2351);
nor U2412 (N_2412,N_2372,N_2378);
or U2413 (N_2413,N_2344,N_2343);
nor U2414 (N_2414,N_2391,N_2340);
nand U2415 (N_2415,N_2354,N_2357);
nor U2416 (N_2416,N_2395,N_2367);
and U2417 (N_2417,N_2341,N_2371);
nand U2418 (N_2418,N_2358,N_2350);
and U2419 (N_2419,N_2345,N_2389);
xnor U2420 (N_2420,N_2360,N_2362);
and U2421 (N_2421,N_2359,N_2392);
nor U2422 (N_2422,N_2390,N_2347);
and U2423 (N_2423,N_2363,N_2368);
or U2424 (N_2424,N_2356,N_2388);
nand U2425 (N_2425,N_2346,N_2366);
nor U2426 (N_2426,N_2399,N_2369);
and U2427 (N_2427,N_2365,N_2353);
nor U2428 (N_2428,N_2379,N_2349);
and U2429 (N_2429,N_2394,N_2374);
or U2430 (N_2430,N_2381,N_2393);
or U2431 (N_2431,N_2342,N_2395);
xnor U2432 (N_2432,N_2380,N_2364);
and U2433 (N_2433,N_2367,N_2366);
or U2434 (N_2434,N_2362,N_2390);
and U2435 (N_2435,N_2343,N_2395);
or U2436 (N_2436,N_2398,N_2392);
or U2437 (N_2437,N_2352,N_2363);
nand U2438 (N_2438,N_2361,N_2386);
xor U2439 (N_2439,N_2375,N_2389);
and U2440 (N_2440,N_2375,N_2344);
nand U2441 (N_2441,N_2344,N_2349);
or U2442 (N_2442,N_2386,N_2371);
nor U2443 (N_2443,N_2384,N_2381);
nor U2444 (N_2444,N_2381,N_2392);
or U2445 (N_2445,N_2392,N_2364);
and U2446 (N_2446,N_2368,N_2348);
and U2447 (N_2447,N_2359,N_2367);
nor U2448 (N_2448,N_2357,N_2348);
nand U2449 (N_2449,N_2355,N_2390);
or U2450 (N_2450,N_2351,N_2347);
nand U2451 (N_2451,N_2356,N_2349);
and U2452 (N_2452,N_2361,N_2364);
or U2453 (N_2453,N_2387,N_2341);
nor U2454 (N_2454,N_2358,N_2362);
xnor U2455 (N_2455,N_2369,N_2386);
nor U2456 (N_2456,N_2394,N_2349);
or U2457 (N_2457,N_2370,N_2359);
or U2458 (N_2458,N_2340,N_2351);
nor U2459 (N_2459,N_2397,N_2372);
nand U2460 (N_2460,N_2413,N_2435);
nand U2461 (N_2461,N_2438,N_2400);
nand U2462 (N_2462,N_2419,N_2424);
and U2463 (N_2463,N_2450,N_2452);
and U2464 (N_2464,N_2421,N_2451);
xor U2465 (N_2465,N_2448,N_2412);
and U2466 (N_2466,N_2404,N_2427);
nand U2467 (N_2467,N_2447,N_2439);
or U2468 (N_2468,N_2416,N_2426);
nor U2469 (N_2469,N_2443,N_2414);
xor U2470 (N_2470,N_2455,N_2402);
nand U2471 (N_2471,N_2429,N_2406);
nand U2472 (N_2472,N_2434,N_2446);
xnor U2473 (N_2473,N_2449,N_2411);
and U2474 (N_2474,N_2433,N_2401);
nand U2475 (N_2475,N_2437,N_2407);
nand U2476 (N_2476,N_2417,N_2408);
and U2477 (N_2477,N_2405,N_2425);
nor U2478 (N_2478,N_2432,N_2440);
nand U2479 (N_2479,N_2454,N_2436);
nor U2480 (N_2480,N_2420,N_2458);
or U2481 (N_2481,N_2453,N_2409);
or U2482 (N_2482,N_2415,N_2431);
and U2483 (N_2483,N_2456,N_2428);
and U2484 (N_2484,N_2403,N_2423);
or U2485 (N_2485,N_2422,N_2444);
xor U2486 (N_2486,N_2457,N_2459);
or U2487 (N_2487,N_2430,N_2442);
nor U2488 (N_2488,N_2445,N_2441);
or U2489 (N_2489,N_2410,N_2418);
nor U2490 (N_2490,N_2404,N_2456);
or U2491 (N_2491,N_2444,N_2458);
nor U2492 (N_2492,N_2423,N_2445);
nand U2493 (N_2493,N_2418,N_2446);
or U2494 (N_2494,N_2415,N_2445);
and U2495 (N_2495,N_2417,N_2428);
nor U2496 (N_2496,N_2451,N_2401);
and U2497 (N_2497,N_2424,N_2430);
or U2498 (N_2498,N_2433,N_2400);
and U2499 (N_2499,N_2442,N_2435);
or U2500 (N_2500,N_2448,N_2447);
or U2501 (N_2501,N_2416,N_2423);
and U2502 (N_2502,N_2422,N_2440);
nand U2503 (N_2503,N_2456,N_2424);
and U2504 (N_2504,N_2402,N_2440);
or U2505 (N_2505,N_2443,N_2416);
or U2506 (N_2506,N_2446,N_2435);
nand U2507 (N_2507,N_2431,N_2418);
nor U2508 (N_2508,N_2432,N_2422);
nor U2509 (N_2509,N_2421,N_2416);
and U2510 (N_2510,N_2457,N_2400);
nor U2511 (N_2511,N_2405,N_2416);
and U2512 (N_2512,N_2420,N_2417);
or U2513 (N_2513,N_2446,N_2449);
and U2514 (N_2514,N_2453,N_2415);
or U2515 (N_2515,N_2412,N_2431);
and U2516 (N_2516,N_2435,N_2434);
nand U2517 (N_2517,N_2425,N_2449);
and U2518 (N_2518,N_2405,N_2451);
and U2519 (N_2519,N_2446,N_2454);
xor U2520 (N_2520,N_2506,N_2462);
and U2521 (N_2521,N_2516,N_2499);
and U2522 (N_2522,N_2480,N_2510);
and U2523 (N_2523,N_2467,N_2503);
or U2524 (N_2524,N_2519,N_2509);
and U2525 (N_2525,N_2495,N_2496);
xnor U2526 (N_2526,N_2490,N_2483);
nand U2527 (N_2527,N_2476,N_2484);
and U2528 (N_2528,N_2511,N_2488);
and U2529 (N_2529,N_2517,N_2507);
or U2530 (N_2530,N_2508,N_2486);
or U2531 (N_2531,N_2482,N_2471);
xor U2532 (N_2532,N_2470,N_2489);
or U2533 (N_2533,N_2463,N_2493);
nand U2534 (N_2534,N_2504,N_2513);
nor U2535 (N_2535,N_2485,N_2492);
nor U2536 (N_2536,N_2465,N_2475);
and U2537 (N_2537,N_2461,N_2501);
nand U2538 (N_2538,N_2518,N_2515);
or U2539 (N_2539,N_2474,N_2494);
nand U2540 (N_2540,N_2468,N_2472);
and U2541 (N_2541,N_2469,N_2464);
nor U2542 (N_2542,N_2466,N_2481);
nand U2543 (N_2543,N_2512,N_2479);
xnor U2544 (N_2544,N_2498,N_2497);
xnor U2545 (N_2545,N_2460,N_2478);
nand U2546 (N_2546,N_2514,N_2487);
or U2547 (N_2547,N_2473,N_2500);
and U2548 (N_2548,N_2505,N_2477);
nor U2549 (N_2549,N_2502,N_2491);
and U2550 (N_2550,N_2514,N_2517);
or U2551 (N_2551,N_2511,N_2484);
nand U2552 (N_2552,N_2513,N_2496);
nor U2553 (N_2553,N_2479,N_2464);
or U2554 (N_2554,N_2508,N_2488);
and U2555 (N_2555,N_2507,N_2486);
nand U2556 (N_2556,N_2477,N_2486);
xnor U2557 (N_2557,N_2485,N_2478);
nand U2558 (N_2558,N_2513,N_2478);
or U2559 (N_2559,N_2518,N_2477);
or U2560 (N_2560,N_2464,N_2501);
and U2561 (N_2561,N_2480,N_2498);
xnor U2562 (N_2562,N_2490,N_2482);
nand U2563 (N_2563,N_2513,N_2516);
nor U2564 (N_2564,N_2489,N_2495);
or U2565 (N_2565,N_2469,N_2499);
or U2566 (N_2566,N_2491,N_2511);
nor U2567 (N_2567,N_2487,N_2468);
nor U2568 (N_2568,N_2507,N_2510);
xnor U2569 (N_2569,N_2470,N_2498);
nor U2570 (N_2570,N_2489,N_2490);
or U2571 (N_2571,N_2463,N_2483);
nand U2572 (N_2572,N_2497,N_2475);
and U2573 (N_2573,N_2467,N_2485);
and U2574 (N_2574,N_2498,N_2516);
nor U2575 (N_2575,N_2491,N_2500);
and U2576 (N_2576,N_2500,N_2518);
nor U2577 (N_2577,N_2517,N_2497);
nor U2578 (N_2578,N_2461,N_2477);
nor U2579 (N_2579,N_2485,N_2498);
xor U2580 (N_2580,N_2559,N_2552);
nor U2581 (N_2581,N_2523,N_2532);
nand U2582 (N_2582,N_2525,N_2531);
and U2583 (N_2583,N_2535,N_2571);
or U2584 (N_2584,N_2529,N_2564);
and U2585 (N_2585,N_2544,N_2577);
nand U2586 (N_2586,N_2574,N_2536);
and U2587 (N_2587,N_2537,N_2573);
or U2588 (N_2588,N_2527,N_2576);
nor U2589 (N_2589,N_2548,N_2561);
nand U2590 (N_2590,N_2566,N_2547);
nor U2591 (N_2591,N_2538,N_2560);
xnor U2592 (N_2592,N_2558,N_2540);
nor U2593 (N_2593,N_2579,N_2550);
nor U2594 (N_2594,N_2554,N_2524);
nand U2595 (N_2595,N_2575,N_2562);
or U2596 (N_2596,N_2521,N_2534);
nand U2597 (N_2597,N_2549,N_2556);
nor U2598 (N_2598,N_2563,N_2545);
and U2599 (N_2599,N_2569,N_2551);
nand U2600 (N_2600,N_2565,N_2570);
nor U2601 (N_2601,N_2557,N_2528);
and U2602 (N_2602,N_2542,N_2522);
and U2603 (N_2603,N_2578,N_2568);
and U2604 (N_2604,N_2572,N_2567);
xor U2605 (N_2605,N_2533,N_2553);
or U2606 (N_2606,N_2539,N_2520);
and U2607 (N_2607,N_2541,N_2530);
xnor U2608 (N_2608,N_2555,N_2526);
nor U2609 (N_2609,N_2543,N_2546);
nor U2610 (N_2610,N_2544,N_2574);
nor U2611 (N_2611,N_2543,N_2540);
or U2612 (N_2612,N_2564,N_2570);
nor U2613 (N_2613,N_2521,N_2535);
or U2614 (N_2614,N_2563,N_2578);
and U2615 (N_2615,N_2575,N_2558);
or U2616 (N_2616,N_2537,N_2520);
and U2617 (N_2617,N_2535,N_2572);
xor U2618 (N_2618,N_2561,N_2556);
or U2619 (N_2619,N_2555,N_2537);
xnor U2620 (N_2620,N_2543,N_2542);
and U2621 (N_2621,N_2569,N_2562);
and U2622 (N_2622,N_2532,N_2574);
nand U2623 (N_2623,N_2574,N_2533);
nand U2624 (N_2624,N_2559,N_2524);
or U2625 (N_2625,N_2559,N_2564);
nand U2626 (N_2626,N_2543,N_2557);
nor U2627 (N_2627,N_2568,N_2556);
nor U2628 (N_2628,N_2575,N_2531);
and U2629 (N_2629,N_2552,N_2562);
nand U2630 (N_2630,N_2553,N_2523);
and U2631 (N_2631,N_2527,N_2522);
and U2632 (N_2632,N_2565,N_2532);
and U2633 (N_2633,N_2561,N_2539);
and U2634 (N_2634,N_2547,N_2575);
nand U2635 (N_2635,N_2572,N_2524);
nand U2636 (N_2636,N_2569,N_2528);
nand U2637 (N_2637,N_2574,N_2535);
nor U2638 (N_2638,N_2548,N_2555);
nor U2639 (N_2639,N_2528,N_2530);
or U2640 (N_2640,N_2622,N_2597);
nand U2641 (N_2641,N_2616,N_2637);
or U2642 (N_2642,N_2606,N_2625);
or U2643 (N_2643,N_2627,N_2582);
nor U2644 (N_2644,N_2594,N_2611);
nand U2645 (N_2645,N_2595,N_2619);
nand U2646 (N_2646,N_2588,N_2598);
nand U2647 (N_2647,N_2609,N_2618);
or U2648 (N_2648,N_2602,N_2634);
or U2649 (N_2649,N_2633,N_2613);
nor U2650 (N_2650,N_2638,N_2585);
and U2651 (N_2651,N_2580,N_2621);
or U2652 (N_2652,N_2614,N_2636);
nor U2653 (N_2653,N_2632,N_2629);
xor U2654 (N_2654,N_2583,N_2612);
and U2655 (N_2655,N_2605,N_2635);
xnor U2656 (N_2656,N_2615,N_2599);
nor U2657 (N_2657,N_2586,N_2610);
nand U2658 (N_2658,N_2601,N_2600);
and U2659 (N_2659,N_2630,N_2608);
nand U2660 (N_2660,N_2617,N_2596);
and U2661 (N_2661,N_2607,N_2589);
and U2662 (N_2662,N_2624,N_2592);
and U2663 (N_2663,N_2591,N_2623);
or U2664 (N_2664,N_2587,N_2593);
and U2665 (N_2665,N_2604,N_2631);
or U2666 (N_2666,N_2639,N_2581);
nor U2667 (N_2667,N_2626,N_2620);
nand U2668 (N_2668,N_2603,N_2590);
xnor U2669 (N_2669,N_2584,N_2628);
and U2670 (N_2670,N_2634,N_2619);
or U2671 (N_2671,N_2607,N_2585);
nand U2672 (N_2672,N_2624,N_2586);
nand U2673 (N_2673,N_2602,N_2621);
nor U2674 (N_2674,N_2586,N_2616);
and U2675 (N_2675,N_2587,N_2629);
and U2676 (N_2676,N_2595,N_2639);
or U2677 (N_2677,N_2614,N_2596);
nand U2678 (N_2678,N_2583,N_2639);
or U2679 (N_2679,N_2619,N_2584);
nor U2680 (N_2680,N_2608,N_2625);
and U2681 (N_2681,N_2623,N_2635);
nor U2682 (N_2682,N_2599,N_2601);
nand U2683 (N_2683,N_2631,N_2615);
and U2684 (N_2684,N_2633,N_2623);
and U2685 (N_2685,N_2630,N_2589);
or U2686 (N_2686,N_2609,N_2583);
xnor U2687 (N_2687,N_2619,N_2624);
or U2688 (N_2688,N_2590,N_2623);
or U2689 (N_2689,N_2627,N_2611);
or U2690 (N_2690,N_2591,N_2617);
or U2691 (N_2691,N_2580,N_2624);
xnor U2692 (N_2692,N_2623,N_2580);
nor U2693 (N_2693,N_2609,N_2589);
or U2694 (N_2694,N_2606,N_2580);
xor U2695 (N_2695,N_2601,N_2611);
nand U2696 (N_2696,N_2606,N_2639);
nor U2697 (N_2697,N_2629,N_2612);
or U2698 (N_2698,N_2600,N_2589);
and U2699 (N_2699,N_2596,N_2600);
and U2700 (N_2700,N_2656,N_2668);
or U2701 (N_2701,N_2661,N_2681);
and U2702 (N_2702,N_2657,N_2673);
or U2703 (N_2703,N_2685,N_2692);
and U2704 (N_2704,N_2658,N_2675);
xnor U2705 (N_2705,N_2671,N_2697);
nand U2706 (N_2706,N_2699,N_2660);
and U2707 (N_2707,N_2651,N_2647);
xnor U2708 (N_2708,N_2683,N_2687);
and U2709 (N_2709,N_2643,N_2677);
nor U2710 (N_2710,N_2640,N_2649);
nor U2711 (N_2711,N_2672,N_2652);
nor U2712 (N_2712,N_2642,N_2644);
and U2713 (N_2713,N_2665,N_2648);
and U2714 (N_2714,N_2662,N_2689);
nor U2715 (N_2715,N_2663,N_2688);
and U2716 (N_2716,N_2694,N_2674);
nor U2717 (N_2717,N_2670,N_2696);
nor U2718 (N_2718,N_2679,N_2669);
and U2719 (N_2719,N_2682,N_2686);
and U2720 (N_2720,N_2650,N_2693);
and U2721 (N_2721,N_2680,N_2654);
and U2722 (N_2722,N_2676,N_2684);
nor U2723 (N_2723,N_2678,N_2664);
nand U2724 (N_2724,N_2645,N_2666);
and U2725 (N_2725,N_2659,N_2646);
xor U2726 (N_2726,N_2655,N_2641);
and U2727 (N_2727,N_2695,N_2653);
xnor U2728 (N_2728,N_2667,N_2698);
and U2729 (N_2729,N_2690,N_2691);
and U2730 (N_2730,N_2668,N_2697);
nand U2731 (N_2731,N_2664,N_2658);
and U2732 (N_2732,N_2643,N_2644);
or U2733 (N_2733,N_2688,N_2697);
nor U2734 (N_2734,N_2695,N_2680);
or U2735 (N_2735,N_2647,N_2658);
nor U2736 (N_2736,N_2692,N_2682);
and U2737 (N_2737,N_2673,N_2671);
nand U2738 (N_2738,N_2655,N_2659);
nor U2739 (N_2739,N_2652,N_2699);
or U2740 (N_2740,N_2672,N_2670);
nand U2741 (N_2741,N_2659,N_2688);
or U2742 (N_2742,N_2673,N_2659);
nand U2743 (N_2743,N_2686,N_2683);
xnor U2744 (N_2744,N_2660,N_2657);
nand U2745 (N_2745,N_2664,N_2666);
and U2746 (N_2746,N_2652,N_2641);
nand U2747 (N_2747,N_2671,N_2666);
xnor U2748 (N_2748,N_2697,N_2659);
or U2749 (N_2749,N_2673,N_2649);
nand U2750 (N_2750,N_2680,N_2649);
and U2751 (N_2751,N_2675,N_2662);
nor U2752 (N_2752,N_2645,N_2696);
or U2753 (N_2753,N_2665,N_2659);
or U2754 (N_2754,N_2698,N_2682);
nand U2755 (N_2755,N_2658,N_2698);
nor U2756 (N_2756,N_2665,N_2641);
and U2757 (N_2757,N_2652,N_2654);
nor U2758 (N_2758,N_2685,N_2651);
or U2759 (N_2759,N_2652,N_2643);
or U2760 (N_2760,N_2704,N_2701);
nand U2761 (N_2761,N_2732,N_2757);
xor U2762 (N_2762,N_2733,N_2756);
nor U2763 (N_2763,N_2758,N_2739);
nor U2764 (N_2764,N_2721,N_2720);
nor U2765 (N_2765,N_2755,N_2700);
nand U2766 (N_2766,N_2729,N_2745);
xor U2767 (N_2767,N_2746,N_2708);
xnor U2768 (N_2768,N_2703,N_2741);
and U2769 (N_2769,N_2743,N_2725);
nor U2770 (N_2770,N_2734,N_2705);
or U2771 (N_2771,N_2710,N_2717);
and U2772 (N_2772,N_2707,N_2711);
and U2773 (N_2773,N_2722,N_2753);
xor U2774 (N_2774,N_2728,N_2714);
nor U2775 (N_2775,N_2747,N_2738);
or U2776 (N_2776,N_2713,N_2706);
nand U2777 (N_2777,N_2727,N_2742);
nor U2778 (N_2778,N_2759,N_2736);
or U2779 (N_2779,N_2735,N_2715);
nor U2780 (N_2780,N_2716,N_2752);
nor U2781 (N_2781,N_2730,N_2702);
or U2782 (N_2782,N_2749,N_2744);
and U2783 (N_2783,N_2709,N_2751);
nor U2784 (N_2784,N_2731,N_2748);
xor U2785 (N_2785,N_2750,N_2740);
or U2786 (N_2786,N_2724,N_2712);
or U2787 (N_2787,N_2754,N_2726);
nor U2788 (N_2788,N_2737,N_2718);
nand U2789 (N_2789,N_2719,N_2723);
nand U2790 (N_2790,N_2758,N_2707);
or U2791 (N_2791,N_2730,N_2741);
xor U2792 (N_2792,N_2708,N_2729);
and U2793 (N_2793,N_2715,N_2730);
nor U2794 (N_2794,N_2739,N_2707);
and U2795 (N_2795,N_2700,N_2750);
and U2796 (N_2796,N_2718,N_2709);
nand U2797 (N_2797,N_2757,N_2723);
nand U2798 (N_2798,N_2731,N_2756);
nand U2799 (N_2799,N_2723,N_2724);
and U2800 (N_2800,N_2728,N_2743);
and U2801 (N_2801,N_2705,N_2723);
and U2802 (N_2802,N_2742,N_2718);
nor U2803 (N_2803,N_2722,N_2746);
or U2804 (N_2804,N_2754,N_2746);
nand U2805 (N_2805,N_2707,N_2728);
and U2806 (N_2806,N_2700,N_2754);
or U2807 (N_2807,N_2731,N_2721);
nand U2808 (N_2808,N_2712,N_2730);
nand U2809 (N_2809,N_2759,N_2740);
nor U2810 (N_2810,N_2716,N_2738);
nand U2811 (N_2811,N_2713,N_2742);
or U2812 (N_2812,N_2717,N_2703);
and U2813 (N_2813,N_2707,N_2721);
xor U2814 (N_2814,N_2723,N_2734);
nor U2815 (N_2815,N_2713,N_2715);
nor U2816 (N_2816,N_2758,N_2752);
or U2817 (N_2817,N_2700,N_2725);
nand U2818 (N_2818,N_2754,N_2731);
and U2819 (N_2819,N_2752,N_2712);
or U2820 (N_2820,N_2772,N_2764);
and U2821 (N_2821,N_2777,N_2766);
or U2822 (N_2822,N_2769,N_2760);
or U2823 (N_2823,N_2795,N_2797);
nor U2824 (N_2824,N_2773,N_2801);
nor U2825 (N_2825,N_2806,N_2793);
nor U2826 (N_2826,N_2816,N_2812);
nand U2827 (N_2827,N_2788,N_2819);
and U2828 (N_2828,N_2810,N_2778);
nor U2829 (N_2829,N_2790,N_2799);
nor U2830 (N_2830,N_2805,N_2798);
nor U2831 (N_2831,N_2817,N_2802);
or U2832 (N_2832,N_2784,N_2783);
xor U2833 (N_2833,N_2779,N_2780);
and U2834 (N_2834,N_2813,N_2811);
nand U2835 (N_2835,N_2762,N_2808);
nor U2836 (N_2836,N_2765,N_2770);
xnor U2837 (N_2837,N_2767,N_2796);
or U2838 (N_2838,N_2818,N_2792);
or U2839 (N_2839,N_2785,N_2782);
or U2840 (N_2840,N_2803,N_2776);
and U2841 (N_2841,N_2787,N_2794);
nand U2842 (N_2842,N_2804,N_2789);
and U2843 (N_2843,N_2781,N_2815);
or U2844 (N_2844,N_2807,N_2771);
nand U2845 (N_2845,N_2800,N_2814);
and U2846 (N_2846,N_2786,N_2761);
nand U2847 (N_2847,N_2763,N_2768);
nor U2848 (N_2848,N_2791,N_2774);
or U2849 (N_2849,N_2775,N_2809);
or U2850 (N_2850,N_2784,N_2765);
nand U2851 (N_2851,N_2797,N_2801);
xor U2852 (N_2852,N_2778,N_2773);
nand U2853 (N_2853,N_2794,N_2789);
or U2854 (N_2854,N_2771,N_2767);
xnor U2855 (N_2855,N_2762,N_2805);
nand U2856 (N_2856,N_2803,N_2815);
nand U2857 (N_2857,N_2772,N_2799);
nor U2858 (N_2858,N_2794,N_2816);
nand U2859 (N_2859,N_2763,N_2774);
or U2860 (N_2860,N_2789,N_2780);
nor U2861 (N_2861,N_2798,N_2789);
nor U2862 (N_2862,N_2795,N_2772);
and U2863 (N_2863,N_2799,N_2773);
nor U2864 (N_2864,N_2810,N_2790);
nor U2865 (N_2865,N_2770,N_2767);
and U2866 (N_2866,N_2769,N_2810);
nand U2867 (N_2867,N_2785,N_2766);
nor U2868 (N_2868,N_2769,N_2818);
xor U2869 (N_2869,N_2790,N_2785);
nor U2870 (N_2870,N_2775,N_2801);
or U2871 (N_2871,N_2771,N_2797);
nor U2872 (N_2872,N_2804,N_2791);
nor U2873 (N_2873,N_2801,N_2782);
and U2874 (N_2874,N_2764,N_2783);
nand U2875 (N_2875,N_2796,N_2770);
and U2876 (N_2876,N_2804,N_2801);
nand U2877 (N_2877,N_2793,N_2784);
xor U2878 (N_2878,N_2791,N_2811);
and U2879 (N_2879,N_2763,N_2767);
and U2880 (N_2880,N_2838,N_2856);
nor U2881 (N_2881,N_2869,N_2872);
and U2882 (N_2882,N_2822,N_2834);
nor U2883 (N_2883,N_2868,N_2875);
xnor U2884 (N_2884,N_2845,N_2852);
and U2885 (N_2885,N_2820,N_2837);
or U2886 (N_2886,N_2859,N_2843);
nand U2887 (N_2887,N_2836,N_2844);
nand U2888 (N_2888,N_2867,N_2840);
xnor U2889 (N_2889,N_2832,N_2825);
nor U2890 (N_2890,N_2871,N_2828);
xnor U2891 (N_2891,N_2874,N_2841);
nand U2892 (N_2892,N_2830,N_2864);
nand U2893 (N_2893,N_2849,N_2865);
and U2894 (N_2894,N_2846,N_2863);
nor U2895 (N_2895,N_2824,N_2833);
and U2896 (N_2896,N_2857,N_2821);
nor U2897 (N_2897,N_2879,N_2877);
nand U2898 (N_2898,N_2870,N_2866);
nor U2899 (N_2899,N_2873,N_2839);
and U2900 (N_2900,N_2829,N_2858);
and U2901 (N_2901,N_2831,N_2855);
and U2902 (N_2902,N_2861,N_2842);
nand U2903 (N_2903,N_2876,N_2862);
or U2904 (N_2904,N_2854,N_2823);
and U2905 (N_2905,N_2826,N_2827);
nor U2906 (N_2906,N_2850,N_2878);
xnor U2907 (N_2907,N_2851,N_2853);
nor U2908 (N_2908,N_2848,N_2847);
or U2909 (N_2909,N_2835,N_2860);
nand U2910 (N_2910,N_2853,N_2843);
nor U2911 (N_2911,N_2823,N_2860);
and U2912 (N_2912,N_2822,N_2868);
nand U2913 (N_2913,N_2875,N_2822);
and U2914 (N_2914,N_2837,N_2877);
nor U2915 (N_2915,N_2838,N_2874);
nand U2916 (N_2916,N_2836,N_2860);
nand U2917 (N_2917,N_2821,N_2829);
and U2918 (N_2918,N_2821,N_2861);
nor U2919 (N_2919,N_2850,N_2879);
xnor U2920 (N_2920,N_2853,N_2865);
and U2921 (N_2921,N_2874,N_2827);
and U2922 (N_2922,N_2831,N_2878);
or U2923 (N_2923,N_2851,N_2848);
nor U2924 (N_2924,N_2866,N_2838);
nand U2925 (N_2925,N_2825,N_2838);
xnor U2926 (N_2926,N_2853,N_2845);
nand U2927 (N_2927,N_2845,N_2829);
xnor U2928 (N_2928,N_2863,N_2825);
or U2929 (N_2929,N_2871,N_2855);
nand U2930 (N_2930,N_2849,N_2879);
or U2931 (N_2931,N_2824,N_2829);
or U2932 (N_2932,N_2869,N_2861);
xor U2933 (N_2933,N_2852,N_2835);
xnor U2934 (N_2934,N_2875,N_2866);
xor U2935 (N_2935,N_2858,N_2843);
or U2936 (N_2936,N_2831,N_2877);
or U2937 (N_2937,N_2858,N_2828);
or U2938 (N_2938,N_2833,N_2874);
and U2939 (N_2939,N_2840,N_2830);
nand U2940 (N_2940,N_2891,N_2899);
nor U2941 (N_2941,N_2937,N_2922);
and U2942 (N_2942,N_2886,N_2906);
and U2943 (N_2943,N_2909,N_2910);
nor U2944 (N_2944,N_2926,N_2883);
xnor U2945 (N_2945,N_2908,N_2880);
or U2946 (N_2946,N_2912,N_2914);
and U2947 (N_2947,N_2901,N_2931);
nor U2948 (N_2948,N_2920,N_2885);
xor U2949 (N_2949,N_2896,N_2933);
or U2950 (N_2950,N_2915,N_2924);
or U2951 (N_2951,N_2928,N_2929);
or U2952 (N_2952,N_2923,N_2903);
and U2953 (N_2953,N_2918,N_2888);
nor U2954 (N_2954,N_2889,N_2893);
nand U2955 (N_2955,N_2904,N_2936);
or U2956 (N_2956,N_2881,N_2900);
nand U2957 (N_2957,N_2887,N_2917);
and U2958 (N_2958,N_2921,N_2882);
and U2959 (N_2959,N_2897,N_2925);
or U2960 (N_2960,N_2895,N_2902);
nand U2961 (N_2961,N_2892,N_2930);
and U2962 (N_2962,N_2894,N_2898);
or U2963 (N_2963,N_2907,N_2932);
nor U2964 (N_2964,N_2911,N_2884);
or U2965 (N_2965,N_2905,N_2938);
nand U2966 (N_2966,N_2935,N_2934);
and U2967 (N_2967,N_2919,N_2927);
and U2968 (N_2968,N_2890,N_2939);
or U2969 (N_2969,N_2913,N_2916);
nand U2970 (N_2970,N_2881,N_2888);
nand U2971 (N_2971,N_2929,N_2915);
nand U2972 (N_2972,N_2886,N_2896);
and U2973 (N_2973,N_2902,N_2912);
xnor U2974 (N_2974,N_2921,N_2908);
or U2975 (N_2975,N_2918,N_2912);
and U2976 (N_2976,N_2901,N_2911);
nor U2977 (N_2977,N_2907,N_2924);
and U2978 (N_2978,N_2904,N_2931);
nor U2979 (N_2979,N_2914,N_2890);
nor U2980 (N_2980,N_2894,N_2913);
nand U2981 (N_2981,N_2882,N_2930);
or U2982 (N_2982,N_2899,N_2900);
nor U2983 (N_2983,N_2938,N_2891);
nand U2984 (N_2984,N_2917,N_2924);
and U2985 (N_2985,N_2883,N_2901);
nor U2986 (N_2986,N_2916,N_2880);
nor U2987 (N_2987,N_2905,N_2923);
nand U2988 (N_2988,N_2934,N_2913);
and U2989 (N_2989,N_2907,N_2893);
or U2990 (N_2990,N_2892,N_2927);
and U2991 (N_2991,N_2906,N_2900);
and U2992 (N_2992,N_2898,N_2903);
and U2993 (N_2993,N_2936,N_2885);
and U2994 (N_2994,N_2880,N_2890);
nor U2995 (N_2995,N_2882,N_2889);
nand U2996 (N_2996,N_2927,N_2884);
nand U2997 (N_2997,N_2897,N_2923);
xnor U2998 (N_2998,N_2933,N_2892);
nor U2999 (N_2999,N_2917,N_2880);
nand UO_0 (O_0,N_2966,N_2962);
nor UO_1 (O_1,N_2985,N_2965);
nor UO_2 (O_2,N_2947,N_2954);
and UO_3 (O_3,N_2998,N_2968);
xor UO_4 (O_4,N_2997,N_2990);
nor UO_5 (O_5,N_2956,N_2958);
and UO_6 (O_6,N_2957,N_2941);
or UO_7 (O_7,N_2953,N_2963);
nand UO_8 (O_8,N_2959,N_2971);
or UO_9 (O_9,N_2942,N_2949);
xor UO_10 (O_10,N_2960,N_2994);
and UO_11 (O_11,N_2979,N_2993);
or UO_12 (O_12,N_2977,N_2951);
and UO_13 (O_13,N_2986,N_2964);
or UO_14 (O_14,N_2972,N_2982);
nor UO_15 (O_15,N_2944,N_2999);
and UO_16 (O_16,N_2984,N_2983);
nor UO_17 (O_17,N_2940,N_2961);
nor UO_18 (O_18,N_2980,N_2987);
and UO_19 (O_19,N_2952,N_2981);
nand UO_20 (O_20,N_2973,N_2969);
nor UO_21 (O_21,N_2974,N_2946);
nor UO_22 (O_22,N_2976,N_2988);
nand UO_23 (O_23,N_2943,N_2996);
nand UO_24 (O_24,N_2975,N_2955);
nand UO_25 (O_25,N_2978,N_2967);
or UO_26 (O_26,N_2992,N_2948);
nor UO_27 (O_27,N_2970,N_2991);
and UO_28 (O_28,N_2945,N_2950);
and UO_29 (O_29,N_2995,N_2989);
xor UO_30 (O_30,N_2973,N_2994);
nand UO_31 (O_31,N_2963,N_2979);
and UO_32 (O_32,N_2975,N_2982);
nor UO_33 (O_33,N_2975,N_2986);
nor UO_34 (O_34,N_2951,N_2942);
nor UO_35 (O_35,N_2999,N_2986);
and UO_36 (O_36,N_2948,N_2969);
and UO_37 (O_37,N_2981,N_2987);
nor UO_38 (O_38,N_2940,N_2967);
and UO_39 (O_39,N_2972,N_2992);
xor UO_40 (O_40,N_2988,N_2945);
or UO_41 (O_41,N_2943,N_2993);
nor UO_42 (O_42,N_2998,N_2955);
nand UO_43 (O_43,N_2962,N_2982);
and UO_44 (O_44,N_2963,N_2976);
nor UO_45 (O_45,N_2978,N_2946);
nand UO_46 (O_46,N_2977,N_2968);
nand UO_47 (O_47,N_2945,N_2973);
and UO_48 (O_48,N_2966,N_2968);
nand UO_49 (O_49,N_2960,N_2984);
xor UO_50 (O_50,N_2952,N_2960);
xor UO_51 (O_51,N_2955,N_2995);
or UO_52 (O_52,N_2961,N_2952);
nand UO_53 (O_53,N_2941,N_2977);
and UO_54 (O_54,N_2984,N_2972);
nand UO_55 (O_55,N_2962,N_2972);
or UO_56 (O_56,N_2964,N_2974);
nand UO_57 (O_57,N_2973,N_2991);
or UO_58 (O_58,N_2970,N_2950);
nor UO_59 (O_59,N_2955,N_2963);
xor UO_60 (O_60,N_2976,N_2967);
and UO_61 (O_61,N_2970,N_2997);
nor UO_62 (O_62,N_2978,N_2953);
nor UO_63 (O_63,N_2962,N_2968);
nand UO_64 (O_64,N_2991,N_2993);
and UO_65 (O_65,N_2991,N_2944);
nor UO_66 (O_66,N_2941,N_2943);
xnor UO_67 (O_67,N_2965,N_2992);
and UO_68 (O_68,N_2985,N_2953);
or UO_69 (O_69,N_2993,N_2998);
and UO_70 (O_70,N_2983,N_2979);
nand UO_71 (O_71,N_2971,N_2957);
nand UO_72 (O_72,N_2985,N_2995);
xnor UO_73 (O_73,N_2967,N_2953);
nor UO_74 (O_74,N_2986,N_2942);
nand UO_75 (O_75,N_2971,N_2976);
and UO_76 (O_76,N_2960,N_2974);
and UO_77 (O_77,N_2966,N_2967);
and UO_78 (O_78,N_2943,N_2962);
nor UO_79 (O_79,N_2959,N_2947);
xor UO_80 (O_80,N_2950,N_2975);
nor UO_81 (O_81,N_2982,N_2940);
and UO_82 (O_82,N_2969,N_2985);
and UO_83 (O_83,N_2962,N_2960);
nand UO_84 (O_84,N_2999,N_2991);
nand UO_85 (O_85,N_2955,N_2950);
and UO_86 (O_86,N_2960,N_2961);
xnor UO_87 (O_87,N_2949,N_2967);
nor UO_88 (O_88,N_2986,N_2941);
or UO_89 (O_89,N_2995,N_2958);
or UO_90 (O_90,N_2994,N_2949);
and UO_91 (O_91,N_2992,N_2995);
and UO_92 (O_92,N_2971,N_2960);
or UO_93 (O_93,N_2989,N_2988);
and UO_94 (O_94,N_2987,N_2971);
xor UO_95 (O_95,N_2982,N_2950);
or UO_96 (O_96,N_2979,N_2962);
and UO_97 (O_97,N_2945,N_2983);
and UO_98 (O_98,N_2975,N_2992);
nand UO_99 (O_99,N_2978,N_2954);
or UO_100 (O_100,N_2944,N_2956);
and UO_101 (O_101,N_2979,N_2948);
and UO_102 (O_102,N_2941,N_2976);
and UO_103 (O_103,N_2949,N_2956);
xor UO_104 (O_104,N_2953,N_2960);
nor UO_105 (O_105,N_2950,N_2963);
nor UO_106 (O_106,N_2990,N_2944);
nand UO_107 (O_107,N_2941,N_2944);
nor UO_108 (O_108,N_2987,N_2969);
nor UO_109 (O_109,N_2990,N_2982);
nor UO_110 (O_110,N_2994,N_2947);
xor UO_111 (O_111,N_2995,N_2991);
nor UO_112 (O_112,N_2968,N_2976);
nand UO_113 (O_113,N_2993,N_2953);
or UO_114 (O_114,N_2970,N_2963);
nand UO_115 (O_115,N_2990,N_2992);
and UO_116 (O_116,N_2985,N_2971);
or UO_117 (O_117,N_2966,N_2947);
nand UO_118 (O_118,N_2947,N_2973);
nand UO_119 (O_119,N_2991,N_2959);
nor UO_120 (O_120,N_2960,N_2999);
and UO_121 (O_121,N_2961,N_2992);
or UO_122 (O_122,N_2971,N_2945);
nand UO_123 (O_123,N_2952,N_2999);
nor UO_124 (O_124,N_2987,N_2986);
and UO_125 (O_125,N_2995,N_2943);
nand UO_126 (O_126,N_2957,N_2983);
nor UO_127 (O_127,N_2982,N_2960);
and UO_128 (O_128,N_2944,N_2966);
or UO_129 (O_129,N_2996,N_2970);
or UO_130 (O_130,N_2974,N_2966);
nand UO_131 (O_131,N_2961,N_2954);
and UO_132 (O_132,N_2981,N_2994);
xor UO_133 (O_133,N_2971,N_2988);
and UO_134 (O_134,N_2963,N_2961);
or UO_135 (O_135,N_2956,N_2975);
and UO_136 (O_136,N_2952,N_2969);
nor UO_137 (O_137,N_2962,N_2985);
or UO_138 (O_138,N_2973,N_2950);
or UO_139 (O_139,N_2989,N_2940);
xor UO_140 (O_140,N_2951,N_2967);
xor UO_141 (O_141,N_2975,N_2996);
and UO_142 (O_142,N_2969,N_2949);
or UO_143 (O_143,N_2981,N_2959);
and UO_144 (O_144,N_2955,N_2964);
xnor UO_145 (O_145,N_2983,N_2982);
nor UO_146 (O_146,N_2994,N_2943);
xor UO_147 (O_147,N_2988,N_2981);
and UO_148 (O_148,N_2993,N_2994);
xnor UO_149 (O_149,N_2973,N_2940);
or UO_150 (O_150,N_2984,N_2951);
or UO_151 (O_151,N_2958,N_2954);
and UO_152 (O_152,N_2966,N_2951);
nor UO_153 (O_153,N_2975,N_2993);
nor UO_154 (O_154,N_2943,N_2972);
and UO_155 (O_155,N_2988,N_2958);
or UO_156 (O_156,N_2966,N_2981);
nand UO_157 (O_157,N_2955,N_2997);
nor UO_158 (O_158,N_2977,N_2953);
xor UO_159 (O_159,N_2962,N_2989);
nand UO_160 (O_160,N_2984,N_2978);
and UO_161 (O_161,N_2978,N_2981);
or UO_162 (O_162,N_2956,N_2973);
or UO_163 (O_163,N_2965,N_2982);
or UO_164 (O_164,N_2981,N_2991);
nor UO_165 (O_165,N_2970,N_2959);
nor UO_166 (O_166,N_2958,N_2989);
and UO_167 (O_167,N_2948,N_2961);
and UO_168 (O_168,N_2987,N_2972);
nand UO_169 (O_169,N_2940,N_2963);
nor UO_170 (O_170,N_2944,N_2963);
nand UO_171 (O_171,N_2952,N_2941);
nand UO_172 (O_172,N_2991,N_2953);
nor UO_173 (O_173,N_2950,N_2957);
xor UO_174 (O_174,N_2979,N_2991);
nor UO_175 (O_175,N_2971,N_2977);
or UO_176 (O_176,N_2959,N_2950);
or UO_177 (O_177,N_2995,N_2966);
nand UO_178 (O_178,N_2980,N_2944);
nand UO_179 (O_179,N_2987,N_2945);
and UO_180 (O_180,N_2985,N_2990);
nand UO_181 (O_181,N_2991,N_2978);
xor UO_182 (O_182,N_2999,N_2974);
nor UO_183 (O_183,N_2985,N_2966);
or UO_184 (O_184,N_2953,N_2980);
or UO_185 (O_185,N_2953,N_2951);
xor UO_186 (O_186,N_2956,N_2979);
and UO_187 (O_187,N_2948,N_2959);
nand UO_188 (O_188,N_2974,N_2951);
or UO_189 (O_189,N_2944,N_2973);
nor UO_190 (O_190,N_2985,N_2959);
and UO_191 (O_191,N_2940,N_2977);
and UO_192 (O_192,N_2996,N_2990);
nand UO_193 (O_193,N_2957,N_2953);
nand UO_194 (O_194,N_2940,N_2960);
nor UO_195 (O_195,N_2995,N_2967);
nor UO_196 (O_196,N_2953,N_2950);
xor UO_197 (O_197,N_2989,N_2945);
nand UO_198 (O_198,N_2943,N_2998);
nor UO_199 (O_199,N_2990,N_2952);
nand UO_200 (O_200,N_2976,N_2961);
and UO_201 (O_201,N_2972,N_2970);
or UO_202 (O_202,N_2992,N_2940);
nor UO_203 (O_203,N_2963,N_2943);
or UO_204 (O_204,N_2972,N_2997);
and UO_205 (O_205,N_2962,N_2990);
nand UO_206 (O_206,N_2965,N_2943);
nand UO_207 (O_207,N_2994,N_2989);
nand UO_208 (O_208,N_2997,N_2987);
nand UO_209 (O_209,N_2959,N_2983);
and UO_210 (O_210,N_2945,N_2999);
and UO_211 (O_211,N_2941,N_2988);
or UO_212 (O_212,N_2990,N_2989);
and UO_213 (O_213,N_2973,N_2996);
nor UO_214 (O_214,N_2984,N_2995);
nand UO_215 (O_215,N_2982,N_2998);
nand UO_216 (O_216,N_2941,N_2974);
nand UO_217 (O_217,N_2969,N_2986);
nor UO_218 (O_218,N_2986,N_2997);
nand UO_219 (O_219,N_2952,N_2963);
and UO_220 (O_220,N_2947,N_2941);
and UO_221 (O_221,N_2947,N_2980);
nand UO_222 (O_222,N_2989,N_2977);
nand UO_223 (O_223,N_2947,N_2982);
or UO_224 (O_224,N_2989,N_2976);
nand UO_225 (O_225,N_2951,N_2945);
and UO_226 (O_226,N_2950,N_2951);
or UO_227 (O_227,N_2946,N_2973);
or UO_228 (O_228,N_2972,N_2961);
or UO_229 (O_229,N_2999,N_2987);
or UO_230 (O_230,N_2955,N_2948);
and UO_231 (O_231,N_2940,N_2966);
nand UO_232 (O_232,N_2972,N_2952);
nor UO_233 (O_233,N_2972,N_2993);
or UO_234 (O_234,N_2991,N_2988);
nor UO_235 (O_235,N_2977,N_2961);
nand UO_236 (O_236,N_2999,N_2981);
and UO_237 (O_237,N_2998,N_2985);
xnor UO_238 (O_238,N_2972,N_2996);
nand UO_239 (O_239,N_2978,N_2943);
xnor UO_240 (O_240,N_2969,N_2978);
nor UO_241 (O_241,N_2961,N_2991);
nand UO_242 (O_242,N_2941,N_2982);
and UO_243 (O_243,N_2994,N_2942);
or UO_244 (O_244,N_2948,N_2954);
or UO_245 (O_245,N_2947,N_2942);
nand UO_246 (O_246,N_2940,N_2947);
xnor UO_247 (O_247,N_2964,N_2994);
and UO_248 (O_248,N_2992,N_2982);
nor UO_249 (O_249,N_2940,N_2956);
nor UO_250 (O_250,N_2981,N_2974);
nand UO_251 (O_251,N_2973,N_2967);
nand UO_252 (O_252,N_2989,N_2991);
nor UO_253 (O_253,N_2947,N_2968);
nor UO_254 (O_254,N_2996,N_2994);
nand UO_255 (O_255,N_2991,N_2965);
and UO_256 (O_256,N_2957,N_2952);
nand UO_257 (O_257,N_2988,N_2986);
nand UO_258 (O_258,N_2984,N_2961);
or UO_259 (O_259,N_2942,N_2962);
or UO_260 (O_260,N_2962,N_2992);
nor UO_261 (O_261,N_2968,N_2941);
or UO_262 (O_262,N_2981,N_2948);
nor UO_263 (O_263,N_2973,N_2990);
nand UO_264 (O_264,N_2963,N_2982);
and UO_265 (O_265,N_2969,N_2995);
nor UO_266 (O_266,N_2947,N_2964);
xor UO_267 (O_267,N_2941,N_2949);
nor UO_268 (O_268,N_2960,N_2968);
nand UO_269 (O_269,N_2942,N_2960);
or UO_270 (O_270,N_2996,N_2958);
nand UO_271 (O_271,N_2987,N_2991);
and UO_272 (O_272,N_2945,N_2960);
nor UO_273 (O_273,N_2951,N_2946);
nor UO_274 (O_274,N_2961,N_2943);
nor UO_275 (O_275,N_2984,N_2996);
xnor UO_276 (O_276,N_2994,N_2992);
or UO_277 (O_277,N_2962,N_2975);
nor UO_278 (O_278,N_2981,N_2992);
and UO_279 (O_279,N_2946,N_2972);
or UO_280 (O_280,N_2958,N_2999);
and UO_281 (O_281,N_2982,N_2969);
nand UO_282 (O_282,N_2986,N_2972);
nor UO_283 (O_283,N_2988,N_2963);
nand UO_284 (O_284,N_2985,N_2946);
nor UO_285 (O_285,N_2955,N_2985);
nand UO_286 (O_286,N_2978,N_2979);
xnor UO_287 (O_287,N_2986,N_2992);
or UO_288 (O_288,N_2969,N_2946);
nor UO_289 (O_289,N_2998,N_2989);
xnor UO_290 (O_290,N_2976,N_2946);
or UO_291 (O_291,N_2956,N_2992);
and UO_292 (O_292,N_2951,N_2975);
xnor UO_293 (O_293,N_2994,N_2984);
nor UO_294 (O_294,N_2989,N_2966);
nor UO_295 (O_295,N_2961,N_2944);
nand UO_296 (O_296,N_2968,N_2944);
or UO_297 (O_297,N_2983,N_2965);
nand UO_298 (O_298,N_2956,N_2994);
xor UO_299 (O_299,N_2946,N_2952);
or UO_300 (O_300,N_2970,N_2953);
or UO_301 (O_301,N_2995,N_2983);
and UO_302 (O_302,N_2974,N_2992);
and UO_303 (O_303,N_2969,N_2968);
and UO_304 (O_304,N_2984,N_2985);
or UO_305 (O_305,N_2967,N_2991);
nand UO_306 (O_306,N_2948,N_2963);
and UO_307 (O_307,N_2993,N_2940);
nor UO_308 (O_308,N_2950,N_2965);
nand UO_309 (O_309,N_2981,N_2956);
and UO_310 (O_310,N_2953,N_2994);
nor UO_311 (O_311,N_2988,N_2972);
and UO_312 (O_312,N_2991,N_2962);
nand UO_313 (O_313,N_2980,N_2976);
and UO_314 (O_314,N_2982,N_2997);
nand UO_315 (O_315,N_2983,N_2997);
nor UO_316 (O_316,N_2966,N_2972);
or UO_317 (O_317,N_2957,N_2988);
or UO_318 (O_318,N_2999,N_2943);
and UO_319 (O_319,N_2996,N_2998);
and UO_320 (O_320,N_2983,N_2980);
and UO_321 (O_321,N_2951,N_2997);
nor UO_322 (O_322,N_2975,N_2944);
xor UO_323 (O_323,N_2945,N_2968);
and UO_324 (O_324,N_2989,N_2969);
xnor UO_325 (O_325,N_2953,N_2952);
or UO_326 (O_326,N_2943,N_2967);
nand UO_327 (O_327,N_2992,N_2955);
or UO_328 (O_328,N_2952,N_2989);
nand UO_329 (O_329,N_2952,N_2998);
xor UO_330 (O_330,N_2957,N_2990);
nor UO_331 (O_331,N_2977,N_2983);
nor UO_332 (O_332,N_2948,N_2990);
nand UO_333 (O_333,N_2968,N_2995);
nand UO_334 (O_334,N_2964,N_2973);
nor UO_335 (O_335,N_2963,N_2959);
or UO_336 (O_336,N_2949,N_2979);
xor UO_337 (O_337,N_2958,N_2976);
nand UO_338 (O_338,N_2985,N_2972);
nor UO_339 (O_339,N_2995,N_2986);
and UO_340 (O_340,N_2980,N_2961);
and UO_341 (O_341,N_2986,N_2965);
nand UO_342 (O_342,N_2993,N_2976);
nor UO_343 (O_343,N_2963,N_2995);
or UO_344 (O_344,N_2944,N_2950);
nand UO_345 (O_345,N_2966,N_2986);
nor UO_346 (O_346,N_2989,N_2987);
or UO_347 (O_347,N_2979,N_2996);
nand UO_348 (O_348,N_2960,N_2946);
and UO_349 (O_349,N_2941,N_2958);
nor UO_350 (O_350,N_2968,N_2985);
nor UO_351 (O_351,N_2997,N_2959);
and UO_352 (O_352,N_2995,N_2949);
nor UO_353 (O_353,N_2944,N_2974);
or UO_354 (O_354,N_2951,N_2980);
nor UO_355 (O_355,N_2980,N_2940);
nand UO_356 (O_356,N_2966,N_2983);
or UO_357 (O_357,N_2952,N_2977);
nand UO_358 (O_358,N_2978,N_2996);
or UO_359 (O_359,N_2963,N_2969);
nor UO_360 (O_360,N_2960,N_2948);
nor UO_361 (O_361,N_2984,N_2982);
nor UO_362 (O_362,N_2980,N_2960);
nor UO_363 (O_363,N_2987,N_2990);
or UO_364 (O_364,N_2987,N_2940);
nor UO_365 (O_365,N_2994,N_2986);
xor UO_366 (O_366,N_2954,N_2979);
and UO_367 (O_367,N_2969,N_2962);
nand UO_368 (O_368,N_2972,N_2964);
xnor UO_369 (O_369,N_2978,N_2942);
or UO_370 (O_370,N_2993,N_2971);
and UO_371 (O_371,N_2983,N_2990);
and UO_372 (O_372,N_2970,N_2987);
nand UO_373 (O_373,N_2973,N_2979);
nand UO_374 (O_374,N_2945,N_2953);
or UO_375 (O_375,N_2969,N_2958);
or UO_376 (O_376,N_2965,N_2981);
and UO_377 (O_377,N_2950,N_2972);
and UO_378 (O_378,N_2941,N_2956);
and UO_379 (O_379,N_2974,N_2965);
and UO_380 (O_380,N_2985,N_2956);
nor UO_381 (O_381,N_2943,N_2949);
nand UO_382 (O_382,N_2973,N_2942);
nand UO_383 (O_383,N_2998,N_2949);
nand UO_384 (O_384,N_2980,N_2943);
and UO_385 (O_385,N_2966,N_2950);
and UO_386 (O_386,N_2978,N_2948);
or UO_387 (O_387,N_2943,N_2986);
or UO_388 (O_388,N_2994,N_2982);
or UO_389 (O_389,N_2991,N_2960);
or UO_390 (O_390,N_2959,N_2946);
nand UO_391 (O_391,N_2941,N_2951);
xor UO_392 (O_392,N_2946,N_2950);
nor UO_393 (O_393,N_2942,N_2956);
or UO_394 (O_394,N_2967,N_2998);
and UO_395 (O_395,N_2980,N_2993);
nand UO_396 (O_396,N_2987,N_2983);
nor UO_397 (O_397,N_2966,N_2961);
nor UO_398 (O_398,N_2971,N_2952);
nand UO_399 (O_399,N_2993,N_2981);
or UO_400 (O_400,N_2994,N_2970);
or UO_401 (O_401,N_2961,N_2974);
and UO_402 (O_402,N_2965,N_2945);
nand UO_403 (O_403,N_2946,N_2943);
and UO_404 (O_404,N_2989,N_2983);
and UO_405 (O_405,N_2950,N_2942);
or UO_406 (O_406,N_2996,N_2967);
and UO_407 (O_407,N_2957,N_2993);
or UO_408 (O_408,N_2948,N_2985);
or UO_409 (O_409,N_2982,N_2966);
and UO_410 (O_410,N_2992,N_2947);
or UO_411 (O_411,N_2997,N_2963);
nand UO_412 (O_412,N_2951,N_2959);
and UO_413 (O_413,N_2951,N_2952);
nor UO_414 (O_414,N_2967,N_2954);
nand UO_415 (O_415,N_2997,N_2975);
nand UO_416 (O_416,N_2990,N_2984);
and UO_417 (O_417,N_2945,N_2991);
nand UO_418 (O_418,N_2976,N_2978);
or UO_419 (O_419,N_2944,N_2945);
nand UO_420 (O_420,N_2947,N_2993);
or UO_421 (O_421,N_2946,N_2999);
nand UO_422 (O_422,N_2943,N_2979);
or UO_423 (O_423,N_2974,N_2980);
nand UO_424 (O_424,N_2955,N_2989);
and UO_425 (O_425,N_2970,N_2966);
nor UO_426 (O_426,N_2965,N_2998);
and UO_427 (O_427,N_2945,N_2984);
nand UO_428 (O_428,N_2974,N_2977);
nand UO_429 (O_429,N_2989,N_2947);
nor UO_430 (O_430,N_2985,N_2945);
and UO_431 (O_431,N_2960,N_2990);
nor UO_432 (O_432,N_2994,N_2954);
nand UO_433 (O_433,N_2974,N_2956);
and UO_434 (O_434,N_2955,N_2971);
and UO_435 (O_435,N_2965,N_2975);
or UO_436 (O_436,N_2986,N_2963);
and UO_437 (O_437,N_2952,N_2997);
nor UO_438 (O_438,N_2957,N_2959);
nor UO_439 (O_439,N_2945,N_2957);
and UO_440 (O_440,N_2979,N_2946);
nand UO_441 (O_441,N_2979,N_2989);
nand UO_442 (O_442,N_2995,N_2978);
or UO_443 (O_443,N_2980,N_2946);
and UO_444 (O_444,N_2986,N_2978);
or UO_445 (O_445,N_2964,N_2999);
nand UO_446 (O_446,N_2976,N_2981);
and UO_447 (O_447,N_2984,N_2940);
or UO_448 (O_448,N_2972,N_2955);
nand UO_449 (O_449,N_2999,N_2963);
and UO_450 (O_450,N_2944,N_2949);
nand UO_451 (O_451,N_2998,N_2994);
or UO_452 (O_452,N_2949,N_2946);
and UO_453 (O_453,N_2971,N_2944);
and UO_454 (O_454,N_2997,N_2977);
xor UO_455 (O_455,N_2951,N_2954);
or UO_456 (O_456,N_2982,N_2956);
and UO_457 (O_457,N_2952,N_2991);
and UO_458 (O_458,N_2941,N_2962);
xnor UO_459 (O_459,N_2991,N_2976);
nand UO_460 (O_460,N_2975,N_2979);
nand UO_461 (O_461,N_2987,N_2943);
nand UO_462 (O_462,N_2991,N_2975);
nor UO_463 (O_463,N_2996,N_2956);
or UO_464 (O_464,N_2976,N_2957);
and UO_465 (O_465,N_2977,N_2999);
or UO_466 (O_466,N_2961,N_2978);
nand UO_467 (O_467,N_2945,N_2977);
or UO_468 (O_468,N_2942,N_2964);
or UO_469 (O_469,N_2989,N_2953);
or UO_470 (O_470,N_2945,N_2956);
nand UO_471 (O_471,N_2981,N_2945);
or UO_472 (O_472,N_2960,N_2998);
or UO_473 (O_473,N_2962,N_2988);
and UO_474 (O_474,N_2990,N_2998);
nand UO_475 (O_475,N_2990,N_2979);
nor UO_476 (O_476,N_2980,N_2949);
or UO_477 (O_477,N_2955,N_2942);
nor UO_478 (O_478,N_2948,N_2966);
or UO_479 (O_479,N_2965,N_2951);
or UO_480 (O_480,N_2950,N_2947);
xnor UO_481 (O_481,N_2972,N_2945);
nor UO_482 (O_482,N_2989,N_2997);
or UO_483 (O_483,N_2950,N_2967);
or UO_484 (O_484,N_2988,N_2967);
nand UO_485 (O_485,N_2980,N_2969);
and UO_486 (O_486,N_2947,N_2943);
or UO_487 (O_487,N_2944,N_2983);
nand UO_488 (O_488,N_2971,N_2986);
xor UO_489 (O_489,N_2951,N_2973);
or UO_490 (O_490,N_2945,N_2941);
nor UO_491 (O_491,N_2947,N_2948);
and UO_492 (O_492,N_2961,N_2970);
or UO_493 (O_493,N_2954,N_2949);
or UO_494 (O_494,N_2943,N_2988);
xnor UO_495 (O_495,N_2952,N_2956);
or UO_496 (O_496,N_2948,N_2982);
nand UO_497 (O_497,N_2961,N_2945);
nand UO_498 (O_498,N_2946,N_2958);
nand UO_499 (O_499,N_2952,N_2980);
endmodule