module basic_1500_15000_2000_5_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xor U0 (N_0,In_1057,In_583);
xor U1 (N_1,In_743,In_1432);
and U2 (N_2,In_98,In_1451);
xor U3 (N_3,In_578,In_99);
or U4 (N_4,In_1472,In_808);
nand U5 (N_5,In_279,In_892);
xor U6 (N_6,In_1207,In_1397);
and U7 (N_7,In_1026,In_1493);
and U8 (N_8,In_1134,In_947);
xor U9 (N_9,In_931,In_1232);
nor U10 (N_10,In_829,In_24);
or U11 (N_11,In_684,In_122);
xnor U12 (N_12,In_955,In_486);
or U13 (N_13,In_1117,In_591);
and U14 (N_14,In_1238,In_354);
or U15 (N_15,In_1306,In_139);
and U16 (N_16,In_1019,In_960);
and U17 (N_17,In_538,In_1132);
xor U18 (N_18,In_225,In_864);
or U19 (N_19,In_1103,In_1473);
and U20 (N_20,In_910,In_360);
and U21 (N_21,In_235,In_537);
nor U22 (N_22,In_803,In_36);
nand U23 (N_23,In_232,In_1190);
nor U24 (N_24,In_316,In_1070);
and U25 (N_25,In_1205,In_293);
nor U26 (N_26,In_795,In_698);
nor U27 (N_27,In_938,In_985);
and U28 (N_28,In_824,In_1258);
or U29 (N_29,In_541,In_677);
nand U30 (N_30,In_1387,In_1046);
nor U31 (N_31,In_718,In_1227);
and U32 (N_32,In_30,In_7);
and U33 (N_33,In_468,In_1083);
nand U34 (N_34,In_1310,In_475);
or U35 (N_35,In_593,In_1374);
nor U36 (N_36,In_791,In_635);
or U37 (N_37,In_618,In_1085);
nor U38 (N_38,In_3,In_1330);
or U39 (N_39,In_1120,In_870);
or U40 (N_40,In_1112,In_1436);
nor U41 (N_41,In_556,In_245);
and U42 (N_42,In_847,In_1323);
nor U43 (N_43,In_57,In_775);
or U44 (N_44,In_118,In_564);
xor U45 (N_45,In_776,In_18);
nand U46 (N_46,In_798,In_1253);
or U47 (N_47,In_372,In_333);
nor U48 (N_48,In_877,In_391);
and U49 (N_49,In_171,In_692);
nand U50 (N_50,In_315,In_309);
and U51 (N_51,In_432,In_143);
nand U52 (N_52,In_220,In_1101);
or U53 (N_53,In_975,In_859);
nand U54 (N_54,In_597,In_5);
nand U55 (N_55,In_280,In_1402);
nor U56 (N_56,In_1452,In_1140);
or U57 (N_57,In_147,In_828);
or U58 (N_58,In_1005,In_262);
nor U59 (N_59,In_444,In_1293);
xnor U60 (N_60,In_1437,In_230);
and U61 (N_61,In_346,In_1089);
and U62 (N_62,In_21,In_1218);
nor U63 (N_63,In_1006,In_277);
and U64 (N_64,In_336,In_1462);
or U65 (N_65,In_901,In_952);
and U66 (N_66,In_1059,In_196);
and U67 (N_67,In_519,In_325);
nand U68 (N_68,In_103,In_160);
nand U69 (N_69,In_1484,In_956);
nand U70 (N_70,In_76,In_1408);
or U71 (N_71,In_375,In_204);
or U72 (N_72,In_484,In_663);
or U73 (N_73,In_886,In_893);
nand U74 (N_74,In_1195,In_80);
xnor U75 (N_75,In_1197,In_1298);
nand U76 (N_76,In_31,In_249);
and U77 (N_77,In_1001,In_1339);
xor U78 (N_78,In_530,In_1318);
nor U79 (N_79,In_800,In_897);
or U80 (N_80,In_634,In_335);
or U81 (N_81,In_1098,In_157);
nor U82 (N_82,In_1248,In_347);
nor U83 (N_83,In_1435,In_550);
xnor U84 (N_84,In_906,In_380);
nand U85 (N_85,In_620,In_959);
nand U86 (N_86,In_883,In_894);
nand U87 (N_87,In_54,In_108);
and U88 (N_88,In_1284,In_457);
or U89 (N_89,In_744,In_246);
nor U90 (N_90,In_1349,In_650);
or U91 (N_91,In_1210,In_382);
nand U92 (N_92,In_546,In_1237);
nand U93 (N_93,In_345,In_281);
nor U94 (N_94,In_505,In_1077);
nor U95 (N_95,In_876,In_533);
nor U96 (N_96,In_481,In_926);
xnor U97 (N_97,In_1440,In_754);
or U98 (N_98,In_693,In_1350);
and U99 (N_99,In_502,In_882);
or U100 (N_100,In_1477,In_1383);
or U101 (N_101,In_1201,In_221);
or U102 (N_102,In_1406,In_804);
nor U103 (N_103,In_1217,In_788);
or U104 (N_104,In_1376,In_848);
nor U105 (N_105,In_590,In_446);
xnor U106 (N_106,In_781,In_855);
and U107 (N_107,In_1388,In_1476);
or U108 (N_108,In_39,In_762);
nand U109 (N_109,In_286,In_1495);
or U110 (N_110,In_951,In_95);
or U111 (N_111,In_1222,In_266);
or U112 (N_112,In_1076,In_1186);
or U113 (N_113,In_168,In_396);
nand U114 (N_114,In_1461,In_945);
nand U115 (N_115,In_615,In_77);
nor U116 (N_116,In_764,In_1123);
nand U117 (N_117,In_717,In_162);
and U118 (N_118,In_227,In_1173);
and U119 (N_119,In_1420,In_67);
nor U120 (N_120,In_254,In_87);
nor U121 (N_121,In_158,In_950);
nand U122 (N_122,In_422,In_374);
or U123 (N_123,In_19,In_154);
nor U124 (N_124,In_1028,In_1147);
nand U125 (N_125,In_362,In_265);
xnor U126 (N_126,In_837,In_469);
nor U127 (N_127,In_1039,In_708);
and U128 (N_128,In_1414,In_1290);
nor U129 (N_129,In_439,In_756);
or U130 (N_130,In_201,In_278);
xnor U131 (N_131,In_1131,In_987);
and U132 (N_132,In_202,In_657);
nand U133 (N_133,In_145,In_23);
and U134 (N_134,In_1268,In_133);
or U135 (N_135,In_1171,In_1417);
or U136 (N_136,In_988,In_236);
and U137 (N_137,In_150,In_1394);
nand U138 (N_138,In_121,In_995);
nor U139 (N_139,In_779,In_1381);
xnor U140 (N_140,In_1271,In_1266);
and U141 (N_141,In_701,In_1000);
nor U142 (N_142,In_1278,In_2);
nor U143 (N_143,In_400,In_734);
nor U144 (N_144,In_1463,In_441);
nand U145 (N_145,In_1304,In_1347);
nor U146 (N_146,In_1482,In_130);
or U147 (N_147,In_1149,In_915);
nand U148 (N_148,In_451,In_177);
nand U149 (N_149,In_120,In_1288);
nand U150 (N_150,In_1092,In_1105);
and U151 (N_151,In_367,In_416);
nor U152 (N_152,In_393,In_517);
nand U153 (N_153,In_330,In_193);
or U154 (N_154,In_102,In_1121);
and U155 (N_155,In_14,In_1024);
xor U156 (N_156,In_1236,In_1246);
nor U157 (N_157,In_211,In_1108);
or U158 (N_158,In_1273,In_1301);
nor U159 (N_159,In_482,In_1294);
or U160 (N_160,In_506,In_1165);
or U161 (N_161,In_1459,In_1156);
nand U162 (N_162,In_1254,In_17);
nand U163 (N_163,In_470,In_96);
nand U164 (N_164,In_182,In_1068);
nor U165 (N_165,In_1229,In_598);
nor U166 (N_166,In_405,In_426);
nor U167 (N_167,In_126,In_531);
and U168 (N_168,In_875,In_888);
and U169 (N_169,In_190,In_369);
xnor U170 (N_170,In_1371,In_799);
nand U171 (N_171,In_737,In_337);
or U172 (N_172,In_664,In_914);
or U173 (N_173,In_106,In_128);
and U174 (N_174,In_704,In_305);
nand U175 (N_175,In_79,In_1355);
and U176 (N_176,In_243,In_794);
xor U177 (N_177,In_332,In_71);
and U178 (N_178,In_689,In_260);
or U179 (N_179,In_1263,In_529);
nand U180 (N_180,In_1145,In_624);
nor U181 (N_181,In_1152,In_1007);
nand U182 (N_182,In_199,In_1021);
and U183 (N_183,In_408,In_1353);
nor U184 (N_184,In_1255,In_324);
and U185 (N_185,In_272,In_480);
nand U186 (N_186,In_739,In_142);
nand U187 (N_187,In_1321,In_1022);
nand U188 (N_188,In_47,In_1429);
nor U189 (N_189,In_215,In_288);
xnor U190 (N_190,In_423,In_1043);
nand U191 (N_191,In_231,In_703);
nand U192 (N_192,In_1176,In_561);
nor U193 (N_193,In_270,In_436);
or U194 (N_194,In_603,In_302);
and U195 (N_195,In_184,In_413);
nor U196 (N_196,In_1133,In_86);
or U197 (N_197,In_1390,In_1471);
or U198 (N_198,In_1213,In_290);
and U199 (N_199,In_0,In_1464);
or U200 (N_200,In_1413,In_1109);
nor U201 (N_201,In_329,In_1483);
and U202 (N_202,In_849,In_805);
nand U203 (N_203,In_666,In_760);
or U204 (N_204,In_844,In_1409);
or U205 (N_205,In_963,In_1069);
and U206 (N_206,In_1469,In_296);
nor U207 (N_207,In_746,In_429);
and U208 (N_208,In_1431,In_9);
or U209 (N_209,In_412,In_726);
or U210 (N_210,In_322,In_358);
or U211 (N_211,In_751,In_1220);
and U212 (N_212,In_6,In_180);
and U213 (N_213,In_247,In_109);
nand U214 (N_214,In_806,In_777);
xor U215 (N_215,In_1300,In_8);
xnor U216 (N_216,In_932,In_939);
and U217 (N_217,In_1317,In_474);
nand U218 (N_218,In_811,In_411);
and U219 (N_219,In_835,In_871);
nor U220 (N_220,In_1136,In_865);
or U221 (N_221,In_796,In_389);
or U222 (N_222,In_1163,In_588);
or U223 (N_223,In_169,In_729);
nor U224 (N_224,In_1179,In_1100);
nand U225 (N_225,In_673,In_1138);
or U226 (N_226,In_56,In_1322);
or U227 (N_227,In_91,In_1426);
and U228 (N_228,In_1282,In_355);
nand U229 (N_229,In_920,In_1419);
or U230 (N_230,In_1286,In_797);
and U231 (N_231,In_1257,In_1096);
or U232 (N_232,In_226,In_459);
and U233 (N_233,In_763,In_283);
nor U234 (N_234,In_287,In_404);
nor U235 (N_235,In_850,In_904);
or U236 (N_236,In_1319,In_114);
nor U237 (N_237,In_999,In_179);
nor U238 (N_238,In_818,In_579);
nand U239 (N_239,In_622,In_890);
and U240 (N_240,In_465,In_1219);
or U241 (N_241,In_1478,In_513);
and U242 (N_242,In_688,In_1392);
and U243 (N_243,In_757,In_1407);
nand U244 (N_244,In_195,In_52);
or U245 (N_245,In_802,In_267);
nand U246 (N_246,In_1405,In_364);
nand U247 (N_247,In_1428,In_532);
or U248 (N_248,In_968,In_935);
or U249 (N_249,In_617,In_881);
nor U250 (N_250,In_297,In_1228);
nor U251 (N_251,In_1211,In_1081);
nor U252 (N_252,In_1017,In_394);
nor U253 (N_253,In_826,In_1249);
nand U254 (N_254,In_1265,In_789);
or U255 (N_255,In_1256,In_1474);
nor U256 (N_256,In_725,In_420);
nor U257 (N_257,In_845,In_823);
and U258 (N_258,In_858,In_1325);
nand U259 (N_259,In_736,In_908);
and U260 (N_260,In_813,In_586);
nor U261 (N_261,In_1303,In_543);
xor U262 (N_262,In_759,In_1328);
nor U263 (N_263,In_878,In_1497);
or U264 (N_264,In_868,In_285);
nor U265 (N_265,In_1343,In_351);
nor U266 (N_266,In_239,In_210);
and U267 (N_267,In_242,In_445);
nor U268 (N_268,In_311,In_1345);
and U269 (N_269,In_765,In_275);
nand U270 (N_270,In_515,In_750);
or U271 (N_271,In_65,In_1240);
nand U272 (N_272,In_1172,In_253);
nor U273 (N_273,In_721,In_1250);
nor U274 (N_274,In_326,In_1155);
nand U275 (N_275,In_1127,In_1358);
or U276 (N_276,In_1275,In_641);
nand U277 (N_277,In_501,In_1276);
or U278 (N_278,In_705,In_790);
nand U279 (N_279,In_857,In_1455);
or U280 (N_280,In_973,In_1267);
nand U281 (N_281,In_1094,In_292);
nand U282 (N_282,In_830,In_1157);
nor U283 (N_283,In_553,In_483);
nor U284 (N_284,In_1193,In_33);
xor U285 (N_285,In_252,In_1074);
and U286 (N_286,In_1078,In_323);
nand U287 (N_287,In_496,In_1044);
and U288 (N_288,In_1064,In_1184);
and U289 (N_289,In_83,In_377);
and U290 (N_290,In_390,In_560);
and U291 (N_291,In_319,In_774);
nand U292 (N_292,In_1457,In_707);
and U293 (N_293,In_1468,In_172);
and U294 (N_294,In_1487,In_1324);
and U295 (N_295,In_499,In_25);
or U296 (N_296,In_206,In_566);
or U297 (N_297,In_584,In_1291);
nor U298 (N_298,In_646,In_152);
or U299 (N_299,In_656,In_403);
nor U300 (N_300,In_1072,In_727);
nand U301 (N_301,In_1245,In_327);
and U302 (N_302,In_58,In_846);
nand U303 (N_303,In_488,In_633);
and U304 (N_304,In_738,In_630);
and U305 (N_305,In_60,In_1456);
and U306 (N_306,In_1332,In_1490);
or U307 (N_307,In_508,In_151);
nor U308 (N_308,In_1233,In_933);
or U309 (N_309,In_214,In_385);
xnor U310 (N_310,In_820,In_1445);
nand U311 (N_311,In_32,In_148);
or U312 (N_312,In_1334,In_643);
nand U313 (N_313,In_1143,In_647);
nor U314 (N_314,In_1223,In_1385);
or U315 (N_315,In_414,In_1460);
and U316 (N_316,In_29,In_902);
or U317 (N_317,In_898,In_175);
or U318 (N_318,In_131,In_1346);
xor U319 (N_319,In_923,In_536);
nor U320 (N_320,In_417,In_1247);
or U321 (N_321,In_1041,In_683);
or U322 (N_322,In_1139,In_1354);
and U323 (N_323,In_907,In_284);
nand U324 (N_324,In_606,In_339);
nand U325 (N_325,In_1488,In_1423);
nor U326 (N_326,In_1329,In_268);
or U327 (N_327,In_1299,In_140);
nand U328 (N_328,In_318,In_1391);
nand U329 (N_329,In_1049,In_608);
nand U330 (N_330,In_1191,In_100);
or U331 (N_331,In_40,In_1313);
or U332 (N_332,In_589,In_887);
nand U333 (N_333,In_163,In_437);
or U334 (N_334,In_1104,In_1055);
and U335 (N_335,In_1002,In_1335);
or U336 (N_336,In_856,In_188);
nand U337 (N_337,In_49,In_1314);
nand U338 (N_338,In_942,In_37);
nor U339 (N_339,In_792,In_1439);
nand U340 (N_340,In_716,In_1187);
nand U341 (N_341,In_1181,In_551);
nand U342 (N_342,In_10,In_4);
nor U343 (N_343,In_1351,In_687);
nor U344 (N_344,In_1088,In_350);
nand U345 (N_345,In_1262,In_782);
and U346 (N_346,In_1344,In_982);
nand U347 (N_347,In_1090,In_16);
or U348 (N_348,In_640,In_625);
nor U349 (N_349,In_383,In_609);
and U350 (N_350,In_900,In_836);
nand U351 (N_351,In_472,In_1020);
xor U352 (N_352,In_1,In_357);
and U353 (N_353,In_1337,In_20);
or U354 (N_354,In_447,In_261);
or U355 (N_355,In_1158,In_771);
nor U356 (N_356,In_812,In_425);
nor U357 (N_357,In_809,In_1422);
nor U358 (N_358,In_395,In_338);
and U359 (N_359,In_974,In_185);
nand U360 (N_360,In_521,In_448);
nand U361 (N_361,In_768,In_922);
or U362 (N_362,In_1242,In_954);
and U363 (N_363,In_548,In_406);
nand U364 (N_364,In_569,In_1012);
and U365 (N_365,In_545,In_632);
nand U366 (N_366,In_682,In_1367);
nor U367 (N_367,In_863,In_710);
or U368 (N_368,In_753,In_219);
and U369 (N_369,In_670,In_1062);
or U370 (N_370,In_282,In_217);
nand U371 (N_371,In_1114,In_653);
and U372 (N_372,In_35,In_1489);
or U373 (N_373,In_317,In_1073);
nand U374 (N_374,In_75,In_1342);
and U375 (N_375,In_1356,In_574);
nand U376 (N_376,In_473,In_917);
or U377 (N_377,In_735,In_507);
nand U378 (N_378,In_1393,In_307);
nor U379 (N_379,In_418,In_119);
or U380 (N_380,In_1175,In_969);
and U381 (N_381,In_658,In_1368);
nor U382 (N_382,In_113,In_549);
and U383 (N_383,In_1033,In_331);
xor U384 (N_384,In_353,In_957);
and U385 (N_385,In_38,In_626);
nand U386 (N_386,In_1183,In_709);
and U387 (N_387,In_1214,In_1159);
nor U388 (N_388,In_1065,In_11);
nand U389 (N_389,In_450,In_112);
nand U390 (N_390,In_368,In_159);
nand U391 (N_391,In_758,In_471);
or U392 (N_392,In_1182,In_1365);
or U393 (N_393,In_466,In_1448);
xor U394 (N_394,In_1360,In_966);
xor U395 (N_395,In_925,In_607);
nand U396 (N_396,In_1167,In_510);
nor U397 (N_397,In_921,In_1038);
or U398 (N_398,In_1162,In_652);
xnor U399 (N_399,In_748,In_1425);
or U400 (N_400,In_415,In_853);
and U401 (N_401,In_341,In_1305);
nor U402 (N_402,In_276,In_526);
nand U403 (N_403,In_1264,In_299);
and U404 (N_404,In_174,In_1142);
and U405 (N_405,In_520,In_238);
and U406 (N_406,In_1225,In_137);
or U407 (N_407,In_1277,In_387);
nor U408 (N_408,In_1341,In_1010);
nand U409 (N_409,In_1285,In_1106);
nor U410 (N_410,In_1434,In_1169);
or U411 (N_411,In_572,In_399);
and U412 (N_412,In_460,In_685);
nor U413 (N_413,In_205,In_66);
nor U414 (N_414,In_376,In_909);
nand U415 (N_415,In_340,In_455);
nor U416 (N_416,In_1035,In_138);
xor U417 (N_417,In_117,In_594);
xnor U418 (N_418,In_321,In_134);
nand U419 (N_419,In_570,In_1308);
and U420 (N_420,In_1202,In_535);
nor U421 (N_421,In_81,In_453);
nor U422 (N_422,In_1260,In_1144);
or U423 (N_423,In_1153,In_1164);
nand U424 (N_424,In_639,In_1221);
nand U425 (N_425,In_1011,In_1364);
and U426 (N_426,In_500,In_752);
and U427 (N_427,In_1485,In_628);
nor U428 (N_428,In_613,In_841);
nor U429 (N_429,In_72,In_1036);
nand U430 (N_430,In_627,In_241);
nor U431 (N_431,In_313,In_493);
or U432 (N_432,In_1087,In_587);
or U433 (N_433,In_344,In_1058);
xnor U434 (N_434,In_554,In_248);
and U435 (N_435,In_977,In_124);
and U436 (N_436,In_69,In_310);
and U437 (N_437,In_911,In_786);
nand U438 (N_438,In_132,In_787);
nand U439 (N_439,In_73,In_967);
and U440 (N_440,In_381,In_479);
nand U441 (N_441,In_192,In_348);
nand U442 (N_442,In_378,In_741);
nand U443 (N_443,In_861,In_107);
nand U444 (N_444,In_919,In_104);
and U445 (N_445,In_306,In_294);
nor U446 (N_446,In_834,In_873);
and U447 (N_447,In_706,In_63);
or U448 (N_448,In_1018,In_880);
xnor U449 (N_449,In_1261,In_509);
nand U450 (N_450,In_300,In_50);
and U451 (N_451,In_1375,In_15);
and U452 (N_452,In_723,In_843);
xor U453 (N_453,In_821,In_662);
or U454 (N_454,In_366,In_101);
and U455 (N_455,In_438,In_623);
nor U456 (N_456,In_478,In_90);
and U457 (N_457,In_1444,In_1494);
nor U458 (N_458,In_793,In_930);
nor U459 (N_459,In_610,In_867);
nor U460 (N_460,In_1234,In_189);
nand U461 (N_461,In_116,In_714);
or U462 (N_462,In_540,In_562);
nand U463 (N_463,In_1251,In_1052);
or U464 (N_464,In_45,In_392);
and U465 (N_465,In_672,In_1185);
and U466 (N_466,In_712,In_636);
and U467 (N_467,In_962,In_251);
and U468 (N_468,In_218,In_976);
nor U469 (N_469,In_229,In_631);
nand U470 (N_470,In_1230,In_1326);
nand U471 (N_471,In_314,In_1194);
and U472 (N_472,In_1124,In_851);
and U473 (N_473,In_1411,In_523);
nor U474 (N_474,In_645,In_994);
nor U475 (N_475,In_492,In_94);
and U476 (N_476,In_233,In_839);
nand U477 (N_477,In_1281,In_720);
nor U478 (N_478,In_905,In_992);
nand U479 (N_479,In_398,In_1166);
or U480 (N_480,In_1309,In_1209);
and U481 (N_481,In_1380,In_1384);
or U482 (N_482,In_815,In_934);
or U483 (N_483,In_386,In_702);
xnor U484 (N_484,In_1279,In_1259);
xnor U485 (N_485,In_181,In_1032);
or U486 (N_486,In_1198,In_1361);
nor U487 (N_487,In_667,In_755);
or U488 (N_488,In_1453,In_1352);
xor U489 (N_489,In_53,In_1366);
nor U490 (N_490,In_141,In_1034);
or U491 (N_491,In_1216,In_518);
and U492 (N_492,In_833,In_200);
or U493 (N_493,In_485,In_495);
nand U494 (N_494,In_567,In_402);
nand U495 (N_495,In_349,In_1243);
xnor U496 (N_496,In_1446,In_1084);
nand U497 (N_497,In_884,In_660);
and U498 (N_498,In_724,In_487);
nor U499 (N_499,In_1244,In_668);
nand U500 (N_500,In_419,In_986);
nand U501 (N_501,In_832,In_1458);
or U502 (N_502,In_989,In_528);
nand U503 (N_503,In_1061,In_840);
xnor U504 (N_504,In_1091,In_749);
nand U505 (N_505,In_222,In_860);
or U506 (N_506,In_409,In_431);
nor U507 (N_507,In_504,In_649);
nand U508 (N_508,In_1292,In_1327);
xor U509 (N_509,In_105,In_780);
xnor U510 (N_510,In_70,In_213);
or U511 (N_511,In_555,In_694);
and U512 (N_512,In_715,In_170);
nand U513 (N_513,In_659,In_1315);
nand U514 (N_514,In_1016,In_223);
nand U515 (N_515,In_770,In_477);
nor U516 (N_516,In_42,In_165);
nor U517 (N_517,In_89,In_1377);
or U518 (N_518,In_454,In_494);
or U519 (N_519,In_250,In_1196);
and U520 (N_520,In_1130,In_946);
and U521 (N_521,In_12,In_971);
or U522 (N_522,In_512,In_84);
nor U523 (N_523,In_82,In_733);
nand U524 (N_524,In_123,In_810);
nand U525 (N_525,In_1421,In_642);
and U526 (N_526,In_1014,In_328);
and U527 (N_527,In_1239,In_912);
xnor U528 (N_528,In_1424,In_1369);
or U529 (N_529,In_822,In_371);
or U530 (N_530,In_48,In_1154);
or U531 (N_531,In_1302,In_1097);
and U532 (N_532,In_1080,In_1031);
xor U533 (N_533,In_879,In_1151);
and U534 (N_534,In_983,In_234);
xnor U535 (N_535,In_1280,In_1336);
or U536 (N_536,In_1045,In_690);
and U537 (N_537,In_173,In_1340);
nand U538 (N_538,In_937,In_1119);
and U539 (N_539,In_719,In_295);
xnor U540 (N_540,In_842,In_1470);
and U541 (N_541,In_604,In_612);
and U542 (N_542,In_961,In_1118);
or U543 (N_543,In_352,In_1150);
xor U544 (N_544,In_1443,In_342);
and U545 (N_545,In_22,In_435);
nand U546 (N_546,In_365,In_1148);
xnor U547 (N_547,In_237,In_1067);
nor U548 (N_548,In_581,In_1189);
and U549 (N_549,In_216,In_434);
nand U550 (N_550,In_1480,In_1466);
nor U551 (N_551,In_552,In_916);
nand U552 (N_552,In_203,In_363);
or U553 (N_553,In_1208,In_370);
nor U554 (N_554,In_427,In_452);
and U555 (N_555,In_301,In_949);
or U556 (N_556,In_1054,In_896);
or U557 (N_557,In_644,In_410);
nor U558 (N_558,In_359,In_1235);
and U559 (N_559,In_1126,In_1027);
and U560 (N_560,In_669,In_958);
nand U561 (N_561,In_699,In_259);
or U562 (N_562,In_944,In_637);
nand U563 (N_563,In_1427,In_224);
nor U564 (N_564,In_936,In_862);
or U565 (N_565,In_700,In_34);
nand U566 (N_566,In_1499,In_1295);
and U567 (N_567,In_558,In_197);
nand U568 (N_568,In_675,In_1204);
nor U569 (N_569,In_489,In_676);
and U570 (N_570,In_621,In_1177);
or U571 (N_571,In_461,In_1396);
nand U572 (N_572,In_442,In_1498);
or U573 (N_573,In_1060,In_990);
nor U574 (N_574,In_674,In_686);
xor U575 (N_575,In_979,In_577);
nor U576 (N_576,In_783,In_428);
or U577 (N_577,In_527,In_430);
nand U578 (N_578,In_1079,In_998);
or U579 (N_579,In_943,In_544);
and U580 (N_580,In_524,In_1357);
and U581 (N_581,In_1141,In_308);
and U582 (N_582,In_1316,In_655);
nor U583 (N_583,In_891,In_476);
nand U584 (N_584,In_1224,In_1200);
xor U585 (N_585,In_722,In_88);
nor U586 (N_586,In_1015,In_997);
and U587 (N_587,In_993,In_1447);
and U588 (N_588,In_186,In_1430);
xnor U589 (N_589,In_1122,In_605);
xnor U590 (N_590,In_304,In_1496);
nand U591 (N_591,In_695,In_1296);
nand U592 (N_592,In_766,In_1433);
and U593 (N_593,In_1192,In_740);
nor U594 (N_594,In_866,In_490);
and U595 (N_595,In_1491,In_547);
nor U596 (N_596,In_885,In_1215);
and U597 (N_597,In_1030,In_212);
nand U598 (N_598,In_563,In_64);
and U599 (N_599,In_1379,In_953);
nor U600 (N_600,In_592,In_827);
nor U601 (N_601,In_388,In_1231);
nor U602 (N_602,In_1442,In_464);
nand U603 (N_603,In_1331,In_1113);
xor U604 (N_604,In_59,In_43);
xnor U605 (N_605,In_149,In_1128);
and U606 (N_606,In_178,In_767);
and U607 (N_607,In_831,In_568);
nor U608 (N_608,In_1050,In_924);
nand U609 (N_609,In_616,In_742);
or U610 (N_610,In_580,In_312);
and U611 (N_611,In_773,In_273);
or U612 (N_612,In_209,In_1178);
or U613 (N_613,In_343,In_449);
nand U614 (N_614,In_1403,In_874);
or U615 (N_615,In_244,In_334);
xor U616 (N_616,In_463,In_852);
nand U617 (N_617,In_1370,In_697);
and U618 (N_618,In_373,In_838);
or U619 (N_619,In_1226,In_28);
or U620 (N_620,In_27,In_198);
nor U621 (N_621,In_497,In_1107);
and U622 (N_622,In_511,In_13);
nor U623 (N_623,In_747,In_731);
nand U624 (N_624,In_41,In_1013);
nor U625 (N_625,In_1135,In_256);
and U626 (N_626,In_361,In_240);
nor U627 (N_627,In_525,In_320);
and U628 (N_628,In_582,In_1082);
and U629 (N_629,In_1206,In_1362);
nor U630 (N_630,In_462,In_379);
and U631 (N_631,In_1212,In_1075);
nor U632 (N_632,In_778,In_1363);
nand U633 (N_633,In_1274,In_671);
or U634 (N_634,In_1137,In_146);
or U635 (N_635,In_611,In_1398);
nand U636 (N_636,In_85,In_1320);
nand U637 (N_637,In_74,In_1481);
nand U638 (N_638,In_421,In_1378);
and U639 (N_639,In_440,In_1146);
and U640 (N_640,In_651,In_565);
nand U641 (N_641,In_51,In_255);
or U642 (N_642,In_228,In_1025);
and U643 (N_643,In_1047,In_1372);
nand U644 (N_644,In_965,In_1241);
nor U645 (N_645,In_903,In_1056);
and U646 (N_646,In_1289,In_274);
nand U647 (N_647,In_424,In_522);
and U648 (N_648,In_1008,In_110);
or U649 (N_649,In_941,In_600);
nor U650 (N_650,In_1199,In_732);
or U651 (N_651,In_44,In_135);
and U652 (N_652,In_1386,In_654);
or U653 (N_653,In_166,In_772);
nor U654 (N_654,In_691,In_978);
nor U655 (N_655,In_984,In_1051);
nand U656 (N_656,In_1111,In_384);
or U657 (N_657,In_1270,In_918);
and U658 (N_658,In_1283,In_401);
or U659 (N_659,In_769,In_1252);
or U660 (N_660,In_129,In_542);
or U661 (N_661,In_1095,In_940);
or U662 (N_662,In_1174,In_356);
nand U663 (N_663,In_1441,In_136);
and U664 (N_664,In_1023,In_55);
nand U665 (N_665,In_1311,In_711);
nor U666 (N_666,In_407,In_125);
or U667 (N_667,In_1272,In_648);
and U668 (N_668,In_1053,In_869);
xor U669 (N_669,In_981,In_68);
nor U670 (N_670,In_257,In_1269);
or U671 (N_671,In_1438,In_534);
and U672 (N_672,In_872,In_176);
and U673 (N_673,In_696,In_1382);
and U674 (N_674,In_1003,In_1099);
nor U675 (N_675,In_1004,In_1063);
and U676 (N_676,In_596,In_1467);
nor U677 (N_677,In_1029,In_539);
or U678 (N_678,In_571,In_498);
nand U679 (N_679,In_1203,In_1359);
and U680 (N_680,In_557,In_1093);
or U681 (N_681,In_97,In_187);
and U682 (N_682,In_1066,In_745);
nand U683 (N_683,In_601,In_785);
xor U684 (N_684,In_913,In_153);
and U685 (N_685,In_614,In_289);
xor U686 (N_686,In_155,In_1418);
nand U687 (N_687,In_996,In_728);
nor U688 (N_688,In_1454,In_680);
and U689 (N_689,In_1415,In_1129);
nor U690 (N_690,In_164,In_1401);
and U691 (N_691,In_467,In_929);
and U692 (N_692,In_1180,In_127);
or U693 (N_693,In_807,In_1188);
and U694 (N_694,In_678,In_1287);
or U695 (N_695,In_1416,In_26);
and U696 (N_696,In_62,In_1042);
and U697 (N_697,In_1116,In_111);
nor U698 (N_698,In_1399,In_1160);
xnor U699 (N_699,In_269,In_1170);
nor U700 (N_700,In_514,In_258);
or U701 (N_701,In_599,In_681);
or U702 (N_702,In_491,In_661);
and U703 (N_703,In_264,In_1479);
xnor U704 (N_704,In_1115,In_576);
and U705 (N_705,In_207,In_208);
nand U706 (N_706,In_602,In_730);
or U707 (N_707,In_1338,In_1475);
nor U708 (N_708,In_825,In_115);
nor U709 (N_709,In_1373,In_629);
nand U710 (N_710,In_638,In_1110);
nand U711 (N_711,In_298,In_1404);
and U712 (N_712,In_1333,In_1410);
and U713 (N_713,In_156,In_816);
or U714 (N_714,In_303,In_61);
nor U715 (N_715,In_948,In_713);
nand U716 (N_716,In_1297,In_619);
nor U717 (N_717,In_443,In_585);
nor U718 (N_718,In_1009,In_263);
or U719 (N_719,In_679,In_1048);
nand U720 (N_720,In_1037,In_1450);
and U721 (N_721,In_1348,In_819);
xor U722 (N_722,In_397,In_194);
xnor U723 (N_723,In_991,In_970);
and U724 (N_724,In_899,In_665);
or U725 (N_725,In_1389,In_1168);
nor U726 (N_726,In_575,In_1449);
nor U727 (N_727,In_516,In_817);
or U728 (N_728,In_1307,In_503);
or U729 (N_729,In_761,In_1125);
xnor U730 (N_730,In_573,In_801);
or U731 (N_731,In_191,In_1492);
nor U732 (N_732,In_1312,In_972);
or U733 (N_733,In_167,In_895);
and U734 (N_734,In_1465,In_1486);
or U735 (N_735,In_814,In_433);
nand U736 (N_736,In_92,In_144);
nor U737 (N_737,In_980,In_889);
and U738 (N_738,In_93,In_784);
nand U739 (N_739,In_458,In_1102);
or U740 (N_740,In_964,In_78);
and U741 (N_741,In_1412,In_854);
nor U742 (N_742,In_927,In_183);
nand U743 (N_743,In_559,In_291);
nand U744 (N_744,In_1086,In_1395);
nor U745 (N_745,In_595,In_456);
and U746 (N_746,In_1071,In_928);
and U747 (N_747,In_46,In_271);
and U748 (N_748,In_161,In_1161);
nand U749 (N_749,In_1040,In_1400);
and U750 (N_750,In_1358,In_884);
or U751 (N_751,In_1456,In_786);
and U752 (N_752,In_280,In_1291);
or U753 (N_753,In_387,In_20);
or U754 (N_754,In_285,In_1393);
nand U755 (N_755,In_18,In_990);
nor U756 (N_756,In_677,In_1427);
nand U757 (N_757,In_926,In_51);
and U758 (N_758,In_803,In_295);
xor U759 (N_759,In_33,In_1408);
nand U760 (N_760,In_656,In_732);
and U761 (N_761,In_1471,In_121);
xnor U762 (N_762,In_663,In_1209);
or U763 (N_763,In_718,In_474);
nand U764 (N_764,In_1350,In_1295);
nor U765 (N_765,In_466,In_1255);
nand U766 (N_766,In_1257,In_1095);
nor U767 (N_767,In_99,In_249);
or U768 (N_768,In_16,In_607);
nor U769 (N_769,In_1029,In_387);
xnor U770 (N_770,In_944,In_27);
nor U771 (N_771,In_948,In_628);
nor U772 (N_772,In_1384,In_930);
nand U773 (N_773,In_1284,In_330);
or U774 (N_774,In_655,In_1411);
or U775 (N_775,In_154,In_162);
nand U776 (N_776,In_1267,In_111);
xnor U777 (N_777,In_94,In_449);
and U778 (N_778,In_45,In_52);
or U779 (N_779,In_132,In_136);
nor U780 (N_780,In_824,In_219);
or U781 (N_781,In_750,In_826);
nand U782 (N_782,In_931,In_1272);
or U783 (N_783,In_1221,In_202);
nand U784 (N_784,In_680,In_734);
nand U785 (N_785,In_1357,In_783);
nand U786 (N_786,In_571,In_425);
and U787 (N_787,In_1450,In_426);
nor U788 (N_788,In_368,In_1450);
or U789 (N_789,In_1405,In_34);
nand U790 (N_790,In_670,In_1446);
xnor U791 (N_791,In_759,In_767);
and U792 (N_792,In_1422,In_1427);
nor U793 (N_793,In_1299,In_1032);
and U794 (N_794,In_953,In_1036);
nand U795 (N_795,In_957,In_844);
nor U796 (N_796,In_45,In_165);
or U797 (N_797,In_292,In_732);
xor U798 (N_798,In_1207,In_149);
and U799 (N_799,In_768,In_583);
and U800 (N_800,In_348,In_371);
and U801 (N_801,In_211,In_914);
or U802 (N_802,In_294,In_995);
and U803 (N_803,In_932,In_1125);
xor U804 (N_804,In_1030,In_1332);
or U805 (N_805,In_949,In_145);
nor U806 (N_806,In_489,In_492);
xnor U807 (N_807,In_819,In_1021);
and U808 (N_808,In_423,In_1158);
and U809 (N_809,In_401,In_104);
nor U810 (N_810,In_90,In_257);
and U811 (N_811,In_1369,In_1147);
nor U812 (N_812,In_224,In_660);
nand U813 (N_813,In_1481,In_1497);
nand U814 (N_814,In_1188,In_936);
or U815 (N_815,In_780,In_850);
nor U816 (N_816,In_1445,In_23);
and U817 (N_817,In_1448,In_1389);
and U818 (N_818,In_1481,In_766);
nor U819 (N_819,In_283,In_10);
xnor U820 (N_820,In_670,In_46);
or U821 (N_821,In_236,In_235);
nor U822 (N_822,In_1284,In_1371);
nand U823 (N_823,In_584,In_726);
nand U824 (N_824,In_1266,In_355);
nand U825 (N_825,In_1107,In_41);
or U826 (N_826,In_67,In_258);
nand U827 (N_827,In_828,In_113);
or U828 (N_828,In_491,In_354);
or U829 (N_829,In_566,In_406);
nor U830 (N_830,In_177,In_1086);
or U831 (N_831,In_897,In_1301);
or U832 (N_832,In_43,In_354);
nand U833 (N_833,In_697,In_380);
nor U834 (N_834,In_1319,In_174);
nand U835 (N_835,In_1163,In_279);
and U836 (N_836,In_627,In_1388);
or U837 (N_837,In_992,In_1049);
nand U838 (N_838,In_1006,In_617);
or U839 (N_839,In_310,In_1449);
nand U840 (N_840,In_734,In_1143);
xnor U841 (N_841,In_335,In_891);
and U842 (N_842,In_1393,In_923);
nand U843 (N_843,In_1444,In_461);
and U844 (N_844,In_804,In_1413);
or U845 (N_845,In_1190,In_249);
xnor U846 (N_846,In_619,In_674);
and U847 (N_847,In_396,In_1215);
nand U848 (N_848,In_357,In_1417);
xor U849 (N_849,In_1225,In_815);
or U850 (N_850,In_1456,In_484);
nor U851 (N_851,In_462,In_470);
nor U852 (N_852,In_914,In_140);
nand U853 (N_853,In_606,In_711);
nor U854 (N_854,In_339,In_643);
nor U855 (N_855,In_834,In_401);
nand U856 (N_856,In_246,In_237);
xnor U857 (N_857,In_1240,In_377);
nor U858 (N_858,In_736,In_641);
or U859 (N_859,In_1498,In_345);
and U860 (N_860,In_1055,In_1299);
or U861 (N_861,In_1343,In_552);
and U862 (N_862,In_806,In_677);
nand U863 (N_863,In_869,In_416);
or U864 (N_864,In_963,In_736);
xor U865 (N_865,In_1194,In_199);
or U866 (N_866,In_1132,In_1301);
or U867 (N_867,In_1057,In_519);
and U868 (N_868,In_651,In_637);
nand U869 (N_869,In_1048,In_756);
and U870 (N_870,In_987,In_86);
nand U871 (N_871,In_472,In_870);
and U872 (N_872,In_767,In_1370);
xor U873 (N_873,In_156,In_1239);
nor U874 (N_874,In_78,In_1213);
xnor U875 (N_875,In_926,In_678);
or U876 (N_876,In_374,In_363);
nor U877 (N_877,In_1400,In_442);
nand U878 (N_878,In_1496,In_796);
nor U879 (N_879,In_610,In_11);
or U880 (N_880,In_101,In_1288);
nor U881 (N_881,In_1227,In_172);
nand U882 (N_882,In_1238,In_1017);
or U883 (N_883,In_584,In_1048);
xnor U884 (N_884,In_624,In_676);
nor U885 (N_885,In_361,In_1385);
and U886 (N_886,In_1496,In_42);
and U887 (N_887,In_1378,In_1211);
and U888 (N_888,In_1045,In_1103);
nand U889 (N_889,In_1462,In_319);
and U890 (N_890,In_895,In_1153);
or U891 (N_891,In_265,In_1092);
or U892 (N_892,In_1133,In_1407);
nor U893 (N_893,In_574,In_89);
and U894 (N_894,In_639,In_267);
nor U895 (N_895,In_1383,In_90);
nor U896 (N_896,In_671,In_807);
nor U897 (N_897,In_1306,In_1193);
or U898 (N_898,In_1232,In_1083);
or U899 (N_899,In_1266,In_922);
and U900 (N_900,In_871,In_417);
xor U901 (N_901,In_602,In_1290);
xnor U902 (N_902,In_1008,In_119);
nand U903 (N_903,In_1197,In_890);
or U904 (N_904,In_281,In_777);
nand U905 (N_905,In_221,In_956);
nand U906 (N_906,In_1052,In_1492);
nor U907 (N_907,In_939,In_1007);
nor U908 (N_908,In_890,In_818);
or U909 (N_909,In_883,In_92);
nor U910 (N_910,In_1312,In_1417);
nand U911 (N_911,In_490,In_143);
nand U912 (N_912,In_975,In_1122);
nor U913 (N_913,In_289,In_1001);
xnor U914 (N_914,In_690,In_281);
and U915 (N_915,In_342,In_373);
xor U916 (N_916,In_977,In_1226);
and U917 (N_917,In_578,In_919);
nand U918 (N_918,In_1468,In_717);
or U919 (N_919,In_158,In_52);
nor U920 (N_920,In_677,In_253);
nand U921 (N_921,In_1284,In_12);
xnor U922 (N_922,In_1449,In_694);
and U923 (N_923,In_755,In_1115);
nand U924 (N_924,In_871,In_1406);
and U925 (N_925,In_802,In_777);
or U926 (N_926,In_937,In_696);
and U927 (N_927,In_1418,In_825);
or U928 (N_928,In_760,In_659);
xor U929 (N_929,In_167,In_84);
and U930 (N_930,In_976,In_98);
nor U931 (N_931,In_674,In_59);
or U932 (N_932,In_500,In_513);
or U933 (N_933,In_644,In_721);
or U934 (N_934,In_1399,In_742);
and U935 (N_935,In_1336,In_143);
and U936 (N_936,In_1478,In_955);
or U937 (N_937,In_1201,In_753);
and U938 (N_938,In_19,In_763);
and U939 (N_939,In_924,In_580);
or U940 (N_940,In_276,In_1183);
or U941 (N_941,In_894,In_1351);
and U942 (N_942,In_582,In_504);
nor U943 (N_943,In_1275,In_419);
or U944 (N_944,In_664,In_969);
and U945 (N_945,In_1033,In_421);
or U946 (N_946,In_186,In_1237);
xnor U947 (N_947,In_587,In_594);
and U948 (N_948,In_1374,In_1100);
or U949 (N_949,In_1057,In_1001);
nor U950 (N_950,In_1180,In_1348);
or U951 (N_951,In_1216,In_612);
nor U952 (N_952,In_225,In_1110);
and U953 (N_953,In_99,In_375);
nor U954 (N_954,In_1110,In_319);
nand U955 (N_955,In_296,In_1398);
nor U956 (N_956,In_1429,In_527);
nand U957 (N_957,In_995,In_829);
and U958 (N_958,In_315,In_669);
nor U959 (N_959,In_491,In_1317);
and U960 (N_960,In_1425,In_980);
or U961 (N_961,In_1038,In_1386);
nor U962 (N_962,In_222,In_255);
and U963 (N_963,In_966,In_431);
or U964 (N_964,In_998,In_400);
nand U965 (N_965,In_812,In_593);
nor U966 (N_966,In_995,In_787);
or U967 (N_967,In_544,In_1370);
or U968 (N_968,In_1347,In_581);
and U969 (N_969,In_736,In_1174);
nor U970 (N_970,In_180,In_418);
nand U971 (N_971,In_1048,In_712);
nand U972 (N_972,In_66,In_1259);
nand U973 (N_973,In_1280,In_469);
or U974 (N_974,In_478,In_464);
nor U975 (N_975,In_71,In_189);
and U976 (N_976,In_891,In_636);
nand U977 (N_977,In_1104,In_458);
and U978 (N_978,In_225,In_304);
nor U979 (N_979,In_1181,In_343);
or U980 (N_980,In_982,In_378);
or U981 (N_981,In_322,In_227);
nor U982 (N_982,In_70,In_915);
and U983 (N_983,In_307,In_732);
and U984 (N_984,In_715,In_455);
and U985 (N_985,In_369,In_516);
nand U986 (N_986,In_1311,In_763);
xnor U987 (N_987,In_244,In_510);
xor U988 (N_988,In_804,In_90);
xnor U989 (N_989,In_635,In_1224);
and U990 (N_990,In_77,In_875);
nor U991 (N_991,In_1025,In_498);
nand U992 (N_992,In_1022,In_377);
and U993 (N_993,In_1491,In_10);
and U994 (N_994,In_402,In_736);
or U995 (N_995,In_197,In_884);
nor U996 (N_996,In_1155,In_1030);
nand U997 (N_997,In_455,In_510);
and U998 (N_998,In_1483,In_425);
or U999 (N_999,In_430,In_1299);
and U1000 (N_1000,In_754,In_251);
nor U1001 (N_1001,In_500,In_1320);
nand U1002 (N_1002,In_531,In_839);
and U1003 (N_1003,In_1303,In_99);
nand U1004 (N_1004,In_82,In_393);
and U1005 (N_1005,In_1277,In_836);
nor U1006 (N_1006,In_151,In_340);
or U1007 (N_1007,In_922,In_974);
nor U1008 (N_1008,In_1388,In_131);
or U1009 (N_1009,In_420,In_1379);
xnor U1010 (N_1010,In_1159,In_226);
xnor U1011 (N_1011,In_395,In_434);
nand U1012 (N_1012,In_1489,In_408);
or U1013 (N_1013,In_983,In_325);
or U1014 (N_1014,In_791,In_1080);
or U1015 (N_1015,In_1081,In_780);
nor U1016 (N_1016,In_1245,In_1025);
nor U1017 (N_1017,In_552,In_682);
nor U1018 (N_1018,In_813,In_1215);
and U1019 (N_1019,In_1084,In_769);
or U1020 (N_1020,In_906,In_860);
nor U1021 (N_1021,In_106,In_417);
and U1022 (N_1022,In_610,In_314);
and U1023 (N_1023,In_1492,In_583);
nor U1024 (N_1024,In_1274,In_439);
or U1025 (N_1025,In_744,In_823);
xnor U1026 (N_1026,In_1119,In_240);
or U1027 (N_1027,In_1239,In_1250);
xor U1028 (N_1028,In_225,In_606);
nand U1029 (N_1029,In_998,In_1155);
and U1030 (N_1030,In_792,In_1096);
nand U1031 (N_1031,In_783,In_884);
and U1032 (N_1032,In_1164,In_1224);
nor U1033 (N_1033,In_39,In_1397);
or U1034 (N_1034,In_464,In_1130);
nor U1035 (N_1035,In_178,In_458);
nor U1036 (N_1036,In_1295,In_615);
nor U1037 (N_1037,In_446,In_1435);
and U1038 (N_1038,In_1305,In_304);
nand U1039 (N_1039,In_28,In_1452);
or U1040 (N_1040,In_243,In_762);
nand U1041 (N_1041,In_1322,In_377);
or U1042 (N_1042,In_1049,In_1470);
nor U1043 (N_1043,In_79,In_536);
xor U1044 (N_1044,In_804,In_483);
and U1045 (N_1045,In_1006,In_117);
xnor U1046 (N_1046,In_144,In_455);
or U1047 (N_1047,In_520,In_232);
or U1048 (N_1048,In_703,In_332);
nor U1049 (N_1049,In_533,In_1081);
nor U1050 (N_1050,In_702,In_371);
nand U1051 (N_1051,In_1279,In_344);
xnor U1052 (N_1052,In_459,In_141);
nand U1053 (N_1053,In_1201,In_871);
or U1054 (N_1054,In_168,In_1484);
or U1055 (N_1055,In_207,In_348);
or U1056 (N_1056,In_1451,In_636);
and U1057 (N_1057,In_371,In_215);
nand U1058 (N_1058,In_1271,In_1415);
or U1059 (N_1059,In_1102,In_150);
or U1060 (N_1060,In_1183,In_195);
nand U1061 (N_1061,In_815,In_943);
nand U1062 (N_1062,In_524,In_1234);
xnor U1063 (N_1063,In_356,In_803);
nand U1064 (N_1064,In_634,In_1491);
and U1065 (N_1065,In_112,In_841);
nand U1066 (N_1066,In_1075,In_1177);
nor U1067 (N_1067,In_702,In_925);
xor U1068 (N_1068,In_750,In_127);
or U1069 (N_1069,In_220,In_152);
nand U1070 (N_1070,In_1409,In_107);
nand U1071 (N_1071,In_1407,In_274);
nand U1072 (N_1072,In_1059,In_470);
and U1073 (N_1073,In_1067,In_1317);
or U1074 (N_1074,In_392,In_221);
nand U1075 (N_1075,In_1314,In_429);
or U1076 (N_1076,In_115,In_694);
nor U1077 (N_1077,In_371,In_114);
nand U1078 (N_1078,In_314,In_446);
and U1079 (N_1079,In_1475,In_699);
nand U1080 (N_1080,In_1041,In_1295);
nor U1081 (N_1081,In_183,In_312);
or U1082 (N_1082,In_393,In_1060);
or U1083 (N_1083,In_495,In_523);
or U1084 (N_1084,In_1243,In_1497);
or U1085 (N_1085,In_1334,In_712);
nor U1086 (N_1086,In_856,In_154);
nand U1087 (N_1087,In_236,In_1386);
xor U1088 (N_1088,In_897,In_463);
xnor U1089 (N_1089,In_1411,In_911);
and U1090 (N_1090,In_1190,In_744);
xor U1091 (N_1091,In_1315,In_728);
or U1092 (N_1092,In_860,In_793);
and U1093 (N_1093,In_1440,In_895);
nand U1094 (N_1094,In_1051,In_343);
or U1095 (N_1095,In_122,In_80);
and U1096 (N_1096,In_1109,In_1011);
or U1097 (N_1097,In_1211,In_937);
or U1098 (N_1098,In_748,In_1323);
and U1099 (N_1099,In_554,In_1463);
or U1100 (N_1100,In_891,In_617);
and U1101 (N_1101,In_183,In_900);
nor U1102 (N_1102,In_857,In_1047);
nand U1103 (N_1103,In_893,In_927);
and U1104 (N_1104,In_1198,In_641);
nand U1105 (N_1105,In_650,In_173);
or U1106 (N_1106,In_1172,In_888);
nand U1107 (N_1107,In_5,In_1154);
xnor U1108 (N_1108,In_1428,In_494);
nor U1109 (N_1109,In_744,In_1452);
nand U1110 (N_1110,In_1432,In_1372);
or U1111 (N_1111,In_128,In_1112);
xnor U1112 (N_1112,In_1288,In_180);
nand U1113 (N_1113,In_23,In_107);
nor U1114 (N_1114,In_1103,In_990);
or U1115 (N_1115,In_535,In_295);
or U1116 (N_1116,In_398,In_156);
nor U1117 (N_1117,In_917,In_36);
xnor U1118 (N_1118,In_157,In_182);
nand U1119 (N_1119,In_332,In_1295);
nand U1120 (N_1120,In_598,In_555);
and U1121 (N_1121,In_1341,In_178);
and U1122 (N_1122,In_318,In_561);
and U1123 (N_1123,In_938,In_698);
and U1124 (N_1124,In_1139,In_1091);
xor U1125 (N_1125,In_83,In_1262);
nor U1126 (N_1126,In_850,In_981);
or U1127 (N_1127,In_184,In_869);
nand U1128 (N_1128,In_1378,In_411);
nor U1129 (N_1129,In_919,In_949);
nand U1130 (N_1130,In_1409,In_857);
or U1131 (N_1131,In_1197,In_1173);
and U1132 (N_1132,In_107,In_781);
or U1133 (N_1133,In_370,In_309);
nor U1134 (N_1134,In_67,In_926);
and U1135 (N_1135,In_31,In_556);
or U1136 (N_1136,In_1201,In_596);
and U1137 (N_1137,In_956,In_972);
and U1138 (N_1138,In_1108,In_1149);
or U1139 (N_1139,In_277,In_428);
or U1140 (N_1140,In_84,In_1032);
or U1141 (N_1141,In_753,In_804);
or U1142 (N_1142,In_244,In_1234);
and U1143 (N_1143,In_877,In_1167);
and U1144 (N_1144,In_1477,In_158);
nand U1145 (N_1145,In_1179,In_1201);
or U1146 (N_1146,In_772,In_787);
nor U1147 (N_1147,In_612,In_566);
nand U1148 (N_1148,In_760,In_533);
and U1149 (N_1149,In_704,In_98);
or U1150 (N_1150,In_496,In_932);
and U1151 (N_1151,In_294,In_879);
or U1152 (N_1152,In_1180,In_679);
nand U1153 (N_1153,In_1098,In_837);
nand U1154 (N_1154,In_22,In_1013);
nand U1155 (N_1155,In_873,In_609);
nor U1156 (N_1156,In_635,In_274);
nand U1157 (N_1157,In_1131,In_244);
or U1158 (N_1158,In_79,In_74);
or U1159 (N_1159,In_1479,In_1387);
nor U1160 (N_1160,In_144,In_1034);
nand U1161 (N_1161,In_523,In_633);
or U1162 (N_1162,In_566,In_1363);
or U1163 (N_1163,In_1320,In_688);
nor U1164 (N_1164,In_709,In_1011);
xnor U1165 (N_1165,In_1450,In_602);
nor U1166 (N_1166,In_1034,In_1307);
nor U1167 (N_1167,In_836,In_671);
or U1168 (N_1168,In_152,In_652);
and U1169 (N_1169,In_47,In_638);
nor U1170 (N_1170,In_1259,In_1330);
nor U1171 (N_1171,In_605,In_929);
xnor U1172 (N_1172,In_1159,In_672);
and U1173 (N_1173,In_862,In_607);
nand U1174 (N_1174,In_117,In_497);
and U1175 (N_1175,In_172,In_419);
nor U1176 (N_1176,In_305,In_96);
nand U1177 (N_1177,In_585,In_1262);
and U1178 (N_1178,In_714,In_133);
or U1179 (N_1179,In_890,In_1450);
nor U1180 (N_1180,In_601,In_1455);
and U1181 (N_1181,In_847,In_1150);
nand U1182 (N_1182,In_1043,In_0);
or U1183 (N_1183,In_607,In_1250);
or U1184 (N_1184,In_1445,In_1418);
nor U1185 (N_1185,In_410,In_440);
nor U1186 (N_1186,In_10,In_1390);
and U1187 (N_1187,In_515,In_935);
or U1188 (N_1188,In_367,In_1216);
and U1189 (N_1189,In_1409,In_78);
nand U1190 (N_1190,In_1237,In_4);
and U1191 (N_1191,In_1082,In_145);
nand U1192 (N_1192,In_293,In_377);
and U1193 (N_1193,In_149,In_926);
xor U1194 (N_1194,In_424,In_83);
or U1195 (N_1195,In_554,In_1452);
xor U1196 (N_1196,In_660,In_739);
nor U1197 (N_1197,In_251,In_316);
nor U1198 (N_1198,In_1019,In_612);
nand U1199 (N_1199,In_886,In_1434);
nor U1200 (N_1200,In_1380,In_635);
or U1201 (N_1201,In_1241,In_312);
and U1202 (N_1202,In_1075,In_307);
nor U1203 (N_1203,In_590,In_1155);
nor U1204 (N_1204,In_208,In_715);
or U1205 (N_1205,In_1135,In_1154);
and U1206 (N_1206,In_1461,In_67);
nor U1207 (N_1207,In_648,In_1103);
nor U1208 (N_1208,In_857,In_152);
and U1209 (N_1209,In_667,In_625);
xor U1210 (N_1210,In_1253,In_329);
nor U1211 (N_1211,In_1496,In_1331);
and U1212 (N_1212,In_819,In_49);
and U1213 (N_1213,In_781,In_469);
or U1214 (N_1214,In_276,In_1264);
nor U1215 (N_1215,In_169,In_652);
nor U1216 (N_1216,In_217,In_604);
nor U1217 (N_1217,In_975,In_854);
or U1218 (N_1218,In_157,In_1215);
and U1219 (N_1219,In_1266,In_1054);
xnor U1220 (N_1220,In_1226,In_618);
or U1221 (N_1221,In_844,In_1024);
or U1222 (N_1222,In_756,In_1395);
nand U1223 (N_1223,In_1230,In_977);
and U1224 (N_1224,In_1307,In_431);
nor U1225 (N_1225,In_284,In_1042);
nand U1226 (N_1226,In_46,In_1450);
nor U1227 (N_1227,In_1372,In_485);
or U1228 (N_1228,In_782,In_1205);
nand U1229 (N_1229,In_1148,In_781);
or U1230 (N_1230,In_943,In_1368);
xor U1231 (N_1231,In_237,In_295);
nand U1232 (N_1232,In_905,In_1339);
nor U1233 (N_1233,In_387,In_573);
nor U1234 (N_1234,In_48,In_246);
nor U1235 (N_1235,In_1017,In_762);
or U1236 (N_1236,In_863,In_1220);
or U1237 (N_1237,In_1309,In_623);
and U1238 (N_1238,In_512,In_881);
or U1239 (N_1239,In_455,In_493);
nor U1240 (N_1240,In_1206,In_301);
nor U1241 (N_1241,In_62,In_499);
and U1242 (N_1242,In_223,In_701);
nand U1243 (N_1243,In_45,In_216);
nor U1244 (N_1244,In_766,In_1424);
and U1245 (N_1245,In_1036,In_358);
and U1246 (N_1246,In_554,In_706);
nor U1247 (N_1247,In_846,In_1089);
nor U1248 (N_1248,In_360,In_1145);
nand U1249 (N_1249,In_475,In_1052);
nor U1250 (N_1250,In_437,In_587);
nor U1251 (N_1251,In_992,In_816);
and U1252 (N_1252,In_1089,In_470);
and U1253 (N_1253,In_104,In_820);
and U1254 (N_1254,In_570,In_1313);
nand U1255 (N_1255,In_620,In_52);
nand U1256 (N_1256,In_876,In_203);
nor U1257 (N_1257,In_1194,In_752);
nor U1258 (N_1258,In_515,In_96);
nor U1259 (N_1259,In_817,In_813);
xnor U1260 (N_1260,In_1414,In_443);
and U1261 (N_1261,In_149,In_1083);
nor U1262 (N_1262,In_171,In_864);
or U1263 (N_1263,In_1261,In_1221);
and U1264 (N_1264,In_278,In_1040);
and U1265 (N_1265,In_16,In_409);
or U1266 (N_1266,In_40,In_272);
nand U1267 (N_1267,In_214,In_942);
or U1268 (N_1268,In_20,In_1460);
or U1269 (N_1269,In_779,In_856);
and U1270 (N_1270,In_710,In_299);
nand U1271 (N_1271,In_409,In_1091);
nor U1272 (N_1272,In_151,In_134);
and U1273 (N_1273,In_838,In_826);
or U1274 (N_1274,In_986,In_469);
nand U1275 (N_1275,In_1482,In_799);
and U1276 (N_1276,In_772,In_815);
nand U1277 (N_1277,In_209,In_687);
or U1278 (N_1278,In_1499,In_108);
xnor U1279 (N_1279,In_743,In_286);
nand U1280 (N_1280,In_107,In_1317);
and U1281 (N_1281,In_1030,In_622);
and U1282 (N_1282,In_467,In_63);
and U1283 (N_1283,In_1154,In_918);
or U1284 (N_1284,In_1280,In_1096);
nor U1285 (N_1285,In_1182,In_1210);
nand U1286 (N_1286,In_1307,In_1065);
nand U1287 (N_1287,In_236,In_222);
nor U1288 (N_1288,In_216,In_1041);
and U1289 (N_1289,In_525,In_701);
or U1290 (N_1290,In_1449,In_753);
and U1291 (N_1291,In_0,In_531);
nand U1292 (N_1292,In_1145,In_1021);
and U1293 (N_1293,In_347,In_304);
or U1294 (N_1294,In_118,In_1132);
nor U1295 (N_1295,In_1463,In_843);
or U1296 (N_1296,In_348,In_550);
xor U1297 (N_1297,In_1126,In_1108);
and U1298 (N_1298,In_321,In_1347);
and U1299 (N_1299,In_557,In_1353);
and U1300 (N_1300,In_467,In_722);
nand U1301 (N_1301,In_165,In_413);
and U1302 (N_1302,In_425,In_317);
or U1303 (N_1303,In_361,In_595);
nor U1304 (N_1304,In_241,In_910);
and U1305 (N_1305,In_201,In_287);
or U1306 (N_1306,In_358,In_294);
or U1307 (N_1307,In_888,In_321);
nor U1308 (N_1308,In_1252,In_915);
or U1309 (N_1309,In_351,In_1359);
or U1310 (N_1310,In_1253,In_197);
nand U1311 (N_1311,In_934,In_530);
and U1312 (N_1312,In_353,In_40);
nor U1313 (N_1313,In_610,In_1269);
or U1314 (N_1314,In_585,In_796);
or U1315 (N_1315,In_1124,In_465);
xnor U1316 (N_1316,In_540,In_370);
xnor U1317 (N_1317,In_810,In_1034);
nand U1318 (N_1318,In_320,In_40);
nor U1319 (N_1319,In_1469,In_520);
and U1320 (N_1320,In_1392,In_125);
and U1321 (N_1321,In_1110,In_1186);
nand U1322 (N_1322,In_672,In_970);
nor U1323 (N_1323,In_64,In_861);
nor U1324 (N_1324,In_1294,In_241);
and U1325 (N_1325,In_1131,In_77);
nand U1326 (N_1326,In_810,In_846);
nor U1327 (N_1327,In_1235,In_1421);
nand U1328 (N_1328,In_237,In_32);
and U1329 (N_1329,In_457,In_744);
or U1330 (N_1330,In_649,In_703);
xor U1331 (N_1331,In_517,In_816);
and U1332 (N_1332,In_572,In_725);
or U1333 (N_1333,In_522,In_945);
or U1334 (N_1334,In_1303,In_279);
nand U1335 (N_1335,In_635,In_333);
or U1336 (N_1336,In_1173,In_166);
and U1337 (N_1337,In_778,In_1178);
nand U1338 (N_1338,In_636,In_118);
nand U1339 (N_1339,In_962,In_494);
nand U1340 (N_1340,In_587,In_1424);
and U1341 (N_1341,In_594,In_967);
and U1342 (N_1342,In_70,In_696);
nor U1343 (N_1343,In_443,In_1009);
xor U1344 (N_1344,In_370,In_400);
nor U1345 (N_1345,In_842,In_764);
and U1346 (N_1346,In_319,In_971);
or U1347 (N_1347,In_104,In_860);
nor U1348 (N_1348,In_344,In_782);
or U1349 (N_1349,In_184,In_671);
xnor U1350 (N_1350,In_1009,In_194);
or U1351 (N_1351,In_401,In_763);
and U1352 (N_1352,In_1434,In_494);
and U1353 (N_1353,In_466,In_881);
xnor U1354 (N_1354,In_1018,In_1468);
nand U1355 (N_1355,In_158,In_1257);
nor U1356 (N_1356,In_1397,In_638);
nand U1357 (N_1357,In_842,In_1339);
nand U1358 (N_1358,In_550,In_599);
and U1359 (N_1359,In_785,In_857);
nand U1360 (N_1360,In_1258,In_847);
and U1361 (N_1361,In_1378,In_860);
xnor U1362 (N_1362,In_406,In_763);
and U1363 (N_1363,In_1080,In_334);
or U1364 (N_1364,In_1417,In_1405);
or U1365 (N_1365,In_745,In_1452);
or U1366 (N_1366,In_144,In_245);
and U1367 (N_1367,In_1391,In_958);
nand U1368 (N_1368,In_284,In_908);
nor U1369 (N_1369,In_3,In_45);
or U1370 (N_1370,In_209,In_325);
nand U1371 (N_1371,In_31,In_1129);
nand U1372 (N_1372,In_1299,In_1382);
nand U1373 (N_1373,In_1204,In_1094);
xnor U1374 (N_1374,In_898,In_1261);
nor U1375 (N_1375,In_1119,In_335);
and U1376 (N_1376,In_242,In_821);
and U1377 (N_1377,In_1306,In_1276);
or U1378 (N_1378,In_1403,In_345);
nor U1379 (N_1379,In_883,In_856);
nand U1380 (N_1380,In_1232,In_1272);
nor U1381 (N_1381,In_592,In_838);
xor U1382 (N_1382,In_203,In_334);
nor U1383 (N_1383,In_433,In_200);
xnor U1384 (N_1384,In_1147,In_547);
and U1385 (N_1385,In_118,In_691);
nand U1386 (N_1386,In_26,In_449);
or U1387 (N_1387,In_574,In_860);
nand U1388 (N_1388,In_914,In_5);
and U1389 (N_1389,In_1212,In_1286);
xnor U1390 (N_1390,In_73,In_494);
nand U1391 (N_1391,In_1342,In_1382);
nand U1392 (N_1392,In_1284,In_1253);
nor U1393 (N_1393,In_860,In_1254);
xor U1394 (N_1394,In_531,In_40);
or U1395 (N_1395,In_1211,In_408);
nor U1396 (N_1396,In_1276,In_882);
nor U1397 (N_1397,In_1466,In_273);
nand U1398 (N_1398,In_777,In_260);
and U1399 (N_1399,In_929,In_1390);
or U1400 (N_1400,In_1427,In_11);
or U1401 (N_1401,In_640,In_227);
and U1402 (N_1402,In_465,In_676);
nand U1403 (N_1403,In_874,In_528);
nor U1404 (N_1404,In_1003,In_1155);
nor U1405 (N_1405,In_488,In_629);
nand U1406 (N_1406,In_747,In_537);
nand U1407 (N_1407,In_1220,In_26);
or U1408 (N_1408,In_1466,In_1157);
or U1409 (N_1409,In_523,In_453);
nor U1410 (N_1410,In_286,In_914);
and U1411 (N_1411,In_1325,In_1483);
and U1412 (N_1412,In_1318,In_368);
xnor U1413 (N_1413,In_1215,In_235);
nand U1414 (N_1414,In_1199,In_1399);
or U1415 (N_1415,In_610,In_494);
nor U1416 (N_1416,In_864,In_496);
or U1417 (N_1417,In_275,In_912);
nor U1418 (N_1418,In_528,In_747);
nor U1419 (N_1419,In_243,In_611);
and U1420 (N_1420,In_873,In_355);
and U1421 (N_1421,In_1387,In_1495);
nor U1422 (N_1422,In_230,In_291);
nand U1423 (N_1423,In_816,In_789);
or U1424 (N_1424,In_209,In_1240);
xnor U1425 (N_1425,In_897,In_1222);
and U1426 (N_1426,In_1496,In_415);
or U1427 (N_1427,In_725,In_1201);
xor U1428 (N_1428,In_840,In_838);
and U1429 (N_1429,In_302,In_166);
or U1430 (N_1430,In_684,In_972);
nand U1431 (N_1431,In_639,In_1303);
nor U1432 (N_1432,In_1203,In_422);
nor U1433 (N_1433,In_389,In_272);
or U1434 (N_1434,In_218,In_486);
or U1435 (N_1435,In_387,In_1303);
nand U1436 (N_1436,In_1493,In_1288);
nand U1437 (N_1437,In_842,In_234);
or U1438 (N_1438,In_1287,In_1068);
nand U1439 (N_1439,In_1458,In_1017);
and U1440 (N_1440,In_1099,In_188);
and U1441 (N_1441,In_878,In_1140);
nor U1442 (N_1442,In_757,In_355);
xnor U1443 (N_1443,In_1290,In_30);
or U1444 (N_1444,In_1176,In_184);
or U1445 (N_1445,In_244,In_1017);
and U1446 (N_1446,In_157,In_1150);
nand U1447 (N_1447,In_850,In_168);
nor U1448 (N_1448,In_507,In_436);
and U1449 (N_1449,In_1248,In_514);
nand U1450 (N_1450,In_812,In_627);
nand U1451 (N_1451,In_1184,In_683);
or U1452 (N_1452,In_1449,In_1062);
nand U1453 (N_1453,In_1400,In_296);
nor U1454 (N_1454,In_1056,In_842);
nand U1455 (N_1455,In_1387,In_1164);
nor U1456 (N_1456,In_222,In_1103);
nor U1457 (N_1457,In_683,In_233);
or U1458 (N_1458,In_1388,In_274);
nor U1459 (N_1459,In_1332,In_1247);
or U1460 (N_1460,In_44,In_1438);
nand U1461 (N_1461,In_909,In_1244);
xor U1462 (N_1462,In_1027,In_56);
nor U1463 (N_1463,In_210,In_1493);
nor U1464 (N_1464,In_1213,In_572);
and U1465 (N_1465,In_146,In_947);
or U1466 (N_1466,In_1386,In_1227);
nand U1467 (N_1467,In_589,In_822);
nor U1468 (N_1468,In_412,In_997);
and U1469 (N_1469,In_693,In_343);
nand U1470 (N_1470,In_1084,In_667);
nor U1471 (N_1471,In_796,In_676);
nand U1472 (N_1472,In_204,In_1014);
and U1473 (N_1473,In_1287,In_66);
and U1474 (N_1474,In_1245,In_161);
and U1475 (N_1475,In_616,In_1329);
nand U1476 (N_1476,In_421,In_782);
nor U1477 (N_1477,In_262,In_655);
xor U1478 (N_1478,In_226,In_34);
nor U1479 (N_1479,In_946,In_795);
or U1480 (N_1480,In_1030,In_26);
and U1481 (N_1481,In_1339,In_771);
or U1482 (N_1482,In_1302,In_966);
or U1483 (N_1483,In_915,In_238);
nand U1484 (N_1484,In_926,In_786);
nand U1485 (N_1485,In_751,In_1241);
nand U1486 (N_1486,In_1092,In_1283);
and U1487 (N_1487,In_1038,In_1207);
or U1488 (N_1488,In_282,In_981);
or U1489 (N_1489,In_423,In_743);
nand U1490 (N_1490,In_274,In_456);
nor U1491 (N_1491,In_988,In_261);
nor U1492 (N_1492,In_1074,In_206);
and U1493 (N_1493,In_239,In_1129);
and U1494 (N_1494,In_1457,In_844);
nand U1495 (N_1495,In_1431,In_619);
and U1496 (N_1496,In_1397,In_239);
and U1497 (N_1497,In_416,In_1064);
and U1498 (N_1498,In_858,In_1141);
xor U1499 (N_1499,In_1441,In_1298);
or U1500 (N_1500,In_1412,In_827);
or U1501 (N_1501,In_1180,In_792);
nor U1502 (N_1502,In_45,In_118);
nand U1503 (N_1503,In_1047,In_337);
or U1504 (N_1504,In_116,In_196);
nand U1505 (N_1505,In_85,In_844);
and U1506 (N_1506,In_84,In_105);
nor U1507 (N_1507,In_388,In_801);
or U1508 (N_1508,In_1105,In_248);
nor U1509 (N_1509,In_1404,In_1199);
and U1510 (N_1510,In_1264,In_730);
xnor U1511 (N_1511,In_275,In_1221);
nor U1512 (N_1512,In_719,In_632);
nand U1513 (N_1513,In_1336,In_578);
and U1514 (N_1514,In_676,In_854);
and U1515 (N_1515,In_75,In_139);
nand U1516 (N_1516,In_1230,In_189);
and U1517 (N_1517,In_1435,In_111);
or U1518 (N_1518,In_1347,In_767);
and U1519 (N_1519,In_963,In_758);
nor U1520 (N_1520,In_429,In_974);
nor U1521 (N_1521,In_1456,In_1136);
and U1522 (N_1522,In_686,In_1022);
nand U1523 (N_1523,In_29,In_95);
nor U1524 (N_1524,In_1303,In_1496);
or U1525 (N_1525,In_1373,In_346);
or U1526 (N_1526,In_1171,In_891);
and U1527 (N_1527,In_671,In_497);
nand U1528 (N_1528,In_1042,In_831);
xnor U1529 (N_1529,In_1446,In_1406);
nor U1530 (N_1530,In_1216,In_139);
and U1531 (N_1531,In_1474,In_1153);
or U1532 (N_1532,In_1196,In_668);
nand U1533 (N_1533,In_554,In_609);
and U1534 (N_1534,In_1226,In_172);
nand U1535 (N_1535,In_850,In_1201);
or U1536 (N_1536,In_82,In_333);
xnor U1537 (N_1537,In_925,In_677);
or U1538 (N_1538,In_507,In_464);
or U1539 (N_1539,In_1322,In_798);
and U1540 (N_1540,In_915,In_77);
nor U1541 (N_1541,In_105,In_681);
and U1542 (N_1542,In_588,In_1397);
and U1543 (N_1543,In_399,In_1412);
or U1544 (N_1544,In_499,In_672);
xor U1545 (N_1545,In_785,In_1257);
nand U1546 (N_1546,In_572,In_48);
or U1547 (N_1547,In_1429,In_185);
nand U1548 (N_1548,In_521,In_418);
or U1549 (N_1549,In_1381,In_1123);
and U1550 (N_1550,In_228,In_80);
and U1551 (N_1551,In_552,In_730);
nor U1552 (N_1552,In_973,In_1037);
xnor U1553 (N_1553,In_1376,In_541);
or U1554 (N_1554,In_985,In_1450);
nand U1555 (N_1555,In_379,In_66);
and U1556 (N_1556,In_1276,In_217);
and U1557 (N_1557,In_991,In_536);
nand U1558 (N_1558,In_550,In_650);
and U1559 (N_1559,In_870,In_1367);
or U1560 (N_1560,In_1245,In_1114);
and U1561 (N_1561,In_398,In_849);
nor U1562 (N_1562,In_498,In_1134);
nand U1563 (N_1563,In_1189,In_994);
or U1564 (N_1564,In_1233,In_1012);
nand U1565 (N_1565,In_216,In_859);
nor U1566 (N_1566,In_984,In_756);
or U1567 (N_1567,In_246,In_937);
and U1568 (N_1568,In_411,In_88);
or U1569 (N_1569,In_794,In_1475);
and U1570 (N_1570,In_52,In_521);
nand U1571 (N_1571,In_198,In_829);
xor U1572 (N_1572,In_1380,In_532);
and U1573 (N_1573,In_1051,In_798);
or U1574 (N_1574,In_977,In_647);
xnor U1575 (N_1575,In_500,In_48);
or U1576 (N_1576,In_990,In_1230);
nand U1577 (N_1577,In_892,In_474);
and U1578 (N_1578,In_852,In_1114);
and U1579 (N_1579,In_901,In_500);
and U1580 (N_1580,In_470,In_99);
and U1581 (N_1581,In_252,In_1092);
and U1582 (N_1582,In_145,In_917);
nor U1583 (N_1583,In_1214,In_146);
and U1584 (N_1584,In_534,In_124);
nand U1585 (N_1585,In_182,In_770);
nor U1586 (N_1586,In_1381,In_1474);
nand U1587 (N_1587,In_203,In_370);
or U1588 (N_1588,In_1176,In_389);
nand U1589 (N_1589,In_1481,In_706);
nor U1590 (N_1590,In_1440,In_53);
or U1591 (N_1591,In_569,In_322);
nor U1592 (N_1592,In_601,In_457);
or U1593 (N_1593,In_72,In_42);
and U1594 (N_1594,In_43,In_647);
nand U1595 (N_1595,In_1437,In_1419);
nor U1596 (N_1596,In_844,In_681);
xor U1597 (N_1597,In_1132,In_1055);
or U1598 (N_1598,In_321,In_630);
and U1599 (N_1599,In_1470,In_128);
xor U1600 (N_1600,In_1273,In_434);
nor U1601 (N_1601,In_438,In_885);
or U1602 (N_1602,In_590,In_949);
and U1603 (N_1603,In_487,In_915);
and U1604 (N_1604,In_921,In_903);
and U1605 (N_1605,In_581,In_1002);
xnor U1606 (N_1606,In_133,In_799);
nand U1607 (N_1607,In_1251,In_1426);
or U1608 (N_1608,In_114,In_929);
and U1609 (N_1609,In_247,In_110);
nand U1610 (N_1610,In_1343,In_2);
nand U1611 (N_1611,In_1034,In_317);
nor U1612 (N_1612,In_41,In_449);
or U1613 (N_1613,In_127,In_79);
and U1614 (N_1614,In_631,In_76);
nor U1615 (N_1615,In_119,In_454);
nand U1616 (N_1616,In_1419,In_299);
nor U1617 (N_1617,In_293,In_1280);
nand U1618 (N_1618,In_1406,In_168);
and U1619 (N_1619,In_522,In_1401);
or U1620 (N_1620,In_338,In_913);
and U1621 (N_1621,In_1005,In_362);
and U1622 (N_1622,In_1173,In_182);
nand U1623 (N_1623,In_279,In_1328);
nor U1624 (N_1624,In_1224,In_1456);
nand U1625 (N_1625,In_1069,In_708);
and U1626 (N_1626,In_291,In_897);
nor U1627 (N_1627,In_340,In_1251);
and U1628 (N_1628,In_1279,In_903);
nor U1629 (N_1629,In_1216,In_1135);
nor U1630 (N_1630,In_160,In_311);
and U1631 (N_1631,In_1158,In_419);
and U1632 (N_1632,In_1471,In_756);
nand U1633 (N_1633,In_614,In_259);
and U1634 (N_1634,In_161,In_881);
and U1635 (N_1635,In_609,In_1173);
nand U1636 (N_1636,In_1281,In_1);
nand U1637 (N_1637,In_1343,In_1402);
nor U1638 (N_1638,In_1396,In_1454);
or U1639 (N_1639,In_932,In_115);
or U1640 (N_1640,In_68,In_1171);
and U1641 (N_1641,In_29,In_1107);
xnor U1642 (N_1642,In_1,In_218);
and U1643 (N_1643,In_979,In_303);
and U1644 (N_1644,In_939,In_629);
or U1645 (N_1645,In_1285,In_586);
and U1646 (N_1646,In_849,In_1317);
xor U1647 (N_1647,In_577,In_1351);
nand U1648 (N_1648,In_148,In_1029);
or U1649 (N_1649,In_23,In_1172);
and U1650 (N_1650,In_1078,In_746);
xor U1651 (N_1651,In_683,In_1008);
nor U1652 (N_1652,In_1033,In_522);
or U1653 (N_1653,In_1421,In_1231);
nand U1654 (N_1654,In_618,In_187);
nand U1655 (N_1655,In_1321,In_620);
and U1656 (N_1656,In_428,In_946);
nor U1657 (N_1657,In_681,In_670);
and U1658 (N_1658,In_275,In_1441);
and U1659 (N_1659,In_479,In_1232);
nand U1660 (N_1660,In_503,In_815);
or U1661 (N_1661,In_1239,In_1206);
nand U1662 (N_1662,In_124,In_706);
nand U1663 (N_1663,In_1355,In_627);
nor U1664 (N_1664,In_1015,In_283);
nor U1665 (N_1665,In_712,In_1141);
xor U1666 (N_1666,In_336,In_1473);
nand U1667 (N_1667,In_330,In_1462);
or U1668 (N_1668,In_236,In_1043);
nor U1669 (N_1669,In_713,In_126);
nand U1670 (N_1670,In_97,In_288);
nor U1671 (N_1671,In_1343,In_1001);
and U1672 (N_1672,In_720,In_361);
nor U1673 (N_1673,In_462,In_799);
nor U1674 (N_1674,In_1225,In_1477);
xnor U1675 (N_1675,In_7,In_537);
and U1676 (N_1676,In_163,In_756);
or U1677 (N_1677,In_889,In_1309);
xor U1678 (N_1678,In_422,In_365);
and U1679 (N_1679,In_455,In_1482);
and U1680 (N_1680,In_1301,In_666);
nor U1681 (N_1681,In_228,In_866);
nor U1682 (N_1682,In_85,In_655);
nand U1683 (N_1683,In_1203,In_1);
or U1684 (N_1684,In_1352,In_332);
or U1685 (N_1685,In_534,In_260);
nor U1686 (N_1686,In_1052,In_590);
nor U1687 (N_1687,In_1282,In_1359);
nand U1688 (N_1688,In_1352,In_1208);
nand U1689 (N_1689,In_1124,In_1442);
nand U1690 (N_1690,In_126,In_332);
xnor U1691 (N_1691,In_1091,In_979);
and U1692 (N_1692,In_770,In_749);
or U1693 (N_1693,In_1089,In_74);
nor U1694 (N_1694,In_779,In_496);
nor U1695 (N_1695,In_933,In_128);
nor U1696 (N_1696,In_951,In_1315);
and U1697 (N_1697,In_392,In_1276);
or U1698 (N_1698,In_72,In_743);
or U1699 (N_1699,In_1351,In_592);
nand U1700 (N_1700,In_971,In_888);
or U1701 (N_1701,In_194,In_965);
nand U1702 (N_1702,In_1453,In_1435);
and U1703 (N_1703,In_1040,In_256);
nand U1704 (N_1704,In_550,In_1038);
and U1705 (N_1705,In_1155,In_289);
or U1706 (N_1706,In_518,In_138);
and U1707 (N_1707,In_633,In_376);
or U1708 (N_1708,In_306,In_1059);
nand U1709 (N_1709,In_403,In_411);
nor U1710 (N_1710,In_147,In_473);
nor U1711 (N_1711,In_1465,In_974);
nor U1712 (N_1712,In_1386,In_1408);
nand U1713 (N_1713,In_1178,In_510);
nor U1714 (N_1714,In_1002,In_89);
xnor U1715 (N_1715,In_116,In_145);
xor U1716 (N_1716,In_1221,In_1251);
or U1717 (N_1717,In_928,In_745);
xor U1718 (N_1718,In_25,In_379);
xor U1719 (N_1719,In_1421,In_588);
nand U1720 (N_1720,In_60,In_943);
nor U1721 (N_1721,In_213,In_1376);
nand U1722 (N_1722,In_62,In_140);
and U1723 (N_1723,In_291,In_352);
xor U1724 (N_1724,In_1061,In_127);
and U1725 (N_1725,In_1135,In_1414);
or U1726 (N_1726,In_1204,In_1085);
or U1727 (N_1727,In_196,In_427);
xnor U1728 (N_1728,In_1219,In_1377);
and U1729 (N_1729,In_1373,In_524);
nand U1730 (N_1730,In_669,In_884);
and U1731 (N_1731,In_59,In_1085);
xor U1732 (N_1732,In_1364,In_1062);
and U1733 (N_1733,In_699,In_1145);
nand U1734 (N_1734,In_151,In_600);
nand U1735 (N_1735,In_1098,In_324);
nand U1736 (N_1736,In_604,In_1055);
nor U1737 (N_1737,In_663,In_350);
and U1738 (N_1738,In_569,In_515);
and U1739 (N_1739,In_1484,In_603);
nor U1740 (N_1740,In_413,In_242);
and U1741 (N_1741,In_1212,In_1375);
nand U1742 (N_1742,In_211,In_68);
nand U1743 (N_1743,In_0,In_1238);
nand U1744 (N_1744,In_697,In_1019);
nor U1745 (N_1745,In_647,In_291);
nor U1746 (N_1746,In_340,In_1016);
xnor U1747 (N_1747,In_1020,In_279);
nand U1748 (N_1748,In_721,In_1263);
or U1749 (N_1749,In_694,In_872);
nor U1750 (N_1750,In_1439,In_503);
or U1751 (N_1751,In_1150,In_1265);
and U1752 (N_1752,In_753,In_957);
xor U1753 (N_1753,In_1448,In_500);
and U1754 (N_1754,In_1087,In_1252);
nand U1755 (N_1755,In_981,In_852);
and U1756 (N_1756,In_107,In_775);
or U1757 (N_1757,In_74,In_1492);
and U1758 (N_1758,In_452,In_799);
nor U1759 (N_1759,In_439,In_1167);
xor U1760 (N_1760,In_180,In_61);
or U1761 (N_1761,In_895,In_662);
or U1762 (N_1762,In_941,In_178);
and U1763 (N_1763,In_827,In_1404);
nor U1764 (N_1764,In_781,In_588);
nand U1765 (N_1765,In_331,In_48);
or U1766 (N_1766,In_1362,In_1349);
and U1767 (N_1767,In_803,In_995);
nor U1768 (N_1768,In_843,In_631);
nor U1769 (N_1769,In_1375,In_417);
or U1770 (N_1770,In_574,In_33);
nor U1771 (N_1771,In_701,In_357);
nor U1772 (N_1772,In_638,In_680);
and U1773 (N_1773,In_1172,In_1142);
or U1774 (N_1774,In_1076,In_441);
nor U1775 (N_1775,In_1219,In_1007);
nor U1776 (N_1776,In_1388,In_352);
or U1777 (N_1777,In_128,In_276);
or U1778 (N_1778,In_1139,In_1234);
and U1779 (N_1779,In_925,In_1371);
nand U1780 (N_1780,In_317,In_1444);
nand U1781 (N_1781,In_226,In_913);
and U1782 (N_1782,In_606,In_1249);
or U1783 (N_1783,In_1103,In_549);
nand U1784 (N_1784,In_1005,In_70);
and U1785 (N_1785,In_152,In_865);
or U1786 (N_1786,In_39,In_1125);
nand U1787 (N_1787,In_343,In_358);
and U1788 (N_1788,In_1016,In_519);
and U1789 (N_1789,In_1462,In_721);
nand U1790 (N_1790,In_767,In_1114);
or U1791 (N_1791,In_1023,In_1152);
nor U1792 (N_1792,In_907,In_521);
or U1793 (N_1793,In_1078,In_118);
and U1794 (N_1794,In_679,In_356);
or U1795 (N_1795,In_177,In_179);
and U1796 (N_1796,In_1373,In_570);
nand U1797 (N_1797,In_429,In_919);
nand U1798 (N_1798,In_1311,In_326);
nor U1799 (N_1799,In_968,In_1336);
nand U1800 (N_1800,In_1497,In_1213);
nor U1801 (N_1801,In_767,In_574);
and U1802 (N_1802,In_1077,In_602);
nand U1803 (N_1803,In_869,In_381);
and U1804 (N_1804,In_1232,In_1475);
and U1805 (N_1805,In_223,In_977);
and U1806 (N_1806,In_1425,In_1125);
nor U1807 (N_1807,In_622,In_493);
xor U1808 (N_1808,In_553,In_1339);
and U1809 (N_1809,In_996,In_1155);
nand U1810 (N_1810,In_299,In_885);
or U1811 (N_1811,In_1034,In_575);
nor U1812 (N_1812,In_1276,In_26);
or U1813 (N_1813,In_883,In_524);
or U1814 (N_1814,In_827,In_148);
nor U1815 (N_1815,In_463,In_702);
nand U1816 (N_1816,In_857,In_742);
or U1817 (N_1817,In_887,In_489);
and U1818 (N_1818,In_354,In_1331);
nor U1819 (N_1819,In_1496,In_1089);
nand U1820 (N_1820,In_330,In_1249);
or U1821 (N_1821,In_1047,In_1338);
xor U1822 (N_1822,In_1349,In_679);
nand U1823 (N_1823,In_420,In_541);
nand U1824 (N_1824,In_247,In_77);
and U1825 (N_1825,In_1333,In_1027);
nor U1826 (N_1826,In_480,In_543);
nand U1827 (N_1827,In_62,In_792);
or U1828 (N_1828,In_129,In_604);
or U1829 (N_1829,In_1085,In_208);
or U1830 (N_1830,In_783,In_1424);
xnor U1831 (N_1831,In_490,In_680);
nand U1832 (N_1832,In_116,In_282);
nor U1833 (N_1833,In_812,In_389);
nor U1834 (N_1834,In_338,In_1310);
nand U1835 (N_1835,In_1012,In_125);
or U1836 (N_1836,In_801,In_259);
nand U1837 (N_1837,In_980,In_1250);
xor U1838 (N_1838,In_585,In_1057);
nand U1839 (N_1839,In_175,In_364);
nor U1840 (N_1840,In_26,In_519);
nor U1841 (N_1841,In_897,In_549);
nor U1842 (N_1842,In_681,In_993);
or U1843 (N_1843,In_1018,In_960);
and U1844 (N_1844,In_1360,In_1352);
nand U1845 (N_1845,In_204,In_1345);
xnor U1846 (N_1846,In_1452,In_823);
and U1847 (N_1847,In_901,In_313);
and U1848 (N_1848,In_766,In_610);
xor U1849 (N_1849,In_146,In_577);
nor U1850 (N_1850,In_807,In_757);
or U1851 (N_1851,In_546,In_790);
and U1852 (N_1852,In_81,In_1437);
and U1853 (N_1853,In_657,In_1184);
nor U1854 (N_1854,In_1132,In_489);
nand U1855 (N_1855,In_683,In_355);
or U1856 (N_1856,In_1156,In_252);
xor U1857 (N_1857,In_153,In_975);
nor U1858 (N_1858,In_139,In_1100);
nor U1859 (N_1859,In_379,In_222);
or U1860 (N_1860,In_175,In_261);
and U1861 (N_1861,In_379,In_1029);
or U1862 (N_1862,In_1431,In_530);
and U1863 (N_1863,In_1207,In_1065);
and U1864 (N_1864,In_877,In_496);
nand U1865 (N_1865,In_167,In_721);
nand U1866 (N_1866,In_1465,In_398);
or U1867 (N_1867,In_381,In_1212);
xnor U1868 (N_1868,In_773,In_596);
nand U1869 (N_1869,In_1149,In_111);
and U1870 (N_1870,In_710,In_1056);
and U1871 (N_1871,In_891,In_937);
nand U1872 (N_1872,In_327,In_889);
nand U1873 (N_1873,In_679,In_1016);
or U1874 (N_1874,In_1059,In_333);
nor U1875 (N_1875,In_264,In_35);
xor U1876 (N_1876,In_841,In_1256);
and U1877 (N_1877,In_483,In_41);
nand U1878 (N_1878,In_126,In_544);
or U1879 (N_1879,In_188,In_1123);
nand U1880 (N_1880,In_1256,In_700);
and U1881 (N_1881,In_995,In_450);
nand U1882 (N_1882,In_475,In_1339);
or U1883 (N_1883,In_521,In_1238);
xnor U1884 (N_1884,In_319,In_477);
and U1885 (N_1885,In_987,In_690);
and U1886 (N_1886,In_234,In_1187);
nor U1887 (N_1887,In_759,In_1445);
or U1888 (N_1888,In_979,In_1048);
nor U1889 (N_1889,In_328,In_1033);
or U1890 (N_1890,In_549,In_58);
and U1891 (N_1891,In_1082,In_1374);
and U1892 (N_1892,In_982,In_465);
or U1893 (N_1893,In_652,In_1402);
and U1894 (N_1894,In_805,In_823);
nand U1895 (N_1895,In_224,In_36);
and U1896 (N_1896,In_1475,In_575);
and U1897 (N_1897,In_96,In_544);
or U1898 (N_1898,In_197,In_488);
nand U1899 (N_1899,In_648,In_240);
and U1900 (N_1900,In_1054,In_230);
nor U1901 (N_1901,In_1423,In_382);
and U1902 (N_1902,In_1148,In_1271);
nand U1903 (N_1903,In_898,In_442);
xor U1904 (N_1904,In_502,In_3);
nand U1905 (N_1905,In_1286,In_471);
nand U1906 (N_1906,In_745,In_774);
or U1907 (N_1907,In_600,In_1342);
nand U1908 (N_1908,In_217,In_1377);
nand U1909 (N_1909,In_845,In_95);
nand U1910 (N_1910,In_680,In_1158);
nor U1911 (N_1911,In_1411,In_1377);
or U1912 (N_1912,In_898,In_428);
nor U1913 (N_1913,In_1418,In_452);
nand U1914 (N_1914,In_541,In_1013);
and U1915 (N_1915,In_264,In_1227);
nand U1916 (N_1916,In_464,In_119);
nand U1917 (N_1917,In_209,In_139);
nor U1918 (N_1918,In_542,In_217);
xnor U1919 (N_1919,In_875,In_1111);
and U1920 (N_1920,In_329,In_1383);
or U1921 (N_1921,In_50,In_1186);
and U1922 (N_1922,In_712,In_1283);
or U1923 (N_1923,In_1032,In_1349);
or U1924 (N_1924,In_474,In_637);
xnor U1925 (N_1925,In_1410,In_1429);
nor U1926 (N_1926,In_1016,In_1336);
nand U1927 (N_1927,In_851,In_692);
nand U1928 (N_1928,In_748,In_1469);
xor U1929 (N_1929,In_1374,In_1235);
or U1930 (N_1930,In_138,In_1142);
nand U1931 (N_1931,In_359,In_1344);
nand U1932 (N_1932,In_1146,In_628);
and U1933 (N_1933,In_298,In_514);
nand U1934 (N_1934,In_949,In_882);
or U1935 (N_1935,In_153,In_1428);
and U1936 (N_1936,In_693,In_1209);
and U1937 (N_1937,In_405,In_455);
and U1938 (N_1938,In_1128,In_436);
and U1939 (N_1939,In_1183,In_670);
or U1940 (N_1940,In_821,In_250);
nor U1941 (N_1941,In_74,In_1194);
nand U1942 (N_1942,In_292,In_895);
nor U1943 (N_1943,In_1001,In_1300);
and U1944 (N_1944,In_470,In_61);
nor U1945 (N_1945,In_1005,In_874);
nor U1946 (N_1946,In_1439,In_149);
nand U1947 (N_1947,In_817,In_126);
nor U1948 (N_1948,In_23,In_1007);
and U1949 (N_1949,In_414,In_1134);
xnor U1950 (N_1950,In_1497,In_1273);
nand U1951 (N_1951,In_1210,In_754);
or U1952 (N_1952,In_366,In_1425);
or U1953 (N_1953,In_70,In_368);
nand U1954 (N_1954,In_1321,In_1192);
and U1955 (N_1955,In_128,In_1378);
or U1956 (N_1956,In_428,In_1069);
and U1957 (N_1957,In_1192,In_1418);
nand U1958 (N_1958,In_1230,In_1294);
and U1959 (N_1959,In_999,In_979);
nand U1960 (N_1960,In_960,In_553);
and U1961 (N_1961,In_314,In_218);
nand U1962 (N_1962,In_1089,In_1179);
nor U1963 (N_1963,In_1060,In_302);
or U1964 (N_1964,In_1484,In_1079);
and U1965 (N_1965,In_764,In_1444);
and U1966 (N_1966,In_628,In_560);
and U1967 (N_1967,In_106,In_219);
xor U1968 (N_1968,In_539,In_78);
nand U1969 (N_1969,In_1379,In_698);
and U1970 (N_1970,In_1453,In_1032);
nor U1971 (N_1971,In_482,In_754);
or U1972 (N_1972,In_305,In_472);
nand U1973 (N_1973,In_327,In_1174);
nor U1974 (N_1974,In_1278,In_1149);
nand U1975 (N_1975,In_919,In_834);
or U1976 (N_1976,In_120,In_461);
or U1977 (N_1977,In_441,In_67);
or U1978 (N_1978,In_1169,In_825);
xor U1979 (N_1979,In_1167,In_1176);
and U1980 (N_1980,In_1358,In_1218);
or U1981 (N_1981,In_669,In_1003);
and U1982 (N_1982,In_229,In_1419);
nand U1983 (N_1983,In_624,In_1124);
nor U1984 (N_1984,In_464,In_261);
nor U1985 (N_1985,In_526,In_71);
nor U1986 (N_1986,In_963,In_131);
nand U1987 (N_1987,In_84,In_1303);
xor U1988 (N_1988,In_1175,In_312);
and U1989 (N_1989,In_748,In_972);
and U1990 (N_1990,In_1497,In_469);
and U1991 (N_1991,In_361,In_581);
and U1992 (N_1992,In_37,In_1060);
and U1993 (N_1993,In_426,In_128);
nand U1994 (N_1994,In_1438,In_1489);
or U1995 (N_1995,In_5,In_1138);
nand U1996 (N_1996,In_667,In_1135);
and U1997 (N_1997,In_830,In_558);
and U1998 (N_1998,In_213,In_525);
nand U1999 (N_1999,In_1371,In_819);
nand U2000 (N_2000,In_688,In_482);
nand U2001 (N_2001,In_435,In_21);
xnor U2002 (N_2002,In_838,In_241);
xor U2003 (N_2003,In_1306,In_716);
nor U2004 (N_2004,In_744,In_209);
and U2005 (N_2005,In_946,In_47);
or U2006 (N_2006,In_559,In_1096);
nand U2007 (N_2007,In_389,In_874);
or U2008 (N_2008,In_1012,In_133);
or U2009 (N_2009,In_875,In_509);
nand U2010 (N_2010,In_328,In_665);
xor U2011 (N_2011,In_128,In_910);
nand U2012 (N_2012,In_600,In_1269);
nor U2013 (N_2013,In_279,In_8);
nor U2014 (N_2014,In_996,In_834);
nand U2015 (N_2015,In_1268,In_317);
and U2016 (N_2016,In_468,In_575);
xnor U2017 (N_2017,In_1140,In_451);
nor U2018 (N_2018,In_551,In_1333);
and U2019 (N_2019,In_1173,In_1100);
or U2020 (N_2020,In_1481,In_1260);
or U2021 (N_2021,In_1417,In_1479);
nand U2022 (N_2022,In_767,In_394);
xnor U2023 (N_2023,In_119,In_444);
and U2024 (N_2024,In_383,In_480);
xor U2025 (N_2025,In_933,In_203);
nand U2026 (N_2026,In_1118,In_1429);
or U2027 (N_2027,In_367,In_667);
or U2028 (N_2028,In_1293,In_71);
nand U2029 (N_2029,In_802,In_852);
xor U2030 (N_2030,In_468,In_510);
xor U2031 (N_2031,In_800,In_434);
nor U2032 (N_2032,In_245,In_405);
and U2033 (N_2033,In_841,In_1430);
and U2034 (N_2034,In_686,In_627);
nand U2035 (N_2035,In_1235,In_55);
nor U2036 (N_2036,In_151,In_987);
nor U2037 (N_2037,In_985,In_802);
or U2038 (N_2038,In_736,In_1236);
nor U2039 (N_2039,In_1255,In_1304);
or U2040 (N_2040,In_1081,In_1427);
xor U2041 (N_2041,In_550,In_299);
nor U2042 (N_2042,In_1287,In_778);
nor U2043 (N_2043,In_546,In_528);
xnor U2044 (N_2044,In_86,In_211);
xor U2045 (N_2045,In_229,In_449);
nand U2046 (N_2046,In_1132,In_505);
xnor U2047 (N_2047,In_1206,In_48);
xor U2048 (N_2048,In_68,In_419);
nand U2049 (N_2049,In_812,In_1002);
nor U2050 (N_2050,In_689,In_1159);
nor U2051 (N_2051,In_219,In_733);
nor U2052 (N_2052,In_1423,In_1417);
and U2053 (N_2053,In_34,In_254);
xnor U2054 (N_2054,In_692,In_38);
nand U2055 (N_2055,In_486,In_136);
nand U2056 (N_2056,In_1308,In_524);
nor U2057 (N_2057,In_235,In_1325);
and U2058 (N_2058,In_69,In_1195);
and U2059 (N_2059,In_436,In_366);
xnor U2060 (N_2060,In_960,In_199);
nor U2061 (N_2061,In_622,In_149);
and U2062 (N_2062,In_1353,In_796);
or U2063 (N_2063,In_58,In_727);
or U2064 (N_2064,In_235,In_1490);
and U2065 (N_2065,In_870,In_10);
nor U2066 (N_2066,In_450,In_934);
or U2067 (N_2067,In_1034,In_427);
or U2068 (N_2068,In_555,In_249);
nand U2069 (N_2069,In_998,In_146);
and U2070 (N_2070,In_1117,In_1039);
xor U2071 (N_2071,In_906,In_123);
xnor U2072 (N_2072,In_359,In_1380);
xnor U2073 (N_2073,In_1210,In_397);
xnor U2074 (N_2074,In_988,In_578);
or U2075 (N_2075,In_763,In_1240);
xnor U2076 (N_2076,In_1129,In_991);
and U2077 (N_2077,In_876,In_1478);
nand U2078 (N_2078,In_331,In_262);
nand U2079 (N_2079,In_179,In_1158);
or U2080 (N_2080,In_1364,In_794);
nor U2081 (N_2081,In_629,In_194);
nor U2082 (N_2082,In_858,In_1455);
nand U2083 (N_2083,In_484,In_1218);
nand U2084 (N_2084,In_420,In_1141);
nand U2085 (N_2085,In_1053,In_363);
nor U2086 (N_2086,In_1441,In_672);
and U2087 (N_2087,In_1294,In_1338);
nand U2088 (N_2088,In_482,In_414);
or U2089 (N_2089,In_274,In_864);
or U2090 (N_2090,In_1083,In_1279);
or U2091 (N_2091,In_862,In_1302);
xor U2092 (N_2092,In_1460,In_1061);
nor U2093 (N_2093,In_1303,In_437);
nor U2094 (N_2094,In_1266,In_613);
and U2095 (N_2095,In_1178,In_1137);
nor U2096 (N_2096,In_31,In_420);
nand U2097 (N_2097,In_1151,In_1192);
nor U2098 (N_2098,In_337,In_770);
or U2099 (N_2099,In_1350,In_119);
xor U2100 (N_2100,In_713,In_1422);
nor U2101 (N_2101,In_17,In_1499);
and U2102 (N_2102,In_465,In_1096);
and U2103 (N_2103,In_1196,In_1145);
nor U2104 (N_2104,In_153,In_1238);
xor U2105 (N_2105,In_1090,In_815);
nor U2106 (N_2106,In_1095,In_808);
nor U2107 (N_2107,In_574,In_49);
or U2108 (N_2108,In_250,In_1151);
nor U2109 (N_2109,In_88,In_311);
nand U2110 (N_2110,In_259,In_1264);
nor U2111 (N_2111,In_308,In_578);
and U2112 (N_2112,In_564,In_1073);
nand U2113 (N_2113,In_1030,In_10);
nand U2114 (N_2114,In_832,In_243);
or U2115 (N_2115,In_602,In_1465);
xor U2116 (N_2116,In_913,In_33);
nand U2117 (N_2117,In_686,In_180);
or U2118 (N_2118,In_1040,In_962);
nor U2119 (N_2119,In_237,In_495);
nor U2120 (N_2120,In_163,In_610);
nor U2121 (N_2121,In_1262,In_1156);
nor U2122 (N_2122,In_9,In_1486);
xor U2123 (N_2123,In_1061,In_1247);
xor U2124 (N_2124,In_443,In_779);
and U2125 (N_2125,In_4,In_921);
nor U2126 (N_2126,In_899,In_223);
nor U2127 (N_2127,In_707,In_1214);
nor U2128 (N_2128,In_631,In_1369);
or U2129 (N_2129,In_607,In_999);
nor U2130 (N_2130,In_1298,In_13);
nand U2131 (N_2131,In_1345,In_41);
nand U2132 (N_2132,In_705,In_128);
and U2133 (N_2133,In_531,In_944);
nor U2134 (N_2134,In_1319,In_683);
and U2135 (N_2135,In_744,In_965);
or U2136 (N_2136,In_1126,In_8);
nor U2137 (N_2137,In_298,In_1420);
nor U2138 (N_2138,In_438,In_859);
nand U2139 (N_2139,In_228,In_506);
nand U2140 (N_2140,In_1374,In_485);
or U2141 (N_2141,In_599,In_1280);
nand U2142 (N_2142,In_320,In_826);
xnor U2143 (N_2143,In_792,In_432);
and U2144 (N_2144,In_730,In_277);
and U2145 (N_2145,In_718,In_351);
and U2146 (N_2146,In_525,In_236);
nand U2147 (N_2147,In_1287,In_945);
xnor U2148 (N_2148,In_743,In_574);
and U2149 (N_2149,In_1416,In_1456);
nor U2150 (N_2150,In_1297,In_1086);
nor U2151 (N_2151,In_7,In_96);
xnor U2152 (N_2152,In_1389,In_366);
nand U2153 (N_2153,In_925,In_272);
nor U2154 (N_2154,In_1245,In_1376);
nand U2155 (N_2155,In_949,In_717);
nor U2156 (N_2156,In_739,In_1378);
nor U2157 (N_2157,In_1338,In_523);
nand U2158 (N_2158,In_414,In_1424);
nor U2159 (N_2159,In_819,In_454);
or U2160 (N_2160,In_1031,In_966);
and U2161 (N_2161,In_37,In_944);
xnor U2162 (N_2162,In_1150,In_1363);
or U2163 (N_2163,In_1462,In_15);
and U2164 (N_2164,In_1234,In_1016);
and U2165 (N_2165,In_1059,In_1074);
nor U2166 (N_2166,In_920,In_1331);
and U2167 (N_2167,In_847,In_1279);
or U2168 (N_2168,In_98,In_300);
nor U2169 (N_2169,In_335,In_515);
nor U2170 (N_2170,In_290,In_1487);
nor U2171 (N_2171,In_736,In_268);
nor U2172 (N_2172,In_415,In_184);
xnor U2173 (N_2173,In_996,In_154);
and U2174 (N_2174,In_136,In_1478);
nor U2175 (N_2175,In_1391,In_901);
xor U2176 (N_2176,In_1322,In_738);
and U2177 (N_2177,In_684,In_590);
nand U2178 (N_2178,In_505,In_1142);
nand U2179 (N_2179,In_359,In_1024);
nor U2180 (N_2180,In_589,In_136);
nand U2181 (N_2181,In_506,In_280);
nor U2182 (N_2182,In_1373,In_759);
or U2183 (N_2183,In_1246,In_1062);
and U2184 (N_2184,In_1079,In_872);
nor U2185 (N_2185,In_53,In_949);
nand U2186 (N_2186,In_830,In_852);
and U2187 (N_2187,In_1210,In_4);
and U2188 (N_2188,In_775,In_203);
and U2189 (N_2189,In_357,In_1181);
nand U2190 (N_2190,In_237,In_244);
nand U2191 (N_2191,In_867,In_1431);
or U2192 (N_2192,In_393,In_645);
nand U2193 (N_2193,In_390,In_252);
xnor U2194 (N_2194,In_483,In_458);
nor U2195 (N_2195,In_161,In_703);
nand U2196 (N_2196,In_444,In_1373);
xor U2197 (N_2197,In_462,In_130);
and U2198 (N_2198,In_678,In_538);
nor U2199 (N_2199,In_1264,In_1252);
nor U2200 (N_2200,In_82,In_765);
or U2201 (N_2201,In_436,In_929);
nor U2202 (N_2202,In_774,In_909);
or U2203 (N_2203,In_756,In_953);
or U2204 (N_2204,In_984,In_624);
or U2205 (N_2205,In_1158,In_928);
nor U2206 (N_2206,In_253,In_1383);
and U2207 (N_2207,In_1147,In_610);
or U2208 (N_2208,In_800,In_561);
or U2209 (N_2209,In_491,In_245);
and U2210 (N_2210,In_938,In_812);
and U2211 (N_2211,In_29,In_510);
nand U2212 (N_2212,In_575,In_533);
nand U2213 (N_2213,In_52,In_787);
and U2214 (N_2214,In_499,In_594);
nor U2215 (N_2215,In_1358,In_611);
nor U2216 (N_2216,In_1108,In_500);
nor U2217 (N_2217,In_315,In_741);
xnor U2218 (N_2218,In_1220,In_918);
nand U2219 (N_2219,In_488,In_984);
nand U2220 (N_2220,In_1130,In_373);
xnor U2221 (N_2221,In_855,In_929);
and U2222 (N_2222,In_37,In_1292);
nor U2223 (N_2223,In_929,In_485);
nand U2224 (N_2224,In_791,In_1333);
and U2225 (N_2225,In_501,In_834);
or U2226 (N_2226,In_1343,In_1303);
and U2227 (N_2227,In_505,In_1356);
nor U2228 (N_2228,In_1132,In_1430);
or U2229 (N_2229,In_614,In_952);
nor U2230 (N_2230,In_1461,In_909);
xor U2231 (N_2231,In_493,In_332);
or U2232 (N_2232,In_1418,In_1044);
nand U2233 (N_2233,In_528,In_620);
nor U2234 (N_2234,In_1383,In_842);
nor U2235 (N_2235,In_656,In_765);
or U2236 (N_2236,In_323,In_13);
and U2237 (N_2237,In_1456,In_1220);
nand U2238 (N_2238,In_772,In_706);
and U2239 (N_2239,In_1463,In_1392);
and U2240 (N_2240,In_731,In_514);
nor U2241 (N_2241,In_690,In_1283);
and U2242 (N_2242,In_461,In_860);
xor U2243 (N_2243,In_193,In_756);
nand U2244 (N_2244,In_210,In_815);
and U2245 (N_2245,In_338,In_1324);
xnor U2246 (N_2246,In_730,In_829);
nand U2247 (N_2247,In_964,In_1104);
nand U2248 (N_2248,In_1294,In_293);
nor U2249 (N_2249,In_457,In_1334);
xnor U2250 (N_2250,In_771,In_1257);
nand U2251 (N_2251,In_812,In_103);
and U2252 (N_2252,In_422,In_958);
and U2253 (N_2253,In_1046,In_507);
nor U2254 (N_2254,In_713,In_944);
and U2255 (N_2255,In_1374,In_305);
nand U2256 (N_2256,In_13,In_1208);
nor U2257 (N_2257,In_692,In_1205);
or U2258 (N_2258,In_962,In_1259);
or U2259 (N_2259,In_122,In_558);
xnor U2260 (N_2260,In_1023,In_1054);
and U2261 (N_2261,In_1140,In_666);
nand U2262 (N_2262,In_956,In_252);
and U2263 (N_2263,In_794,In_374);
nor U2264 (N_2264,In_1256,In_1498);
and U2265 (N_2265,In_1396,In_181);
and U2266 (N_2266,In_869,In_256);
or U2267 (N_2267,In_743,In_193);
or U2268 (N_2268,In_241,In_1056);
nand U2269 (N_2269,In_1339,In_829);
and U2270 (N_2270,In_949,In_93);
xnor U2271 (N_2271,In_1173,In_1231);
and U2272 (N_2272,In_401,In_428);
nor U2273 (N_2273,In_1160,In_1273);
nand U2274 (N_2274,In_1448,In_1142);
nand U2275 (N_2275,In_591,In_45);
nand U2276 (N_2276,In_480,In_1469);
or U2277 (N_2277,In_687,In_334);
nor U2278 (N_2278,In_1037,In_403);
or U2279 (N_2279,In_1246,In_930);
and U2280 (N_2280,In_1107,In_1454);
and U2281 (N_2281,In_67,In_1057);
nand U2282 (N_2282,In_964,In_1374);
and U2283 (N_2283,In_877,In_197);
and U2284 (N_2284,In_483,In_627);
xnor U2285 (N_2285,In_1157,In_978);
xor U2286 (N_2286,In_1013,In_1107);
or U2287 (N_2287,In_1049,In_1333);
or U2288 (N_2288,In_1162,In_358);
nor U2289 (N_2289,In_719,In_1156);
or U2290 (N_2290,In_262,In_917);
and U2291 (N_2291,In_729,In_1376);
nand U2292 (N_2292,In_1304,In_1270);
and U2293 (N_2293,In_1121,In_1414);
nand U2294 (N_2294,In_347,In_1268);
and U2295 (N_2295,In_1110,In_98);
xor U2296 (N_2296,In_1285,In_157);
nand U2297 (N_2297,In_1355,In_846);
or U2298 (N_2298,In_1267,In_1338);
or U2299 (N_2299,In_28,In_750);
xor U2300 (N_2300,In_1401,In_1109);
or U2301 (N_2301,In_201,In_197);
or U2302 (N_2302,In_1482,In_1377);
xor U2303 (N_2303,In_565,In_56);
nand U2304 (N_2304,In_134,In_629);
nand U2305 (N_2305,In_1254,In_794);
nand U2306 (N_2306,In_459,In_935);
nor U2307 (N_2307,In_382,In_252);
nor U2308 (N_2308,In_716,In_244);
nand U2309 (N_2309,In_213,In_46);
xor U2310 (N_2310,In_920,In_875);
or U2311 (N_2311,In_524,In_370);
and U2312 (N_2312,In_1152,In_336);
nand U2313 (N_2313,In_268,In_237);
nor U2314 (N_2314,In_657,In_700);
xor U2315 (N_2315,In_599,In_93);
nor U2316 (N_2316,In_165,In_277);
nand U2317 (N_2317,In_1496,In_567);
nor U2318 (N_2318,In_273,In_717);
and U2319 (N_2319,In_415,In_1282);
nand U2320 (N_2320,In_558,In_533);
or U2321 (N_2321,In_1013,In_339);
or U2322 (N_2322,In_281,In_811);
and U2323 (N_2323,In_886,In_172);
nor U2324 (N_2324,In_827,In_585);
xor U2325 (N_2325,In_619,In_105);
nor U2326 (N_2326,In_1205,In_395);
xnor U2327 (N_2327,In_571,In_494);
and U2328 (N_2328,In_1413,In_555);
and U2329 (N_2329,In_797,In_109);
nor U2330 (N_2330,In_352,In_1246);
nor U2331 (N_2331,In_304,In_1131);
nor U2332 (N_2332,In_235,In_63);
or U2333 (N_2333,In_1000,In_1046);
and U2334 (N_2334,In_142,In_308);
nor U2335 (N_2335,In_737,In_1051);
nand U2336 (N_2336,In_1336,In_1236);
or U2337 (N_2337,In_227,In_790);
nand U2338 (N_2338,In_984,In_788);
nor U2339 (N_2339,In_1070,In_32);
and U2340 (N_2340,In_1097,In_1409);
nand U2341 (N_2341,In_16,In_244);
nand U2342 (N_2342,In_72,In_1029);
or U2343 (N_2343,In_155,In_1155);
and U2344 (N_2344,In_1417,In_355);
nor U2345 (N_2345,In_826,In_1383);
and U2346 (N_2346,In_419,In_119);
nor U2347 (N_2347,In_891,In_35);
or U2348 (N_2348,In_451,In_462);
nor U2349 (N_2349,In_1194,In_1291);
nor U2350 (N_2350,In_1020,In_1041);
nand U2351 (N_2351,In_965,In_1415);
or U2352 (N_2352,In_1125,In_400);
xor U2353 (N_2353,In_1425,In_274);
or U2354 (N_2354,In_1239,In_19);
nand U2355 (N_2355,In_1342,In_903);
nand U2356 (N_2356,In_779,In_1467);
and U2357 (N_2357,In_517,In_227);
and U2358 (N_2358,In_931,In_524);
xnor U2359 (N_2359,In_570,In_780);
nand U2360 (N_2360,In_862,In_194);
and U2361 (N_2361,In_1262,In_293);
nor U2362 (N_2362,In_903,In_96);
nand U2363 (N_2363,In_869,In_705);
nor U2364 (N_2364,In_622,In_823);
nor U2365 (N_2365,In_1188,In_269);
or U2366 (N_2366,In_1254,In_1273);
nor U2367 (N_2367,In_1367,In_250);
nor U2368 (N_2368,In_17,In_422);
and U2369 (N_2369,In_1005,In_503);
nor U2370 (N_2370,In_1017,In_247);
nor U2371 (N_2371,In_686,In_123);
nor U2372 (N_2372,In_261,In_1177);
xnor U2373 (N_2373,In_1120,In_61);
nor U2374 (N_2374,In_1109,In_1241);
nor U2375 (N_2375,In_776,In_72);
and U2376 (N_2376,In_96,In_552);
xor U2377 (N_2377,In_133,In_782);
nor U2378 (N_2378,In_944,In_958);
and U2379 (N_2379,In_993,In_763);
and U2380 (N_2380,In_1292,In_1013);
nand U2381 (N_2381,In_890,In_126);
or U2382 (N_2382,In_230,In_383);
and U2383 (N_2383,In_1,In_31);
nor U2384 (N_2384,In_1013,In_1168);
nand U2385 (N_2385,In_686,In_1010);
nor U2386 (N_2386,In_154,In_791);
or U2387 (N_2387,In_659,In_745);
nor U2388 (N_2388,In_162,In_0);
nor U2389 (N_2389,In_487,In_218);
nor U2390 (N_2390,In_112,In_318);
nand U2391 (N_2391,In_1038,In_604);
xor U2392 (N_2392,In_258,In_38);
xnor U2393 (N_2393,In_1386,In_355);
nand U2394 (N_2394,In_1152,In_149);
or U2395 (N_2395,In_160,In_454);
and U2396 (N_2396,In_138,In_1194);
or U2397 (N_2397,In_286,In_1135);
nand U2398 (N_2398,In_1499,In_764);
nand U2399 (N_2399,In_622,In_145);
nand U2400 (N_2400,In_454,In_285);
xor U2401 (N_2401,In_826,In_390);
or U2402 (N_2402,In_1484,In_570);
nand U2403 (N_2403,In_983,In_291);
nor U2404 (N_2404,In_125,In_811);
nand U2405 (N_2405,In_734,In_505);
nand U2406 (N_2406,In_579,In_8);
nor U2407 (N_2407,In_5,In_878);
nand U2408 (N_2408,In_1480,In_1342);
nand U2409 (N_2409,In_230,In_197);
xnor U2410 (N_2410,In_1400,In_616);
nor U2411 (N_2411,In_1263,In_565);
and U2412 (N_2412,In_756,In_1248);
nor U2413 (N_2413,In_1471,In_778);
nand U2414 (N_2414,In_301,In_441);
nand U2415 (N_2415,In_716,In_86);
nor U2416 (N_2416,In_795,In_263);
and U2417 (N_2417,In_1332,In_111);
nor U2418 (N_2418,In_529,In_205);
xor U2419 (N_2419,In_892,In_803);
nand U2420 (N_2420,In_629,In_720);
and U2421 (N_2421,In_750,In_98);
and U2422 (N_2422,In_1213,In_983);
xor U2423 (N_2423,In_1450,In_513);
nor U2424 (N_2424,In_974,In_1082);
or U2425 (N_2425,In_268,In_748);
nand U2426 (N_2426,In_967,In_965);
nand U2427 (N_2427,In_912,In_811);
or U2428 (N_2428,In_696,In_222);
or U2429 (N_2429,In_841,In_1393);
or U2430 (N_2430,In_1007,In_81);
nor U2431 (N_2431,In_203,In_225);
and U2432 (N_2432,In_883,In_341);
and U2433 (N_2433,In_1420,In_409);
nand U2434 (N_2434,In_159,In_274);
xnor U2435 (N_2435,In_1264,In_1491);
or U2436 (N_2436,In_619,In_178);
and U2437 (N_2437,In_1486,In_1189);
nand U2438 (N_2438,In_260,In_246);
or U2439 (N_2439,In_1412,In_1186);
and U2440 (N_2440,In_361,In_379);
and U2441 (N_2441,In_79,In_481);
or U2442 (N_2442,In_791,In_123);
or U2443 (N_2443,In_1441,In_978);
nor U2444 (N_2444,In_353,In_695);
nand U2445 (N_2445,In_1359,In_878);
or U2446 (N_2446,In_1198,In_670);
nor U2447 (N_2447,In_224,In_237);
nor U2448 (N_2448,In_952,In_506);
nor U2449 (N_2449,In_797,In_265);
nand U2450 (N_2450,In_130,In_272);
or U2451 (N_2451,In_1,In_1381);
nor U2452 (N_2452,In_55,In_173);
or U2453 (N_2453,In_415,In_377);
nand U2454 (N_2454,In_1018,In_1062);
nand U2455 (N_2455,In_936,In_787);
nand U2456 (N_2456,In_1437,In_705);
nand U2457 (N_2457,In_1178,In_315);
or U2458 (N_2458,In_337,In_235);
nand U2459 (N_2459,In_165,In_307);
nor U2460 (N_2460,In_542,In_975);
nor U2461 (N_2461,In_212,In_568);
nor U2462 (N_2462,In_510,In_1336);
or U2463 (N_2463,In_1384,In_968);
or U2464 (N_2464,In_1243,In_1088);
xnor U2465 (N_2465,In_1439,In_349);
or U2466 (N_2466,In_1201,In_92);
and U2467 (N_2467,In_182,In_604);
xnor U2468 (N_2468,In_1227,In_1205);
nand U2469 (N_2469,In_517,In_1439);
nand U2470 (N_2470,In_545,In_845);
nand U2471 (N_2471,In_1459,In_1218);
or U2472 (N_2472,In_1204,In_961);
and U2473 (N_2473,In_1050,In_1297);
and U2474 (N_2474,In_160,In_1249);
nand U2475 (N_2475,In_919,In_1257);
or U2476 (N_2476,In_245,In_1437);
nand U2477 (N_2477,In_1157,In_1068);
nor U2478 (N_2478,In_638,In_780);
nor U2479 (N_2479,In_708,In_1492);
nor U2480 (N_2480,In_896,In_1009);
nand U2481 (N_2481,In_261,In_173);
nor U2482 (N_2482,In_772,In_49);
nor U2483 (N_2483,In_911,In_1243);
nand U2484 (N_2484,In_539,In_1224);
and U2485 (N_2485,In_1295,In_1470);
nor U2486 (N_2486,In_1110,In_1381);
nand U2487 (N_2487,In_518,In_80);
nand U2488 (N_2488,In_1407,In_238);
nand U2489 (N_2489,In_457,In_807);
and U2490 (N_2490,In_815,In_113);
nor U2491 (N_2491,In_160,In_61);
nand U2492 (N_2492,In_574,In_692);
nand U2493 (N_2493,In_258,In_14);
and U2494 (N_2494,In_948,In_1173);
nor U2495 (N_2495,In_1362,In_904);
and U2496 (N_2496,In_350,In_964);
or U2497 (N_2497,In_618,In_984);
or U2498 (N_2498,In_347,In_1155);
or U2499 (N_2499,In_1282,In_491);
xnor U2500 (N_2500,In_1170,In_954);
nand U2501 (N_2501,In_545,In_732);
nand U2502 (N_2502,In_941,In_1307);
or U2503 (N_2503,In_638,In_272);
nor U2504 (N_2504,In_111,In_708);
nor U2505 (N_2505,In_1086,In_874);
nand U2506 (N_2506,In_1094,In_1401);
or U2507 (N_2507,In_24,In_415);
xor U2508 (N_2508,In_1490,In_31);
nor U2509 (N_2509,In_989,In_380);
and U2510 (N_2510,In_833,In_894);
and U2511 (N_2511,In_1000,In_1193);
xnor U2512 (N_2512,In_177,In_170);
nand U2513 (N_2513,In_192,In_861);
and U2514 (N_2514,In_612,In_621);
nor U2515 (N_2515,In_1274,In_905);
or U2516 (N_2516,In_618,In_697);
and U2517 (N_2517,In_273,In_1343);
and U2518 (N_2518,In_812,In_69);
and U2519 (N_2519,In_299,In_147);
or U2520 (N_2520,In_213,In_195);
nand U2521 (N_2521,In_537,In_401);
and U2522 (N_2522,In_649,In_175);
or U2523 (N_2523,In_222,In_1369);
xnor U2524 (N_2524,In_181,In_1363);
xor U2525 (N_2525,In_1014,In_610);
and U2526 (N_2526,In_937,In_960);
nand U2527 (N_2527,In_433,In_1426);
and U2528 (N_2528,In_791,In_1437);
or U2529 (N_2529,In_853,In_625);
or U2530 (N_2530,In_454,In_1160);
or U2531 (N_2531,In_881,In_817);
nor U2532 (N_2532,In_1305,In_751);
or U2533 (N_2533,In_303,In_400);
or U2534 (N_2534,In_544,In_38);
xor U2535 (N_2535,In_604,In_1465);
and U2536 (N_2536,In_1004,In_375);
or U2537 (N_2537,In_903,In_1423);
xor U2538 (N_2538,In_933,In_1286);
nand U2539 (N_2539,In_473,In_1240);
nand U2540 (N_2540,In_420,In_230);
nand U2541 (N_2541,In_475,In_65);
nand U2542 (N_2542,In_1231,In_211);
and U2543 (N_2543,In_806,In_305);
nand U2544 (N_2544,In_755,In_87);
nand U2545 (N_2545,In_898,In_6);
nand U2546 (N_2546,In_717,In_31);
and U2547 (N_2547,In_814,In_656);
nor U2548 (N_2548,In_416,In_764);
and U2549 (N_2549,In_1008,In_814);
nand U2550 (N_2550,In_35,In_1260);
or U2551 (N_2551,In_1185,In_501);
nand U2552 (N_2552,In_122,In_1329);
and U2553 (N_2553,In_258,In_1353);
nor U2554 (N_2554,In_1362,In_856);
xor U2555 (N_2555,In_1167,In_817);
nand U2556 (N_2556,In_885,In_161);
nand U2557 (N_2557,In_23,In_871);
and U2558 (N_2558,In_1084,In_733);
and U2559 (N_2559,In_854,In_444);
and U2560 (N_2560,In_1358,In_446);
and U2561 (N_2561,In_847,In_897);
and U2562 (N_2562,In_597,In_398);
nand U2563 (N_2563,In_689,In_417);
or U2564 (N_2564,In_963,In_916);
nor U2565 (N_2565,In_1286,In_1095);
nand U2566 (N_2566,In_651,In_339);
or U2567 (N_2567,In_1467,In_894);
nor U2568 (N_2568,In_981,In_939);
and U2569 (N_2569,In_1289,In_723);
nand U2570 (N_2570,In_946,In_476);
and U2571 (N_2571,In_390,In_272);
xor U2572 (N_2572,In_980,In_592);
and U2573 (N_2573,In_1203,In_221);
and U2574 (N_2574,In_640,In_1256);
or U2575 (N_2575,In_1309,In_1015);
and U2576 (N_2576,In_349,In_1012);
nor U2577 (N_2577,In_251,In_832);
and U2578 (N_2578,In_1495,In_12);
and U2579 (N_2579,In_674,In_739);
and U2580 (N_2580,In_1040,In_1212);
nor U2581 (N_2581,In_1153,In_686);
nand U2582 (N_2582,In_1312,In_539);
nand U2583 (N_2583,In_1145,In_461);
and U2584 (N_2584,In_764,In_1417);
nor U2585 (N_2585,In_1161,In_107);
or U2586 (N_2586,In_265,In_746);
nor U2587 (N_2587,In_1086,In_1);
nor U2588 (N_2588,In_1293,In_120);
or U2589 (N_2589,In_69,In_500);
or U2590 (N_2590,In_1296,In_717);
nand U2591 (N_2591,In_1059,In_1282);
nand U2592 (N_2592,In_639,In_349);
or U2593 (N_2593,In_923,In_633);
nand U2594 (N_2594,In_544,In_1134);
or U2595 (N_2595,In_969,In_1227);
or U2596 (N_2596,In_30,In_502);
or U2597 (N_2597,In_626,In_696);
nor U2598 (N_2598,In_676,In_295);
nand U2599 (N_2599,In_965,In_176);
nand U2600 (N_2600,In_224,In_1180);
or U2601 (N_2601,In_228,In_679);
or U2602 (N_2602,In_447,In_1206);
nor U2603 (N_2603,In_824,In_417);
nand U2604 (N_2604,In_774,In_1470);
nand U2605 (N_2605,In_281,In_718);
xor U2606 (N_2606,In_1455,In_853);
nor U2607 (N_2607,In_1184,In_210);
or U2608 (N_2608,In_1399,In_843);
xor U2609 (N_2609,In_1458,In_1366);
or U2610 (N_2610,In_568,In_620);
nand U2611 (N_2611,In_574,In_593);
and U2612 (N_2612,In_392,In_423);
or U2613 (N_2613,In_49,In_942);
xor U2614 (N_2614,In_1494,In_346);
nand U2615 (N_2615,In_337,In_440);
nor U2616 (N_2616,In_793,In_1392);
and U2617 (N_2617,In_26,In_745);
nand U2618 (N_2618,In_61,In_1459);
nand U2619 (N_2619,In_393,In_1036);
or U2620 (N_2620,In_1354,In_31);
nand U2621 (N_2621,In_1266,In_1076);
nor U2622 (N_2622,In_793,In_992);
nor U2623 (N_2623,In_1163,In_321);
and U2624 (N_2624,In_36,In_518);
and U2625 (N_2625,In_816,In_122);
and U2626 (N_2626,In_249,In_414);
nand U2627 (N_2627,In_965,In_844);
nor U2628 (N_2628,In_364,In_130);
nor U2629 (N_2629,In_747,In_1275);
or U2630 (N_2630,In_874,In_885);
nor U2631 (N_2631,In_601,In_685);
nand U2632 (N_2632,In_1379,In_38);
or U2633 (N_2633,In_372,In_509);
nor U2634 (N_2634,In_973,In_592);
and U2635 (N_2635,In_210,In_809);
nor U2636 (N_2636,In_699,In_77);
xnor U2637 (N_2637,In_285,In_534);
or U2638 (N_2638,In_654,In_3);
xnor U2639 (N_2639,In_141,In_393);
nand U2640 (N_2640,In_837,In_341);
and U2641 (N_2641,In_929,In_524);
or U2642 (N_2642,In_806,In_997);
and U2643 (N_2643,In_1279,In_646);
and U2644 (N_2644,In_995,In_563);
nand U2645 (N_2645,In_126,In_399);
nand U2646 (N_2646,In_927,In_236);
nor U2647 (N_2647,In_1309,In_1431);
nor U2648 (N_2648,In_1242,In_168);
nand U2649 (N_2649,In_904,In_1466);
nor U2650 (N_2650,In_66,In_1381);
xnor U2651 (N_2651,In_591,In_539);
nand U2652 (N_2652,In_1331,In_1131);
or U2653 (N_2653,In_796,In_132);
or U2654 (N_2654,In_252,In_812);
nor U2655 (N_2655,In_952,In_499);
nand U2656 (N_2656,In_1392,In_673);
and U2657 (N_2657,In_305,In_1122);
or U2658 (N_2658,In_1296,In_402);
xor U2659 (N_2659,In_340,In_1288);
nor U2660 (N_2660,In_1399,In_1046);
xor U2661 (N_2661,In_344,In_144);
xnor U2662 (N_2662,In_257,In_1144);
or U2663 (N_2663,In_768,In_446);
and U2664 (N_2664,In_1058,In_37);
or U2665 (N_2665,In_851,In_811);
nand U2666 (N_2666,In_383,In_177);
nand U2667 (N_2667,In_1058,In_368);
nand U2668 (N_2668,In_491,In_1277);
nand U2669 (N_2669,In_556,In_891);
nor U2670 (N_2670,In_778,In_890);
xnor U2671 (N_2671,In_459,In_277);
and U2672 (N_2672,In_923,In_344);
nor U2673 (N_2673,In_1328,In_412);
and U2674 (N_2674,In_1357,In_422);
or U2675 (N_2675,In_1140,In_959);
or U2676 (N_2676,In_1390,In_638);
or U2677 (N_2677,In_1375,In_628);
xnor U2678 (N_2678,In_1404,In_647);
nand U2679 (N_2679,In_574,In_178);
xor U2680 (N_2680,In_582,In_805);
nand U2681 (N_2681,In_74,In_396);
xor U2682 (N_2682,In_250,In_865);
and U2683 (N_2683,In_1356,In_304);
or U2684 (N_2684,In_1202,In_745);
or U2685 (N_2685,In_923,In_634);
or U2686 (N_2686,In_433,In_628);
or U2687 (N_2687,In_1201,In_1112);
or U2688 (N_2688,In_1137,In_1390);
nand U2689 (N_2689,In_572,In_1040);
nand U2690 (N_2690,In_821,In_324);
nand U2691 (N_2691,In_645,In_550);
xnor U2692 (N_2692,In_1101,In_49);
xor U2693 (N_2693,In_1152,In_1429);
and U2694 (N_2694,In_820,In_942);
xor U2695 (N_2695,In_1270,In_604);
nor U2696 (N_2696,In_333,In_1382);
nor U2697 (N_2697,In_493,In_232);
and U2698 (N_2698,In_14,In_1028);
xor U2699 (N_2699,In_877,In_224);
nor U2700 (N_2700,In_559,In_967);
nor U2701 (N_2701,In_1243,In_885);
or U2702 (N_2702,In_453,In_575);
and U2703 (N_2703,In_1067,In_1439);
or U2704 (N_2704,In_1262,In_50);
nor U2705 (N_2705,In_1282,In_879);
or U2706 (N_2706,In_174,In_15);
xnor U2707 (N_2707,In_725,In_783);
or U2708 (N_2708,In_1440,In_579);
nor U2709 (N_2709,In_1462,In_1414);
and U2710 (N_2710,In_558,In_193);
or U2711 (N_2711,In_1181,In_335);
xnor U2712 (N_2712,In_486,In_110);
or U2713 (N_2713,In_688,In_634);
or U2714 (N_2714,In_816,In_443);
nor U2715 (N_2715,In_1257,In_559);
and U2716 (N_2716,In_901,In_1337);
xor U2717 (N_2717,In_217,In_955);
and U2718 (N_2718,In_292,In_1136);
xor U2719 (N_2719,In_1201,In_273);
nor U2720 (N_2720,In_239,In_871);
nand U2721 (N_2721,In_17,In_403);
nor U2722 (N_2722,In_394,In_226);
and U2723 (N_2723,In_127,In_1490);
nor U2724 (N_2724,In_1423,In_764);
and U2725 (N_2725,In_1064,In_1310);
or U2726 (N_2726,In_158,In_564);
nand U2727 (N_2727,In_1192,In_111);
and U2728 (N_2728,In_283,In_594);
nand U2729 (N_2729,In_76,In_271);
xor U2730 (N_2730,In_229,In_294);
nor U2731 (N_2731,In_190,In_974);
xnor U2732 (N_2732,In_545,In_397);
nor U2733 (N_2733,In_817,In_956);
nor U2734 (N_2734,In_1236,In_1494);
nand U2735 (N_2735,In_12,In_1416);
nand U2736 (N_2736,In_425,In_1154);
nor U2737 (N_2737,In_723,In_680);
nand U2738 (N_2738,In_474,In_699);
nand U2739 (N_2739,In_1041,In_1343);
and U2740 (N_2740,In_863,In_1080);
xnor U2741 (N_2741,In_1130,In_1434);
and U2742 (N_2742,In_1289,In_120);
xnor U2743 (N_2743,In_1404,In_660);
or U2744 (N_2744,In_1158,In_1390);
or U2745 (N_2745,In_1006,In_91);
xor U2746 (N_2746,In_914,In_1006);
xor U2747 (N_2747,In_70,In_246);
nor U2748 (N_2748,In_1456,In_915);
or U2749 (N_2749,In_272,In_576);
nand U2750 (N_2750,In_390,In_1040);
nor U2751 (N_2751,In_1343,In_432);
nand U2752 (N_2752,In_1478,In_121);
xor U2753 (N_2753,In_1240,In_1133);
or U2754 (N_2754,In_1099,In_1200);
xor U2755 (N_2755,In_647,In_992);
or U2756 (N_2756,In_1293,In_1413);
nand U2757 (N_2757,In_559,In_1083);
nor U2758 (N_2758,In_419,In_1349);
and U2759 (N_2759,In_457,In_1120);
or U2760 (N_2760,In_1421,In_1096);
nor U2761 (N_2761,In_418,In_1190);
nand U2762 (N_2762,In_630,In_1264);
xor U2763 (N_2763,In_132,In_1134);
and U2764 (N_2764,In_454,In_96);
or U2765 (N_2765,In_433,In_840);
or U2766 (N_2766,In_315,In_90);
nand U2767 (N_2767,In_112,In_89);
or U2768 (N_2768,In_202,In_9);
or U2769 (N_2769,In_1093,In_1247);
or U2770 (N_2770,In_737,In_707);
and U2771 (N_2771,In_414,In_1098);
xor U2772 (N_2772,In_480,In_689);
nor U2773 (N_2773,In_1222,In_1404);
or U2774 (N_2774,In_309,In_618);
nand U2775 (N_2775,In_997,In_392);
and U2776 (N_2776,In_1410,In_1455);
or U2777 (N_2777,In_153,In_642);
or U2778 (N_2778,In_1347,In_1375);
and U2779 (N_2779,In_626,In_1373);
nand U2780 (N_2780,In_325,In_52);
nand U2781 (N_2781,In_175,In_93);
xnor U2782 (N_2782,In_169,In_1036);
nand U2783 (N_2783,In_1073,In_1031);
xor U2784 (N_2784,In_649,In_1064);
nand U2785 (N_2785,In_472,In_991);
nor U2786 (N_2786,In_409,In_1018);
and U2787 (N_2787,In_174,In_752);
or U2788 (N_2788,In_66,In_1206);
nand U2789 (N_2789,In_974,In_1459);
and U2790 (N_2790,In_1450,In_488);
or U2791 (N_2791,In_139,In_35);
or U2792 (N_2792,In_1126,In_1488);
xnor U2793 (N_2793,In_816,In_1040);
and U2794 (N_2794,In_1198,In_932);
and U2795 (N_2795,In_1144,In_1170);
nor U2796 (N_2796,In_237,In_608);
xnor U2797 (N_2797,In_789,In_901);
and U2798 (N_2798,In_675,In_425);
nand U2799 (N_2799,In_1342,In_531);
nand U2800 (N_2800,In_1397,In_1024);
and U2801 (N_2801,In_571,In_1188);
and U2802 (N_2802,In_337,In_1255);
nand U2803 (N_2803,In_1318,In_1462);
nor U2804 (N_2804,In_1369,In_1417);
nor U2805 (N_2805,In_387,In_114);
nor U2806 (N_2806,In_1183,In_1223);
and U2807 (N_2807,In_1175,In_882);
or U2808 (N_2808,In_330,In_705);
nor U2809 (N_2809,In_178,In_64);
nor U2810 (N_2810,In_587,In_529);
nand U2811 (N_2811,In_154,In_304);
nor U2812 (N_2812,In_160,In_896);
and U2813 (N_2813,In_812,In_655);
or U2814 (N_2814,In_247,In_155);
nand U2815 (N_2815,In_348,In_201);
nand U2816 (N_2816,In_1132,In_1297);
or U2817 (N_2817,In_1054,In_611);
nand U2818 (N_2818,In_413,In_1141);
nor U2819 (N_2819,In_138,In_1184);
or U2820 (N_2820,In_1252,In_477);
xor U2821 (N_2821,In_1273,In_1175);
or U2822 (N_2822,In_367,In_897);
nand U2823 (N_2823,In_753,In_1280);
and U2824 (N_2824,In_1327,In_480);
or U2825 (N_2825,In_1426,In_990);
or U2826 (N_2826,In_367,In_513);
nand U2827 (N_2827,In_227,In_457);
and U2828 (N_2828,In_786,In_1311);
and U2829 (N_2829,In_185,In_1384);
nand U2830 (N_2830,In_944,In_186);
nor U2831 (N_2831,In_1197,In_1449);
nand U2832 (N_2832,In_261,In_896);
nand U2833 (N_2833,In_950,In_251);
nand U2834 (N_2834,In_500,In_53);
or U2835 (N_2835,In_1138,In_760);
and U2836 (N_2836,In_1091,In_1348);
nor U2837 (N_2837,In_154,In_1447);
or U2838 (N_2838,In_524,In_121);
nand U2839 (N_2839,In_951,In_732);
and U2840 (N_2840,In_1315,In_302);
xnor U2841 (N_2841,In_736,In_1212);
and U2842 (N_2842,In_1172,In_1090);
or U2843 (N_2843,In_1090,In_758);
nand U2844 (N_2844,In_1343,In_68);
or U2845 (N_2845,In_1150,In_354);
nor U2846 (N_2846,In_944,In_75);
or U2847 (N_2847,In_1489,In_1407);
nor U2848 (N_2848,In_1197,In_922);
nand U2849 (N_2849,In_301,In_1072);
and U2850 (N_2850,In_446,In_1003);
and U2851 (N_2851,In_361,In_709);
or U2852 (N_2852,In_1208,In_1093);
or U2853 (N_2853,In_170,In_686);
and U2854 (N_2854,In_128,In_966);
and U2855 (N_2855,In_947,In_1316);
or U2856 (N_2856,In_1328,In_1339);
nor U2857 (N_2857,In_1039,In_761);
xor U2858 (N_2858,In_56,In_1232);
and U2859 (N_2859,In_164,In_894);
and U2860 (N_2860,In_903,In_808);
and U2861 (N_2861,In_1442,In_1185);
nand U2862 (N_2862,In_930,In_176);
nor U2863 (N_2863,In_878,In_590);
or U2864 (N_2864,In_13,In_606);
nand U2865 (N_2865,In_1358,In_1126);
nor U2866 (N_2866,In_432,In_1379);
and U2867 (N_2867,In_302,In_1433);
nor U2868 (N_2868,In_622,In_906);
or U2869 (N_2869,In_933,In_1051);
nand U2870 (N_2870,In_929,In_556);
nor U2871 (N_2871,In_644,In_325);
nor U2872 (N_2872,In_1381,In_1205);
nand U2873 (N_2873,In_1261,In_1106);
or U2874 (N_2874,In_523,In_1146);
xnor U2875 (N_2875,In_1343,In_1049);
nor U2876 (N_2876,In_366,In_1180);
or U2877 (N_2877,In_1260,In_722);
and U2878 (N_2878,In_1374,In_363);
or U2879 (N_2879,In_124,In_1136);
nor U2880 (N_2880,In_430,In_704);
nor U2881 (N_2881,In_787,In_135);
nor U2882 (N_2882,In_1400,In_1280);
or U2883 (N_2883,In_921,In_522);
nand U2884 (N_2884,In_533,In_1061);
and U2885 (N_2885,In_741,In_623);
nand U2886 (N_2886,In_892,In_1367);
nand U2887 (N_2887,In_21,In_860);
and U2888 (N_2888,In_771,In_1387);
nor U2889 (N_2889,In_210,In_1472);
nand U2890 (N_2890,In_774,In_854);
xor U2891 (N_2891,In_1205,In_429);
or U2892 (N_2892,In_193,In_266);
nor U2893 (N_2893,In_1022,In_526);
nand U2894 (N_2894,In_695,In_185);
nor U2895 (N_2895,In_1019,In_1246);
or U2896 (N_2896,In_340,In_1436);
nor U2897 (N_2897,In_1309,In_450);
and U2898 (N_2898,In_1310,In_94);
nand U2899 (N_2899,In_1390,In_1240);
and U2900 (N_2900,In_716,In_468);
or U2901 (N_2901,In_1087,In_342);
and U2902 (N_2902,In_1022,In_958);
and U2903 (N_2903,In_1234,In_1265);
or U2904 (N_2904,In_1080,In_1442);
nand U2905 (N_2905,In_564,In_298);
nand U2906 (N_2906,In_770,In_649);
or U2907 (N_2907,In_821,In_290);
nor U2908 (N_2908,In_490,In_220);
and U2909 (N_2909,In_543,In_709);
nand U2910 (N_2910,In_973,In_884);
or U2911 (N_2911,In_1233,In_535);
nand U2912 (N_2912,In_1023,In_1354);
nand U2913 (N_2913,In_802,In_868);
nor U2914 (N_2914,In_1159,In_516);
nand U2915 (N_2915,In_1046,In_767);
nor U2916 (N_2916,In_185,In_956);
or U2917 (N_2917,In_1159,In_1139);
and U2918 (N_2918,In_282,In_1041);
nor U2919 (N_2919,In_718,In_226);
or U2920 (N_2920,In_1382,In_934);
and U2921 (N_2921,In_478,In_1244);
nor U2922 (N_2922,In_1014,In_1197);
and U2923 (N_2923,In_847,In_912);
or U2924 (N_2924,In_1206,In_705);
or U2925 (N_2925,In_446,In_1273);
or U2926 (N_2926,In_1355,In_1232);
or U2927 (N_2927,In_250,In_336);
xor U2928 (N_2928,In_1190,In_342);
nor U2929 (N_2929,In_550,In_12);
nand U2930 (N_2930,In_1009,In_848);
nand U2931 (N_2931,In_1035,In_1314);
nor U2932 (N_2932,In_515,In_694);
xor U2933 (N_2933,In_722,In_533);
nand U2934 (N_2934,In_484,In_979);
nor U2935 (N_2935,In_297,In_303);
or U2936 (N_2936,In_1318,In_417);
nor U2937 (N_2937,In_1187,In_531);
or U2938 (N_2938,In_758,In_164);
xnor U2939 (N_2939,In_177,In_860);
nor U2940 (N_2940,In_802,In_147);
or U2941 (N_2941,In_736,In_1004);
nor U2942 (N_2942,In_1259,In_172);
xor U2943 (N_2943,In_291,In_917);
and U2944 (N_2944,In_1028,In_799);
nand U2945 (N_2945,In_153,In_943);
and U2946 (N_2946,In_758,In_296);
and U2947 (N_2947,In_692,In_469);
xnor U2948 (N_2948,In_1274,In_1015);
nor U2949 (N_2949,In_1050,In_633);
or U2950 (N_2950,In_988,In_1190);
or U2951 (N_2951,In_1404,In_332);
and U2952 (N_2952,In_947,In_1037);
nor U2953 (N_2953,In_476,In_374);
and U2954 (N_2954,In_627,In_10);
and U2955 (N_2955,In_444,In_1483);
and U2956 (N_2956,In_263,In_689);
nand U2957 (N_2957,In_734,In_1457);
nor U2958 (N_2958,In_691,In_1270);
nor U2959 (N_2959,In_965,In_544);
xor U2960 (N_2960,In_235,In_188);
and U2961 (N_2961,In_1131,In_1497);
nand U2962 (N_2962,In_800,In_1298);
and U2963 (N_2963,In_565,In_26);
and U2964 (N_2964,In_1320,In_885);
nand U2965 (N_2965,In_220,In_304);
nor U2966 (N_2966,In_1406,In_359);
nand U2967 (N_2967,In_458,In_1143);
nor U2968 (N_2968,In_467,In_627);
nor U2969 (N_2969,In_1186,In_88);
nor U2970 (N_2970,In_609,In_993);
nand U2971 (N_2971,In_1203,In_375);
nand U2972 (N_2972,In_869,In_868);
xor U2973 (N_2973,In_715,In_603);
or U2974 (N_2974,In_90,In_1043);
or U2975 (N_2975,In_867,In_363);
xnor U2976 (N_2976,In_1445,In_148);
and U2977 (N_2977,In_1476,In_593);
or U2978 (N_2978,In_902,In_80);
nor U2979 (N_2979,In_1101,In_28);
and U2980 (N_2980,In_504,In_1236);
nor U2981 (N_2981,In_659,In_612);
nor U2982 (N_2982,In_626,In_377);
nor U2983 (N_2983,In_329,In_1259);
or U2984 (N_2984,In_677,In_585);
and U2985 (N_2985,In_1170,In_1461);
and U2986 (N_2986,In_996,In_1358);
nand U2987 (N_2987,In_603,In_928);
and U2988 (N_2988,In_868,In_1306);
and U2989 (N_2989,In_737,In_340);
nor U2990 (N_2990,In_1174,In_653);
or U2991 (N_2991,In_675,In_1483);
nand U2992 (N_2992,In_1293,In_1393);
or U2993 (N_2993,In_637,In_270);
or U2994 (N_2994,In_821,In_423);
or U2995 (N_2995,In_767,In_1400);
and U2996 (N_2996,In_1372,In_543);
nor U2997 (N_2997,In_109,In_633);
nand U2998 (N_2998,In_382,In_1106);
nand U2999 (N_2999,In_111,In_69);
or U3000 (N_3000,N_2898,N_289);
xnor U3001 (N_3001,N_361,N_2836);
nor U3002 (N_3002,N_169,N_2246);
or U3003 (N_3003,N_399,N_1954);
nand U3004 (N_3004,N_1583,N_2143);
and U3005 (N_3005,N_1675,N_1771);
or U3006 (N_3006,N_731,N_852);
nor U3007 (N_3007,N_373,N_1429);
nor U3008 (N_3008,N_796,N_1461);
nand U3009 (N_3009,N_1054,N_2659);
nand U3010 (N_3010,N_1229,N_52);
nor U3011 (N_3011,N_2779,N_1252);
or U3012 (N_3012,N_131,N_204);
nand U3013 (N_3013,N_1802,N_1581);
xnor U3014 (N_3014,N_2690,N_2451);
nor U3015 (N_3015,N_1761,N_700);
xnor U3016 (N_3016,N_2834,N_1957);
or U3017 (N_3017,N_2676,N_1361);
nand U3018 (N_3018,N_759,N_819);
nor U3019 (N_3019,N_19,N_1371);
nand U3020 (N_3020,N_2635,N_2383);
nor U3021 (N_3021,N_1791,N_562);
nand U3022 (N_3022,N_133,N_83);
and U3023 (N_3023,N_2430,N_1166);
and U3024 (N_3024,N_1551,N_2101);
and U3025 (N_3025,N_942,N_2213);
and U3026 (N_3026,N_2996,N_2128);
or U3027 (N_3027,N_2726,N_839);
or U3028 (N_3028,N_32,N_2298);
or U3029 (N_3029,N_1159,N_733);
or U3030 (N_3030,N_1576,N_111);
and U3031 (N_3031,N_2619,N_246);
and U3032 (N_3032,N_1622,N_2134);
nand U3033 (N_3033,N_656,N_1860);
or U3034 (N_3034,N_1413,N_1094);
xor U3035 (N_3035,N_2950,N_481);
nand U3036 (N_3036,N_2174,N_2548);
and U3037 (N_3037,N_1187,N_647);
or U3038 (N_3038,N_1378,N_2867);
nand U3039 (N_3039,N_2640,N_1731);
nand U3040 (N_3040,N_1018,N_2400);
and U3041 (N_3041,N_2471,N_1686);
nand U3042 (N_3042,N_87,N_846);
and U3043 (N_3043,N_322,N_1818);
nor U3044 (N_3044,N_869,N_2569);
nand U3045 (N_3045,N_2670,N_371);
nor U3046 (N_3046,N_150,N_2324);
or U3047 (N_3047,N_2194,N_777);
or U3048 (N_3048,N_1082,N_1477);
or U3049 (N_3049,N_2654,N_2853);
nand U3050 (N_3050,N_2695,N_2012);
nor U3051 (N_3051,N_1634,N_2292);
nand U3052 (N_3052,N_2064,N_1584);
nand U3053 (N_3053,N_884,N_2010);
nand U3054 (N_3054,N_1379,N_2166);
nand U3055 (N_3055,N_2500,N_2328);
nand U3056 (N_3056,N_2508,N_2109);
and U3057 (N_3057,N_2335,N_2436);
nand U3058 (N_3058,N_383,N_1782);
nor U3059 (N_3059,N_2655,N_27);
nor U3060 (N_3060,N_527,N_2503);
nor U3061 (N_3061,N_734,N_422);
nor U3062 (N_3062,N_1036,N_2389);
nor U3063 (N_3063,N_1130,N_1568);
xnor U3064 (N_3064,N_2744,N_1198);
and U3065 (N_3065,N_1876,N_1455);
and U3066 (N_3066,N_2602,N_1918);
and U3067 (N_3067,N_482,N_2790);
nor U3068 (N_3068,N_2320,N_1299);
xnor U3069 (N_3069,N_1964,N_646);
and U3070 (N_3070,N_924,N_202);
or U3071 (N_3071,N_2886,N_2939);
nor U3072 (N_3072,N_7,N_2050);
nand U3073 (N_3073,N_735,N_847);
xor U3074 (N_3074,N_2276,N_1640);
and U3075 (N_3075,N_597,N_2986);
or U3076 (N_3076,N_959,N_2678);
and U3077 (N_3077,N_2582,N_1269);
nor U3078 (N_3078,N_2259,N_1137);
nor U3079 (N_3079,N_2813,N_854);
or U3080 (N_3080,N_196,N_2756);
or U3081 (N_3081,N_2881,N_521);
nand U3082 (N_3082,N_1631,N_2578);
or U3083 (N_3083,N_761,N_2282);
or U3084 (N_3084,N_2597,N_2700);
nand U3085 (N_3085,N_2421,N_2423);
and U3086 (N_3086,N_2065,N_485);
or U3087 (N_3087,N_214,N_1750);
and U3088 (N_3088,N_1365,N_312);
nor U3089 (N_3089,N_1265,N_1146);
or U3090 (N_3090,N_2888,N_1796);
and U3091 (N_3091,N_2146,N_2802);
or U3092 (N_3092,N_44,N_810);
nor U3093 (N_3093,N_1523,N_126);
nor U3094 (N_3094,N_2549,N_1868);
nand U3095 (N_3095,N_222,N_327);
or U3096 (N_3096,N_2752,N_2434);
nor U3097 (N_3097,N_2971,N_1110);
and U3098 (N_3098,N_2793,N_1266);
nand U3099 (N_3099,N_14,N_1104);
and U3100 (N_3100,N_1232,N_66);
nor U3101 (N_3101,N_1904,N_173);
or U3102 (N_3102,N_1138,N_424);
and U3103 (N_3103,N_79,N_2369);
nand U3104 (N_3104,N_1960,N_108);
nand U3105 (N_3105,N_1069,N_2673);
or U3106 (N_3106,N_2804,N_139);
nor U3107 (N_3107,N_2754,N_1778);
xnor U3108 (N_3108,N_1692,N_1925);
xor U3109 (N_3109,N_2186,N_2225);
nand U3110 (N_3110,N_1617,N_2869);
nand U3111 (N_3111,N_895,N_1126);
nand U3112 (N_3112,N_1784,N_532);
nor U3113 (N_3113,N_1596,N_2532);
nand U3114 (N_3114,N_353,N_2788);
nor U3115 (N_3115,N_99,N_51);
nand U3116 (N_3116,N_1204,N_1698);
xnor U3117 (N_3117,N_711,N_1812);
nor U3118 (N_3118,N_189,N_2585);
and U3119 (N_3119,N_1518,N_314);
and U3120 (N_3120,N_364,N_2505);
nor U3121 (N_3121,N_2830,N_929);
xnor U3122 (N_3122,N_2658,N_1517);
or U3123 (N_3123,N_467,N_1522);
or U3124 (N_3124,N_2543,N_2637);
nor U3125 (N_3125,N_750,N_1);
nor U3126 (N_3126,N_720,N_1820);
or U3127 (N_3127,N_511,N_1873);
and U3128 (N_3128,N_2047,N_1756);
and U3129 (N_3129,N_2171,N_2835);
or U3130 (N_3130,N_1096,N_1380);
nand U3131 (N_3131,N_1403,N_2590);
nand U3132 (N_3132,N_2734,N_1079);
and U3133 (N_3133,N_1641,N_661);
xor U3134 (N_3134,N_1907,N_1469);
or U3135 (N_3135,N_2284,N_1383);
nor U3136 (N_3136,N_2561,N_1453);
or U3137 (N_3137,N_1884,N_1608);
nand U3138 (N_3138,N_2714,N_881);
xor U3139 (N_3139,N_1277,N_1938);
or U3140 (N_3140,N_172,N_198);
nor U3141 (N_3141,N_1047,N_1373);
nand U3142 (N_3142,N_1430,N_2475);
and U3143 (N_3143,N_2182,N_2237);
nor U3144 (N_3144,N_2603,N_1512);
nand U3145 (N_3145,N_678,N_1890);
and U3146 (N_3146,N_542,N_1537);
or U3147 (N_3147,N_872,N_1892);
and U3148 (N_3148,N_1670,N_1111);
xnor U3149 (N_3149,N_69,N_226);
and U3150 (N_3150,N_821,N_2220);
and U3151 (N_3151,N_441,N_830);
and U3152 (N_3152,N_921,N_2405);
and U3153 (N_3153,N_2795,N_4);
and U3154 (N_3154,N_698,N_402);
nand U3155 (N_3155,N_1226,N_899);
and U3156 (N_3156,N_2008,N_1411);
xnor U3157 (N_3157,N_1943,N_59);
nand U3158 (N_3158,N_2534,N_2078);
and U3159 (N_3159,N_2643,N_2183);
xnor U3160 (N_3160,N_1899,N_1118);
xnor U3161 (N_3161,N_1959,N_119);
xor U3162 (N_3162,N_2859,N_2583);
nor U3163 (N_3163,N_2350,N_2621);
or U3164 (N_3164,N_2469,N_2573);
nor U3165 (N_3165,N_1627,N_1149);
or U3166 (N_3166,N_291,N_1431);
nand U3167 (N_3167,N_2222,N_2392);
nand U3168 (N_3168,N_102,N_706);
or U3169 (N_3169,N_1835,N_2862);
xor U3170 (N_3170,N_128,N_1224);
or U3171 (N_3171,N_339,N_1950);
or U3172 (N_3172,N_2223,N_1789);
or U3173 (N_3173,N_2185,N_1292);
and U3174 (N_3174,N_2150,N_982);
nand U3175 (N_3175,N_2336,N_181);
or U3176 (N_3176,N_55,N_822);
nor U3177 (N_3177,N_2656,N_1081);
or U3178 (N_3178,N_2495,N_1356);
xor U3179 (N_3179,N_2825,N_1471);
xor U3180 (N_3180,N_1632,N_1560);
and U3181 (N_3181,N_265,N_2079);
nand U3182 (N_3182,N_394,N_815);
and U3183 (N_3183,N_687,N_2506);
nand U3184 (N_3184,N_638,N_376);
nor U3185 (N_3185,N_1780,N_785);
and U3186 (N_3186,N_1309,N_89);
or U3187 (N_3187,N_1170,N_1473);
nor U3188 (N_3188,N_2168,N_2196);
or U3189 (N_3189,N_1769,N_2059);
nand U3190 (N_3190,N_2646,N_2488);
nand U3191 (N_3191,N_1688,N_671);
nor U3192 (N_3192,N_874,N_2195);
and U3193 (N_3193,N_776,N_2293);
nand U3194 (N_3194,N_271,N_1434);
nor U3195 (N_3195,N_2342,N_753);
nor U3196 (N_3196,N_1690,N_231);
or U3197 (N_3197,N_1474,N_875);
or U3198 (N_3198,N_2786,N_2021);
xor U3199 (N_3199,N_2896,N_2904);
nand U3200 (N_3200,N_1019,N_1445);
and U3201 (N_3201,N_2753,N_2227);
nor U3202 (N_3202,N_2990,N_1157);
xor U3203 (N_3203,N_2016,N_2340);
or U3204 (N_3204,N_857,N_1150);
xor U3205 (N_3205,N_1888,N_1586);
nor U3206 (N_3206,N_1107,N_1412);
or U3207 (N_3207,N_2061,N_1003);
nand U3208 (N_3208,N_2466,N_1303);
or U3209 (N_3209,N_1946,N_1867);
nand U3210 (N_3210,N_1822,N_1462);
nand U3211 (N_3211,N_1452,N_1020);
nor U3212 (N_3212,N_333,N_2188);
xnor U3213 (N_3213,N_405,N_2901);
and U3214 (N_3214,N_516,N_1768);
nand U3215 (N_3215,N_2210,N_205);
or U3216 (N_3216,N_1465,N_2147);
nor U3217 (N_3217,N_1311,N_252);
and U3218 (N_3218,N_971,N_2450);
nand U3219 (N_3219,N_2811,N_2402);
nand U3220 (N_3220,N_555,N_630);
or U3221 (N_3221,N_1405,N_2628);
nor U3222 (N_3222,N_667,N_1664);
or U3223 (N_3223,N_1031,N_166);
and U3224 (N_3224,N_417,N_596);
xnor U3225 (N_3225,N_805,N_911);
nand U3226 (N_3226,N_756,N_1597);
nand U3227 (N_3227,N_1382,N_2837);
and U3228 (N_3228,N_1760,N_9);
nor U3229 (N_3229,N_1005,N_1589);
or U3230 (N_3230,N_2663,N_2133);
xnor U3231 (N_3231,N_790,N_581);
nor U3232 (N_3232,N_285,N_378);
and U3233 (N_3233,N_2262,N_451);
and U3234 (N_3234,N_2002,N_154);
or U3235 (N_3235,N_1209,N_744);
or U3236 (N_3236,N_628,N_195);
nor U3237 (N_3237,N_2040,N_2018);
nor U3238 (N_3238,N_1933,N_1024);
and U3239 (N_3239,N_709,N_1934);
nor U3240 (N_3240,N_2415,N_325);
nand U3241 (N_3241,N_640,N_966);
or U3242 (N_3242,N_2121,N_174);
nand U3243 (N_3243,N_1416,N_2544);
and U3244 (N_3244,N_918,N_2871);
and U3245 (N_3245,N_2992,N_1994);
nor U3246 (N_3246,N_786,N_273);
and U3247 (N_3247,N_2317,N_307);
nor U3248 (N_3248,N_389,N_122);
or U3249 (N_3249,N_2445,N_1499);
or U3250 (N_3250,N_2954,N_2374);
nand U3251 (N_3251,N_2080,N_1359);
and U3252 (N_3252,N_2420,N_1786);
and U3253 (N_3253,N_2562,N_1273);
nand U3254 (N_3254,N_1353,N_2789);
and U3255 (N_3255,N_2189,N_2920);
and U3256 (N_3256,N_943,N_685);
xnor U3257 (N_3257,N_1563,N_1775);
and U3258 (N_3258,N_1603,N_100);
nand U3259 (N_3259,N_103,N_2085);
or U3260 (N_3260,N_680,N_136);
nor U3261 (N_3261,N_1801,N_1655);
and U3262 (N_3262,N_2232,N_2046);
nor U3263 (N_3263,N_2709,N_2748);
nor U3264 (N_3264,N_2907,N_1004);
and U3265 (N_3265,N_2899,N_1975);
and U3266 (N_3266,N_2941,N_2448);
or U3267 (N_3267,N_2806,N_1279);
nor U3268 (N_3268,N_1553,N_1259);
and U3269 (N_3269,N_639,N_679);
nand U3270 (N_3270,N_708,N_86);
and U3271 (N_3271,N_845,N_1401);
xor U3272 (N_3272,N_829,N_2208);
xnor U3273 (N_3273,N_1013,N_922);
or U3274 (N_3274,N_408,N_401);
or U3275 (N_3275,N_2918,N_835);
nor U3276 (N_3276,N_2615,N_2666);
and U3277 (N_3277,N_1857,N_856);
nand U3278 (N_3278,N_1438,N_989);
xor U3279 (N_3279,N_374,N_2257);
nor U3280 (N_3280,N_2801,N_358);
or U3281 (N_3281,N_2791,N_1202);
nand U3282 (N_3282,N_876,N_2279);
and U3283 (N_3283,N_572,N_904);
or U3284 (N_3284,N_2880,N_2359);
and U3285 (N_3285,N_1425,N_1908);
and U3286 (N_3286,N_283,N_2604);
nor U3287 (N_3287,N_2401,N_1949);
nor U3288 (N_3288,N_1962,N_964);
nor U3289 (N_3289,N_1487,N_2672);
nor U3290 (N_3290,N_331,N_3);
and U3291 (N_3291,N_1856,N_2936);
or U3292 (N_3292,N_2798,N_2140);
xor U3293 (N_3293,N_1263,N_2349);
nor U3294 (N_3294,N_2942,N_1881);
and U3295 (N_3295,N_2390,N_2281);
nor U3296 (N_3296,N_1703,N_1637);
nand U3297 (N_3297,N_2757,N_2381);
xor U3298 (N_3298,N_676,N_728);
xor U3299 (N_3299,N_2647,N_984);
nand U3300 (N_3300,N_2775,N_57);
or U3301 (N_3301,N_2139,N_2152);
or U3302 (N_3302,N_2538,N_2158);
xnor U3303 (N_3303,N_972,N_1776);
nand U3304 (N_3304,N_2641,N_1956);
or U3305 (N_3305,N_1552,N_1321);
and U3306 (N_3306,N_1395,N_2119);
nor U3307 (N_3307,N_2125,N_2329);
xnor U3308 (N_3308,N_2073,N_2872);
or U3309 (N_3309,N_192,N_1101);
or U3310 (N_3310,N_2832,N_2600);
nor U3311 (N_3311,N_213,N_797);
and U3312 (N_3312,N_293,N_1239);
and U3313 (N_3313,N_1351,N_18);
nor U3314 (N_3314,N_2129,N_336);
nand U3315 (N_3315,N_575,N_1814);
and U3316 (N_3316,N_2307,N_945);
or U3317 (N_3317,N_1996,N_1609);
and U3318 (N_3318,N_1056,N_120);
and U3319 (N_3319,N_326,N_266);
and U3320 (N_3320,N_1065,N_2737);
nor U3321 (N_3321,N_1807,N_1175);
nand U3322 (N_3322,N_2787,N_831);
and U3323 (N_3323,N_2393,N_1642);
xnor U3324 (N_3324,N_1834,N_428);
nor U3325 (N_3325,N_2566,N_2740);
nor U3326 (N_3326,N_563,N_1725);
nor U3327 (N_3327,N_690,N_2706);
nor U3328 (N_3328,N_20,N_2919);
nand U3329 (N_3329,N_443,N_1720);
or U3330 (N_3330,N_80,N_1532);
or U3331 (N_3331,N_2060,N_249);
or U3332 (N_3332,N_863,N_2197);
nand U3333 (N_3333,N_1183,N_2481);
and U3334 (N_3334,N_1852,N_694);
xor U3335 (N_3335,N_1457,N_1237);
and U3336 (N_3336,N_324,N_2);
and U3337 (N_3337,N_2441,N_10);
nand U3338 (N_3338,N_1488,N_2226);
or U3339 (N_3339,N_520,N_1932);
nand U3340 (N_3340,N_2122,N_2153);
xnor U3341 (N_3341,N_2325,N_2199);
and U3342 (N_3342,N_1489,N_435);
and U3343 (N_3343,N_159,N_2945);
nand U3344 (N_3344,N_741,N_560);
nand U3345 (N_3345,N_223,N_2033);
or U3346 (N_3346,N_2090,N_557);
nor U3347 (N_3347,N_2092,N_1143);
nand U3348 (N_3348,N_2989,N_1008);
or U3349 (N_3349,N_714,N_2537);
nor U3350 (N_3350,N_2531,N_1386);
and U3351 (N_3351,N_632,N_2219);
nor U3352 (N_3352,N_689,N_592);
and U3353 (N_3353,N_2413,N_270);
xor U3354 (N_3354,N_2498,N_2493);
nor U3355 (N_3355,N_470,N_2960);
nor U3356 (N_3356,N_788,N_2854);
xnor U3357 (N_3357,N_1078,N_968);
nor U3358 (N_3358,N_713,N_2499);
or U3359 (N_3359,N_2574,N_299);
and U3360 (N_3360,N_1774,N_2053);
nand U3361 (N_3361,N_431,N_2394);
nand U3362 (N_3362,N_682,N_1038);
or U3363 (N_3363,N_1506,N_965);
or U3364 (N_3364,N_2269,N_1555);
nand U3365 (N_3365,N_323,N_188);
nor U3366 (N_3366,N_828,N_1828);
or U3367 (N_3367,N_660,N_93);
nor U3368 (N_3368,N_721,N_1995);
xor U3369 (N_3369,N_1805,N_2797);
nand U3370 (N_3370,N_1449,N_276);
and U3371 (N_3371,N_2003,N_1712);
nand U3372 (N_3372,N_2444,N_2912);
nand U3373 (N_3373,N_263,N_1976);
nor U3374 (N_3374,N_877,N_2844);
nand U3375 (N_3375,N_739,N_2617);
nand U3376 (N_3376,N_937,N_110);
and U3377 (N_3377,N_1220,N_356);
nand U3378 (N_3378,N_2925,N_2418);
nand U3379 (N_3379,N_200,N_1501);
nand U3380 (N_3380,N_2684,N_1313);
and U3381 (N_3381,N_1119,N_433);
xor U3382 (N_3382,N_701,N_2686);
and U3383 (N_3383,N_920,N_1635);
and U3384 (N_3384,N_382,N_794);
and U3385 (N_3385,N_1402,N_2831);
and U3386 (N_3386,N_1582,N_2841);
xor U3387 (N_3387,N_1875,N_1257);
or U3388 (N_3388,N_981,N_2652);
nand U3389 (N_3389,N_1192,N_1874);
or U3390 (N_3390,N_1677,N_2360);
nand U3391 (N_3391,N_1646,N_1314);
xnor U3392 (N_3392,N_2967,N_1973);
and U3393 (N_3393,N_343,N_502);
and U3394 (N_3394,N_1645,N_880);
or U3395 (N_3395,N_1838,N_1441);
nand U3396 (N_3396,N_658,N_2978);
and U3397 (N_3397,N_1320,N_490);
or U3398 (N_3398,N_2198,N_2042);
and U3399 (N_3399,N_269,N_344);
nand U3400 (N_3400,N_2395,N_454);
nor U3401 (N_3401,N_951,N_107);
or U3402 (N_3402,N_2963,N_1840);
nand U3403 (N_3403,N_1729,N_2497);
or U3404 (N_3404,N_1007,N_2368);
nor U3405 (N_3405,N_157,N_760);
nor U3406 (N_3406,N_1034,N_894);
nor U3407 (N_3407,N_2765,N_1979);
nand U3408 (N_3408,N_1318,N_864);
nor U3409 (N_3409,N_235,N_729);
or U3410 (N_3410,N_1590,N_915);
nand U3411 (N_3411,N_509,N_1951);
xnor U3412 (N_3412,N_2406,N_2792);
xnor U3413 (N_3413,N_1194,N_611);
nand U3414 (N_3414,N_445,N_180);
and U3415 (N_3415,N_257,N_523);
or U3416 (N_3416,N_2771,N_2345);
nand U3417 (N_3417,N_54,N_2149);
and U3418 (N_3418,N_1666,N_1030);
and U3419 (N_3419,N_2723,N_2034);
nor U3420 (N_3420,N_2275,N_2087);
or U3421 (N_3421,N_2929,N_1606);
nand U3422 (N_3422,N_610,N_472);
or U3423 (N_3423,N_2037,N_97);
and U3424 (N_3424,N_1284,N_2591);
nor U3425 (N_3425,N_2849,N_1837);
and U3426 (N_3426,N_2162,N_812);
xor U3427 (N_3427,N_2234,N_1832);
nor U3428 (N_3428,N_418,N_2738);
xor U3429 (N_3429,N_397,N_1173);
nand U3430 (N_3430,N_2218,N_1495);
nand U3431 (N_3431,N_1375,N_2358);
nand U3432 (N_3432,N_1540,N_2852);
or U3433 (N_3433,N_2411,N_462);
nor U3434 (N_3434,N_1432,N_2427);
nand U3435 (N_3435,N_2554,N_2766);
nand U3436 (N_3436,N_2217,N_295);
nor U3437 (N_3437,N_1508,N_1022);
nand U3438 (N_3438,N_1861,N_140);
xnor U3439 (N_3439,N_987,N_416);
xnor U3440 (N_3440,N_738,N_1562);
nand U3441 (N_3441,N_758,N_2005);
nand U3442 (N_3442,N_953,N_1573);
or U3443 (N_3443,N_2306,N_1671);
and U3444 (N_3444,N_912,N_1121);
and U3445 (N_3445,N_142,N_1058);
nand U3446 (N_3446,N_2961,N_859);
nand U3447 (N_3447,N_294,N_71);
nor U3448 (N_3448,N_2995,N_2823);
nor U3449 (N_3449,N_550,N_2127);
and U3450 (N_3450,N_2523,N_1390);
xor U3451 (N_3451,N_2557,N_221);
or U3452 (N_3452,N_2386,N_994);
or U3453 (N_3453,N_2860,N_691);
xnor U3454 (N_3454,N_1307,N_1737);
and U3455 (N_3455,N_840,N_199);
nand U3456 (N_3456,N_407,N_2161);
xor U3457 (N_3457,N_1792,N_2858);
and U3458 (N_3458,N_1850,N_64);
and U3459 (N_3459,N_1798,N_2202);
nor U3460 (N_3460,N_2327,N_1733);
xnor U3461 (N_3461,N_260,N_2482);
and U3462 (N_3462,N_2951,N_2568);
nor U3463 (N_3463,N_1944,N_2058);
xor U3464 (N_3464,N_537,N_1804);
nor U3465 (N_3465,N_1577,N_747);
or U3466 (N_3466,N_1913,N_2045);
and U3467 (N_3467,N_2755,N_1859);
xnor U3468 (N_3468,N_732,N_348);
and U3469 (N_3469,N_372,N_2409);
nor U3470 (N_3470,N_2923,N_1542);
nand U3471 (N_3471,N_896,N_2533);
or U3472 (N_3472,N_2843,N_2593);
xor U3473 (N_3473,N_775,N_2252);
nand U3474 (N_3474,N_2922,N_1770);
nor U3475 (N_3475,N_1358,N_1485);
and U3476 (N_3476,N_156,N_392);
nand U3477 (N_3477,N_1345,N_1773);
and U3478 (N_3478,N_1526,N_2464);
xnor U3479 (N_3479,N_352,N_1088);
and U3480 (N_3480,N_2746,N_2052);
and U3481 (N_3481,N_2253,N_1335);
nor U3482 (N_3482,N_564,N_1463);
or U3483 (N_3483,N_185,N_1135);
or U3484 (N_3484,N_2135,N_1855);
xnor U3485 (N_3485,N_673,N_1963);
or U3486 (N_3486,N_106,N_1601);
nor U3487 (N_3487,N_2560,N_1765);
and U3488 (N_3488,N_1419,N_187);
or U3489 (N_3489,N_2370,N_2728);
nor U3490 (N_3490,N_1529,N_2838);
nand U3491 (N_3491,N_2577,N_2627);
nand U3492 (N_3492,N_2710,N_838);
and U3493 (N_3493,N_1258,N_385);
nor U3494 (N_3494,N_1754,N_1988);
xor U3495 (N_3495,N_1986,N_2962);
and U3496 (N_3496,N_146,N_1743);
nand U3497 (N_3497,N_704,N_2030);
nor U3498 (N_3498,N_1710,N_2887);
nand U3499 (N_3499,N_2072,N_1283);
or U3500 (N_3500,N_580,N_1521);
nor U3501 (N_3501,N_1695,N_1514);
or U3502 (N_3502,N_2081,N_1657);
nor U3503 (N_3503,N_2879,N_1217);
nor U3504 (N_3504,N_1851,N_2776);
and U3505 (N_3505,N_2366,N_388);
xnor U3506 (N_3506,N_791,N_566);
nand U3507 (N_3507,N_1447,N_1251);
or U3508 (N_3508,N_594,N_137);
nand U3509 (N_3509,N_2476,N_740);
nor U3510 (N_3510,N_447,N_2249);
nor U3511 (N_3511,N_1153,N_1315);
xnor U3512 (N_3512,N_1684,N_193);
nand U3513 (N_3513,N_1227,N_936);
nand U3514 (N_3514,N_1997,N_1682);
and U3515 (N_3515,N_1700,N_1559);
nand U3516 (N_3516,N_1410,N_1006);
nor U3517 (N_3517,N_2020,N_1696);
or U3518 (N_3518,N_238,N_1691);
or U3519 (N_3519,N_1060,N_589);
and U3520 (N_3520,N_1140,N_278);
nor U3521 (N_3521,N_251,N_1162);
or U3522 (N_3522,N_403,N_827);
nor U3523 (N_3523,N_225,N_2644);
and U3524 (N_3524,N_1879,N_2172);
or U3525 (N_3525,N_1228,N_2458);
or U3526 (N_3526,N_190,N_316);
or U3527 (N_3527,N_2032,N_947);
nand U3528 (N_3528,N_1528,N_917);
or U3529 (N_3529,N_783,N_0);
xnor U3530 (N_3530,N_1628,N_2535);
or U3531 (N_3531,N_547,N_2772);
nand U3532 (N_3532,N_1970,N_1923);
and U3533 (N_3533,N_1978,N_1945);
or U3534 (N_3534,N_1163,N_889);
nand U3535 (N_3535,N_1880,N_2067);
nand U3536 (N_3536,N_306,N_404);
nand U3537 (N_3537,N_387,N_1511);
or U3538 (N_3538,N_1530,N_1539);
nor U3539 (N_3539,N_147,N_2556);
xor U3540 (N_3540,N_524,N_2006);
xnor U3541 (N_3541,N_1824,N_2283);
nor U3542 (N_3542,N_124,N_2680);
and U3543 (N_3543,N_1811,N_280);
or U3544 (N_3544,N_2618,N_2868);
or U3545 (N_3545,N_662,N_1249);
or U3546 (N_3546,N_500,N_579);
or U3547 (N_3547,N_642,N_1316);
nand U3548 (N_3548,N_825,N_1293);
or U3549 (N_3549,N_568,N_2541);
nor U3550 (N_3550,N_1993,N_218);
or U3551 (N_3551,N_2759,N_1862);
nor U3552 (N_3552,N_1337,N_2611);
xnor U3553 (N_3553,N_816,N_1406);
and U3554 (N_3554,N_368,N_300);
nand U3555 (N_3555,N_1721,N_923);
nand U3556 (N_3556,N_2391,N_396);
and U3557 (N_3557,N_1866,N_2993);
or U3558 (N_3558,N_2850,N_2935);
nor U3559 (N_3559,N_2367,N_2552);
or U3560 (N_3560,N_2976,N_540);
and U3561 (N_3561,N_1484,N_1600);
nor U3562 (N_3562,N_2312,N_1830);
nand U3563 (N_3563,N_2988,N_2595);
nor U3564 (N_3564,N_1123,N_2302);
and U3565 (N_3565,N_807,N_1052);
xnor U3566 (N_3566,N_2522,N_234);
nand U3567 (N_3567,N_2422,N_2014);
and U3568 (N_3568,N_478,N_1362);
nor U3569 (N_3569,N_2808,N_1678);
nand U3570 (N_3570,N_134,N_461);
nor U3571 (N_3571,N_1388,N_1909);
nor U3572 (N_3572,N_2169,N_1254);
and U3573 (N_3573,N_2657,N_897);
and U3574 (N_3574,N_2818,N_2536);
or U3575 (N_3575,N_1400,N_224);
nand U3576 (N_3576,N_1387,N_1887);
or U3577 (N_3577,N_2287,N_2446);
nand U3578 (N_3578,N_939,N_230);
xor U3579 (N_3579,N_2979,N_1057);
nand U3580 (N_3580,N_2289,N_1706);
nor U3581 (N_3581,N_1077,N_2623);
or U3582 (N_3582,N_1207,N_2118);
nor U3583 (N_3583,N_1418,N_1225);
nand U3584 (N_3584,N_2187,N_1360);
nor U3585 (N_3585,N_2530,N_1290);
or U3586 (N_3586,N_2510,N_535);
nor U3587 (N_3587,N_2846,N_1399);
or U3588 (N_3588,N_2236,N_2731);
and U3589 (N_3589,N_553,N_2084);
and U3590 (N_3590,N_2665,N_2699);
nor U3591 (N_3591,N_1865,N_941);
nor U3592 (N_3592,N_1442,N_2780);
or U3593 (N_3593,N_2473,N_2364);
and U3594 (N_3594,N_1165,N_8);
and U3595 (N_3595,N_891,N_1492);
nand U3596 (N_3596,N_2201,N_1347);
nor U3597 (N_3597,N_1342,N_2460);
or U3598 (N_3598,N_2952,N_1294);
xnor U3599 (N_3599,N_1547,N_1940);
nand U3600 (N_3600,N_2586,N_2035);
nand U3601 (N_3601,N_2958,N_1730);
or U3602 (N_3602,N_552,N_1714);
or U3603 (N_3603,N_530,N_25);
and U3604 (N_3604,N_2751,N_622);
nand U3605 (N_3605,N_724,N_6);
or U3606 (N_3606,N_366,N_1930);
or U3607 (N_3607,N_456,N_1133);
or U3608 (N_3608,N_702,N_1061);
and U3609 (N_3609,N_842,N_850);
xor U3610 (N_3610,N_1305,N_1992);
nor U3611 (N_3611,N_2612,N_2909);
and U3612 (N_3612,N_1331,N_2730);
nand U3613 (N_3613,N_395,N_132);
or U3614 (N_3614,N_1389,N_882);
nand U3615 (N_3615,N_1012,N_303);
and U3616 (N_3616,N_210,N_1667);
nor U3617 (N_3617,N_2428,N_1561);
nor U3618 (N_3618,N_2449,N_2159);
and U3619 (N_3619,N_1203,N_2719);
xnor U3620 (N_3620,N_1687,N_244);
or U3621 (N_3621,N_650,N_1894);
xnor U3622 (N_3622,N_2524,N_77);
nand U3623 (N_3623,N_1800,N_2563);
nand U3624 (N_3624,N_1877,N_1112);
xnor U3625 (N_3625,N_2365,N_2459);
nand U3626 (N_3626,N_161,N_567);
or U3627 (N_3627,N_1039,N_2900);
and U3628 (N_3628,N_1980,N_985);
nand U3629 (N_3629,N_2192,N_1394);
or U3630 (N_3630,N_1724,N_811);
xor U3631 (N_3631,N_179,N_430);
or U3632 (N_3632,N_888,N_2605);
nor U3633 (N_3633,N_2086,N_2204);
nand U3634 (N_3634,N_1736,N_268);
and U3635 (N_3635,N_2540,N_390);
or U3636 (N_3636,N_229,N_26);
xnor U3637 (N_3637,N_2068,N_1417);
xor U3638 (N_3638,N_2036,N_1565);
nand U3639 (N_3639,N_1336,N_1397);
nand U3640 (N_3640,N_2403,N_534);
and U3641 (N_3641,N_2555,N_1167);
and U3642 (N_3642,N_2521,N_2947);
nor U3643 (N_3643,N_696,N_2826);
xor U3644 (N_3644,N_212,N_617);
nand U3645 (N_3645,N_1145,N_604);
nor U3646 (N_3646,N_1242,N_1497);
and U3647 (N_3647,N_991,N_2074);
nand U3648 (N_3648,N_2270,N_420);
nand U3649 (N_3649,N_643,N_1364);
nand U3650 (N_3650,N_1500,N_2991);
and U3651 (N_3651,N_2083,N_1639);
or U3652 (N_3652,N_1989,N_2483);
and U3653 (N_3653,N_778,N_2903);
or U3654 (N_3654,N_1864,N_2144);
nor U3655 (N_3655,N_2847,N_1067);
nand U3656 (N_3656,N_2969,N_2462);
nand U3657 (N_3657,N_2761,N_1593);
and U3658 (N_3658,N_2517,N_2741);
and U3659 (N_3659,N_1424,N_2321);
or U3660 (N_3660,N_561,N_2051);
xnor U3661 (N_3661,N_2994,N_2764);
xnor U3662 (N_3662,N_693,N_967);
and U3663 (N_3663,N_1028,N_2877);
nor U3664 (N_3664,N_1604,N_1470);
or U3665 (N_3665,N_384,N_1393);
or U3666 (N_3666,N_2906,N_518);
or U3667 (N_3667,N_1803,N_554);
nor U3668 (N_3668,N_2981,N_2468);
or U3669 (N_3669,N_22,N_2433);
nor U3670 (N_3670,N_2478,N_298);
and U3671 (N_3671,N_910,N_2376);
nand U3672 (N_3672,N_488,N_1089);
nor U3673 (N_3673,N_240,N_1329);
nand U3674 (N_3674,N_1799,N_665);
and U3675 (N_3675,N_2120,N_2645);
nand U3676 (N_3676,N_1624,N_2272);
nand U3677 (N_3677,N_2944,N_38);
nand U3678 (N_3678,N_1264,N_474);
nor U3679 (N_3679,N_2890,N_1548);
or U3680 (N_3680,N_1817,N_1186);
or U3681 (N_3681,N_1826,N_873);
and U3682 (N_3682,N_506,N_2096);
and U3683 (N_3683,N_2897,N_1212);
or U3684 (N_3684,N_577,N_2519);
nor U3685 (N_3685,N_2875,N_498);
nor U3686 (N_3686,N_1179,N_1809);
xor U3687 (N_3687,N_837,N_495);
or U3688 (N_3688,N_2845,N_2309);
or U3689 (N_3689,N_39,N_2528);
or U3690 (N_3690,N_183,N_2231);
nand U3691 (N_3691,N_457,N_1190);
nor U3692 (N_3692,N_615,N_2239);
nand U3693 (N_3693,N_620,N_905);
nand U3694 (N_3694,N_1325,N_1340);
and U3695 (N_3695,N_2492,N_1048);
and U3696 (N_3696,N_1755,N_1633);
nor U3697 (N_3697,N_513,N_1618);
or U3698 (N_3698,N_1063,N_1569);
nor U3699 (N_3699,N_2864,N_233);
or U3700 (N_3700,N_1070,N_2416);
xor U3701 (N_3701,N_1233,N_804);
xor U3702 (N_3702,N_855,N_1611);
nor U3703 (N_3703,N_2653,N_258);
and U3704 (N_3704,N_878,N_41);
and U3705 (N_3705,N_2207,N_2915);
and U3706 (N_3706,N_1055,N_250);
xor U3707 (N_3707,N_2633,N_1787);
xor U3708 (N_3708,N_2529,N_2822);
nand U3709 (N_3709,N_1948,N_453);
nor U3710 (N_3710,N_1966,N_725);
and U3711 (N_3711,N_2763,N_784);
or U3712 (N_3712,N_16,N_946);
nor U3713 (N_3713,N_1716,N_1437);
nand U3714 (N_3714,N_1607,N_46);
nand U3715 (N_3715,N_2894,N_2727);
nand U3716 (N_3716,N_1240,N_2550);
nor U3717 (N_3717,N_1377,N_1043);
nand U3718 (N_3718,N_1422,N_2514);
nand U3719 (N_3719,N_1545,N_1046);
and U3720 (N_3720,N_2203,N_1459);
or U3721 (N_3721,N_2426,N_2974);
and U3722 (N_3722,N_74,N_1981);
nor U3723 (N_3723,N_219,N_2634);
and U3724 (N_3724,N_1467,N_2661);
and U3725 (N_3725,N_1092,N_207);
or U3726 (N_3726,N_2477,N_2639);
nand U3727 (N_3727,N_1587,N_1669);
and U3728 (N_3728,N_1426,N_1189);
and U3729 (N_3729,N_2398,N_302);
or U3730 (N_3730,N_543,N_901);
nand U3731 (N_3731,N_1598,N_2296);
or U3732 (N_3732,N_2333,N_2334);
and U3733 (N_3733,N_1556,N_528);
and U3734 (N_3734,N_719,N_2688);
nor U3735 (N_3735,N_365,N_1027);
nor U3736 (N_3736,N_115,N_950);
or U3737 (N_3737,N_1408,N_1797);
nor U3738 (N_3738,N_860,N_1969);
nor U3739 (N_3739,N_155,N_2013);
and U3740 (N_3740,N_1282,N_2683);
nor U3741 (N_3741,N_637,N_2778);
nor U3742 (N_3742,N_2480,N_2902);
xnor U3743 (N_3743,N_2608,N_2457);
nor U3744 (N_3744,N_1781,N_2882);
nor U3745 (N_3745,N_2148,N_319);
xnor U3746 (N_3746,N_1017,N_1087);
and U3747 (N_3747,N_2380,N_935);
nor U3748 (N_3748,N_914,N_931);
xor U3749 (N_3749,N_95,N_2807);
nand U3750 (N_3750,N_2304,N_1333);
and U3751 (N_3751,N_1235,N_1652);
or U3752 (N_3752,N_927,N_1793);
nor U3753 (N_3753,N_571,N_669);
xnor U3754 (N_3754,N_2933,N_1160);
xor U3755 (N_3755,N_1653,N_2895);
or U3756 (N_3756,N_1673,N_1747);
and U3757 (N_3757,N_1738,N_480);
or U3758 (N_3758,N_1326,N_593);
nor U3759 (N_3759,N_1922,N_606);
and U3760 (N_3760,N_11,N_2908);
nor U3761 (N_3761,N_33,N_105);
xnor U3762 (N_3762,N_1509,N_317);
or U3763 (N_3763,N_56,N_1102);
xnor U3764 (N_3764,N_259,N_2581);
or U3765 (N_3765,N_491,N_85);
and U3766 (N_3766,N_2362,N_1201);
and U3767 (N_3767,N_2905,N_2762);
and U3768 (N_3768,N_410,N_802);
or U3769 (N_3769,N_2104,N_1621);
or U3770 (N_3770,N_1086,N_1114);
nor U3771 (N_3771,N_145,N_1001);
or U3772 (N_3772,N_2917,N_1914);
or U3773 (N_3773,N_1958,N_2355);
xor U3774 (N_3774,N_442,N_2484);
nor U3775 (N_3775,N_2660,N_1766);
nand U3776 (N_3776,N_861,N_1141);
or U3777 (N_3777,N_2163,N_2774);
nand U3778 (N_3778,N_1739,N_381);
or U3779 (N_3779,N_814,N_2322);
and U3780 (N_3780,N_2267,N_254);
nor U3781 (N_3781,N_2520,N_2648);
xnor U3782 (N_3782,N_2378,N_1374);
and U3783 (N_3783,N_2375,N_1161);
nor U3784 (N_3784,N_2011,N_695);
nand U3785 (N_3785,N_688,N_151);
nand U3786 (N_3786,N_1810,N_976);
and U3787 (N_3787,N_1767,N_2876);
and U3788 (N_3788,N_2742,N_2432);
nor U3789 (N_3789,N_1836,N_1953);
nor U3790 (N_3790,N_350,N_2551);
xor U3791 (N_3791,N_1128,N_1363);
xor U3792 (N_3792,N_1965,N_391);
and U3793 (N_3793,N_2810,N_2255);
nand U3794 (N_3794,N_2662,N_81);
or U3795 (N_3795,N_1898,N_718);
and U3796 (N_3796,N_2579,N_2175);
xnor U3797 (N_3797,N_1790,N_742);
and U3798 (N_3798,N_2970,N_1156);
or U3799 (N_3799,N_808,N_2689);
and U3800 (N_3800,N_2539,N_2443);
nand U3801 (N_3801,N_2509,N_1435);
xnor U3802 (N_3802,N_2260,N_2141);
nand U3803 (N_3803,N_206,N_1349);
or U3804 (N_3804,N_1045,N_1764);
nand U3805 (N_3805,N_1241,N_1456);
nand U3806 (N_3806,N_879,N_2100);
nand U3807 (N_3807,N_573,N_2485);
and U3808 (N_3808,N_2702,N_1295);
nor U3809 (N_3809,N_979,N_332);
nand U3810 (N_3810,N_2733,N_1541);
or U3811 (N_3811,N_304,N_697);
nand U3812 (N_3812,N_2842,N_1032);
nand U3813 (N_3813,N_2697,N_1843);
nand U3814 (N_3814,N_328,N_613);
and U3815 (N_3815,N_82,N_309);
and U3816 (N_3816,N_357,N_2397);
xor U3817 (N_3817,N_1846,N_2982);
nor U3818 (N_3818,N_514,N_138);
or U3819 (N_3819,N_67,N_275);
nor U3820 (N_3820,N_1719,N_177);
nand U3821 (N_3821,N_208,N_2038);
nor U3822 (N_3822,N_2614,N_2610);
xor U3823 (N_3823,N_2910,N_1446);
nand U3824 (N_3824,N_1910,N_618);
and U3825 (N_3825,N_2474,N_1234);
xnor U3826 (N_3826,N_1693,N_282);
and U3827 (N_3827,N_2596,N_787);
and U3828 (N_3828,N_538,N_1699);
nand U3829 (N_3829,N_1842,N_2681);
xnor U3830 (N_3830,N_2829,N_1064);
or U3831 (N_3831,N_1496,N_2799);
nor U3832 (N_3832,N_2587,N_1211);
nand U3833 (N_3833,N_672,N_598);
or U3834 (N_3834,N_477,N_1580);
and U3835 (N_3835,N_393,N_2372);
or U3836 (N_3836,N_1924,N_2009);
nand U3837 (N_3837,N_858,N_1327);
and U3838 (N_3838,N_1991,N_1074);
or U3839 (N_3839,N_507,N_722);
nor U3840 (N_3840,N_1176,N_1520);
nand U3841 (N_3841,N_907,N_616);
and U3842 (N_3842,N_2973,N_335);
nand U3843 (N_3843,N_633,N_2525);
or U3844 (N_3844,N_1011,N_436);
and U3845 (N_3845,N_239,N_466);
nor U3846 (N_3846,N_2332,N_1080);
or U3847 (N_3847,N_584,N_1466);
or U3848 (N_3848,N_1097,N_2044);
nor U3849 (N_3849,N_2650,N_2290);
nor U3850 (N_3850,N_1343,N_1158);
and U3851 (N_3851,N_1872,N_1103);
nand U3852 (N_3852,N_2440,N_1505);
or U3853 (N_3853,N_1722,N_1735);
nor U3854 (N_3854,N_1777,N_957);
nand U3855 (N_3855,N_88,N_723);
xnor U3856 (N_3856,N_426,N_2705);
nand U3857 (N_3857,N_237,N_1275);
or U3858 (N_3858,N_2082,N_1367);
and U3859 (N_3859,N_746,N_969);
nor U3860 (N_3860,N_1831,N_771);
nand U3861 (N_3861,N_2572,N_1460);
or U3862 (N_3862,N_1660,N_940);
nor U3863 (N_3863,N_2773,N_2711);
or U3864 (N_3864,N_1659,N_1023);
and U3865 (N_3865,N_129,N_2347);
and U3866 (N_3866,N_1238,N_23);
nor U3867 (N_3867,N_2720,N_2063);
or U3868 (N_3868,N_37,N_1250);
and U3869 (N_3869,N_712,N_253);
xnor U3870 (N_3870,N_2708,N_2693);
nor U3871 (N_3871,N_2352,N_2571);
or U3872 (N_3872,N_1368,N_2419);
nor U3873 (N_3873,N_1125,N_1718);
or U3874 (N_3874,N_101,N_2233);
and U3875 (N_3875,N_1296,N_1745);
or U3876 (N_3876,N_334,N_998);
or U3877 (N_3877,N_1255,N_2075);
or U3878 (N_3878,N_1599,N_2512);
nand U3879 (N_3879,N_2851,N_2518);
nand U3880 (N_3880,N_853,N_2138);
or U3881 (N_3881,N_2339,N_1795);
or U3882 (N_3882,N_1701,N_2893);
nand U3883 (N_3883,N_2244,N_539);
or U3884 (N_3884,N_1734,N_1244);
and U3885 (N_3885,N_886,N_1658);
nand U3886 (N_3886,N_2297,N_2351);
nor U3887 (N_3887,N_2721,N_2089);
nand U3888 (N_3888,N_1906,N_1131);
nand U3889 (N_3889,N_1051,N_681);
and U3890 (N_3890,N_1071,N_2399);
or U3891 (N_3891,N_2745,N_163);
and U3892 (N_3892,N_715,N_2314);
xor U3893 (N_3893,N_2354,N_2268);
nand U3894 (N_3894,N_826,N_125);
and U3895 (N_3895,N_933,N_1262);
nand U3896 (N_3896,N_2463,N_160);
nor U3897 (N_3897,N_1813,N_1588);
nand U3898 (N_3898,N_1683,N_2687);
and U3899 (N_3899,N_764,N_2004);
nor U3900 (N_3900,N_2964,N_1191);
nor U3901 (N_3901,N_2927,N_546);
or U3902 (N_3902,N_1376,N_12);
and U3903 (N_3903,N_1815,N_2911);
nor U3904 (N_3904,N_1661,N_2410);
nand U3905 (N_3905,N_2624,N_1116);
xor U3906 (N_3906,N_2630,N_2725);
or U3907 (N_3907,N_494,N_1483);
nand U3908 (N_3908,N_517,N_1816);
nand U3909 (N_3909,N_1536,N_1648);
xor U3910 (N_3910,N_1972,N_2261);
and U3911 (N_3911,N_113,N_409);
and U3912 (N_3912,N_1450,N_1935);
and U3913 (N_3913,N_2953,N_2631);
and U3914 (N_3914,N_1221,N_707);
and U3915 (N_3915,N_1544,N_870);
and U3916 (N_3916,N_1829,N_958);
or U3917 (N_3917,N_2414,N_948);
xnor U3918 (N_3918,N_2884,N_1955);
nand U3919 (N_3919,N_2323,N_2770);
or U3920 (N_3920,N_2997,N_2921);
and U3921 (N_3921,N_1939,N_913);
nor U3922 (N_3922,N_168,N_686);
and U3923 (N_3923,N_2212,N_774);
or U3924 (N_3924,N_1304,N_2948);
nor U3925 (N_3925,N_2692,N_1214);
nand U3926 (N_3926,N_1905,N_834);
or U3927 (N_3927,N_703,N_2273);
and U3928 (N_3928,N_1439,N_162);
or U3929 (N_3929,N_1016,N_2265);
xnor U3930 (N_3930,N_117,N_2636);
nand U3931 (N_3931,N_489,N_2592);
nand U3932 (N_3932,N_726,N_996);
nor U3933 (N_3933,N_2928,N_308);
nor U3934 (N_3934,N_2490,N_820);
and U3935 (N_3935,N_2805,N_2266);
nand U3936 (N_3936,N_2224,N_413);
or U3937 (N_3937,N_2885,N_909);
nand U3938 (N_3938,N_800,N_1115);
or U3939 (N_3939,N_2968,N_841);
or U3940 (N_3940,N_1538,N_1180);
or U3941 (N_3941,N_2337,N_2564);
nand U3942 (N_3942,N_1595,N_1276);
nor U3943 (N_3943,N_1285,N_347);
nor U3944 (N_3944,N_60,N_2863);
and U3945 (N_3945,N_2229,N_1727);
and U3946 (N_3946,N_1533,N_118);
or U3947 (N_3947,N_1281,N_1106);
and U3948 (N_3948,N_2452,N_608);
xor U3949 (N_3949,N_1398,N_1585);
nor U3950 (N_3950,N_536,N_2931);
and U3951 (N_3951,N_2816,N_1848);
nor U3952 (N_3952,N_1053,N_792);
or U3953 (N_3953,N_1821,N_1168);
nor U3954 (N_3954,N_342,N_1346);
and U3955 (N_3955,N_1921,N_2914);
nor U3956 (N_3956,N_2515,N_866);
or U3957 (N_3957,N_526,N_2999);
or U3958 (N_3958,N_1494,N_2248);
xor U3959 (N_3959,N_1172,N_1075);
nor U3960 (N_3960,N_2472,N_1668);
and U3961 (N_3961,N_1679,N_2179);
nor U3962 (N_3962,N_1708,N_1381);
and U3963 (N_3963,N_2206,N_1223);
and U3964 (N_3964,N_2496,N_930);
nand U3965 (N_3965,N_215,N_627);
nand U3966 (N_3966,N_476,N_657);
xnor U3967 (N_3967,N_605,N_2527);
nor U3968 (N_3968,N_2076,N_2965);
nor U3969 (N_3969,N_1122,N_684);
or U3970 (N_3970,N_2071,N_799);
nand U3971 (N_3971,N_503,N_2767);
nor U3972 (N_3972,N_902,N_1344);
nand U3973 (N_3973,N_1644,N_379);
and U3974 (N_3974,N_607,N_1694);
and U3975 (N_3975,N_1109,N_2388);
and U3976 (N_3976,N_1260,N_245);
nand U3977 (N_3977,N_1147,N_1849);
nor U3978 (N_3978,N_2055,N_2820);
and U3979 (N_3979,N_1182,N_29);
nor U3980 (N_3980,N_45,N_1142);
and U3981 (N_3981,N_1564,N_1947);
or U3982 (N_3982,N_868,N_2238);
or U3983 (N_3983,N_2724,N_439);
or U3984 (N_3984,N_1744,N_806);
nor U3985 (N_3985,N_153,N_848);
nand U3986 (N_3986,N_782,N_414);
or U3987 (N_3987,N_623,N_459);
or U3988 (N_3988,N_2247,N_1218);
nor U3989 (N_3989,N_980,N_1546);
and U3990 (N_3990,N_2300,N_452);
nor U3991 (N_3991,N_823,N_2110);
or U3992 (N_3992,N_890,N_121);
nor U3993 (N_3993,N_1654,N_429);
or U3994 (N_3994,N_1154,N_1261);
nor U3995 (N_3995,N_2679,N_2387);
and U3996 (N_3996,N_315,N_1863);
and U3997 (N_3997,N_484,N_832);
nand U3998 (N_3998,N_421,N_375);
nand U3999 (N_3999,N_1093,N_2157);
and U4000 (N_4000,N_652,N_1740);
or U4001 (N_4001,N_2889,N_2115);
or U4002 (N_4002,N_2299,N_1748);
nor U4003 (N_4003,N_2256,N_1298);
and U4004 (N_4004,N_341,N_2768);
xor U4005 (N_4005,N_2308,N_1164);
nor U4006 (N_4006,N_2817,N_228);
or U4007 (N_4007,N_1680,N_127);
nor U4008 (N_4008,N_1310,N_1579);
nand U4009 (N_4009,N_227,N_1709);
or U4010 (N_4010,N_599,N_1984);
nand U4011 (N_4011,N_1853,N_1746);
and U4012 (N_4012,N_2274,N_2447);
and U4013 (N_4013,N_2924,N_2465);
xor U4014 (N_4014,N_898,N_2305);
nand U4015 (N_4015,N_400,N_2722);
and U4016 (N_4016,N_1759,N_320);
or U4017 (N_4017,N_2467,N_932);
and U4018 (N_4018,N_256,N_743);
nor U4019 (N_4019,N_2311,N_2865);
or U4020 (N_4020,N_1274,N_2054);
nand U4021 (N_4021,N_1971,N_2396);
nand U4022 (N_4022,N_501,N_96);
or U4023 (N_4023,N_2093,N_582);
or U4024 (N_4024,N_2955,N_2007);
or U4025 (N_4025,N_1384,N_176);
nor U4026 (N_4026,N_2356,N_471);
nor U4027 (N_4027,N_1967,N_1323);
xnor U4028 (N_4028,N_588,N_2216);
and U4029 (N_4029,N_2782,N_836);
xnor U4030 (N_4030,N_2594,N_1833);
nor U4031 (N_4031,N_1099,N_2043);
nor U4032 (N_4032,N_654,N_1985);
or U4033 (N_4033,N_595,N_446);
and U4034 (N_4034,N_1936,N_499);
nor U4035 (N_4035,N_2916,N_2589);
nand U4036 (N_4036,N_1594,N_2112);
and U4037 (N_4037,N_362,N_2584);
xnor U4038 (N_4038,N_1289,N_2489);
nor U4039 (N_4039,N_1717,N_565);
or U4040 (N_4040,N_1482,N_1124);
nor U4041 (N_4041,N_1915,N_2095);
and U4042 (N_4042,N_2783,N_2866);
or U4043 (N_4043,N_2839,N_1614);
or U4044 (N_4044,N_1270,N_1396);
and U4045 (N_4045,N_1288,N_2326);
xnor U4046 (N_4046,N_956,N_2097);
nor U4047 (N_4047,N_1084,N_1650);
and U4048 (N_4048,N_988,N_1136);
xor U4049 (N_4049,N_2442,N_2985);
nor U4050 (N_4050,N_2057,N_201);
and U4051 (N_4051,N_2348,N_2956);
and U4052 (N_4052,N_1616,N_2384);
nand U4053 (N_4053,N_1571,N_1341);
nor U4054 (N_4054,N_745,N_549);
nand U4055 (N_4055,N_1144,N_531);
xnor U4056 (N_4056,N_2099,N_541);
nor U4057 (N_4057,N_570,N_1752);
xnor U4058 (N_4058,N_2039,N_380);
nor U4059 (N_4059,N_2926,N_1372);
and U4060 (N_4060,N_2343,N_444);
nand U4061 (N_4061,N_171,N_2176);
and U4062 (N_4062,N_2622,N_1002);
and U4063 (N_4063,N_1216,N_1468);
nor U4064 (N_4064,N_944,N_651);
or U4065 (N_4065,N_1278,N_2664);
nor U4066 (N_4066,N_1527,N_274);
and U4067 (N_4067,N_2131,N_1723);
nor U4068 (N_4068,N_1982,N_2713);
nand U4069 (N_4069,N_954,N_962);
or U4070 (N_4070,N_1256,N_1912);
and U4071 (N_4071,N_406,N_2155);
or U4072 (N_4072,N_736,N_425);
or U4073 (N_4073,N_1510,N_2116);
xor U4074 (N_4074,N_1073,N_1557);
nor U4075 (N_4075,N_1354,N_2251);
or U4076 (N_4076,N_1324,N_284);
nand U4077 (N_4077,N_1941,N_2856);
xor U4078 (N_4078,N_1444,N_699);
nand U4079 (N_4079,N_197,N_2769);
nand U4080 (N_4080,N_2815,N_2698);
nand U4081 (N_4081,N_2777,N_2701);
nand U4082 (N_4082,N_2966,N_1507);
xor U4083 (N_4083,N_519,N_601);
nor U4084 (N_4084,N_659,N_130);
or U4085 (N_4085,N_2211,N_217);
nand U4086 (N_4086,N_2575,N_1998);
or U4087 (N_4087,N_867,N_1674);
or U4088 (N_4088,N_1741,N_1854);
nor U4089 (N_4089,N_448,N_2743);
and U4090 (N_4090,N_727,N_2930);
xnor U4091 (N_4091,N_1451,N_1369);
nand U4092 (N_4092,N_1197,N_479);
or U4093 (N_4093,N_1575,N_1883);
and U4094 (N_4094,N_903,N_1625);
or U4095 (N_4095,N_1902,N_2453);
or U4096 (N_4096,N_1404,N_411);
nor U4097 (N_4097,N_455,N_2732);
nand U4098 (N_4098,N_2735,N_43);
nor U4099 (N_4099,N_2346,N_1392);
nor U4100 (N_4100,N_1685,N_809);
or U4101 (N_4101,N_31,N_798);
or U4102 (N_4102,N_975,N_2417);
and U4103 (N_4103,N_2435,N_1440);
or U4104 (N_4104,N_585,N_2642);
or U4105 (N_4105,N_2707,N_717);
nand U4106 (N_4106,N_2178,N_2363);
or U4107 (N_4107,N_496,N_2379);
nor U4108 (N_4108,N_1788,N_2455);
nand U4109 (N_4109,N_2957,N_1267);
nand U4110 (N_4110,N_458,N_1847);
nand U4111 (N_4111,N_2280,N_40);
nand U4112 (N_4112,N_1882,N_2001);
or U4113 (N_4113,N_1574,N_551);
and U4114 (N_4114,N_2205,N_2833);
nor U4115 (N_4115,N_2892,N_209);
nor U4116 (N_4116,N_995,N_109);
nor U4117 (N_4117,N_1785,N_243);
or U4118 (N_4118,N_2412,N_1171);
and U4119 (N_4119,N_2516,N_1643);
and U4120 (N_4120,N_2685,N_2156);
nand U4121 (N_4121,N_1480,N_952);
nand U4122 (N_4122,N_98,N_1566);
nand U4123 (N_4123,N_893,N_2861);
nand U4124 (N_4124,N_993,N_1230);
xnor U4125 (N_4125,N_1148,N_1479);
and U4126 (N_4126,N_1707,N_2098);
nand U4127 (N_4127,N_35,N_262);
xnor U4128 (N_4128,N_1592,N_2313);
nor U4129 (N_4129,N_636,N_569);
nand U4130 (N_4130,N_2972,N_510);
nand U4131 (N_4131,N_1014,N_664);
nor U4132 (N_4132,N_591,N_1974);
nor U4133 (N_4133,N_1728,N_287);
nand U4134 (N_4134,N_674,N_2987);
nor U4135 (N_4135,N_1332,N_772);
and U4136 (N_4136,N_17,N_1704);
nor U4137 (N_4137,N_626,N_1236);
xnor U4138 (N_4138,N_2959,N_184);
nand U4139 (N_4139,N_2291,N_13);
or U4140 (N_4140,N_2819,N_556);
nor U4141 (N_4141,N_1300,N_773);
nor U4142 (N_4142,N_1794,N_757);
nor U4143 (N_4143,N_2794,N_2682);
or U4144 (N_4144,N_1026,N_49);
nand U4145 (N_4145,N_449,N_2160);
or U4146 (N_4146,N_15,N_2949);
nor U4147 (N_4147,N_1472,N_1245);
nand U4148 (N_4148,N_1927,N_473);
nor U4149 (N_4149,N_504,N_1370);
and U4150 (N_4150,N_255,N_851);
xor U4151 (N_4151,N_2382,N_2479);
or U4152 (N_4152,N_1715,N_1420);
nor U4153 (N_4153,N_1638,N_2066);
and U4154 (N_4154,N_2357,N_1871);
nor U4155 (N_4155,N_2338,N_1066);
or U4156 (N_4156,N_1476,N_1044);
or U4157 (N_4157,N_1029,N_2062);
xnor U4158 (N_4158,N_2750,N_970);
and U4159 (N_4159,N_1481,N_1901);
nor U4160 (N_4160,N_2456,N_305);
nand U4161 (N_4161,N_1612,N_1033);
nand U4162 (N_4162,N_2629,N_2601);
and U4163 (N_4163,N_2932,N_70);
nor U4164 (N_4164,N_2056,N_2113);
nand U4165 (N_4165,N_1572,N_883);
and U4166 (N_4166,N_1177,N_1322);
or U4167 (N_4167,N_281,N_1042);
xor U4168 (N_4168,N_574,N_90);
nor U4169 (N_4169,N_1742,N_1478);
or U4170 (N_4170,N_1519,N_1098);
nand U4171 (N_4171,N_1891,N_53);
xor U4172 (N_4172,N_2288,N_1895);
nand U4173 (N_4173,N_765,N_505);
and U4174 (N_4174,N_2502,N_2588);
nand U4175 (N_4175,N_1195,N_2570);
and U4176 (N_4176,N_427,N_1391);
nand U4177 (N_4177,N_330,N_2758);
and U4178 (N_4178,N_2937,N_2437);
and U4179 (N_4179,N_123,N_1035);
and U4180 (N_4180,N_1291,N_2848);
and U4181 (N_4181,N_766,N_2353);
or U4182 (N_4182,N_2803,N_1504);
nor U4183 (N_4183,N_2975,N_2840);
nand U4184 (N_4184,N_2855,N_1630);
and U4185 (N_4185,N_1663,N_2632);
xnor U4186 (N_4186,N_1602,N_165);
nor U4187 (N_4187,N_2221,N_2609);
or U4188 (N_4188,N_751,N_76);
nor U4189 (N_4189,N_2407,N_789);
nand U4190 (N_4190,N_916,N_2809);
and U4191 (N_4191,N_1558,N_892);
nor U4192 (N_4192,N_267,N_762);
and U4193 (N_4193,N_297,N_1886);
nor U4194 (N_4194,N_2598,N_655);
xor U4195 (N_4195,N_670,N_2694);
and U4196 (N_4196,N_2230,N_2235);
xor U4197 (N_4197,N_649,N_1762);
or U4198 (N_4198,N_749,N_1059);
nor U4199 (N_4199,N_1049,N_1845);
or U4200 (N_4200,N_2373,N_2669);
nand U4201 (N_4201,N_1550,N_1199);
and U4202 (N_4202,N_1464,N_1113);
xor U4203 (N_4203,N_277,N_1870);
or U4204 (N_4204,N_1050,N_2715);
nor U4205 (N_4205,N_104,N_2264);
nor U4206 (N_4206,N_2031,N_493);
xor U4207 (N_4207,N_2214,N_1626);
nor U4208 (N_4208,N_2181,N_1243);
nor U4209 (N_4209,N_1297,N_2784);
and U4210 (N_4210,N_143,N_602);
nand U4211 (N_4211,N_1219,N_844);
and U4212 (N_4212,N_2404,N_1423);
nor U4213 (N_4213,N_2546,N_2263);
nor U4214 (N_4214,N_2108,N_2547);
nor U4215 (N_4215,N_2511,N_586);
nand U4216 (N_4216,N_438,N_1134);
and U4217 (N_4217,N_2857,N_2027);
nor U4218 (N_4218,N_2878,N_973);
and U4219 (N_4219,N_781,N_1757);
nand U4220 (N_4220,N_1900,N_175);
nand U4221 (N_4221,N_578,N_434);
and U4222 (N_4222,N_1841,N_634);
or U4223 (N_4223,N_2616,N_1286);
or U4224 (N_4224,N_641,N_232);
nand U4225 (N_4225,N_2651,N_1491);
nor U4226 (N_4226,N_1428,N_1328);
and U4227 (N_4227,N_2984,N_2243);
nor U4228 (N_4228,N_1366,N_75);
and U4229 (N_4229,N_2874,N_2946);
nand U4230 (N_4230,N_1210,N_2019);
or U4231 (N_4231,N_1928,N_2760);
nor U4232 (N_4232,N_2696,N_1732);
and U4233 (N_4233,N_2977,N_1037);
or U4234 (N_4234,N_2431,N_705);
and U4235 (N_4235,N_272,N_1352);
and U4236 (N_4236,N_1917,N_1713);
nand U4237 (N_4237,N_2341,N_469);
and U4238 (N_4238,N_2048,N_386);
or U4239 (N_4239,N_68,N_1929);
nor U4240 (N_4240,N_1155,N_296);
and U4241 (N_4241,N_1931,N_2102);
nor U4242 (N_4242,N_1605,N_603);
nand U4243 (N_4243,N_170,N_432);
or U4244 (N_4244,N_2344,N_135);
and U4245 (N_4245,N_236,N_2599);
xor U4246 (N_4246,N_763,N_1253);
nor U4247 (N_4247,N_1897,N_2980);
or U4248 (N_4248,N_925,N_625);
nand U4249 (N_4249,N_2154,N_1531);
xor U4250 (N_4250,N_2821,N_1697);
nor U4251 (N_4251,N_2024,N_900);
nor U4252 (N_4252,N_36,N_1823);
xor U4253 (N_4253,N_1247,N_345);
xor U4254 (N_4254,N_398,N_94);
and U4255 (N_4255,N_1076,N_2377);
and U4256 (N_4256,N_533,N_2254);
nand U4257 (N_4257,N_1613,N_2716);
nand U4258 (N_4258,N_62,N_1083);
nor U4259 (N_4259,N_367,N_2215);
and U4260 (N_4260,N_1196,N_559);
nor U4261 (N_4261,N_310,N_2165);
and U4262 (N_4262,N_1869,N_675);
nor U4263 (N_4263,N_1893,N_2123);
nand U4264 (N_4264,N_1132,N_2691);
xnor U4265 (N_4265,N_288,N_423);
xor U4266 (N_4266,N_817,N_1021);
nor U4267 (N_4267,N_158,N_2241);
and U4268 (N_4268,N_1498,N_2729);
or U4269 (N_4269,N_2164,N_497);
nor U4270 (N_4270,N_683,N_2649);
and U4271 (N_4271,N_1534,N_545);
nand U4272 (N_4272,N_590,N_2180);
nor U4273 (N_4273,N_2285,N_73);
nand U4274 (N_4274,N_1000,N_986);
xor U4275 (N_4275,N_1129,N_2983);
xor U4276 (N_4276,N_1591,N_2712);
nor U4277 (N_4277,N_2209,N_2258);
nor U4278 (N_4278,N_1188,N_2938);
nor U4279 (N_4279,N_2107,N_779);
xnor U4280 (N_4280,N_1178,N_359);
and U4281 (N_4281,N_2828,N_1702);
and U4282 (N_4282,N_492,N_619);
or U4283 (N_4283,N_2132,N_2491);
and U4284 (N_4284,N_1200,N_1977);
nand U4285 (N_4285,N_1105,N_1819);
nor U4286 (N_4286,N_2137,N_116);
nor U4287 (N_4287,N_1968,N_2278);
xnor U4288 (N_4288,N_1827,N_1681);
nor U4289 (N_4289,N_2316,N_1515);
xnor U4290 (N_4290,N_2668,N_2439);
and U4291 (N_4291,N_2934,N_1665);
nor U4292 (N_4292,N_1268,N_1749);
and U4293 (N_4293,N_824,N_1758);
and U4294 (N_4294,N_1726,N_1306);
nand U4295 (N_4295,N_313,N_1301);
and U4296 (N_4296,N_2025,N_141);
and U4297 (N_4297,N_65,N_2173);
and U4298 (N_4298,N_182,N_1525);
nor U4299 (N_4299,N_91,N_1763);
nand U4300 (N_4300,N_92,N_2408);
xor U4301 (N_4301,N_2545,N_216);
nand U4302 (N_4302,N_2184,N_803);
nand U4303 (N_4303,N_1272,N_34);
or U4304 (N_4304,N_849,N_2513);
nor U4305 (N_4305,N_1844,N_1458);
and U4306 (N_4306,N_2667,N_1636);
nand U4307 (N_4307,N_692,N_1248);
or U4308 (N_4308,N_1091,N_938);
nor U4309 (N_4309,N_1753,N_2310);
or U4310 (N_4310,N_1839,N_2607);
nand U4311 (N_4311,N_926,N_2558);
and U4312 (N_4312,N_1317,N_1090);
nand U4313 (N_4313,N_1139,N_2142);
or U4314 (N_4314,N_754,N_292);
xor U4315 (N_4315,N_465,N_1825);
or U4316 (N_4316,N_1193,N_248);
nand U4317 (N_4317,N_522,N_1503);
nand U4318 (N_4318,N_24,N_349);
or U4319 (N_4319,N_47,N_72);
and U4320 (N_4320,N_48,N_1231);
or U4321 (N_4321,N_737,N_377);
or U4322 (N_4322,N_1672,N_1475);
xnor U4323 (N_4323,N_813,N_2286);
or U4324 (N_4324,N_977,N_2739);
nor U4325 (N_4325,N_2105,N_2041);
nor U4326 (N_4326,N_576,N_961);
nand U4327 (N_4327,N_1184,N_1942);
or U4328 (N_4328,N_752,N_1095);
and U4329 (N_4329,N_716,N_2319);
or U4330 (N_4330,N_2167,N_1676);
nand U4331 (N_4331,N_1516,N_1085);
or U4332 (N_4332,N_1952,N_843);
and U4333 (N_4333,N_1570,N_318);
and U4334 (N_4334,N_1647,N_644);
xor U4335 (N_4335,N_614,N_2814);
and U4336 (N_4336,N_2277,N_2385);
nand U4337 (N_4337,N_1937,N_1916);
xnor U4338 (N_4338,N_1421,N_2070);
nor U4339 (N_4339,N_583,N_21);
xor U4340 (N_4340,N_2177,N_311);
or U4341 (N_4341,N_793,N_1549);
and U4342 (N_4342,N_1415,N_1117);
nor U4343 (N_4343,N_1271,N_2747);
nand U4344 (N_4344,N_963,N_1656);
nand U4345 (N_4345,N_61,N_460);
and U4346 (N_4346,N_908,N_949);
nor U4347 (N_4347,N_2303,N_2940);
or U4348 (N_4348,N_1651,N_279);
xnor U4349 (N_4349,N_1806,N_363);
nor U4350 (N_4350,N_261,N_2494);
or U4351 (N_4351,N_548,N_2077);
and U4352 (N_4352,N_955,N_2028);
nor U4353 (N_4353,N_415,N_2913);
and U4354 (N_4354,N_1206,N_755);
nor U4355 (N_4355,N_1567,N_419);
or U4356 (N_4356,N_1490,N_1610);
and U4357 (N_4357,N_2294,N_871);
nand U4358 (N_4358,N_1649,N_1041);
or U4359 (N_4359,N_621,N_1100);
nor U4360 (N_4360,N_1443,N_2017);
nand U4361 (N_4361,N_2796,N_1409);
xor U4362 (N_4362,N_2542,N_770);
or U4363 (N_4363,N_220,N_990);
nand U4364 (N_4364,N_558,N_2736);
nor U4365 (N_4365,N_1174,N_544);
and U4366 (N_4366,N_2429,N_1338);
or U4367 (N_4367,N_2718,N_2576);
nor U4368 (N_4368,N_780,N_1127);
or U4369 (N_4369,N_463,N_1999);
xnor U4370 (N_4370,N_2454,N_2553);
nand U4371 (N_4371,N_2675,N_769);
xnor U4372 (N_4372,N_1334,N_2891);
nand U4373 (N_4373,N_2526,N_286);
or U4374 (N_4374,N_887,N_2103);
xnor U4375 (N_4375,N_42,N_2824);
nand U4376 (N_4376,N_795,N_360);
or U4377 (N_4377,N_437,N_609);
and U4378 (N_4378,N_152,N_241);
or U4379 (N_4379,N_28,N_2151);
and U4380 (N_4380,N_355,N_2870);
or U4381 (N_4381,N_862,N_818);
and U4382 (N_4382,N_450,N_1448);
nor U4383 (N_4383,N_1493,N_2200);
and U4384 (N_4384,N_337,N_1919);
xnor U4385 (N_4385,N_440,N_2567);
nand U4386 (N_4386,N_1513,N_148);
or U4387 (N_4387,N_351,N_612);
nand U4388 (N_4388,N_833,N_2193);
and U4389 (N_4389,N_1987,N_2638);
and U4390 (N_4390,N_2717,N_666);
or U4391 (N_4391,N_2295,N_468);
or U4392 (N_4392,N_629,N_2943);
or U4393 (N_4393,N_748,N_2000);
nor U4394 (N_4394,N_1068,N_508);
nor U4395 (N_4395,N_2470,N_1312);
or U4396 (N_4396,N_631,N_338);
nand U4397 (N_4397,N_321,N_978);
nor U4398 (N_4398,N_1990,N_1427);
or U4399 (N_4399,N_2620,N_203);
nand U4400 (N_4400,N_2507,N_2191);
and U4401 (N_4401,N_2190,N_2271);
nor U4402 (N_4402,N_865,N_1414);
and U4403 (N_4403,N_1615,N_2677);
nand U4404 (N_4404,N_997,N_2704);
or U4405 (N_4405,N_1120,N_112);
or U4406 (N_4406,N_1169,N_1705);
or U4407 (N_4407,N_354,N_919);
nor U4408 (N_4408,N_2318,N_2094);
xor U4409 (N_4409,N_2015,N_5);
nand U4410 (N_4410,N_2111,N_653);
and U4411 (N_4411,N_1578,N_2781);
or U4412 (N_4412,N_149,N_677);
xnor U4413 (N_4413,N_1108,N_1454);
or U4414 (N_4414,N_2330,N_2873);
and U4415 (N_4415,N_730,N_2069);
nor U4416 (N_4416,N_2504,N_1885);
nand U4417 (N_4417,N_1911,N_2331);
nor U4418 (N_4418,N_2625,N_1350);
or U4419 (N_4419,N_2126,N_1205);
xnor U4420 (N_4420,N_2749,N_50);
nor U4421 (N_4421,N_1858,N_515);
nand U4422 (N_4422,N_2361,N_2315);
and U4423 (N_4423,N_600,N_2114);
nand U4424 (N_4424,N_194,N_2228);
or U4425 (N_4425,N_1920,N_1151);
nand U4426 (N_4426,N_635,N_1407);
nand U4427 (N_4427,N_2883,N_2117);
or U4428 (N_4428,N_648,N_885);
or U4429 (N_4429,N_1772,N_264);
or U4430 (N_4430,N_2023,N_486);
nor U4431 (N_4431,N_1015,N_242);
and U4432 (N_4432,N_1903,N_84);
or U4433 (N_4433,N_164,N_1543);
or U4434 (N_4434,N_1554,N_767);
or U4435 (N_4435,N_1213,N_2170);
and U4436 (N_4436,N_529,N_2240);
and U4437 (N_4437,N_2145,N_1302);
nand U4438 (N_4438,N_2487,N_1215);
nor U4439 (N_4439,N_1348,N_999);
and U4440 (N_4440,N_1433,N_2501);
and U4441 (N_4441,N_178,N_1319);
xor U4442 (N_4442,N_1339,N_290);
and U4443 (N_4443,N_487,N_801);
nor U4444 (N_4444,N_983,N_1629);
nand U4445 (N_4445,N_1751,N_369);
nor U4446 (N_4446,N_2106,N_974);
nor U4447 (N_4447,N_475,N_1783);
or U4448 (N_4448,N_2301,N_992);
nand U4449 (N_4449,N_2674,N_1620);
nand U4450 (N_4450,N_2245,N_1025);
and U4451 (N_4451,N_2606,N_114);
nor U4452 (N_4452,N_587,N_2565);
and U4453 (N_4453,N_2029,N_2130);
or U4454 (N_4454,N_668,N_1926);
or U4455 (N_4455,N_624,N_2026);
xnor U4456 (N_4456,N_1040,N_346);
xnor U4457 (N_4457,N_2425,N_30);
and U4458 (N_4458,N_928,N_710);
xnor U4459 (N_4459,N_2998,N_1009);
nand U4460 (N_4460,N_512,N_301);
and U4461 (N_4461,N_2136,N_2371);
or U4462 (N_4462,N_1355,N_186);
and U4463 (N_4463,N_1486,N_2671);
xor U4464 (N_4464,N_1308,N_1152);
nand U4465 (N_4465,N_1779,N_1330);
nand U4466 (N_4466,N_144,N_1072);
or U4467 (N_4467,N_78,N_1287);
nor U4468 (N_4468,N_1208,N_2785);
and U4469 (N_4469,N_1662,N_340);
xnor U4470 (N_4470,N_2424,N_1896);
or U4471 (N_4471,N_412,N_2438);
nand U4472 (N_4472,N_2812,N_1502);
nand U4473 (N_4473,N_2088,N_1983);
and U4474 (N_4474,N_2242,N_167);
or U4475 (N_4475,N_960,N_1385);
or U4476 (N_4476,N_2580,N_247);
nand U4477 (N_4477,N_2091,N_2827);
nand U4478 (N_4478,N_1808,N_2049);
xor U4479 (N_4479,N_1961,N_2800);
and U4480 (N_4480,N_1889,N_2626);
nand U4481 (N_4481,N_1689,N_2559);
or U4482 (N_4482,N_58,N_2461);
nor U4483 (N_4483,N_2022,N_464);
nor U4484 (N_4484,N_2486,N_1185);
or U4485 (N_4485,N_191,N_906);
nor U4486 (N_4486,N_663,N_1623);
and U4487 (N_4487,N_370,N_329);
or U4488 (N_4488,N_1524,N_483);
nor U4489 (N_4489,N_1878,N_1357);
nor U4490 (N_4490,N_768,N_525);
or U4491 (N_4491,N_1181,N_1010);
nand U4492 (N_4492,N_1711,N_934);
xnor U4493 (N_4493,N_2250,N_63);
nor U4494 (N_4494,N_2124,N_1062);
nand U4495 (N_4495,N_645,N_1246);
nand U4496 (N_4496,N_1222,N_1619);
and U4497 (N_4497,N_1535,N_2703);
or U4498 (N_4498,N_1436,N_2613);
or U4499 (N_4499,N_1280,N_211);
nand U4500 (N_4500,N_787,N_2404);
and U4501 (N_4501,N_1738,N_2219);
nor U4502 (N_4502,N_383,N_2561);
nor U4503 (N_4503,N_784,N_2556);
and U4504 (N_4504,N_1827,N_1017);
or U4505 (N_4505,N_239,N_556);
nand U4506 (N_4506,N_1208,N_788);
nor U4507 (N_4507,N_2000,N_1011);
or U4508 (N_4508,N_2416,N_2642);
or U4509 (N_4509,N_2327,N_2941);
nand U4510 (N_4510,N_387,N_44);
nand U4511 (N_4511,N_2940,N_1783);
nor U4512 (N_4512,N_1096,N_2153);
nor U4513 (N_4513,N_2070,N_1731);
nand U4514 (N_4514,N_2677,N_557);
or U4515 (N_4515,N_921,N_2391);
nand U4516 (N_4516,N_628,N_1409);
and U4517 (N_4517,N_75,N_1001);
nand U4518 (N_4518,N_2763,N_1429);
nand U4519 (N_4519,N_2144,N_1761);
nor U4520 (N_4520,N_2468,N_2361);
nor U4521 (N_4521,N_1487,N_2781);
nand U4522 (N_4522,N_2656,N_2259);
nor U4523 (N_4523,N_400,N_2297);
nand U4524 (N_4524,N_1420,N_1133);
or U4525 (N_4525,N_462,N_2211);
or U4526 (N_4526,N_1185,N_2872);
and U4527 (N_4527,N_2546,N_2434);
nor U4528 (N_4528,N_2196,N_1880);
nand U4529 (N_4529,N_2106,N_2357);
and U4530 (N_4530,N_1662,N_1464);
and U4531 (N_4531,N_622,N_1103);
and U4532 (N_4532,N_416,N_524);
and U4533 (N_4533,N_1244,N_1211);
and U4534 (N_4534,N_1000,N_154);
nand U4535 (N_4535,N_940,N_1996);
or U4536 (N_4536,N_331,N_1127);
or U4537 (N_4537,N_2556,N_588);
and U4538 (N_4538,N_1521,N_2312);
or U4539 (N_4539,N_2159,N_1899);
nor U4540 (N_4540,N_2541,N_1772);
nor U4541 (N_4541,N_2150,N_783);
or U4542 (N_4542,N_2348,N_1281);
and U4543 (N_4543,N_1581,N_2619);
nor U4544 (N_4544,N_1834,N_1426);
xor U4545 (N_4545,N_272,N_2694);
or U4546 (N_4546,N_2322,N_1196);
nor U4547 (N_4547,N_139,N_712);
and U4548 (N_4548,N_2100,N_683);
xor U4549 (N_4549,N_699,N_1835);
nor U4550 (N_4550,N_2737,N_2199);
xnor U4551 (N_4551,N_2203,N_2684);
and U4552 (N_4552,N_1379,N_2936);
nor U4553 (N_4553,N_2857,N_1337);
nand U4554 (N_4554,N_483,N_2401);
and U4555 (N_4555,N_2106,N_857);
or U4556 (N_4556,N_1622,N_2847);
nor U4557 (N_4557,N_2691,N_2824);
nand U4558 (N_4558,N_1429,N_2995);
and U4559 (N_4559,N_872,N_1033);
nand U4560 (N_4560,N_1095,N_1274);
or U4561 (N_4561,N_36,N_2934);
nand U4562 (N_4562,N_2881,N_363);
xnor U4563 (N_4563,N_2143,N_1119);
or U4564 (N_4564,N_1269,N_2047);
and U4565 (N_4565,N_2863,N_2039);
or U4566 (N_4566,N_698,N_748);
or U4567 (N_4567,N_849,N_1884);
nand U4568 (N_4568,N_741,N_1902);
or U4569 (N_4569,N_1021,N_895);
and U4570 (N_4570,N_1948,N_30);
nor U4571 (N_4571,N_1270,N_1033);
nor U4572 (N_4572,N_2767,N_815);
or U4573 (N_4573,N_143,N_2947);
nand U4574 (N_4574,N_2916,N_717);
nand U4575 (N_4575,N_2036,N_2714);
nor U4576 (N_4576,N_2954,N_2765);
nor U4577 (N_4577,N_2824,N_1012);
and U4578 (N_4578,N_784,N_303);
or U4579 (N_4579,N_2784,N_305);
nand U4580 (N_4580,N_1571,N_2466);
xor U4581 (N_4581,N_2463,N_2536);
and U4582 (N_4582,N_1488,N_1954);
and U4583 (N_4583,N_176,N_2187);
nand U4584 (N_4584,N_263,N_368);
or U4585 (N_4585,N_1149,N_1907);
or U4586 (N_4586,N_1963,N_2797);
and U4587 (N_4587,N_394,N_575);
and U4588 (N_4588,N_1288,N_1984);
nor U4589 (N_4589,N_1123,N_2314);
or U4590 (N_4590,N_2381,N_149);
nor U4591 (N_4591,N_2515,N_431);
nand U4592 (N_4592,N_2587,N_1631);
xnor U4593 (N_4593,N_1860,N_1141);
nor U4594 (N_4594,N_1072,N_2723);
nand U4595 (N_4595,N_1138,N_1794);
nand U4596 (N_4596,N_885,N_1845);
or U4597 (N_4597,N_1866,N_2526);
nand U4598 (N_4598,N_1278,N_2244);
and U4599 (N_4599,N_2686,N_508);
nand U4600 (N_4600,N_314,N_865);
nand U4601 (N_4601,N_2550,N_1867);
nand U4602 (N_4602,N_1848,N_1054);
xor U4603 (N_4603,N_1366,N_1643);
and U4604 (N_4604,N_935,N_797);
nand U4605 (N_4605,N_2487,N_2881);
nor U4606 (N_4606,N_1257,N_504);
nor U4607 (N_4607,N_2739,N_1516);
and U4608 (N_4608,N_523,N_1709);
and U4609 (N_4609,N_1110,N_728);
or U4610 (N_4610,N_797,N_1379);
or U4611 (N_4611,N_448,N_2997);
xor U4612 (N_4612,N_674,N_1642);
nand U4613 (N_4613,N_174,N_2639);
nor U4614 (N_4614,N_580,N_2477);
and U4615 (N_4615,N_668,N_1809);
nand U4616 (N_4616,N_946,N_1122);
nand U4617 (N_4617,N_2684,N_2044);
or U4618 (N_4618,N_193,N_121);
or U4619 (N_4619,N_1886,N_1759);
and U4620 (N_4620,N_394,N_2631);
nor U4621 (N_4621,N_2990,N_2783);
nor U4622 (N_4622,N_1886,N_1346);
xor U4623 (N_4623,N_2142,N_1116);
xnor U4624 (N_4624,N_595,N_2907);
or U4625 (N_4625,N_555,N_1789);
or U4626 (N_4626,N_2358,N_1310);
nand U4627 (N_4627,N_2997,N_1593);
nand U4628 (N_4628,N_1826,N_1473);
and U4629 (N_4629,N_2181,N_831);
or U4630 (N_4630,N_1990,N_2474);
nand U4631 (N_4631,N_8,N_2419);
nand U4632 (N_4632,N_653,N_1101);
xor U4633 (N_4633,N_2275,N_1835);
and U4634 (N_4634,N_1477,N_400);
nand U4635 (N_4635,N_1361,N_490);
nor U4636 (N_4636,N_19,N_394);
nor U4637 (N_4637,N_2040,N_2030);
nor U4638 (N_4638,N_1752,N_1056);
nor U4639 (N_4639,N_206,N_1388);
nand U4640 (N_4640,N_1033,N_935);
nand U4641 (N_4641,N_2773,N_1213);
nor U4642 (N_4642,N_2881,N_1567);
xnor U4643 (N_4643,N_221,N_1934);
and U4644 (N_4644,N_2300,N_1955);
or U4645 (N_4645,N_2436,N_1441);
xnor U4646 (N_4646,N_1915,N_1441);
or U4647 (N_4647,N_2813,N_73);
nor U4648 (N_4648,N_2955,N_1034);
nor U4649 (N_4649,N_2458,N_2563);
nor U4650 (N_4650,N_220,N_2261);
nor U4651 (N_4651,N_2861,N_2223);
xnor U4652 (N_4652,N_1733,N_929);
or U4653 (N_4653,N_203,N_2316);
and U4654 (N_4654,N_2862,N_149);
nand U4655 (N_4655,N_1313,N_2180);
nor U4656 (N_4656,N_23,N_2648);
nand U4657 (N_4657,N_2141,N_126);
xnor U4658 (N_4658,N_2898,N_173);
or U4659 (N_4659,N_1114,N_175);
nor U4660 (N_4660,N_180,N_2919);
or U4661 (N_4661,N_2440,N_1216);
or U4662 (N_4662,N_1294,N_2853);
and U4663 (N_4663,N_820,N_1991);
nand U4664 (N_4664,N_2862,N_1501);
and U4665 (N_4665,N_2706,N_1504);
or U4666 (N_4666,N_1428,N_1196);
or U4667 (N_4667,N_1874,N_1687);
nand U4668 (N_4668,N_20,N_784);
and U4669 (N_4669,N_1026,N_2904);
xnor U4670 (N_4670,N_2587,N_1682);
nand U4671 (N_4671,N_805,N_717);
nand U4672 (N_4672,N_1587,N_2694);
xor U4673 (N_4673,N_2485,N_1316);
or U4674 (N_4674,N_2357,N_1122);
xor U4675 (N_4675,N_950,N_1144);
or U4676 (N_4676,N_2551,N_449);
xor U4677 (N_4677,N_891,N_1619);
nand U4678 (N_4678,N_2700,N_240);
and U4679 (N_4679,N_180,N_2960);
xor U4680 (N_4680,N_663,N_1893);
or U4681 (N_4681,N_2514,N_1386);
or U4682 (N_4682,N_860,N_2174);
or U4683 (N_4683,N_1913,N_438);
nand U4684 (N_4684,N_693,N_604);
nor U4685 (N_4685,N_275,N_781);
nand U4686 (N_4686,N_988,N_1296);
or U4687 (N_4687,N_2713,N_892);
and U4688 (N_4688,N_244,N_1539);
or U4689 (N_4689,N_2971,N_826);
nand U4690 (N_4690,N_1385,N_828);
or U4691 (N_4691,N_1161,N_479);
nor U4692 (N_4692,N_844,N_59);
and U4693 (N_4693,N_894,N_473);
or U4694 (N_4694,N_360,N_2327);
and U4695 (N_4695,N_2181,N_2614);
xor U4696 (N_4696,N_1573,N_1229);
nand U4697 (N_4697,N_1167,N_1821);
nor U4698 (N_4698,N_122,N_1667);
xnor U4699 (N_4699,N_558,N_1683);
nor U4700 (N_4700,N_1045,N_2683);
and U4701 (N_4701,N_2073,N_2297);
nand U4702 (N_4702,N_2462,N_90);
and U4703 (N_4703,N_916,N_878);
or U4704 (N_4704,N_1167,N_1639);
nor U4705 (N_4705,N_943,N_92);
nand U4706 (N_4706,N_2534,N_2556);
nand U4707 (N_4707,N_312,N_531);
nor U4708 (N_4708,N_2771,N_1995);
xnor U4709 (N_4709,N_1585,N_1809);
or U4710 (N_4710,N_57,N_524);
nor U4711 (N_4711,N_2435,N_627);
and U4712 (N_4712,N_1330,N_2675);
nor U4713 (N_4713,N_312,N_1234);
xnor U4714 (N_4714,N_2973,N_2029);
nor U4715 (N_4715,N_2999,N_1702);
nor U4716 (N_4716,N_1672,N_2643);
and U4717 (N_4717,N_1529,N_1840);
xnor U4718 (N_4718,N_248,N_1003);
nand U4719 (N_4719,N_1706,N_2716);
nor U4720 (N_4720,N_2138,N_84);
nor U4721 (N_4721,N_1154,N_40);
and U4722 (N_4722,N_140,N_2982);
nor U4723 (N_4723,N_2903,N_2007);
nor U4724 (N_4724,N_2159,N_2871);
and U4725 (N_4725,N_2062,N_2212);
and U4726 (N_4726,N_2647,N_1322);
and U4727 (N_4727,N_1804,N_2929);
or U4728 (N_4728,N_1312,N_2411);
nor U4729 (N_4729,N_948,N_530);
nand U4730 (N_4730,N_2213,N_2871);
nor U4731 (N_4731,N_1285,N_884);
and U4732 (N_4732,N_1155,N_2266);
nor U4733 (N_4733,N_2656,N_1674);
or U4734 (N_4734,N_87,N_1666);
nand U4735 (N_4735,N_339,N_2037);
and U4736 (N_4736,N_1998,N_2885);
nand U4737 (N_4737,N_2032,N_2413);
nand U4738 (N_4738,N_975,N_1047);
nor U4739 (N_4739,N_2078,N_1158);
nand U4740 (N_4740,N_1472,N_1596);
or U4741 (N_4741,N_1980,N_2322);
or U4742 (N_4742,N_2936,N_576);
nand U4743 (N_4743,N_1772,N_559);
nor U4744 (N_4744,N_1662,N_2216);
nor U4745 (N_4745,N_2540,N_538);
and U4746 (N_4746,N_1144,N_576);
and U4747 (N_4747,N_1060,N_1705);
nand U4748 (N_4748,N_2870,N_2056);
and U4749 (N_4749,N_2771,N_1045);
xnor U4750 (N_4750,N_2967,N_2653);
or U4751 (N_4751,N_2829,N_1652);
or U4752 (N_4752,N_1876,N_593);
and U4753 (N_4753,N_2933,N_1152);
and U4754 (N_4754,N_926,N_980);
and U4755 (N_4755,N_2139,N_831);
nor U4756 (N_4756,N_2070,N_2233);
xnor U4757 (N_4757,N_1230,N_2869);
nor U4758 (N_4758,N_886,N_1377);
nor U4759 (N_4759,N_1853,N_2047);
and U4760 (N_4760,N_2261,N_531);
xnor U4761 (N_4761,N_798,N_2645);
or U4762 (N_4762,N_450,N_344);
nand U4763 (N_4763,N_2203,N_305);
and U4764 (N_4764,N_2456,N_315);
or U4765 (N_4765,N_1554,N_523);
nor U4766 (N_4766,N_1376,N_1775);
or U4767 (N_4767,N_2434,N_2768);
nand U4768 (N_4768,N_240,N_1523);
and U4769 (N_4769,N_2602,N_625);
nor U4770 (N_4770,N_1705,N_2135);
nand U4771 (N_4771,N_2472,N_918);
nand U4772 (N_4772,N_1056,N_1969);
xnor U4773 (N_4773,N_1012,N_973);
or U4774 (N_4774,N_538,N_114);
and U4775 (N_4775,N_1322,N_1229);
xnor U4776 (N_4776,N_1973,N_2563);
xnor U4777 (N_4777,N_1168,N_1678);
nor U4778 (N_4778,N_1143,N_2264);
or U4779 (N_4779,N_324,N_1539);
and U4780 (N_4780,N_679,N_159);
xnor U4781 (N_4781,N_1166,N_1032);
nor U4782 (N_4782,N_1184,N_1815);
or U4783 (N_4783,N_326,N_680);
and U4784 (N_4784,N_2911,N_2580);
nand U4785 (N_4785,N_2929,N_879);
and U4786 (N_4786,N_2086,N_256);
or U4787 (N_4787,N_919,N_2957);
xnor U4788 (N_4788,N_1964,N_689);
xor U4789 (N_4789,N_1457,N_2366);
nor U4790 (N_4790,N_1767,N_2815);
or U4791 (N_4791,N_749,N_1403);
or U4792 (N_4792,N_2499,N_1939);
or U4793 (N_4793,N_1761,N_1867);
nor U4794 (N_4794,N_2190,N_2696);
nand U4795 (N_4795,N_2802,N_2971);
nand U4796 (N_4796,N_2940,N_1684);
nand U4797 (N_4797,N_1131,N_219);
and U4798 (N_4798,N_2844,N_1471);
nand U4799 (N_4799,N_1135,N_2122);
nand U4800 (N_4800,N_2454,N_593);
and U4801 (N_4801,N_1959,N_2956);
or U4802 (N_4802,N_675,N_630);
xor U4803 (N_4803,N_256,N_2365);
nand U4804 (N_4804,N_793,N_1987);
and U4805 (N_4805,N_604,N_2996);
or U4806 (N_4806,N_2182,N_182);
and U4807 (N_4807,N_1026,N_2118);
or U4808 (N_4808,N_390,N_1053);
nand U4809 (N_4809,N_1408,N_348);
nand U4810 (N_4810,N_2760,N_922);
nor U4811 (N_4811,N_1582,N_2988);
nand U4812 (N_4812,N_127,N_1753);
and U4813 (N_4813,N_1664,N_2994);
and U4814 (N_4814,N_1925,N_2421);
nor U4815 (N_4815,N_1319,N_1704);
nand U4816 (N_4816,N_2712,N_1642);
xor U4817 (N_4817,N_50,N_829);
nor U4818 (N_4818,N_2470,N_2709);
or U4819 (N_4819,N_2715,N_2373);
nand U4820 (N_4820,N_11,N_1898);
nand U4821 (N_4821,N_1899,N_1049);
nor U4822 (N_4822,N_2615,N_1755);
or U4823 (N_4823,N_1283,N_1616);
nor U4824 (N_4824,N_239,N_328);
nor U4825 (N_4825,N_1280,N_1035);
xor U4826 (N_4826,N_556,N_33);
or U4827 (N_4827,N_74,N_1039);
nand U4828 (N_4828,N_974,N_2935);
or U4829 (N_4829,N_1340,N_52);
or U4830 (N_4830,N_2019,N_1159);
or U4831 (N_4831,N_1176,N_255);
or U4832 (N_4832,N_2009,N_1614);
and U4833 (N_4833,N_827,N_2891);
nand U4834 (N_4834,N_1807,N_322);
nand U4835 (N_4835,N_115,N_501);
nor U4836 (N_4836,N_1630,N_86);
and U4837 (N_4837,N_2480,N_1376);
and U4838 (N_4838,N_1895,N_2858);
or U4839 (N_4839,N_2538,N_2072);
nor U4840 (N_4840,N_2099,N_1029);
xnor U4841 (N_4841,N_435,N_898);
or U4842 (N_4842,N_2964,N_2975);
nor U4843 (N_4843,N_674,N_2160);
nand U4844 (N_4844,N_1919,N_2005);
or U4845 (N_4845,N_2170,N_2938);
nor U4846 (N_4846,N_1104,N_1805);
nor U4847 (N_4847,N_870,N_2661);
xor U4848 (N_4848,N_2384,N_361);
nand U4849 (N_4849,N_2215,N_2908);
xnor U4850 (N_4850,N_44,N_1601);
and U4851 (N_4851,N_1620,N_1563);
nor U4852 (N_4852,N_2402,N_1592);
and U4853 (N_4853,N_138,N_973);
and U4854 (N_4854,N_1447,N_2391);
nor U4855 (N_4855,N_2627,N_2626);
xor U4856 (N_4856,N_14,N_1204);
or U4857 (N_4857,N_1351,N_2853);
nor U4858 (N_4858,N_1099,N_1429);
nand U4859 (N_4859,N_403,N_2479);
xor U4860 (N_4860,N_1897,N_403);
xor U4861 (N_4861,N_1439,N_2640);
or U4862 (N_4862,N_2380,N_2827);
xor U4863 (N_4863,N_1158,N_519);
and U4864 (N_4864,N_719,N_2308);
and U4865 (N_4865,N_2735,N_939);
nand U4866 (N_4866,N_1374,N_716);
nor U4867 (N_4867,N_792,N_859);
and U4868 (N_4868,N_531,N_421);
xor U4869 (N_4869,N_1668,N_549);
xor U4870 (N_4870,N_2761,N_992);
nand U4871 (N_4871,N_866,N_2783);
xnor U4872 (N_4872,N_31,N_2981);
and U4873 (N_4873,N_11,N_1228);
nor U4874 (N_4874,N_1948,N_864);
and U4875 (N_4875,N_386,N_1871);
and U4876 (N_4876,N_86,N_2336);
and U4877 (N_4877,N_521,N_105);
nor U4878 (N_4878,N_330,N_2145);
nor U4879 (N_4879,N_2190,N_570);
nor U4880 (N_4880,N_1654,N_2365);
nor U4881 (N_4881,N_1576,N_865);
and U4882 (N_4882,N_887,N_1541);
nand U4883 (N_4883,N_1486,N_2546);
or U4884 (N_4884,N_1941,N_435);
nor U4885 (N_4885,N_2807,N_362);
xor U4886 (N_4886,N_2377,N_2235);
and U4887 (N_4887,N_1057,N_552);
xnor U4888 (N_4888,N_2843,N_1756);
nor U4889 (N_4889,N_2026,N_1916);
xor U4890 (N_4890,N_261,N_2602);
or U4891 (N_4891,N_604,N_546);
and U4892 (N_4892,N_2316,N_317);
or U4893 (N_4893,N_192,N_1900);
nand U4894 (N_4894,N_1883,N_1785);
and U4895 (N_4895,N_1056,N_562);
or U4896 (N_4896,N_611,N_100);
or U4897 (N_4897,N_1054,N_1943);
nand U4898 (N_4898,N_2212,N_310);
xor U4899 (N_4899,N_2619,N_2224);
nand U4900 (N_4900,N_65,N_986);
xor U4901 (N_4901,N_854,N_1818);
xor U4902 (N_4902,N_1561,N_2205);
xnor U4903 (N_4903,N_686,N_1413);
nand U4904 (N_4904,N_2083,N_2745);
and U4905 (N_4905,N_1941,N_1928);
nand U4906 (N_4906,N_2815,N_753);
or U4907 (N_4907,N_1182,N_1250);
or U4908 (N_4908,N_338,N_475);
or U4909 (N_4909,N_978,N_2052);
nand U4910 (N_4910,N_1187,N_2422);
or U4911 (N_4911,N_29,N_1008);
or U4912 (N_4912,N_932,N_516);
or U4913 (N_4913,N_406,N_897);
nand U4914 (N_4914,N_1214,N_2919);
xor U4915 (N_4915,N_2903,N_2984);
and U4916 (N_4916,N_701,N_2411);
nor U4917 (N_4917,N_17,N_2022);
and U4918 (N_4918,N_427,N_2591);
or U4919 (N_4919,N_691,N_1150);
nand U4920 (N_4920,N_2616,N_2126);
and U4921 (N_4921,N_1961,N_1149);
or U4922 (N_4922,N_1922,N_60);
xor U4923 (N_4923,N_1090,N_2037);
or U4924 (N_4924,N_1626,N_2410);
or U4925 (N_4925,N_1406,N_288);
nand U4926 (N_4926,N_383,N_2330);
or U4927 (N_4927,N_52,N_2784);
xnor U4928 (N_4928,N_1438,N_2154);
nand U4929 (N_4929,N_1300,N_1899);
or U4930 (N_4930,N_1759,N_2649);
nor U4931 (N_4931,N_1824,N_2257);
or U4932 (N_4932,N_946,N_143);
or U4933 (N_4933,N_297,N_16);
or U4934 (N_4934,N_24,N_1080);
or U4935 (N_4935,N_756,N_1444);
nor U4936 (N_4936,N_2983,N_697);
nor U4937 (N_4937,N_2833,N_1039);
nand U4938 (N_4938,N_2425,N_905);
and U4939 (N_4939,N_1489,N_2227);
or U4940 (N_4940,N_1444,N_1207);
nor U4941 (N_4941,N_548,N_756);
xor U4942 (N_4942,N_1857,N_1791);
or U4943 (N_4943,N_784,N_1631);
nor U4944 (N_4944,N_2257,N_2907);
nor U4945 (N_4945,N_513,N_1574);
nand U4946 (N_4946,N_1613,N_2182);
or U4947 (N_4947,N_2700,N_1241);
and U4948 (N_4948,N_1935,N_2618);
and U4949 (N_4949,N_795,N_99);
nand U4950 (N_4950,N_1349,N_1809);
nand U4951 (N_4951,N_1440,N_1412);
nand U4952 (N_4952,N_2310,N_1763);
or U4953 (N_4953,N_1054,N_1771);
nand U4954 (N_4954,N_1059,N_1369);
and U4955 (N_4955,N_268,N_473);
or U4956 (N_4956,N_2455,N_2743);
and U4957 (N_4957,N_1500,N_442);
nor U4958 (N_4958,N_2918,N_1514);
and U4959 (N_4959,N_2393,N_2517);
nor U4960 (N_4960,N_2276,N_243);
xor U4961 (N_4961,N_600,N_1829);
and U4962 (N_4962,N_2335,N_423);
nand U4963 (N_4963,N_1182,N_1223);
or U4964 (N_4964,N_731,N_734);
or U4965 (N_4965,N_167,N_1510);
nor U4966 (N_4966,N_951,N_1823);
and U4967 (N_4967,N_425,N_1554);
and U4968 (N_4968,N_2767,N_836);
nand U4969 (N_4969,N_520,N_2541);
and U4970 (N_4970,N_549,N_79);
nand U4971 (N_4971,N_912,N_1824);
nand U4972 (N_4972,N_2995,N_2882);
and U4973 (N_4973,N_1696,N_1264);
nand U4974 (N_4974,N_2296,N_495);
and U4975 (N_4975,N_1223,N_2684);
nor U4976 (N_4976,N_2843,N_1142);
or U4977 (N_4977,N_1471,N_2837);
nor U4978 (N_4978,N_2458,N_1487);
and U4979 (N_4979,N_1844,N_200);
and U4980 (N_4980,N_2816,N_2642);
or U4981 (N_4981,N_1899,N_1952);
or U4982 (N_4982,N_2345,N_272);
xor U4983 (N_4983,N_1885,N_1550);
nand U4984 (N_4984,N_1134,N_2768);
nor U4985 (N_4985,N_264,N_1512);
xor U4986 (N_4986,N_1481,N_1191);
and U4987 (N_4987,N_923,N_1016);
xor U4988 (N_4988,N_2087,N_71);
nand U4989 (N_4989,N_2475,N_2274);
nor U4990 (N_4990,N_1034,N_1674);
and U4991 (N_4991,N_195,N_1510);
nor U4992 (N_4992,N_683,N_2687);
nor U4993 (N_4993,N_1788,N_615);
and U4994 (N_4994,N_666,N_1560);
or U4995 (N_4995,N_443,N_2370);
or U4996 (N_4996,N_2572,N_2991);
and U4997 (N_4997,N_1322,N_1389);
or U4998 (N_4998,N_571,N_511);
and U4999 (N_4999,N_2329,N_156);
nor U5000 (N_5000,N_2882,N_394);
or U5001 (N_5001,N_316,N_199);
nor U5002 (N_5002,N_1515,N_965);
xnor U5003 (N_5003,N_772,N_2198);
nor U5004 (N_5004,N_2837,N_2520);
xor U5005 (N_5005,N_1681,N_2925);
nor U5006 (N_5006,N_2007,N_1041);
and U5007 (N_5007,N_641,N_2792);
nor U5008 (N_5008,N_746,N_1453);
nor U5009 (N_5009,N_2345,N_211);
xnor U5010 (N_5010,N_1209,N_2335);
nand U5011 (N_5011,N_2871,N_746);
xor U5012 (N_5012,N_2643,N_75);
and U5013 (N_5013,N_505,N_1316);
or U5014 (N_5014,N_1883,N_1164);
nand U5015 (N_5015,N_199,N_2669);
and U5016 (N_5016,N_2995,N_1404);
xnor U5017 (N_5017,N_1224,N_1051);
or U5018 (N_5018,N_2021,N_1041);
nor U5019 (N_5019,N_1597,N_2420);
nor U5020 (N_5020,N_2715,N_2271);
or U5021 (N_5021,N_2318,N_709);
or U5022 (N_5022,N_218,N_1566);
nor U5023 (N_5023,N_2637,N_1769);
or U5024 (N_5024,N_2493,N_2883);
nor U5025 (N_5025,N_864,N_2835);
nand U5026 (N_5026,N_762,N_497);
nor U5027 (N_5027,N_1568,N_2238);
and U5028 (N_5028,N_2720,N_2379);
xor U5029 (N_5029,N_2573,N_1488);
nand U5030 (N_5030,N_2116,N_1877);
nand U5031 (N_5031,N_2227,N_2702);
nor U5032 (N_5032,N_2419,N_2652);
or U5033 (N_5033,N_577,N_2552);
and U5034 (N_5034,N_450,N_548);
and U5035 (N_5035,N_444,N_1003);
nor U5036 (N_5036,N_1536,N_2275);
and U5037 (N_5037,N_1646,N_2148);
nand U5038 (N_5038,N_2014,N_1879);
nor U5039 (N_5039,N_2958,N_827);
nand U5040 (N_5040,N_490,N_965);
nand U5041 (N_5041,N_870,N_2371);
xor U5042 (N_5042,N_2525,N_2587);
xor U5043 (N_5043,N_2873,N_299);
nand U5044 (N_5044,N_1701,N_2028);
nand U5045 (N_5045,N_2138,N_523);
nand U5046 (N_5046,N_721,N_1956);
or U5047 (N_5047,N_1943,N_2139);
xnor U5048 (N_5048,N_2044,N_2151);
nor U5049 (N_5049,N_1803,N_1857);
nand U5050 (N_5050,N_2096,N_2305);
xor U5051 (N_5051,N_1308,N_1124);
and U5052 (N_5052,N_895,N_201);
and U5053 (N_5053,N_2939,N_2989);
nand U5054 (N_5054,N_901,N_718);
nor U5055 (N_5055,N_1435,N_2118);
xnor U5056 (N_5056,N_1086,N_2204);
or U5057 (N_5057,N_1627,N_367);
nor U5058 (N_5058,N_78,N_1202);
xnor U5059 (N_5059,N_1899,N_677);
nand U5060 (N_5060,N_268,N_26);
and U5061 (N_5061,N_891,N_2236);
nor U5062 (N_5062,N_2627,N_2838);
or U5063 (N_5063,N_546,N_2613);
nor U5064 (N_5064,N_1287,N_529);
and U5065 (N_5065,N_2957,N_2581);
xor U5066 (N_5066,N_1525,N_2852);
or U5067 (N_5067,N_1619,N_2147);
or U5068 (N_5068,N_405,N_1364);
nand U5069 (N_5069,N_1724,N_963);
nor U5070 (N_5070,N_2469,N_1047);
xnor U5071 (N_5071,N_2776,N_1315);
xor U5072 (N_5072,N_2535,N_1689);
nand U5073 (N_5073,N_2161,N_2311);
nor U5074 (N_5074,N_2183,N_1157);
xnor U5075 (N_5075,N_1457,N_505);
nor U5076 (N_5076,N_1797,N_178);
nor U5077 (N_5077,N_1333,N_2511);
nor U5078 (N_5078,N_409,N_832);
nor U5079 (N_5079,N_2721,N_2030);
nor U5080 (N_5080,N_2338,N_1415);
nor U5081 (N_5081,N_1813,N_1989);
nand U5082 (N_5082,N_481,N_346);
nor U5083 (N_5083,N_2093,N_2200);
or U5084 (N_5084,N_2291,N_543);
or U5085 (N_5085,N_209,N_1220);
nand U5086 (N_5086,N_1739,N_1745);
nand U5087 (N_5087,N_1276,N_284);
xor U5088 (N_5088,N_167,N_377);
and U5089 (N_5089,N_2812,N_2668);
and U5090 (N_5090,N_1629,N_1507);
or U5091 (N_5091,N_258,N_1972);
and U5092 (N_5092,N_2250,N_495);
xor U5093 (N_5093,N_2251,N_1754);
nor U5094 (N_5094,N_1081,N_1345);
nand U5095 (N_5095,N_2968,N_843);
nor U5096 (N_5096,N_1965,N_300);
or U5097 (N_5097,N_930,N_2138);
and U5098 (N_5098,N_1395,N_1972);
or U5099 (N_5099,N_2110,N_397);
nand U5100 (N_5100,N_1979,N_753);
nand U5101 (N_5101,N_1356,N_306);
xor U5102 (N_5102,N_804,N_2387);
or U5103 (N_5103,N_838,N_2715);
nor U5104 (N_5104,N_2636,N_2910);
and U5105 (N_5105,N_936,N_1500);
and U5106 (N_5106,N_730,N_1348);
nor U5107 (N_5107,N_1861,N_2664);
or U5108 (N_5108,N_1476,N_2112);
and U5109 (N_5109,N_2984,N_2713);
nand U5110 (N_5110,N_188,N_1783);
nor U5111 (N_5111,N_2585,N_2776);
xor U5112 (N_5112,N_1637,N_1816);
and U5113 (N_5113,N_433,N_569);
or U5114 (N_5114,N_1519,N_1635);
and U5115 (N_5115,N_2292,N_1718);
or U5116 (N_5116,N_2346,N_662);
and U5117 (N_5117,N_2802,N_2548);
nand U5118 (N_5118,N_1107,N_639);
or U5119 (N_5119,N_1806,N_796);
or U5120 (N_5120,N_894,N_659);
nor U5121 (N_5121,N_2443,N_2826);
and U5122 (N_5122,N_2540,N_399);
xor U5123 (N_5123,N_2473,N_2280);
nor U5124 (N_5124,N_2709,N_614);
nand U5125 (N_5125,N_1937,N_2633);
or U5126 (N_5126,N_1657,N_2826);
nor U5127 (N_5127,N_1951,N_11);
or U5128 (N_5128,N_1666,N_461);
nor U5129 (N_5129,N_2906,N_1508);
xnor U5130 (N_5130,N_828,N_415);
nand U5131 (N_5131,N_1978,N_967);
nor U5132 (N_5132,N_1602,N_978);
nand U5133 (N_5133,N_2291,N_142);
xor U5134 (N_5134,N_1245,N_431);
or U5135 (N_5135,N_97,N_2453);
and U5136 (N_5136,N_1904,N_2450);
nand U5137 (N_5137,N_1972,N_1283);
nor U5138 (N_5138,N_229,N_1765);
and U5139 (N_5139,N_195,N_162);
and U5140 (N_5140,N_1037,N_1165);
nand U5141 (N_5141,N_2425,N_340);
nand U5142 (N_5142,N_1904,N_2141);
nor U5143 (N_5143,N_1819,N_2622);
and U5144 (N_5144,N_2650,N_1086);
nand U5145 (N_5145,N_1899,N_1789);
nand U5146 (N_5146,N_2743,N_2186);
or U5147 (N_5147,N_2586,N_2635);
or U5148 (N_5148,N_2442,N_2188);
nor U5149 (N_5149,N_1712,N_1951);
nor U5150 (N_5150,N_1315,N_2337);
and U5151 (N_5151,N_911,N_360);
nand U5152 (N_5152,N_2431,N_2899);
nor U5153 (N_5153,N_753,N_864);
or U5154 (N_5154,N_2401,N_264);
and U5155 (N_5155,N_2960,N_603);
nand U5156 (N_5156,N_22,N_2126);
nand U5157 (N_5157,N_1600,N_1524);
xor U5158 (N_5158,N_590,N_821);
xor U5159 (N_5159,N_593,N_17);
or U5160 (N_5160,N_6,N_1280);
and U5161 (N_5161,N_2215,N_2429);
nor U5162 (N_5162,N_2947,N_160);
and U5163 (N_5163,N_2946,N_1951);
nor U5164 (N_5164,N_82,N_131);
nor U5165 (N_5165,N_601,N_676);
nor U5166 (N_5166,N_1950,N_2928);
or U5167 (N_5167,N_1106,N_2093);
or U5168 (N_5168,N_656,N_1149);
xor U5169 (N_5169,N_368,N_1878);
xnor U5170 (N_5170,N_1905,N_1951);
xor U5171 (N_5171,N_2215,N_2817);
nand U5172 (N_5172,N_318,N_994);
nand U5173 (N_5173,N_2578,N_1579);
nand U5174 (N_5174,N_359,N_1023);
or U5175 (N_5175,N_877,N_801);
nor U5176 (N_5176,N_431,N_1996);
nor U5177 (N_5177,N_118,N_2817);
and U5178 (N_5178,N_1624,N_301);
xnor U5179 (N_5179,N_236,N_2774);
and U5180 (N_5180,N_1866,N_2916);
and U5181 (N_5181,N_502,N_762);
or U5182 (N_5182,N_2486,N_2485);
nand U5183 (N_5183,N_2064,N_1104);
nor U5184 (N_5184,N_297,N_1665);
nand U5185 (N_5185,N_2876,N_1371);
nor U5186 (N_5186,N_1862,N_857);
xor U5187 (N_5187,N_765,N_963);
and U5188 (N_5188,N_1563,N_2577);
nor U5189 (N_5189,N_2168,N_1692);
nor U5190 (N_5190,N_957,N_1040);
nor U5191 (N_5191,N_2356,N_1815);
nand U5192 (N_5192,N_114,N_2604);
and U5193 (N_5193,N_788,N_2631);
xnor U5194 (N_5194,N_2231,N_1737);
nand U5195 (N_5195,N_1554,N_2522);
or U5196 (N_5196,N_2533,N_2948);
or U5197 (N_5197,N_2377,N_2180);
xnor U5198 (N_5198,N_2089,N_2922);
nand U5199 (N_5199,N_2004,N_486);
and U5200 (N_5200,N_2818,N_753);
and U5201 (N_5201,N_2046,N_1349);
nand U5202 (N_5202,N_2642,N_2814);
nor U5203 (N_5203,N_2405,N_2846);
xor U5204 (N_5204,N_1215,N_2892);
and U5205 (N_5205,N_398,N_1063);
nor U5206 (N_5206,N_1058,N_18);
and U5207 (N_5207,N_774,N_479);
nor U5208 (N_5208,N_2894,N_1103);
nand U5209 (N_5209,N_745,N_202);
nor U5210 (N_5210,N_1476,N_1484);
and U5211 (N_5211,N_1410,N_2885);
nor U5212 (N_5212,N_2419,N_2012);
nand U5213 (N_5213,N_1670,N_2120);
nor U5214 (N_5214,N_414,N_90);
nor U5215 (N_5215,N_25,N_2047);
nand U5216 (N_5216,N_2385,N_889);
nor U5217 (N_5217,N_2455,N_1285);
and U5218 (N_5218,N_1489,N_853);
nor U5219 (N_5219,N_2652,N_1898);
nand U5220 (N_5220,N_123,N_2664);
or U5221 (N_5221,N_1247,N_1905);
or U5222 (N_5222,N_2701,N_678);
and U5223 (N_5223,N_1440,N_2531);
nor U5224 (N_5224,N_1107,N_210);
nor U5225 (N_5225,N_553,N_2440);
and U5226 (N_5226,N_2036,N_60);
nand U5227 (N_5227,N_1735,N_398);
or U5228 (N_5228,N_1062,N_921);
nand U5229 (N_5229,N_2282,N_359);
xor U5230 (N_5230,N_1753,N_582);
or U5231 (N_5231,N_1640,N_330);
or U5232 (N_5232,N_966,N_2851);
and U5233 (N_5233,N_817,N_1334);
nor U5234 (N_5234,N_2191,N_283);
or U5235 (N_5235,N_2308,N_1213);
nor U5236 (N_5236,N_2324,N_1916);
nor U5237 (N_5237,N_1239,N_880);
or U5238 (N_5238,N_2936,N_1913);
nand U5239 (N_5239,N_1413,N_435);
and U5240 (N_5240,N_936,N_2498);
nand U5241 (N_5241,N_1535,N_477);
nor U5242 (N_5242,N_1348,N_1653);
or U5243 (N_5243,N_1050,N_965);
nand U5244 (N_5244,N_312,N_2400);
xor U5245 (N_5245,N_1668,N_724);
or U5246 (N_5246,N_202,N_2563);
and U5247 (N_5247,N_2146,N_1467);
nor U5248 (N_5248,N_2193,N_2078);
and U5249 (N_5249,N_2413,N_1240);
and U5250 (N_5250,N_754,N_1155);
nand U5251 (N_5251,N_1894,N_2551);
xnor U5252 (N_5252,N_529,N_2229);
nand U5253 (N_5253,N_1641,N_2602);
or U5254 (N_5254,N_1390,N_1216);
and U5255 (N_5255,N_2952,N_481);
or U5256 (N_5256,N_1294,N_2807);
nor U5257 (N_5257,N_511,N_2061);
xor U5258 (N_5258,N_630,N_288);
nor U5259 (N_5259,N_636,N_1256);
xor U5260 (N_5260,N_1808,N_1083);
and U5261 (N_5261,N_1566,N_585);
and U5262 (N_5262,N_2332,N_2668);
and U5263 (N_5263,N_584,N_2453);
nor U5264 (N_5264,N_1014,N_2565);
nand U5265 (N_5265,N_1709,N_2723);
xor U5266 (N_5266,N_603,N_717);
nand U5267 (N_5267,N_1179,N_1574);
nand U5268 (N_5268,N_2694,N_1981);
xor U5269 (N_5269,N_1574,N_2330);
xnor U5270 (N_5270,N_2987,N_1773);
nand U5271 (N_5271,N_1129,N_476);
nand U5272 (N_5272,N_2902,N_2581);
or U5273 (N_5273,N_2294,N_1448);
nand U5274 (N_5274,N_1170,N_622);
and U5275 (N_5275,N_244,N_1870);
and U5276 (N_5276,N_851,N_140);
and U5277 (N_5277,N_2969,N_1961);
and U5278 (N_5278,N_1097,N_179);
nor U5279 (N_5279,N_2263,N_2932);
nor U5280 (N_5280,N_535,N_2747);
and U5281 (N_5281,N_2083,N_349);
nand U5282 (N_5282,N_599,N_2707);
nor U5283 (N_5283,N_1306,N_1301);
nor U5284 (N_5284,N_287,N_737);
or U5285 (N_5285,N_1221,N_2125);
or U5286 (N_5286,N_2378,N_607);
and U5287 (N_5287,N_549,N_154);
nand U5288 (N_5288,N_2843,N_2812);
and U5289 (N_5289,N_136,N_2289);
or U5290 (N_5290,N_1777,N_413);
nand U5291 (N_5291,N_1460,N_1395);
and U5292 (N_5292,N_2924,N_2308);
and U5293 (N_5293,N_82,N_826);
nor U5294 (N_5294,N_1048,N_1408);
xnor U5295 (N_5295,N_1723,N_2227);
nor U5296 (N_5296,N_2004,N_2313);
nand U5297 (N_5297,N_2729,N_1654);
or U5298 (N_5298,N_2835,N_278);
nor U5299 (N_5299,N_186,N_1459);
nor U5300 (N_5300,N_1614,N_732);
or U5301 (N_5301,N_2593,N_1800);
or U5302 (N_5302,N_711,N_1838);
nor U5303 (N_5303,N_1477,N_2449);
nor U5304 (N_5304,N_1728,N_2928);
or U5305 (N_5305,N_547,N_15);
nor U5306 (N_5306,N_1432,N_2981);
nand U5307 (N_5307,N_2634,N_239);
nor U5308 (N_5308,N_1931,N_1998);
and U5309 (N_5309,N_2730,N_2568);
or U5310 (N_5310,N_672,N_1028);
nand U5311 (N_5311,N_2896,N_2810);
or U5312 (N_5312,N_2443,N_78);
nand U5313 (N_5313,N_1681,N_736);
nand U5314 (N_5314,N_2568,N_2301);
nand U5315 (N_5315,N_790,N_2283);
nand U5316 (N_5316,N_550,N_219);
nand U5317 (N_5317,N_1384,N_2198);
nor U5318 (N_5318,N_2291,N_1003);
xnor U5319 (N_5319,N_249,N_990);
and U5320 (N_5320,N_2176,N_2334);
or U5321 (N_5321,N_1930,N_1707);
nor U5322 (N_5322,N_1754,N_375);
and U5323 (N_5323,N_1086,N_809);
nor U5324 (N_5324,N_1949,N_843);
nand U5325 (N_5325,N_752,N_2440);
and U5326 (N_5326,N_1676,N_1);
nand U5327 (N_5327,N_2132,N_2303);
nand U5328 (N_5328,N_2716,N_1752);
or U5329 (N_5329,N_1952,N_2283);
and U5330 (N_5330,N_52,N_2421);
and U5331 (N_5331,N_1628,N_468);
or U5332 (N_5332,N_2435,N_1577);
nor U5333 (N_5333,N_2505,N_1582);
nor U5334 (N_5334,N_523,N_1825);
nor U5335 (N_5335,N_1803,N_2125);
or U5336 (N_5336,N_1075,N_2988);
or U5337 (N_5337,N_595,N_431);
or U5338 (N_5338,N_532,N_2406);
and U5339 (N_5339,N_2230,N_230);
nand U5340 (N_5340,N_1032,N_262);
and U5341 (N_5341,N_2718,N_332);
nand U5342 (N_5342,N_2919,N_249);
nand U5343 (N_5343,N_2566,N_1547);
xor U5344 (N_5344,N_1742,N_178);
nand U5345 (N_5345,N_2609,N_1633);
nor U5346 (N_5346,N_2107,N_1601);
nor U5347 (N_5347,N_746,N_2399);
nand U5348 (N_5348,N_2439,N_328);
or U5349 (N_5349,N_1278,N_118);
xor U5350 (N_5350,N_1170,N_2409);
or U5351 (N_5351,N_1348,N_2205);
nand U5352 (N_5352,N_2913,N_737);
xor U5353 (N_5353,N_48,N_2325);
and U5354 (N_5354,N_2855,N_2719);
xnor U5355 (N_5355,N_43,N_2454);
nor U5356 (N_5356,N_2279,N_2005);
and U5357 (N_5357,N_1022,N_2451);
or U5358 (N_5358,N_525,N_2170);
and U5359 (N_5359,N_2054,N_1460);
xor U5360 (N_5360,N_523,N_922);
xnor U5361 (N_5361,N_1175,N_2038);
nand U5362 (N_5362,N_812,N_283);
and U5363 (N_5363,N_2278,N_1553);
nand U5364 (N_5364,N_347,N_1094);
nor U5365 (N_5365,N_428,N_184);
xnor U5366 (N_5366,N_2457,N_2379);
nor U5367 (N_5367,N_2648,N_1372);
nor U5368 (N_5368,N_1898,N_1884);
and U5369 (N_5369,N_1881,N_2613);
nand U5370 (N_5370,N_2792,N_2189);
nor U5371 (N_5371,N_860,N_1315);
and U5372 (N_5372,N_2611,N_974);
and U5373 (N_5373,N_1823,N_522);
and U5374 (N_5374,N_1609,N_547);
nor U5375 (N_5375,N_992,N_303);
nand U5376 (N_5376,N_1199,N_1510);
or U5377 (N_5377,N_924,N_358);
or U5378 (N_5378,N_54,N_631);
nor U5379 (N_5379,N_575,N_2966);
or U5380 (N_5380,N_1076,N_2578);
nand U5381 (N_5381,N_517,N_1894);
nor U5382 (N_5382,N_1707,N_1207);
or U5383 (N_5383,N_243,N_439);
nand U5384 (N_5384,N_2189,N_778);
nand U5385 (N_5385,N_2055,N_454);
and U5386 (N_5386,N_2846,N_2732);
nand U5387 (N_5387,N_1931,N_117);
and U5388 (N_5388,N_2187,N_186);
xor U5389 (N_5389,N_1205,N_2143);
xor U5390 (N_5390,N_2274,N_1770);
and U5391 (N_5391,N_1150,N_2604);
xor U5392 (N_5392,N_2546,N_1239);
xnor U5393 (N_5393,N_1757,N_2094);
and U5394 (N_5394,N_669,N_1219);
nor U5395 (N_5395,N_1603,N_1521);
and U5396 (N_5396,N_517,N_2293);
nor U5397 (N_5397,N_1779,N_1145);
nand U5398 (N_5398,N_1686,N_134);
nand U5399 (N_5399,N_425,N_254);
nand U5400 (N_5400,N_1656,N_443);
nor U5401 (N_5401,N_2228,N_1948);
nor U5402 (N_5402,N_1594,N_2738);
nand U5403 (N_5403,N_2057,N_8);
or U5404 (N_5404,N_1220,N_1694);
nand U5405 (N_5405,N_1093,N_628);
or U5406 (N_5406,N_246,N_275);
xor U5407 (N_5407,N_909,N_1411);
or U5408 (N_5408,N_1669,N_1410);
and U5409 (N_5409,N_1734,N_807);
or U5410 (N_5410,N_1033,N_412);
nor U5411 (N_5411,N_2278,N_2831);
nand U5412 (N_5412,N_1672,N_1684);
xnor U5413 (N_5413,N_671,N_2994);
and U5414 (N_5414,N_2600,N_2855);
nor U5415 (N_5415,N_429,N_774);
and U5416 (N_5416,N_1064,N_1754);
or U5417 (N_5417,N_2727,N_2203);
or U5418 (N_5418,N_2049,N_1933);
nor U5419 (N_5419,N_825,N_2934);
nand U5420 (N_5420,N_2992,N_2934);
nor U5421 (N_5421,N_1892,N_1797);
nand U5422 (N_5422,N_381,N_2347);
nand U5423 (N_5423,N_2881,N_931);
nor U5424 (N_5424,N_2232,N_1993);
and U5425 (N_5425,N_2300,N_738);
and U5426 (N_5426,N_547,N_2964);
nand U5427 (N_5427,N_2494,N_1897);
nor U5428 (N_5428,N_5,N_1592);
or U5429 (N_5429,N_884,N_186);
and U5430 (N_5430,N_2485,N_803);
nand U5431 (N_5431,N_244,N_1202);
xor U5432 (N_5432,N_2302,N_465);
nand U5433 (N_5433,N_652,N_1354);
nand U5434 (N_5434,N_1355,N_2314);
nand U5435 (N_5435,N_182,N_1347);
nor U5436 (N_5436,N_1495,N_231);
xor U5437 (N_5437,N_2209,N_2689);
or U5438 (N_5438,N_2020,N_2892);
nor U5439 (N_5439,N_880,N_641);
nor U5440 (N_5440,N_227,N_2431);
or U5441 (N_5441,N_2524,N_1619);
and U5442 (N_5442,N_2330,N_1072);
xnor U5443 (N_5443,N_611,N_1314);
or U5444 (N_5444,N_776,N_1863);
xor U5445 (N_5445,N_1012,N_1914);
and U5446 (N_5446,N_840,N_656);
or U5447 (N_5447,N_2117,N_827);
and U5448 (N_5448,N_1096,N_2651);
nand U5449 (N_5449,N_1713,N_159);
and U5450 (N_5450,N_211,N_2477);
nor U5451 (N_5451,N_1415,N_611);
or U5452 (N_5452,N_1764,N_1540);
or U5453 (N_5453,N_1342,N_630);
nand U5454 (N_5454,N_1864,N_580);
or U5455 (N_5455,N_2133,N_2522);
and U5456 (N_5456,N_794,N_79);
nand U5457 (N_5457,N_2293,N_2802);
or U5458 (N_5458,N_2227,N_2931);
or U5459 (N_5459,N_1464,N_527);
nand U5460 (N_5460,N_935,N_1156);
and U5461 (N_5461,N_1048,N_515);
and U5462 (N_5462,N_128,N_2290);
nand U5463 (N_5463,N_2748,N_2979);
or U5464 (N_5464,N_2445,N_769);
nand U5465 (N_5465,N_765,N_49);
nor U5466 (N_5466,N_244,N_2766);
and U5467 (N_5467,N_605,N_48);
or U5468 (N_5468,N_1504,N_2889);
nor U5469 (N_5469,N_2341,N_1359);
or U5470 (N_5470,N_2652,N_2276);
nand U5471 (N_5471,N_1536,N_550);
nor U5472 (N_5472,N_2201,N_2215);
or U5473 (N_5473,N_2016,N_1887);
and U5474 (N_5474,N_2710,N_1557);
nor U5475 (N_5475,N_1211,N_2272);
and U5476 (N_5476,N_286,N_308);
or U5477 (N_5477,N_1265,N_1436);
and U5478 (N_5478,N_1376,N_2116);
and U5479 (N_5479,N_1956,N_1940);
nand U5480 (N_5480,N_2588,N_547);
xnor U5481 (N_5481,N_2590,N_491);
or U5482 (N_5482,N_2810,N_2829);
xnor U5483 (N_5483,N_85,N_2129);
or U5484 (N_5484,N_1401,N_2335);
nor U5485 (N_5485,N_1089,N_1327);
nor U5486 (N_5486,N_404,N_1421);
or U5487 (N_5487,N_1333,N_2745);
and U5488 (N_5488,N_612,N_842);
nand U5489 (N_5489,N_2007,N_1575);
nor U5490 (N_5490,N_2570,N_708);
xnor U5491 (N_5491,N_163,N_2676);
or U5492 (N_5492,N_1423,N_2968);
nand U5493 (N_5493,N_1445,N_2515);
or U5494 (N_5494,N_852,N_1609);
and U5495 (N_5495,N_1658,N_914);
and U5496 (N_5496,N_1870,N_2780);
nand U5497 (N_5497,N_1806,N_193);
nor U5498 (N_5498,N_1967,N_2509);
nor U5499 (N_5499,N_647,N_416);
and U5500 (N_5500,N_1138,N_2147);
nor U5501 (N_5501,N_876,N_2878);
xor U5502 (N_5502,N_2913,N_1413);
nor U5503 (N_5503,N_2104,N_7);
nand U5504 (N_5504,N_2496,N_899);
or U5505 (N_5505,N_849,N_919);
and U5506 (N_5506,N_1153,N_2542);
xnor U5507 (N_5507,N_24,N_1970);
and U5508 (N_5508,N_256,N_2788);
xor U5509 (N_5509,N_2338,N_599);
or U5510 (N_5510,N_2452,N_461);
and U5511 (N_5511,N_881,N_174);
xnor U5512 (N_5512,N_2082,N_1678);
and U5513 (N_5513,N_1190,N_2866);
or U5514 (N_5514,N_1840,N_2414);
or U5515 (N_5515,N_2364,N_1829);
xor U5516 (N_5516,N_957,N_2672);
nor U5517 (N_5517,N_1935,N_186);
and U5518 (N_5518,N_2412,N_807);
nand U5519 (N_5519,N_1163,N_84);
xnor U5520 (N_5520,N_1155,N_2778);
nand U5521 (N_5521,N_1352,N_169);
or U5522 (N_5522,N_353,N_1269);
and U5523 (N_5523,N_2816,N_276);
nor U5524 (N_5524,N_2751,N_1955);
nor U5525 (N_5525,N_2527,N_1137);
or U5526 (N_5526,N_1340,N_1100);
and U5527 (N_5527,N_2302,N_1227);
nor U5528 (N_5528,N_2935,N_1716);
nor U5529 (N_5529,N_1025,N_1161);
or U5530 (N_5530,N_367,N_563);
nor U5531 (N_5531,N_1757,N_182);
or U5532 (N_5532,N_1163,N_1225);
and U5533 (N_5533,N_2938,N_2583);
nor U5534 (N_5534,N_1191,N_2798);
or U5535 (N_5535,N_1808,N_2384);
or U5536 (N_5536,N_30,N_1989);
nand U5537 (N_5537,N_482,N_55);
nand U5538 (N_5538,N_1585,N_2851);
nor U5539 (N_5539,N_807,N_1497);
nor U5540 (N_5540,N_1390,N_1262);
nor U5541 (N_5541,N_517,N_425);
nand U5542 (N_5542,N_1845,N_2908);
nand U5543 (N_5543,N_2222,N_2878);
or U5544 (N_5544,N_275,N_2760);
and U5545 (N_5545,N_2418,N_1953);
xor U5546 (N_5546,N_1767,N_1416);
xnor U5547 (N_5547,N_1044,N_2006);
xor U5548 (N_5548,N_156,N_99);
nor U5549 (N_5549,N_1944,N_351);
nor U5550 (N_5550,N_2853,N_1737);
or U5551 (N_5551,N_1266,N_1079);
or U5552 (N_5552,N_1550,N_1946);
xor U5553 (N_5553,N_2897,N_724);
nand U5554 (N_5554,N_2630,N_110);
nand U5555 (N_5555,N_368,N_2862);
xnor U5556 (N_5556,N_1615,N_1227);
nor U5557 (N_5557,N_755,N_83);
nor U5558 (N_5558,N_501,N_1517);
and U5559 (N_5559,N_2821,N_398);
or U5560 (N_5560,N_495,N_2248);
nor U5561 (N_5561,N_989,N_2847);
nor U5562 (N_5562,N_2004,N_208);
nand U5563 (N_5563,N_963,N_415);
and U5564 (N_5564,N_1496,N_2222);
nand U5565 (N_5565,N_2345,N_2105);
and U5566 (N_5566,N_2840,N_1222);
or U5567 (N_5567,N_2840,N_2832);
nor U5568 (N_5568,N_1744,N_1229);
or U5569 (N_5569,N_1950,N_2085);
nand U5570 (N_5570,N_1480,N_299);
or U5571 (N_5571,N_2478,N_835);
nor U5572 (N_5572,N_1846,N_1155);
nor U5573 (N_5573,N_505,N_954);
and U5574 (N_5574,N_2642,N_2226);
or U5575 (N_5575,N_2828,N_2733);
nor U5576 (N_5576,N_2276,N_1201);
nand U5577 (N_5577,N_1206,N_464);
xnor U5578 (N_5578,N_320,N_570);
xor U5579 (N_5579,N_2897,N_1354);
nor U5580 (N_5580,N_2879,N_2536);
or U5581 (N_5581,N_2257,N_2062);
or U5582 (N_5582,N_43,N_2716);
nor U5583 (N_5583,N_2921,N_1764);
nor U5584 (N_5584,N_2308,N_2953);
or U5585 (N_5585,N_353,N_1858);
and U5586 (N_5586,N_426,N_1867);
nand U5587 (N_5587,N_1038,N_1427);
or U5588 (N_5588,N_2272,N_416);
xor U5589 (N_5589,N_1981,N_1567);
or U5590 (N_5590,N_899,N_572);
and U5591 (N_5591,N_5,N_639);
and U5592 (N_5592,N_1644,N_73);
nand U5593 (N_5593,N_2418,N_1700);
and U5594 (N_5594,N_2773,N_2477);
or U5595 (N_5595,N_2788,N_1526);
nand U5596 (N_5596,N_1791,N_1585);
nand U5597 (N_5597,N_1455,N_2102);
or U5598 (N_5598,N_1624,N_2138);
and U5599 (N_5599,N_2983,N_2852);
and U5600 (N_5600,N_2983,N_506);
nand U5601 (N_5601,N_491,N_1805);
xor U5602 (N_5602,N_1292,N_2505);
and U5603 (N_5603,N_796,N_875);
nor U5604 (N_5604,N_760,N_830);
and U5605 (N_5605,N_293,N_1768);
or U5606 (N_5606,N_2096,N_2024);
nand U5607 (N_5607,N_2649,N_929);
or U5608 (N_5608,N_2721,N_2395);
or U5609 (N_5609,N_23,N_2342);
and U5610 (N_5610,N_2224,N_2141);
nor U5611 (N_5611,N_1940,N_2365);
or U5612 (N_5612,N_1480,N_289);
nor U5613 (N_5613,N_2304,N_1078);
nand U5614 (N_5614,N_821,N_1632);
and U5615 (N_5615,N_197,N_2662);
and U5616 (N_5616,N_2023,N_1823);
nand U5617 (N_5617,N_1177,N_1229);
or U5618 (N_5618,N_1298,N_2226);
nand U5619 (N_5619,N_1769,N_879);
or U5620 (N_5620,N_1581,N_703);
or U5621 (N_5621,N_1258,N_2281);
nor U5622 (N_5622,N_1049,N_2602);
nand U5623 (N_5623,N_2246,N_707);
and U5624 (N_5624,N_2472,N_2454);
and U5625 (N_5625,N_157,N_1414);
or U5626 (N_5626,N_1586,N_2035);
and U5627 (N_5627,N_190,N_2367);
nand U5628 (N_5628,N_1367,N_971);
or U5629 (N_5629,N_2239,N_1127);
and U5630 (N_5630,N_108,N_775);
or U5631 (N_5631,N_1363,N_1755);
nand U5632 (N_5632,N_372,N_1162);
nand U5633 (N_5633,N_21,N_1314);
xnor U5634 (N_5634,N_197,N_144);
nand U5635 (N_5635,N_1699,N_965);
or U5636 (N_5636,N_2595,N_1872);
and U5637 (N_5637,N_1316,N_169);
or U5638 (N_5638,N_804,N_1277);
nor U5639 (N_5639,N_1552,N_1484);
xnor U5640 (N_5640,N_2495,N_2110);
or U5641 (N_5641,N_2121,N_339);
nand U5642 (N_5642,N_2136,N_2786);
nand U5643 (N_5643,N_2995,N_1110);
nand U5644 (N_5644,N_1047,N_2250);
nor U5645 (N_5645,N_1917,N_1681);
nor U5646 (N_5646,N_1420,N_367);
or U5647 (N_5647,N_2445,N_627);
nand U5648 (N_5648,N_1586,N_2232);
and U5649 (N_5649,N_457,N_821);
and U5650 (N_5650,N_2736,N_2888);
nor U5651 (N_5651,N_920,N_929);
nor U5652 (N_5652,N_1398,N_305);
nand U5653 (N_5653,N_466,N_1048);
or U5654 (N_5654,N_2143,N_856);
nand U5655 (N_5655,N_1546,N_1458);
and U5656 (N_5656,N_2366,N_1872);
nand U5657 (N_5657,N_2547,N_2603);
xnor U5658 (N_5658,N_1542,N_325);
and U5659 (N_5659,N_177,N_1892);
or U5660 (N_5660,N_1795,N_985);
xnor U5661 (N_5661,N_2663,N_606);
xor U5662 (N_5662,N_300,N_2012);
nor U5663 (N_5663,N_1018,N_439);
nand U5664 (N_5664,N_995,N_1375);
nand U5665 (N_5665,N_2862,N_1272);
or U5666 (N_5666,N_2709,N_2345);
xor U5667 (N_5667,N_2985,N_2636);
nand U5668 (N_5668,N_316,N_1033);
nand U5669 (N_5669,N_153,N_2535);
nor U5670 (N_5670,N_1580,N_1050);
xnor U5671 (N_5671,N_1969,N_1959);
nand U5672 (N_5672,N_2465,N_2967);
or U5673 (N_5673,N_783,N_1241);
nor U5674 (N_5674,N_2864,N_37);
or U5675 (N_5675,N_1877,N_379);
nand U5676 (N_5676,N_1333,N_2110);
nand U5677 (N_5677,N_344,N_1020);
and U5678 (N_5678,N_824,N_871);
nand U5679 (N_5679,N_2573,N_2891);
nor U5680 (N_5680,N_903,N_1729);
nand U5681 (N_5681,N_272,N_58);
or U5682 (N_5682,N_1541,N_837);
and U5683 (N_5683,N_1607,N_2485);
nor U5684 (N_5684,N_1368,N_1061);
or U5685 (N_5685,N_1131,N_2963);
or U5686 (N_5686,N_2505,N_977);
or U5687 (N_5687,N_321,N_2686);
and U5688 (N_5688,N_908,N_1697);
nand U5689 (N_5689,N_1280,N_442);
nand U5690 (N_5690,N_2949,N_175);
nand U5691 (N_5691,N_2400,N_1303);
xor U5692 (N_5692,N_1745,N_156);
nand U5693 (N_5693,N_1141,N_1742);
nor U5694 (N_5694,N_1301,N_932);
nand U5695 (N_5695,N_1460,N_485);
and U5696 (N_5696,N_413,N_2028);
nand U5697 (N_5697,N_1063,N_1957);
nand U5698 (N_5698,N_1373,N_2821);
or U5699 (N_5699,N_1654,N_2134);
nand U5700 (N_5700,N_266,N_2466);
nor U5701 (N_5701,N_274,N_2405);
and U5702 (N_5702,N_1107,N_1710);
and U5703 (N_5703,N_107,N_548);
and U5704 (N_5704,N_1097,N_36);
nand U5705 (N_5705,N_443,N_255);
nand U5706 (N_5706,N_2570,N_53);
nor U5707 (N_5707,N_1538,N_2435);
or U5708 (N_5708,N_2943,N_2822);
nor U5709 (N_5709,N_608,N_1168);
or U5710 (N_5710,N_779,N_454);
nor U5711 (N_5711,N_6,N_2473);
nor U5712 (N_5712,N_2872,N_2782);
xor U5713 (N_5713,N_2760,N_1892);
or U5714 (N_5714,N_168,N_690);
and U5715 (N_5715,N_2438,N_2718);
nand U5716 (N_5716,N_945,N_2091);
nand U5717 (N_5717,N_2223,N_2930);
nand U5718 (N_5718,N_749,N_826);
nor U5719 (N_5719,N_2247,N_2725);
or U5720 (N_5720,N_1320,N_970);
and U5721 (N_5721,N_7,N_474);
nand U5722 (N_5722,N_2170,N_984);
and U5723 (N_5723,N_544,N_2943);
nand U5724 (N_5724,N_1455,N_304);
and U5725 (N_5725,N_1421,N_809);
nand U5726 (N_5726,N_574,N_754);
nor U5727 (N_5727,N_216,N_2250);
xnor U5728 (N_5728,N_573,N_2381);
or U5729 (N_5729,N_1496,N_269);
and U5730 (N_5730,N_759,N_1735);
or U5731 (N_5731,N_2022,N_2119);
xnor U5732 (N_5732,N_1991,N_679);
nor U5733 (N_5733,N_1048,N_440);
xnor U5734 (N_5734,N_1674,N_952);
or U5735 (N_5735,N_2380,N_2779);
nand U5736 (N_5736,N_1490,N_1299);
and U5737 (N_5737,N_2170,N_2205);
xnor U5738 (N_5738,N_998,N_2654);
nor U5739 (N_5739,N_762,N_2698);
nor U5740 (N_5740,N_2424,N_1747);
nand U5741 (N_5741,N_1613,N_1616);
or U5742 (N_5742,N_1792,N_755);
nand U5743 (N_5743,N_614,N_2683);
and U5744 (N_5744,N_83,N_1359);
nor U5745 (N_5745,N_2021,N_2674);
nor U5746 (N_5746,N_1520,N_1617);
and U5747 (N_5747,N_82,N_2976);
nor U5748 (N_5748,N_1574,N_401);
and U5749 (N_5749,N_836,N_2505);
nand U5750 (N_5750,N_127,N_718);
xor U5751 (N_5751,N_2017,N_307);
and U5752 (N_5752,N_1248,N_1849);
xnor U5753 (N_5753,N_689,N_1158);
or U5754 (N_5754,N_722,N_670);
or U5755 (N_5755,N_1027,N_2647);
or U5756 (N_5756,N_282,N_2420);
or U5757 (N_5757,N_25,N_1985);
xor U5758 (N_5758,N_1432,N_506);
nor U5759 (N_5759,N_2550,N_1133);
nor U5760 (N_5760,N_1830,N_1940);
xnor U5761 (N_5761,N_2583,N_314);
nor U5762 (N_5762,N_596,N_240);
nand U5763 (N_5763,N_1369,N_1082);
xnor U5764 (N_5764,N_920,N_2839);
or U5765 (N_5765,N_2490,N_427);
and U5766 (N_5766,N_1198,N_2302);
nor U5767 (N_5767,N_2019,N_2514);
xor U5768 (N_5768,N_2655,N_686);
and U5769 (N_5769,N_2017,N_2987);
or U5770 (N_5770,N_750,N_692);
nand U5771 (N_5771,N_332,N_366);
xor U5772 (N_5772,N_2675,N_169);
xnor U5773 (N_5773,N_1291,N_2813);
nand U5774 (N_5774,N_2681,N_598);
or U5775 (N_5775,N_915,N_1944);
or U5776 (N_5776,N_2162,N_1199);
nand U5777 (N_5777,N_1650,N_1665);
nand U5778 (N_5778,N_1226,N_557);
nand U5779 (N_5779,N_277,N_531);
nor U5780 (N_5780,N_2223,N_962);
and U5781 (N_5781,N_2135,N_1080);
and U5782 (N_5782,N_119,N_2750);
nor U5783 (N_5783,N_1151,N_1649);
xor U5784 (N_5784,N_2945,N_672);
nor U5785 (N_5785,N_2961,N_190);
nand U5786 (N_5786,N_2359,N_2422);
or U5787 (N_5787,N_1334,N_551);
nor U5788 (N_5788,N_2776,N_2229);
and U5789 (N_5789,N_1394,N_1838);
and U5790 (N_5790,N_19,N_834);
or U5791 (N_5791,N_680,N_991);
nand U5792 (N_5792,N_977,N_2188);
or U5793 (N_5793,N_2033,N_2175);
nor U5794 (N_5794,N_925,N_559);
nand U5795 (N_5795,N_2445,N_1793);
and U5796 (N_5796,N_377,N_1736);
nand U5797 (N_5797,N_88,N_2407);
or U5798 (N_5798,N_2337,N_1);
nor U5799 (N_5799,N_1511,N_1282);
nand U5800 (N_5800,N_1139,N_445);
nand U5801 (N_5801,N_14,N_1421);
or U5802 (N_5802,N_2748,N_2364);
nand U5803 (N_5803,N_1843,N_569);
xnor U5804 (N_5804,N_2744,N_1706);
nand U5805 (N_5805,N_2764,N_1168);
xor U5806 (N_5806,N_699,N_1185);
xnor U5807 (N_5807,N_2983,N_925);
nand U5808 (N_5808,N_2728,N_1489);
nor U5809 (N_5809,N_1565,N_1271);
xor U5810 (N_5810,N_2372,N_242);
nand U5811 (N_5811,N_2508,N_530);
or U5812 (N_5812,N_2018,N_1333);
and U5813 (N_5813,N_2387,N_163);
nand U5814 (N_5814,N_245,N_2383);
and U5815 (N_5815,N_2220,N_506);
and U5816 (N_5816,N_334,N_647);
nor U5817 (N_5817,N_2898,N_1153);
xnor U5818 (N_5818,N_1138,N_1859);
nor U5819 (N_5819,N_2291,N_887);
nand U5820 (N_5820,N_2316,N_122);
nor U5821 (N_5821,N_133,N_1336);
nand U5822 (N_5822,N_2572,N_1158);
and U5823 (N_5823,N_2030,N_1978);
nor U5824 (N_5824,N_1105,N_1747);
nand U5825 (N_5825,N_1188,N_254);
nand U5826 (N_5826,N_1793,N_2957);
and U5827 (N_5827,N_665,N_1290);
nor U5828 (N_5828,N_1328,N_1474);
or U5829 (N_5829,N_1077,N_176);
nor U5830 (N_5830,N_2335,N_2120);
or U5831 (N_5831,N_640,N_2284);
nand U5832 (N_5832,N_6,N_2771);
or U5833 (N_5833,N_2409,N_30);
nand U5834 (N_5834,N_202,N_490);
nor U5835 (N_5835,N_2290,N_46);
nand U5836 (N_5836,N_560,N_2777);
or U5837 (N_5837,N_1182,N_1156);
xor U5838 (N_5838,N_2010,N_2739);
nand U5839 (N_5839,N_2104,N_443);
and U5840 (N_5840,N_2093,N_490);
nor U5841 (N_5841,N_1564,N_362);
or U5842 (N_5842,N_1056,N_2834);
and U5843 (N_5843,N_2390,N_2070);
xnor U5844 (N_5844,N_265,N_559);
nand U5845 (N_5845,N_1351,N_2687);
nand U5846 (N_5846,N_1497,N_832);
and U5847 (N_5847,N_83,N_1211);
and U5848 (N_5848,N_2454,N_422);
nand U5849 (N_5849,N_1692,N_2874);
nor U5850 (N_5850,N_649,N_1511);
and U5851 (N_5851,N_2754,N_2716);
or U5852 (N_5852,N_1274,N_85);
nand U5853 (N_5853,N_2635,N_1719);
nor U5854 (N_5854,N_1693,N_578);
xnor U5855 (N_5855,N_2220,N_1838);
or U5856 (N_5856,N_1835,N_1113);
nor U5857 (N_5857,N_1442,N_522);
or U5858 (N_5858,N_2895,N_1496);
or U5859 (N_5859,N_599,N_2107);
nand U5860 (N_5860,N_1575,N_592);
nor U5861 (N_5861,N_2430,N_459);
and U5862 (N_5862,N_2165,N_2901);
or U5863 (N_5863,N_800,N_2329);
nor U5864 (N_5864,N_2431,N_6);
nor U5865 (N_5865,N_869,N_751);
nand U5866 (N_5866,N_1699,N_2305);
nor U5867 (N_5867,N_2936,N_2088);
or U5868 (N_5868,N_352,N_1654);
nand U5869 (N_5869,N_515,N_2361);
nand U5870 (N_5870,N_1196,N_23);
and U5871 (N_5871,N_1944,N_1640);
xnor U5872 (N_5872,N_8,N_2445);
and U5873 (N_5873,N_552,N_1689);
and U5874 (N_5874,N_465,N_2147);
or U5875 (N_5875,N_827,N_634);
xor U5876 (N_5876,N_2967,N_2755);
and U5877 (N_5877,N_1433,N_1993);
nor U5878 (N_5878,N_886,N_1210);
xor U5879 (N_5879,N_2146,N_673);
nor U5880 (N_5880,N_1724,N_1136);
and U5881 (N_5881,N_83,N_2599);
nand U5882 (N_5882,N_843,N_1548);
nand U5883 (N_5883,N_2750,N_2184);
or U5884 (N_5884,N_1640,N_1496);
nand U5885 (N_5885,N_2469,N_1236);
nor U5886 (N_5886,N_2745,N_2620);
nor U5887 (N_5887,N_1504,N_873);
xnor U5888 (N_5888,N_1680,N_452);
nand U5889 (N_5889,N_2998,N_597);
and U5890 (N_5890,N_629,N_1371);
and U5891 (N_5891,N_2802,N_1503);
and U5892 (N_5892,N_1893,N_909);
or U5893 (N_5893,N_2039,N_2461);
nand U5894 (N_5894,N_2641,N_437);
nor U5895 (N_5895,N_352,N_1150);
nor U5896 (N_5896,N_967,N_24);
nor U5897 (N_5897,N_1020,N_2500);
and U5898 (N_5898,N_1711,N_540);
or U5899 (N_5899,N_2391,N_732);
xor U5900 (N_5900,N_1473,N_333);
xor U5901 (N_5901,N_2887,N_2301);
and U5902 (N_5902,N_376,N_2566);
and U5903 (N_5903,N_1098,N_2979);
and U5904 (N_5904,N_1323,N_2586);
and U5905 (N_5905,N_2938,N_2295);
nand U5906 (N_5906,N_1869,N_720);
nand U5907 (N_5907,N_1145,N_1231);
and U5908 (N_5908,N_169,N_1802);
or U5909 (N_5909,N_2153,N_42);
and U5910 (N_5910,N_1318,N_2606);
and U5911 (N_5911,N_2535,N_2307);
or U5912 (N_5912,N_1798,N_426);
or U5913 (N_5913,N_33,N_2157);
nor U5914 (N_5914,N_2556,N_1766);
and U5915 (N_5915,N_1008,N_35);
nand U5916 (N_5916,N_2277,N_1300);
and U5917 (N_5917,N_1901,N_2513);
or U5918 (N_5918,N_2389,N_1080);
nand U5919 (N_5919,N_474,N_2330);
nand U5920 (N_5920,N_314,N_721);
nand U5921 (N_5921,N_2855,N_854);
nor U5922 (N_5922,N_2677,N_80);
nor U5923 (N_5923,N_2092,N_2558);
nor U5924 (N_5924,N_2642,N_1784);
or U5925 (N_5925,N_2546,N_2849);
nor U5926 (N_5926,N_2736,N_2356);
nand U5927 (N_5927,N_1184,N_1049);
or U5928 (N_5928,N_2555,N_416);
nor U5929 (N_5929,N_263,N_116);
nand U5930 (N_5930,N_671,N_1267);
or U5931 (N_5931,N_636,N_1940);
nor U5932 (N_5932,N_1131,N_998);
nand U5933 (N_5933,N_1921,N_1787);
and U5934 (N_5934,N_1527,N_2397);
or U5935 (N_5935,N_941,N_428);
nand U5936 (N_5936,N_1315,N_870);
or U5937 (N_5937,N_1204,N_2467);
or U5938 (N_5938,N_2821,N_1270);
or U5939 (N_5939,N_2369,N_2580);
nand U5940 (N_5940,N_799,N_53);
and U5941 (N_5941,N_1887,N_41);
nand U5942 (N_5942,N_1368,N_1048);
and U5943 (N_5943,N_253,N_2315);
nand U5944 (N_5944,N_873,N_2800);
xnor U5945 (N_5945,N_151,N_992);
and U5946 (N_5946,N_2778,N_1517);
nor U5947 (N_5947,N_2445,N_1446);
or U5948 (N_5948,N_748,N_2312);
nor U5949 (N_5949,N_696,N_2852);
and U5950 (N_5950,N_2251,N_1013);
nand U5951 (N_5951,N_1184,N_2660);
or U5952 (N_5952,N_256,N_935);
or U5953 (N_5953,N_2661,N_2125);
nor U5954 (N_5954,N_663,N_2144);
and U5955 (N_5955,N_883,N_2222);
nor U5956 (N_5956,N_2856,N_2762);
xnor U5957 (N_5957,N_123,N_927);
nand U5958 (N_5958,N_2699,N_2997);
or U5959 (N_5959,N_2951,N_457);
nand U5960 (N_5960,N_1426,N_1314);
nand U5961 (N_5961,N_2447,N_718);
nor U5962 (N_5962,N_1002,N_1186);
and U5963 (N_5963,N_1473,N_76);
nor U5964 (N_5964,N_2073,N_1089);
and U5965 (N_5965,N_2584,N_2886);
nor U5966 (N_5966,N_2967,N_1575);
or U5967 (N_5967,N_1984,N_1580);
xor U5968 (N_5968,N_1648,N_656);
or U5969 (N_5969,N_256,N_1398);
nand U5970 (N_5970,N_2154,N_6);
xor U5971 (N_5971,N_2575,N_2658);
and U5972 (N_5972,N_1656,N_163);
and U5973 (N_5973,N_1284,N_1034);
and U5974 (N_5974,N_20,N_594);
nand U5975 (N_5975,N_1011,N_2962);
or U5976 (N_5976,N_794,N_1190);
or U5977 (N_5977,N_2729,N_1807);
or U5978 (N_5978,N_809,N_1873);
nand U5979 (N_5979,N_1617,N_2880);
nand U5980 (N_5980,N_1183,N_129);
nand U5981 (N_5981,N_469,N_2007);
and U5982 (N_5982,N_2820,N_1501);
nor U5983 (N_5983,N_2338,N_2187);
nor U5984 (N_5984,N_2520,N_942);
nand U5985 (N_5985,N_1851,N_1359);
and U5986 (N_5986,N_562,N_2805);
and U5987 (N_5987,N_1031,N_655);
nand U5988 (N_5988,N_2209,N_1421);
or U5989 (N_5989,N_1749,N_811);
and U5990 (N_5990,N_786,N_178);
nor U5991 (N_5991,N_1907,N_1220);
nor U5992 (N_5992,N_456,N_2902);
nor U5993 (N_5993,N_2643,N_139);
and U5994 (N_5994,N_1537,N_275);
nand U5995 (N_5995,N_2620,N_1826);
nor U5996 (N_5996,N_224,N_708);
or U5997 (N_5997,N_2898,N_258);
and U5998 (N_5998,N_2461,N_2270);
nor U5999 (N_5999,N_61,N_2608);
nor U6000 (N_6000,N_5064,N_4015);
and U6001 (N_6001,N_5724,N_5694);
and U6002 (N_6002,N_5225,N_4953);
and U6003 (N_6003,N_4142,N_3636);
or U6004 (N_6004,N_5433,N_3880);
and U6005 (N_6005,N_4014,N_3143);
nand U6006 (N_6006,N_4501,N_3674);
nor U6007 (N_6007,N_5213,N_5691);
nor U6008 (N_6008,N_4235,N_5012);
and U6009 (N_6009,N_5134,N_4489);
nand U6010 (N_6010,N_3995,N_4960);
and U6011 (N_6011,N_3212,N_4423);
or U6012 (N_6012,N_5574,N_3946);
or U6013 (N_6013,N_4279,N_3399);
nand U6014 (N_6014,N_4356,N_5478);
nor U6015 (N_6015,N_4633,N_5749);
nor U6016 (N_6016,N_4940,N_5952);
or U6017 (N_6017,N_5778,N_3067);
nand U6018 (N_6018,N_4944,N_5455);
nand U6019 (N_6019,N_3698,N_4078);
nor U6020 (N_6020,N_3099,N_5401);
and U6021 (N_6021,N_3232,N_3227);
or U6022 (N_6022,N_5877,N_4867);
nor U6023 (N_6023,N_3510,N_4201);
nand U6024 (N_6024,N_5886,N_3870);
nand U6025 (N_6025,N_3216,N_5775);
nor U6026 (N_6026,N_3779,N_3860);
nor U6027 (N_6027,N_4318,N_4337);
and U6028 (N_6028,N_4568,N_5638);
xor U6029 (N_6029,N_5634,N_3200);
nor U6030 (N_6030,N_3245,N_3097);
nand U6031 (N_6031,N_5677,N_4473);
and U6032 (N_6032,N_5227,N_3693);
nand U6033 (N_6033,N_5828,N_4150);
nand U6034 (N_6034,N_4796,N_3699);
and U6035 (N_6035,N_4663,N_3569);
nor U6036 (N_6036,N_4052,N_3148);
nand U6037 (N_6037,N_5335,N_5649);
and U6038 (N_6038,N_4515,N_5395);
xnor U6039 (N_6039,N_3126,N_5743);
or U6040 (N_6040,N_5562,N_3804);
or U6041 (N_6041,N_4726,N_3061);
nand U6042 (N_6042,N_5945,N_3554);
or U6043 (N_6043,N_3602,N_5275);
and U6044 (N_6044,N_3764,N_3685);
or U6045 (N_6045,N_5827,N_4116);
or U6046 (N_6046,N_3401,N_5757);
nand U6047 (N_6047,N_5417,N_5509);
and U6048 (N_6048,N_4479,N_5760);
nand U6049 (N_6049,N_3701,N_5473);
and U6050 (N_6050,N_4065,N_5390);
nor U6051 (N_6051,N_3335,N_5198);
or U6052 (N_6052,N_5246,N_4163);
nand U6053 (N_6053,N_5502,N_5815);
xor U6054 (N_6054,N_3956,N_5533);
nand U6055 (N_6055,N_5920,N_5072);
or U6056 (N_6056,N_4708,N_4300);
and U6057 (N_6057,N_4781,N_5239);
nor U6058 (N_6058,N_5821,N_3262);
nor U6059 (N_6059,N_3840,N_4918);
and U6060 (N_6060,N_3937,N_3523);
nor U6061 (N_6061,N_4763,N_5273);
or U6062 (N_6062,N_5159,N_5494);
and U6063 (N_6063,N_3219,N_4657);
nand U6064 (N_6064,N_5705,N_4553);
nand U6065 (N_6065,N_4689,N_5863);
nor U6066 (N_6066,N_3953,N_3588);
nor U6067 (N_6067,N_4873,N_3711);
nor U6068 (N_6068,N_3084,N_4248);
xor U6069 (N_6069,N_3958,N_5481);
nor U6070 (N_6070,N_4125,N_4123);
or U6071 (N_6071,N_5497,N_4577);
nand U6072 (N_6072,N_5862,N_5936);
nand U6073 (N_6073,N_3844,N_5950);
nand U6074 (N_6074,N_3120,N_5267);
nand U6075 (N_6075,N_5905,N_3482);
and U6076 (N_6076,N_3154,N_4081);
nor U6077 (N_6077,N_3225,N_3773);
or U6078 (N_6078,N_5324,N_4878);
xnor U6079 (N_6079,N_5105,N_3975);
and U6080 (N_6080,N_5088,N_4244);
nor U6081 (N_6081,N_3119,N_4250);
nand U6082 (N_6082,N_3891,N_4310);
nand U6083 (N_6083,N_4406,N_4897);
nor U6084 (N_6084,N_5908,N_4676);
or U6085 (N_6085,N_4110,N_4358);
nand U6086 (N_6086,N_4634,N_4478);
and U6087 (N_6087,N_3258,N_5291);
or U6088 (N_6088,N_3996,N_3866);
nand U6089 (N_6089,N_4916,N_5600);
or U6090 (N_6090,N_3207,N_3717);
xnor U6091 (N_6091,N_5988,N_5697);
and U6092 (N_6092,N_4542,N_3578);
or U6093 (N_6093,N_5116,N_4044);
or U6094 (N_6094,N_3793,N_5621);
and U6095 (N_6095,N_4107,N_5255);
or U6096 (N_6096,N_5791,N_5445);
nand U6097 (N_6097,N_3352,N_5276);
nor U6098 (N_6098,N_3090,N_4105);
or U6099 (N_6099,N_5949,N_5575);
and U6100 (N_6100,N_5491,N_4359);
and U6101 (N_6101,N_4742,N_5327);
nor U6102 (N_6102,N_5144,N_5178);
or U6103 (N_6103,N_4745,N_4412);
and U6104 (N_6104,N_3679,N_3576);
or U6105 (N_6105,N_5034,N_5103);
and U6106 (N_6106,N_3177,N_3849);
and U6107 (N_6107,N_5293,N_4834);
nand U6108 (N_6108,N_4050,N_3398);
or U6109 (N_6109,N_5939,N_5305);
or U6110 (N_6110,N_4186,N_4367);
nand U6111 (N_6111,N_5850,N_5902);
nor U6112 (N_6112,N_4283,N_5205);
nand U6113 (N_6113,N_5814,N_3312);
and U6114 (N_6114,N_3038,N_4465);
or U6115 (N_6115,N_4270,N_3051);
or U6116 (N_6116,N_4806,N_4573);
nor U6117 (N_6117,N_5471,N_4938);
xor U6118 (N_6118,N_5832,N_5215);
xnor U6119 (N_6119,N_5851,N_5182);
nor U6120 (N_6120,N_4333,N_5256);
nand U6121 (N_6121,N_3281,N_4472);
and U6122 (N_6122,N_5953,N_5216);
or U6123 (N_6123,N_5762,N_4089);
and U6124 (N_6124,N_4626,N_5984);
or U6125 (N_6125,N_3354,N_3323);
nor U6126 (N_6126,N_4994,N_5260);
and U6127 (N_6127,N_5448,N_4240);
and U6128 (N_6128,N_5113,N_3350);
nand U6129 (N_6129,N_5410,N_4450);
or U6130 (N_6130,N_4857,N_5752);
or U6131 (N_6131,N_5517,N_5195);
nor U6132 (N_6132,N_3533,N_4507);
nand U6133 (N_6133,N_5413,N_3722);
nor U6134 (N_6134,N_5641,N_4073);
nand U6135 (N_6135,N_4389,N_3759);
and U6136 (N_6136,N_5364,N_3729);
or U6137 (N_6137,N_4364,N_5929);
nand U6138 (N_6138,N_4332,N_3414);
or U6139 (N_6139,N_3279,N_5711);
and U6140 (N_6140,N_3425,N_5024);
nor U6141 (N_6141,N_5842,N_4809);
and U6142 (N_6142,N_5858,N_5896);
or U6143 (N_6143,N_3089,N_3182);
nand U6144 (N_6144,N_5067,N_5405);
and U6145 (N_6145,N_5015,N_3596);
xor U6146 (N_6146,N_3893,N_5385);
and U6147 (N_6147,N_3696,N_5132);
or U6148 (N_6148,N_3951,N_3978);
or U6149 (N_6149,N_3908,N_3678);
or U6150 (N_6150,N_4481,N_3074);
or U6151 (N_6151,N_4506,N_3430);
xnor U6152 (N_6152,N_4314,N_4509);
or U6153 (N_6153,N_4503,N_3725);
nor U6154 (N_6154,N_4625,N_3771);
or U6155 (N_6155,N_3500,N_5788);
and U6156 (N_6156,N_3303,N_3113);
xnor U6157 (N_6157,N_4870,N_4524);
xor U6158 (N_6158,N_4146,N_4949);
nor U6159 (N_6159,N_4903,N_4339);
and U6160 (N_6160,N_5095,N_4043);
or U6161 (N_6161,N_4579,N_4714);
or U6162 (N_6162,N_3502,N_4609);
nor U6163 (N_6163,N_4425,N_4232);
or U6164 (N_6164,N_3986,N_3364);
xor U6165 (N_6165,N_5716,N_4593);
or U6166 (N_6166,N_3030,N_4414);
and U6167 (N_6167,N_4770,N_3733);
or U6168 (N_6168,N_5152,N_3691);
xnor U6169 (N_6169,N_5767,N_3020);
or U6170 (N_6170,N_3315,N_5874);
and U6171 (N_6171,N_4346,N_3229);
or U6172 (N_6172,N_3540,N_5758);
and U6173 (N_6173,N_4894,N_3230);
nand U6174 (N_6174,N_4914,N_3104);
or U6175 (N_6175,N_3585,N_5895);
or U6176 (N_6176,N_3014,N_5200);
nand U6177 (N_6177,N_5352,N_4119);
and U6178 (N_6178,N_5354,N_4607);
nand U6179 (N_6179,N_5386,N_3651);
nand U6180 (N_6180,N_4212,N_3171);
nand U6181 (N_6181,N_5991,N_3034);
nor U6182 (N_6182,N_4521,N_4302);
xor U6183 (N_6183,N_3121,N_5943);
or U6184 (N_6184,N_4269,N_4145);
xnor U6185 (N_6185,N_3675,N_5302);
xor U6186 (N_6186,N_3170,N_4251);
nor U6187 (N_6187,N_5542,N_4988);
nor U6188 (N_6188,N_3826,N_4736);
nor U6189 (N_6189,N_3606,N_5313);
or U6190 (N_6190,N_5903,N_4608);
nor U6191 (N_6191,N_5438,N_4751);
nand U6192 (N_6192,N_3950,N_4924);
and U6193 (N_6193,N_3663,N_5566);
and U6194 (N_6194,N_5393,N_3314);
nor U6195 (N_6195,N_5681,N_3808);
nor U6196 (N_6196,N_3261,N_5240);
nor U6197 (N_6197,N_5882,N_5613);
xor U6198 (N_6198,N_4945,N_5278);
and U6199 (N_6199,N_5578,N_3235);
or U6200 (N_6200,N_4784,N_5781);
nand U6201 (N_6201,N_5308,N_3457);
or U6202 (N_6202,N_4828,N_3224);
nand U6203 (N_6203,N_3993,N_3254);
or U6204 (N_6204,N_3060,N_3562);
or U6205 (N_6205,N_3484,N_3290);
and U6206 (N_6206,N_5014,N_3057);
and U6207 (N_6207,N_4650,N_4740);
and U6208 (N_6208,N_3647,N_3491);
nor U6209 (N_6209,N_3412,N_5328);
or U6210 (N_6210,N_4586,N_4669);
nand U6211 (N_6211,N_5346,N_5028);
and U6212 (N_6212,N_3183,N_3980);
nand U6213 (N_6213,N_4833,N_4535);
or U6214 (N_6214,N_4243,N_4217);
or U6215 (N_6215,N_5362,N_3496);
or U6216 (N_6216,N_3546,N_5869);
nor U6217 (N_6217,N_3580,N_4651);
and U6218 (N_6218,N_3468,N_5234);
nor U6219 (N_6219,N_3659,N_5114);
nand U6220 (N_6220,N_5338,N_5830);
nor U6221 (N_6221,N_3851,N_3267);
nor U6222 (N_6222,N_3452,N_4816);
nand U6223 (N_6223,N_5204,N_4207);
nor U6224 (N_6224,N_5053,N_3926);
nand U6225 (N_6225,N_4868,N_5996);
and U6226 (N_6226,N_4559,N_5449);
nand U6227 (N_6227,N_3334,N_3861);
or U6228 (N_6228,N_3718,N_5027);
nand U6229 (N_6229,N_3370,N_5763);
or U6230 (N_6230,N_4746,N_4055);
nand U6231 (N_6231,N_4376,N_5564);
nor U6232 (N_6232,N_4200,N_4999);
or U6233 (N_6233,N_3454,N_3018);
xnor U6234 (N_6234,N_3820,N_4848);
and U6235 (N_6235,N_4902,N_4036);
and U6236 (N_6236,N_3048,N_5075);
xnor U6237 (N_6237,N_4812,N_5357);
nor U6238 (N_6238,N_5165,N_5203);
xor U6239 (N_6239,N_4261,N_4645);
nor U6240 (N_6240,N_5639,N_3927);
nor U6241 (N_6241,N_4854,N_5777);
xor U6242 (N_6242,N_4672,N_5056);
nor U6243 (N_6243,N_5129,N_3702);
xnor U6244 (N_6244,N_4908,N_4589);
nand U6245 (N_6245,N_4907,N_4749);
nor U6246 (N_6246,N_3371,N_3758);
and U6247 (N_6247,N_4268,N_4215);
and U6248 (N_6248,N_3406,N_5987);
and U6249 (N_6249,N_5706,N_3260);
and U6250 (N_6250,N_5847,N_3797);
or U6251 (N_6251,N_4785,N_4292);
and U6252 (N_6252,N_5817,N_4305);
nand U6253 (N_6253,N_5373,N_5342);
and U6254 (N_6254,N_3210,N_3932);
nand U6255 (N_6255,N_5212,N_4622);
xnor U6256 (N_6256,N_3710,N_5477);
nor U6257 (N_6257,N_5787,N_3650);
nand U6258 (N_6258,N_3521,N_3742);
and U6259 (N_6259,N_4466,N_4939);
nor U6260 (N_6260,N_5748,N_4952);
or U6261 (N_6261,N_3751,N_5507);
or U6262 (N_6262,N_5859,N_3690);
nand U6263 (N_6263,N_3013,N_3007);
and U6264 (N_6264,N_3150,N_5286);
nand U6265 (N_6265,N_3103,N_4502);
nand U6266 (N_6266,N_4467,N_4344);
nand U6267 (N_6267,N_3041,N_5932);
and U6268 (N_6268,N_3556,N_4071);
or U6269 (N_6269,N_3108,N_5604);
and U6270 (N_6270,N_3242,N_3466);
nor U6271 (N_6271,N_5210,N_4840);
and U6272 (N_6272,N_4104,N_4538);
nand U6273 (N_6273,N_3898,N_4741);
nor U6274 (N_6274,N_3599,N_5661);
nor U6275 (N_6275,N_3786,N_5111);
nor U6276 (N_6276,N_4716,N_5051);
nor U6277 (N_6277,N_3582,N_3577);
nor U6278 (N_6278,N_5321,N_4446);
or U6279 (N_6279,N_5146,N_3363);
or U6280 (N_6280,N_4427,N_4764);
or U6281 (N_6281,N_3351,N_3895);
xnor U6282 (N_6282,N_5675,N_5557);
and U6283 (N_6283,N_5617,N_4169);
or U6284 (N_6284,N_3700,N_3811);
or U6285 (N_6285,N_3519,N_3244);
and U6286 (N_6286,N_5403,N_5538);
or U6287 (N_6287,N_3716,N_3744);
xor U6288 (N_6288,N_3522,N_3823);
or U6289 (N_6289,N_4004,N_5893);
nor U6290 (N_6290,N_5504,N_5214);
or U6291 (N_6291,N_3283,N_5942);
nor U6292 (N_6292,N_3854,N_5539);
nand U6293 (N_6293,N_3903,N_4516);
nor U6294 (N_6294,N_4133,N_5086);
nand U6295 (N_6295,N_4564,N_3324);
or U6296 (N_6296,N_5220,N_4199);
nand U6297 (N_6297,N_4368,N_3667);
and U6298 (N_6298,N_3963,N_4421);
or U6299 (N_6299,N_4101,N_4003);
and U6300 (N_6300,N_3535,N_4881);
or U6301 (N_6301,N_5124,N_3044);
and U6302 (N_6302,N_3465,N_3033);
and U6303 (N_6303,N_3055,N_5732);
and U6304 (N_6304,N_4681,N_4259);
nor U6305 (N_6305,N_4578,N_3257);
nand U6306 (N_6306,N_4852,N_3941);
and U6307 (N_6307,N_5710,N_5516);
nor U6308 (N_6308,N_4748,N_4487);
or U6309 (N_6309,N_4700,N_3217);
or U6310 (N_6310,N_5868,N_3526);
and U6311 (N_6311,N_4449,N_4590);
or U6312 (N_6312,N_4468,N_3876);
or U6313 (N_6313,N_5367,N_3874);
nor U6314 (N_6314,N_5892,N_5599);
xor U6315 (N_6315,N_5148,N_4025);
nand U6316 (N_6316,N_4001,N_3096);
xor U6317 (N_6317,N_3933,N_5805);
or U6318 (N_6318,N_5921,N_4743);
nand U6319 (N_6319,N_5085,N_5699);
nand U6320 (N_6320,N_4866,N_5147);
nand U6321 (N_6321,N_3868,N_4042);
or U6322 (N_6322,N_5059,N_5655);
nor U6323 (N_6323,N_4678,N_3136);
or U6324 (N_6324,N_3991,N_5138);
nor U6325 (N_6325,N_3709,N_3458);
or U6326 (N_6326,N_4188,N_3656);
or U6327 (N_6327,N_3112,N_3648);
and U6328 (N_6328,N_4419,N_4418);
and U6329 (N_6329,N_5684,N_3288);
nor U6330 (N_6330,N_4638,N_4301);
nand U6331 (N_6331,N_3091,N_4992);
and U6332 (N_6332,N_4080,N_3316);
or U6333 (N_6333,N_4532,N_3568);
and U6334 (N_6334,N_5495,N_3552);
xor U6335 (N_6335,N_5126,N_3439);
nor U6336 (N_6336,N_5512,N_3503);
xor U6337 (N_6337,N_4031,N_3271);
and U6338 (N_6338,N_3459,N_5408);
nor U6339 (N_6339,N_4889,N_5443);
nor U6340 (N_6340,N_4263,N_3419);
or U6341 (N_6341,N_4288,N_4216);
and U6342 (N_6342,N_4218,N_3715);
and U6343 (N_6343,N_3138,N_3175);
and U6344 (N_6344,N_5631,N_4159);
or U6345 (N_6345,N_3087,N_5946);
nor U6346 (N_6346,N_4138,N_4331);
or U6347 (N_6347,N_5041,N_5727);
and U6348 (N_6348,N_3997,N_3407);
or U6349 (N_6349,N_5570,N_5174);
nor U6350 (N_6350,N_5796,N_5585);
or U6351 (N_6351,N_5556,N_3449);
nor U6352 (N_6352,N_4006,N_3240);
or U6353 (N_6353,N_5836,N_3118);
nand U6354 (N_6354,N_3321,N_5567);
or U6355 (N_6355,N_3079,N_5436);
and U6356 (N_6356,N_5518,N_3762);
nor U6357 (N_6357,N_4998,N_4082);
xor U6358 (N_6358,N_3536,N_3945);
or U6359 (N_6359,N_3890,N_3174);
or U6360 (N_6360,N_5771,N_5924);
and U6361 (N_6361,N_4238,N_4715);
nand U6362 (N_6362,N_3388,N_4658);
or U6363 (N_6363,N_3539,N_5971);
nor U6364 (N_6364,N_3687,N_5894);
nand U6365 (N_6365,N_4896,N_4893);
nand U6366 (N_6366,N_5843,N_5161);
nor U6367 (N_6367,N_4817,N_5521);
xor U6368 (N_6368,N_5657,N_5573);
nor U6369 (N_6369,N_5972,N_4416);
nand U6370 (N_6370,N_4039,N_3355);
or U6371 (N_6371,N_4758,N_4075);
or U6372 (N_6372,N_4103,N_3389);
nand U6373 (N_6373,N_3551,N_4326);
and U6374 (N_6374,N_5097,N_4347);
or U6375 (N_6375,N_4915,N_5022);
nor U6376 (N_6376,N_5394,N_3830);
xnor U6377 (N_6377,N_4340,N_3251);
or U6378 (N_6378,N_4931,N_5365);
nand U6379 (N_6379,N_4810,N_3515);
or U6380 (N_6380,N_5652,N_4695);
xnor U6381 (N_6381,N_3712,N_4005);
nor U6382 (N_6382,N_5166,N_4253);
nor U6383 (N_6383,N_5602,N_4773);
nor U6384 (N_6384,N_5510,N_4802);
and U6385 (N_6385,N_5044,N_5720);
and U6386 (N_6386,N_4363,N_5180);
or U6387 (N_6387,N_3672,N_4293);
nand U6388 (N_6388,N_3906,N_4160);
nand U6389 (N_6389,N_5363,N_4022);
or U6390 (N_6390,N_3379,N_5849);
nor U6391 (N_6391,N_3329,N_3948);
nand U6392 (N_6392,N_4665,N_5717);
or U6393 (N_6393,N_4691,N_3291);
nor U6394 (N_6394,N_4641,N_3686);
and U6395 (N_6395,N_5962,N_3250);
nor U6396 (N_6396,N_5981,N_4325);
xnor U6397 (N_6397,N_5714,N_5800);
and U6398 (N_6398,N_5558,N_5834);
nor U6399 (N_6399,N_4723,N_3537);
or U6400 (N_6400,N_3435,N_3309);
nand U6401 (N_6401,N_3847,N_5682);
nand U6402 (N_6402,N_4754,N_3477);
nor U6403 (N_6403,N_4179,N_4853);
nor U6404 (N_6404,N_4486,N_3110);
or U6405 (N_6405,N_5531,N_3513);
xnor U6406 (N_6406,N_3828,N_3532);
and U6407 (N_6407,N_4971,N_3151);
and U6408 (N_6408,N_5187,N_5462);
xor U6409 (N_6409,N_4165,N_4835);
nand U6410 (N_6410,N_5783,N_5569);
nor U6411 (N_6411,N_3476,N_3741);
nor U6412 (N_6412,N_3300,N_5961);
and U6413 (N_6413,N_5397,N_5799);
and U6414 (N_6414,N_5208,N_4818);
or U6415 (N_6415,N_4092,N_3272);
nor U6416 (N_6416,N_3015,N_5000);
xnor U6417 (N_6417,N_3620,N_3134);
or U6418 (N_6418,N_5270,N_4555);
or U6419 (N_6419,N_5927,N_4371);
nor U6420 (N_6420,N_4456,N_5446);
xnor U6421 (N_6421,N_4613,N_5460);
and U6422 (N_6422,N_5082,N_3359);
nand U6423 (N_6423,N_3470,N_4137);
nor U6424 (N_6424,N_3509,N_3567);
and U6425 (N_6425,N_4072,N_4192);
or U6426 (N_6426,N_3915,N_5222);
and U6427 (N_6427,N_4699,N_5434);
or U6428 (N_6428,N_5201,N_4826);
or U6429 (N_6429,N_5279,N_5389);
xnor U6430 (N_6430,N_3193,N_3058);
nor U6431 (N_6431,N_4382,N_4122);
and U6432 (N_6432,N_3204,N_4571);
and U6433 (N_6433,N_3127,N_3129);
xor U6434 (N_6434,N_5588,N_3310);
or U6435 (N_6435,N_5820,N_4534);
and U6436 (N_6436,N_5196,N_3117);
nor U6437 (N_6437,N_3481,N_4551);
nand U6438 (N_6438,N_4012,N_4727);
and U6439 (N_6439,N_3787,N_4153);
xor U6440 (N_6440,N_4819,N_3317);
or U6441 (N_6441,N_4531,N_3542);
or U6442 (N_6442,N_3855,N_4321);
nor U6443 (N_6443,N_5125,N_4987);
xor U6444 (N_6444,N_5729,N_4303);
or U6445 (N_6445,N_5190,N_5447);
or U6446 (N_6446,N_3339,N_3128);
or U6447 (N_6447,N_4435,N_3657);
or U6448 (N_6448,N_5316,N_5087);
nor U6449 (N_6449,N_5704,N_5676);
or U6450 (N_6450,N_5311,N_3485);
or U6451 (N_6451,N_4139,N_4522);
nor U6452 (N_6452,N_5548,N_3531);
and U6453 (N_6453,N_5700,N_4846);
or U6454 (N_6454,N_4724,N_4051);
nand U6455 (N_6455,N_4951,N_5741);
and U6456 (N_6456,N_3897,N_3766);
nor U6457 (N_6457,N_4351,N_4102);
or U6458 (N_6458,N_5959,N_3821);
nor U6459 (N_6459,N_4093,N_4281);
and U6460 (N_6460,N_4777,N_5057);
or U6461 (N_6461,N_4211,N_3955);
or U6462 (N_6462,N_3402,N_4757);
and U6463 (N_6463,N_4297,N_4954);
and U6464 (N_6464,N_5751,N_3031);
or U6465 (N_6465,N_3631,N_5326);
nor U6466 (N_6466,N_5254,N_5659);
and U6467 (N_6467,N_3652,N_5848);
and U6468 (N_6468,N_4843,N_5025);
and U6469 (N_6469,N_4229,N_5911);
nor U6470 (N_6470,N_5231,N_3342);
nand U6471 (N_6471,N_5232,N_4287);
and U6472 (N_6472,N_3149,N_4490);
or U6473 (N_6473,N_3440,N_4357);
nand U6474 (N_6474,N_4766,N_5283);
and U6475 (N_6475,N_4654,N_5274);
nand U6476 (N_6476,N_4797,N_4483);
and U6477 (N_6477,N_5992,N_4737);
nand U6478 (N_6478,N_4823,N_3557);
or U6479 (N_6479,N_3116,N_3789);
nand U6480 (N_6480,N_4152,N_3085);
and U6481 (N_6481,N_3069,N_5835);
xnor U6482 (N_6482,N_4631,N_5484);
or U6483 (N_6483,N_5513,N_4824);
and U6484 (N_6484,N_3749,N_4245);
or U6485 (N_6485,N_5090,N_5653);
and U6486 (N_6486,N_4260,N_4045);
xnor U6487 (N_6487,N_3056,N_4230);
or U6488 (N_6488,N_5726,N_5441);
nand U6489 (N_6489,N_5914,N_4920);
and U6490 (N_6490,N_3912,N_3432);
nand U6491 (N_6491,N_3905,N_3021);
nand U6492 (N_6492,N_5437,N_4144);
nand U6493 (N_6493,N_5384,N_5709);
nand U6494 (N_6494,N_5591,N_3624);
nor U6495 (N_6495,N_4910,N_4289);
and U6496 (N_6496,N_5974,N_3009);
or U6497 (N_6497,N_4662,N_4717);
or U6498 (N_6498,N_3424,N_5303);
nor U6499 (N_6499,N_4448,N_5468);
or U6500 (N_6500,N_4943,N_5310);
nor U6501 (N_6501,N_5689,N_4735);
nand U6502 (N_6502,N_4675,N_5789);
or U6503 (N_6503,N_4033,N_3036);
nand U6504 (N_6504,N_5155,N_4401);
or U6505 (N_6505,N_5633,N_5167);
nand U6506 (N_6506,N_5400,N_5170);
nand U6507 (N_6507,N_4610,N_5004);
nor U6508 (N_6508,N_5262,N_3100);
nor U6509 (N_6509,N_5611,N_4202);
and U6510 (N_6510,N_3418,N_4134);
or U6511 (N_6511,N_4296,N_5444);
and U6512 (N_6512,N_5597,N_4247);
or U6513 (N_6513,N_4183,N_4342);
nand U6514 (N_6514,N_3834,N_5546);
and U6515 (N_6515,N_3463,N_5457);
nor U6516 (N_6516,N_5219,N_5353);
nor U6517 (N_6517,N_4927,N_3964);
nand U6518 (N_6518,N_5151,N_5568);
and U6519 (N_6519,N_3688,N_3483);
or U6520 (N_6520,N_5983,N_5292);
and U6521 (N_6521,N_5620,N_3382);
and U6522 (N_6522,N_3810,N_4851);
or U6523 (N_6523,N_5191,N_5046);
or U6524 (N_6524,N_5803,N_3684);
and U6525 (N_6525,N_3892,N_5315);
or U6526 (N_6526,N_4604,N_4554);
and U6527 (N_6527,N_4256,N_5804);
or U6528 (N_6528,N_4863,N_4929);
or U6529 (N_6529,N_4362,N_5233);
nand U6530 (N_6530,N_4632,N_3989);
nand U6531 (N_6531,N_4057,N_5463);
xnor U6532 (N_6532,N_5586,N_3516);
nand U6533 (N_6533,N_5248,N_4860);
and U6534 (N_6534,N_3682,N_3761);
nand U6535 (N_6535,N_3825,N_5982);
xnor U6536 (N_6536,N_4680,N_4606);
nand U6537 (N_6537,N_4827,N_5318);
nand U6538 (N_6538,N_4508,N_5419);
nor U6539 (N_6539,N_4871,N_5524);
nand U6540 (N_6540,N_4009,N_3799);
nor U6541 (N_6541,N_3587,N_5332);
or U6542 (N_6542,N_3486,N_3105);
nand U6543 (N_6543,N_3563,N_3848);
and U6544 (N_6544,N_3899,N_4615);
nor U6545 (N_6545,N_3632,N_4266);
and U6546 (N_6546,N_3158,N_3809);
or U6547 (N_6547,N_5670,N_4966);
nor U6548 (N_6548,N_3203,N_3883);
and U6549 (N_6549,N_5866,N_5637);
nor U6550 (N_6550,N_3367,N_5019);
nor U6551 (N_6551,N_4474,N_3222);
nor U6552 (N_6552,N_3163,N_4290);
or U6553 (N_6553,N_5237,N_4611);
nand U6554 (N_6554,N_4783,N_5461);
and U6555 (N_6555,N_4109,N_5488);
or U6556 (N_6556,N_4782,N_4495);
and U6557 (N_6557,N_4400,N_3822);
or U6558 (N_6558,N_5066,N_5402);
nand U6559 (N_6559,N_3162,N_5740);
nand U6560 (N_6560,N_3697,N_3579);
xnor U6561 (N_6561,N_3059,N_5325);
or U6562 (N_6562,N_4327,N_3653);
nand U6563 (N_6563,N_3658,N_3337);
and U6564 (N_6564,N_5119,N_3086);
or U6565 (N_6565,N_5268,N_5241);
or U6566 (N_6566,N_3421,N_3792);
or U6567 (N_6567,N_5900,N_5723);
or U6568 (N_6568,N_3942,N_5742);
xor U6569 (N_6569,N_5282,N_3180);
and U6570 (N_6570,N_3943,N_4617);
nand U6571 (N_6571,N_3394,N_3547);
nor U6572 (N_6572,N_5052,N_3743);
and U6573 (N_6573,N_4696,N_4729);
and U6574 (N_6574,N_5563,N_4892);
nor U6575 (N_6575,N_3378,N_5145);
nor U6576 (N_6576,N_4900,N_5035);
nor U6577 (N_6577,N_5435,N_4791);
xor U6578 (N_6578,N_3360,N_4086);
nor U6579 (N_6579,N_3548,N_5535);
and U6580 (N_6580,N_5141,N_4580);
or U6581 (N_6581,N_3558,N_5926);
and U6582 (N_6582,N_4013,N_3719);
nand U6583 (N_6583,N_3517,N_3233);
or U6584 (N_6584,N_5825,N_3735);
and U6585 (N_6585,N_4341,N_3001);
nor U6586 (N_6586,N_3405,N_3640);
or U6587 (N_6587,N_5580,N_4690);
and U6588 (N_6588,N_5288,N_5658);
nor U6589 (N_6589,N_4517,N_3153);
nand U6590 (N_6590,N_4989,N_3824);
nand U6591 (N_6591,N_3475,N_4932);
nand U6592 (N_6592,N_5065,N_5404);
and U6593 (N_6593,N_4649,N_5532);
nand U6594 (N_6594,N_3185,N_3800);
or U6595 (N_6595,N_4628,N_3583);
nand U6596 (N_6596,N_3464,N_4068);
nor U6597 (N_6597,N_5150,N_5648);
nor U6598 (N_6598,N_4605,N_3333);
nor U6599 (N_6599,N_4793,N_3520);
and U6600 (N_6600,N_5192,N_5271);
xnor U6601 (N_6601,N_3377,N_3479);
xor U6602 (N_6602,N_5485,N_4032);
and U6603 (N_6603,N_4106,N_4529);
or U6604 (N_6604,N_5467,N_4061);
or U6605 (N_6605,N_3448,N_4112);
nor U6606 (N_6606,N_3011,N_5818);
nor U6607 (N_6607,N_3618,N_4099);
xnor U6608 (N_6608,N_4221,N_5852);
or U6609 (N_6609,N_5544,N_5453);
nor U6610 (N_6610,N_3623,N_3269);
or U6611 (N_6611,N_5218,N_3564);
and U6612 (N_6612,N_3444,N_4469);
nor U6613 (N_6613,N_4493,N_5074);
nand U6614 (N_6614,N_3192,N_4097);
xor U6615 (N_6615,N_4798,N_3282);
nand U6616 (N_6616,N_3480,N_3215);
or U6617 (N_6617,N_3524,N_5931);
and U6618 (N_6618,N_5865,N_5884);
nor U6619 (N_6619,N_4157,N_5142);
or U6620 (N_6620,N_3438,N_4433);
or U6621 (N_6621,N_4258,N_3109);
and U6622 (N_6622,N_4821,N_5543);
nor U6623 (N_6623,N_4755,N_5511);
nand U6624 (N_6624,N_5409,N_4402);
and U6625 (N_6625,N_3092,N_3982);
or U6626 (N_6626,N_5572,N_5654);
and U6627 (N_6627,N_3689,N_3131);
and U6628 (N_6628,N_4702,N_3608);
nand U6629 (N_6629,N_4431,N_4576);
nor U6630 (N_6630,N_3610,N_3088);
xnor U6631 (N_6631,N_5307,N_5380);
nand U6632 (N_6632,N_5160,N_5483);
nor U6633 (N_6633,N_3348,N_4923);
xor U6634 (N_6634,N_5281,N_4761);
and U6635 (N_6635,N_5263,N_4277);
or U6636 (N_6636,N_4038,N_4704);
nor U6637 (N_6637,N_5910,N_3186);
nand U6638 (N_6638,N_3325,N_4278);
and U6639 (N_6639,N_3450,N_4140);
and U6640 (N_6640,N_5236,N_5559);
or U6641 (N_6641,N_5250,N_5412);
nor U6642 (N_6642,N_4679,N_3708);
and U6643 (N_6643,N_3574,N_5582);
nand U6644 (N_6644,N_4510,N_3505);
and U6645 (N_6645,N_4193,N_5526);
nor U6646 (N_6646,N_4659,N_4182);
nand U6647 (N_6647,N_5423,N_3296);
or U6648 (N_6648,N_4588,N_3043);
and U6649 (N_6649,N_3944,N_5043);
nand U6650 (N_6650,N_3169,N_5431);
nor U6651 (N_6651,N_5829,N_4706);
and U6652 (N_6652,N_4213,N_5130);
nor U6653 (N_6653,N_3752,N_3226);
nand U6654 (N_6654,N_3680,N_5486);
and U6655 (N_6655,N_3304,N_4518);
or U6656 (N_6656,N_5173,N_4544);
nand U6657 (N_6657,N_3872,N_4765);
nor U6658 (N_6658,N_5845,N_4505);
nand U6659 (N_6659,N_4066,N_3813);
or U6660 (N_6660,N_5990,N_3952);
nand U6661 (N_6661,N_5098,N_4541);
or U6662 (N_6662,N_5107,N_4637);
and U6663 (N_6663,N_3492,N_3864);
xor U6664 (N_6664,N_5712,N_5944);
and U6665 (N_6665,N_4060,N_3616);
or U6666 (N_6666,N_3487,N_5679);
or U6667 (N_6667,N_3178,N_3772);
and U6668 (N_6668,N_4189,N_3605);
nand U6669 (N_6669,N_3570,N_4830);
nand U6670 (N_6670,N_3970,N_3400);
nor U6671 (N_6671,N_4338,N_3141);
nand U6672 (N_6672,N_3968,N_3504);
or U6673 (N_6673,N_3062,N_4028);
or U6674 (N_6674,N_3376,N_4198);
and U6675 (N_6675,N_3853,N_4636);
nor U6676 (N_6676,N_3586,N_4887);
or U6677 (N_6677,N_4855,N_3173);
or U6678 (N_6678,N_3471,N_4453);
nand U6679 (N_6679,N_4286,N_5765);
nand U6680 (N_6680,N_4734,N_4246);
nand U6681 (N_6681,N_3427,N_4836);
nor U6682 (N_6682,N_4648,N_4614);
nand U6683 (N_6683,N_4890,N_5592);
nor U6684 (N_6684,N_4603,N_3133);
and U6685 (N_6685,N_5430,N_5475);
and U6686 (N_6686,N_4799,N_4563);
nor U6687 (N_6687,N_4720,N_5985);
nand U6688 (N_6688,N_3198,N_3846);
nand U6689 (N_6689,N_4062,N_5696);
or U6690 (N_6690,N_4219,N_4002);
and U6691 (N_6691,N_3130,N_4850);
and U6692 (N_6692,N_4661,N_5211);
or U6693 (N_6693,N_4383,N_5888);
and U6694 (N_6694,N_4760,N_4774);
nor U6695 (N_6695,N_3411,N_3832);
nor U6696 (N_6696,N_5683,N_3529);
or U6697 (N_6697,N_5784,N_3525);
nor U6698 (N_6698,N_5904,N_4807);
and U6699 (N_6699,N_5069,N_3441);
and U6700 (N_6700,N_5080,N_5456);
or U6701 (N_6701,N_5688,N_5169);
nand U6702 (N_6702,N_3683,N_3677);
or U6703 (N_6703,N_5957,N_4323);
nor U6704 (N_6704,N_5377,N_5887);
xnor U6705 (N_6705,N_5425,N_5917);
nor U6706 (N_6706,N_4085,N_3575);
and U6707 (N_6707,N_5493,N_5702);
and U6708 (N_6708,N_4461,N_5429);
nand U6709 (N_6709,N_4778,N_4822);
and U6710 (N_6710,N_4582,N_5674);
nand U6711 (N_6711,N_3012,N_5667);
or U6712 (N_6712,N_5666,N_5003);
nor U6713 (N_6713,N_5707,N_5793);
nand U6714 (N_6714,N_4366,N_3962);
nor U6715 (N_6715,N_3194,N_4149);
and U6716 (N_6716,N_4537,N_4108);
or U6717 (N_6717,N_3231,N_5819);
xnor U6718 (N_6718,N_5356,N_3330);
or U6719 (N_6719,N_3806,N_3984);
nor U6720 (N_6720,N_5120,N_3746);
nor U6721 (N_6721,N_3553,N_4772);
nand U6722 (N_6722,N_5560,N_3446);
nor U6723 (N_6723,N_5623,N_3268);
and U6724 (N_6724,N_4034,N_5109);
nand U6725 (N_6725,N_4904,N_3327);
or U6726 (N_6726,N_5773,N_4594);
or U6727 (N_6727,N_4825,N_4788);
nand U6728 (N_6728,N_4767,N_3886);
or U6729 (N_6729,N_3498,N_4444);
and U6730 (N_6730,N_5645,N_3195);
nand U6731 (N_6731,N_5020,N_5615);
and U6732 (N_6732,N_4935,N_3818);
and U6733 (N_6733,N_3050,N_4898);
or U6734 (N_6734,N_4079,N_4520);
and U6735 (N_6735,N_5603,N_3362);
nand U6736 (N_6736,N_4725,N_3328);
or U6737 (N_6737,N_5379,N_3919);
nand U6738 (N_6738,N_3243,N_4635);
nor U6739 (N_6739,N_3756,N_4174);
nand U6740 (N_6740,N_5770,N_5901);
nand U6741 (N_6741,N_5031,N_3633);
xor U6742 (N_6742,N_5680,N_5965);
and U6743 (N_6743,N_3559,N_5399);
nand U6744 (N_6744,N_3628,N_5008);
nor U6745 (N_6745,N_5206,N_3745);
nor U6746 (N_6746,N_5345,N_5925);
xor U6747 (N_6747,N_3456,N_4167);
nor U6748 (N_6748,N_5011,N_4370);
or U6749 (N_6749,N_5339,N_5371);
nand U6750 (N_6750,N_3278,N_4947);
and U6751 (N_6751,N_5340,N_5854);
and U6752 (N_6752,N_3994,N_3453);
xor U6753 (N_6753,N_3494,N_5047);
nand U6754 (N_6754,N_5989,N_5398);
and U6755 (N_6755,N_5979,N_4452);
nand U6756 (N_6756,N_5768,N_5298);
nand U6757 (N_6757,N_3760,N_5733);
or U6758 (N_6758,N_4859,N_4991);
nand U6759 (N_6759,N_5721,N_5747);
xor U6760 (N_6760,N_3426,N_4977);
and U6761 (N_6761,N_3045,N_4203);
and U6762 (N_6762,N_3434,N_5722);
or U6763 (N_6763,N_5391,N_5855);
or U6764 (N_6764,N_5149,N_5197);
nand U6765 (N_6765,N_4019,N_4917);
nor U6766 (N_6766,N_4879,N_3794);
or U6767 (N_6767,N_3921,N_4178);
nor U6768 (N_6768,N_5411,N_3168);
or U6769 (N_6769,N_3839,N_4454);
nor U6770 (N_6770,N_4842,N_3039);
nor U6771 (N_6771,N_3721,N_4482);
and U6772 (N_6772,N_3064,N_3146);
nand U6773 (N_6773,N_3987,N_3026);
nor U6774 (N_6774,N_5330,N_3369);
and U6775 (N_6775,N_4312,N_3256);
nand U6776 (N_6776,N_5545,N_5744);
nand U6777 (N_6777,N_5692,N_5628);
nor U6778 (N_6778,N_3164,N_5550);
or U6779 (N_6779,N_5156,N_5806);
nand U6780 (N_6780,N_3988,N_4909);
or U6781 (N_6781,N_5223,N_5084);
or U6782 (N_6782,N_5503,N_5651);
and U6783 (N_6783,N_3433,N_4233);
or U6784 (N_6784,N_3107,N_5042);
nor U6785 (N_6785,N_4629,N_4117);
or U6786 (N_6786,N_3755,N_4858);
nand U6787 (N_6787,N_3728,N_3703);
nand U6788 (N_6788,N_4317,N_4705);
or U6789 (N_6789,N_4546,N_5089);
xor U6790 (N_6790,N_4485,N_5994);
and U6791 (N_6791,N_5601,N_3187);
and U6792 (N_6792,N_5351,N_3862);
nand U6793 (N_6793,N_5265,N_4738);
xor U6794 (N_6794,N_4451,N_3139);
and U6795 (N_6795,N_5309,N_3122);
nor U6796 (N_6796,N_3622,N_3417);
xor U6797 (N_6797,N_4115,N_3461);
or U6798 (N_6798,N_3584,N_5551);
and U6799 (N_6799,N_3387,N_3731);
nand U6800 (N_6800,N_3145,N_3904);
nand U6801 (N_6801,N_3859,N_3305);
or U6802 (N_6802,N_3753,N_3842);
or U6803 (N_6803,N_4311,N_3637);
and U6804 (N_6804,N_4392,N_5244);
nor U6805 (N_6805,N_3863,N_5595);
nand U6806 (N_6806,N_3336,N_5331);
nand U6807 (N_6807,N_4335,N_4919);
and U6808 (N_6808,N_5055,N_5314);
or U6809 (N_6809,N_5523,N_4280);
or U6810 (N_6810,N_3197,N_5823);
or U6811 (N_6811,N_5581,N_5063);
or U6812 (N_6812,N_3817,N_5023);
or U6813 (N_6813,N_3416,N_4581);
nor U6814 (N_6814,N_3447,N_3340);
nor U6815 (N_6815,N_3075,N_5506);
or U6816 (N_6816,N_5242,N_3966);
nor U6817 (N_6817,N_4385,N_5499);
or U6818 (N_6818,N_3769,N_4982);
nand U6819 (N_6819,N_5687,N_3971);
nand U6820 (N_6820,N_3879,N_3887);
nor U6821 (N_6821,N_5579,N_3917);
xnor U6822 (N_6822,N_5026,N_5229);
or U6823 (N_6823,N_4262,N_5387);
or U6824 (N_6824,N_3734,N_3101);
xor U6825 (N_6825,N_4921,N_4492);
nor U6826 (N_6826,N_3714,N_3875);
and U6827 (N_6827,N_4619,N_5816);
nand U6828 (N_6828,N_4464,N_3287);
or U6829 (N_6829,N_4861,N_3528);
and U6830 (N_6830,N_4130,N_3008);
or U6831 (N_6831,N_3368,N_4114);
nand U6832 (N_6832,N_4069,N_4187);
nor U6833 (N_6833,N_3420,N_5101);
and U6834 (N_6834,N_5472,N_4728);
or U6835 (N_6835,N_5238,N_4008);
or U6836 (N_6836,N_3206,N_3106);
nand U6837 (N_6837,N_4780,N_4804);
nor U6838 (N_6838,N_5081,N_3992);
nand U6839 (N_6839,N_5624,N_4350);
nand U6840 (N_6840,N_3973,N_3469);
nand U6841 (N_6841,N_3920,N_3455);
nor U6842 (N_6842,N_5049,N_4514);
xor U6843 (N_6843,N_5995,N_5833);
and U6844 (N_6844,N_3176,N_5871);
nand U6845 (N_6845,N_3429,N_3816);
and U6846 (N_6846,N_4841,N_3534);
and U6847 (N_6847,N_5162,N_4888);
nor U6848 (N_6848,N_4667,N_3072);
or U6849 (N_6849,N_5934,N_5415);
nand U6850 (N_6850,N_4970,N_5522);
and U6851 (N_6851,N_3302,N_4417);
xor U6852 (N_6852,N_5913,N_5589);
nor U6853 (N_6853,N_4334,N_3234);
nand U6854 (N_6854,N_3723,N_4721);
nand U6855 (N_6855,N_4602,N_4511);
or U6856 (N_6856,N_3293,N_4127);
and U6857 (N_6857,N_4701,N_5734);
or U6858 (N_6858,N_3437,N_5553);
nand U6859 (N_6859,N_3918,N_4911);
nor U6860 (N_6860,N_4794,N_3313);
xnor U6861 (N_6861,N_4845,N_5422);
and U6862 (N_6862,N_3319,N_4849);
nor U6863 (N_6863,N_4985,N_5690);
and U6864 (N_6864,N_3255,N_5490);
and U6865 (N_6865,N_5737,N_4976);
and U6866 (N_6866,N_3837,N_3029);
nor U6867 (N_6867,N_3473,N_4768);
nor U6868 (N_6868,N_5093,N_4355);
nand U6869 (N_6869,N_3157,N_4972);
xor U6870 (N_6870,N_3396,N_3852);
or U6871 (N_6871,N_3740,N_3082);
and U6872 (N_6872,N_3549,N_5964);
nand U6873 (N_6873,N_4623,N_3544);
nor U6874 (N_6874,N_3032,N_5300);
nand U6875 (N_6875,N_5343,N_3514);
and U6876 (N_6876,N_4697,N_5672);
or U6877 (N_6877,N_4058,N_4353);
and U6878 (N_6878,N_5890,N_5693);
or U6879 (N_6879,N_4204,N_3042);
and U6880 (N_6880,N_5045,N_3527);
nor U6881 (N_6881,N_5844,N_5016);
and U6882 (N_6882,N_5701,N_4070);
nor U6883 (N_6883,N_5414,N_4556);
nor U6884 (N_6884,N_5388,N_3049);
or U6885 (N_6885,N_4498,N_3181);
and U6886 (N_6886,N_3236,N_4208);
and U6887 (N_6887,N_5258,N_4885);
nor U6888 (N_6888,N_4308,N_5476);
nand U6889 (N_6889,N_5956,N_3270);
and U6890 (N_6890,N_4056,N_4963);
nand U6891 (N_6891,N_4621,N_4462);
and U6892 (N_6892,N_4275,N_4143);
or U6893 (N_6893,N_4205,N_4372);
or U6894 (N_6894,N_3869,N_3949);
xnor U6895 (N_6895,N_3990,N_5368);
nand U6896 (N_6896,N_5264,N_5537);
or U6897 (N_6897,N_3322,N_4091);
and U6898 (N_6898,N_4569,N_5245);
and U6899 (N_6899,N_4320,N_4304);
nor U6900 (N_6900,N_4064,N_3393);
nor U6901 (N_6901,N_5698,N_3025);
and U6902 (N_6902,N_3202,N_3617);
nor U6903 (N_6903,N_5966,N_3010);
nor U6904 (N_6904,N_4847,N_3284);
nand U6905 (N_6905,N_5780,N_3221);
nor U6906 (N_6906,N_5663,N_4227);
or U6907 (N_6907,N_5017,N_4561);
or U6908 (N_6908,N_3985,N_3220);
and U6909 (N_6909,N_3778,N_4076);
nor U6910 (N_6910,N_3894,N_5465);
nand U6911 (N_6911,N_5277,N_3654);
or U6912 (N_6912,N_3142,N_4948);
and U6913 (N_6913,N_3277,N_4549);
or U6914 (N_6914,N_5975,N_5750);
nand U6915 (N_6915,N_5735,N_3144);
nor U6916 (N_6916,N_4131,N_4957);
or U6917 (N_6917,N_3784,N_5366);
and U6918 (N_6918,N_4545,N_4397);
or U6919 (N_6919,N_3366,N_5039);
and U6920 (N_6920,N_3318,N_5209);
nand U6921 (N_6921,N_4184,N_5121);
or U6922 (N_6922,N_4922,N_3878);
xor U6923 (N_6923,N_3681,N_3223);
nor U6924 (N_6924,N_4181,N_3783);
xor U6925 (N_6925,N_5665,N_4294);
and U6926 (N_6926,N_4776,N_4040);
or U6927 (N_6927,N_3346,N_3913);
and U6928 (N_6928,N_5587,N_5037);
xor U6929 (N_6929,N_3780,N_3228);
xnor U6930 (N_6930,N_3639,N_3375);
or U6931 (N_6931,N_3209,N_3541);
nand U6932 (N_6932,N_5381,N_4709);
nand U6933 (N_6933,N_3053,N_3738);
nand U6934 (N_6934,N_4525,N_3750);
nand U6935 (N_6935,N_5891,N_3155);
or U6936 (N_6936,N_5635,N_3873);
and U6937 (N_6937,N_3615,N_5505);
xnor U6938 (N_6938,N_4126,N_4961);
nor U6939 (N_6939,N_3662,N_4185);
or U6940 (N_6940,N_4272,N_4234);
nor U6941 (N_6941,N_3156,N_5629);
nor U6942 (N_6942,N_5708,N_4265);
nor U6943 (N_6943,N_3338,N_3098);
nand U6944 (N_6944,N_4771,N_4744);
and U6945 (N_6945,N_5565,N_3353);
nand U6946 (N_6946,N_4415,N_4523);
nor U6947 (N_6947,N_3189,N_4925);
and U6948 (N_6948,N_4054,N_4049);
nand U6949 (N_6949,N_4194,N_5879);
or U6950 (N_6950,N_5664,N_4154);
nor U6951 (N_6951,N_5458,N_4630);
and U6952 (N_6952,N_4378,N_3002);
nor U6953 (N_6953,N_5406,N_4170);
nor U6954 (N_6954,N_3345,N_4113);
nor U6955 (N_6955,N_5135,N_5798);
xor U6956 (N_6956,N_5980,N_4162);
xor U6957 (N_6957,N_4018,N_5459);
nor U6958 (N_6958,N_4801,N_3805);
nand U6959 (N_6959,N_5739,N_3959);
and U6960 (N_6960,N_5669,N_4059);
nand U6961 (N_6961,N_4813,N_5555);
and U6962 (N_6962,N_4295,N_4196);
and U6963 (N_6963,N_4225,N_3403);
and U6964 (N_6964,N_4967,N_5630);
and U6965 (N_6965,N_4644,N_4026);
and U6966 (N_6966,N_5154,N_4548);
nand U6967 (N_6967,N_4365,N_5662);
nor U6968 (N_6968,N_3592,N_4429);
and U6969 (N_6969,N_4550,N_4239);
or U6970 (N_6970,N_5857,N_4098);
nand U6971 (N_6971,N_5091,N_4710);
nor U6972 (N_6972,N_4083,N_4673);
nand U6973 (N_6973,N_3383,N_5421);
or U6974 (N_6974,N_5252,N_4786);
and U6975 (N_6975,N_5998,N_3124);
nand U6976 (N_6976,N_5519,N_5685);
xnor U6977 (N_6977,N_3833,N_4639);
nand U6978 (N_6978,N_5986,N_3881);
or U6979 (N_6979,N_5143,N_3630);
nor U6980 (N_6980,N_4926,N_5715);
nor U6981 (N_6981,N_5703,N_3016);
and U6982 (N_6982,N_4475,N_4158);
nor U6983 (N_6983,N_4360,N_4029);
and U6984 (N_6984,N_4575,N_3843);
and U6985 (N_6985,N_4722,N_5614);
or U6986 (N_6986,N_5374,N_3172);
nor U6987 (N_6987,N_3442,N_3649);
and U6988 (N_6988,N_3093,N_3581);
nand U6989 (N_6989,N_5977,N_3625);
xor U6990 (N_6990,N_3571,N_4624);
nand U6991 (N_6991,N_5334,N_5967);
xor U6992 (N_6992,N_3726,N_3238);
nand U6993 (N_6993,N_5529,N_3409);
or U6994 (N_6994,N_4980,N_3241);
nor U6995 (N_6995,N_4499,N_3770);
and U6996 (N_6996,N_4273,N_4017);
or U6997 (N_6997,N_3263,N_3626);
nand U6998 (N_6998,N_5054,N_3573);
nor U6999 (N_6999,N_4872,N_3923);
or U7000 (N_7000,N_4912,N_3349);
nand U7001 (N_7001,N_3135,N_5794);
or U7002 (N_7002,N_5746,N_4905);
nand U7003 (N_7003,N_4135,N_3812);
nand U7004 (N_7004,N_3957,N_3237);
xor U7005 (N_7005,N_5018,N_3692);
nor U7006 (N_7006,N_3747,N_4195);
and U7007 (N_7007,N_4411,N_3961);
nor U7008 (N_7008,N_4769,N_3507);
and U7009 (N_7009,N_3003,N_3111);
or U7010 (N_7010,N_4504,N_5416);
nand U7011 (N_7011,N_3066,N_4484);
or U7012 (N_7012,N_3070,N_3670);
nor U7013 (N_7013,N_4494,N_5153);
and U7014 (N_7014,N_4132,N_4642);
nor U7015 (N_7015,N_4274,N_5058);
nand U7016 (N_7016,N_3102,N_3775);
and U7017 (N_7017,N_3737,N_3603);
and U7018 (N_7018,N_3478,N_3974);
or U7019 (N_7019,N_5754,N_5469);
and U7020 (N_7020,N_4316,N_4856);
or U7021 (N_7021,N_5514,N_4601);
or U7022 (N_7022,N_5336,N_3598);
nor U7023 (N_7023,N_5736,N_4381);
nand U7024 (N_7024,N_3802,N_5541);
nor U7025 (N_7025,N_4618,N_3909);
or U7026 (N_7026,N_4805,N_5492);
and U7027 (N_7027,N_5033,N_5140);
and U7028 (N_7028,N_3004,N_4792);
nand U7029 (N_7029,N_3977,N_4164);
xor U7030 (N_7030,N_4874,N_4838);
nand U7031 (N_7031,N_5062,N_3023);
nor U7032 (N_7032,N_3972,N_5133);
and U7033 (N_7033,N_3706,N_5297);
nor U7034 (N_7034,N_4739,N_5450);
xnor U7035 (N_7035,N_5348,N_5428);
or U7036 (N_7036,N_5766,N_5452);
or U7037 (N_7037,N_5745,N_4403);
or U7038 (N_7038,N_4913,N_3065);
nor U7039 (N_7039,N_5322,N_3037);
xor U7040 (N_7040,N_3530,N_3704);
and U7041 (N_7041,N_4021,N_4432);
and U7042 (N_7042,N_3597,N_5713);
or U7043 (N_7043,N_3889,N_3838);
nor U7044 (N_7044,N_3068,N_5349);
nand U7045 (N_7045,N_4007,N_3777);
or U7046 (N_7046,N_5813,N_4477);
or U7047 (N_7047,N_3545,N_4790);
and U7048 (N_7048,N_4488,N_4956);
nor U7049 (N_7049,N_3925,N_3292);
nand U7050 (N_7050,N_5922,N_4530);
and U7051 (N_7051,N_5184,N_5073);
nand U7052 (N_7052,N_3911,N_4354);
xor U7053 (N_7053,N_3922,N_3081);
or U7054 (N_7054,N_3815,N_4242);
nand U7055 (N_7055,N_5077,N_4313);
nor U7056 (N_7056,N_5496,N_3115);
and U7057 (N_7057,N_5790,N_5839);
or U7058 (N_7058,N_3397,N_5272);
nor U7059 (N_7059,N_5571,N_4291);
nand U7060 (N_7060,N_4396,N_5915);
nand U7061 (N_7061,N_5840,N_5179);
nor U7062 (N_7062,N_3538,N_5266);
nor U7063 (N_7063,N_3390,N_5188);
nand U7064 (N_7064,N_5360,N_5189);
and U7065 (N_7065,N_3246,N_4282);
nand U7066 (N_7066,N_3644,N_4387);
xor U7067 (N_7067,N_3289,N_5605);
and U7068 (N_7068,N_4443,N_5846);
nor U7069 (N_7069,N_3867,N_4046);
and U7070 (N_7070,N_4175,N_4955);
or U7071 (N_7071,N_4386,N_5104);
or U7072 (N_7072,N_3850,N_3646);
xor U7073 (N_7073,N_5883,N_3358);
xor U7074 (N_7074,N_5369,N_4869);
or U7075 (N_7075,N_3604,N_3474);
xor U7076 (N_7076,N_3512,N_3614);
or U7077 (N_7077,N_3190,N_4787);
and U7078 (N_7078,N_5040,N_3462);
nand U7079 (N_7079,N_5006,N_3410);
and U7080 (N_7080,N_5164,N_3694);
or U7081 (N_7081,N_3591,N_4088);
or U7082 (N_7082,N_4803,N_3910);
nor U7083 (N_7083,N_5916,N_4220);
and U7084 (N_7084,N_3754,N_4377);
xnor U7085 (N_7085,N_5779,N_5359);
and U7086 (N_7086,N_4129,N_3858);
nor U7087 (N_7087,N_4811,N_4686);
and U7088 (N_7088,N_5079,N_3884);
or U7089 (N_7089,N_4352,N_3123);
nor U7090 (N_7090,N_4995,N_4934);
and U7091 (N_7091,N_4016,N_3343);
or U7092 (N_7092,N_5728,N_4329);
and U7093 (N_7093,N_4526,N_4118);
xnor U7094 (N_7094,N_3550,N_3969);
and U7095 (N_7095,N_4997,N_3566);
nor U7096 (N_7096,N_4168,N_4222);
nor U7097 (N_7097,N_4950,N_3979);
or U7098 (N_7098,N_3273,N_4719);
or U7099 (N_7099,N_4373,N_5440);
nand U7100 (N_7100,N_3252,N_3611);
nor U7101 (N_7101,N_3907,N_4682);
nand U7102 (N_7102,N_5341,N_5312);
nand U7103 (N_7103,N_5333,N_5947);
nand U7104 (N_7104,N_3063,N_4420);
and U7105 (N_7105,N_5383,N_4441);
nor U7106 (N_7106,N_5970,N_3071);
nand U7107 (N_7107,N_3311,N_5812);
xnor U7108 (N_7108,N_3589,N_5856);
nor U7109 (N_7109,N_3024,N_4237);
nor U7110 (N_7110,N_4880,N_5479);
nor U7111 (N_7111,N_5163,N_3518);
xor U7112 (N_7112,N_4684,N_4600);
or U7113 (N_7113,N_3600,N_4147);
nor U7114 (N_7114,N_5139,N_3214);
or U7115 (N_7115,N_4528,N_3076);
nand U7116 (N_7116,N_3885,N_4285);
nand U7117 (N_7117,N_4513,N_5940);
and U7118 (N_7118,N_3720,N_4585);
nand U7119 (N_7119,N_3017,N_4560);
and U7120 (N_7120,N_3436,N_3856);
nand U7121 (N_7121,N_4990,N_5897);
and U7122 (N_7122,N_4814,N_4616);
and U7123 (N_7123,N_3497,N_4837);
or U7124 (N_7124,N_4968,N_5172);
xor U7125 (N_7125,N_3595,N_4171);
nor U7126 (N_7126,N_5759,N_4718);
nor U7127 (N_7127,N_5695,N_3308);
or U7128 (N_7128,N_3981,N_4100);
xnor U7129 (N_7129,N_5171,N_4671);
nor U7130 (N_7130,N_5627,N_3073);
and U7131 (N_7131,N_5837,N_5764);
or U7132 (N_7132,N_3841,N_3019);
or U7133 (N_7133,N_4958,N_4674);
nand U7134 (N_7134,N_4228,N_5576);
nand U7135 (N_7135,N_5583,N_4035);
nor U7136 (N_7136,N_3499,N_5873);
or U7137 (N_7137,N_5347,N_4962);
and U7138 (N_7138,N_3976,N_5809);
nand U7139 (N_7139,N_5607,N_4476);
nor U7140 (N_7140,N_3555,N_3934);
or U7141 (N_7141,N_3404,N_4527);
and U7142 (N_7142,N_3167,N_5951);
nand U7143 (N_7143,N_5969,N_5520);
nand U7144 (N_7144,N_3249,N_5731);
xor U7145 (N_7145,N_4688,N_4120);
or U7146 (N_7146,N_5382,N_3052);
nand U7147 (N_7147,N_4343,N_5909);
nor U7148 (N_7148,N_5061,N_4864);
or U7149 (N_7149,N_3836,N_4000);
nand U7150 (N_7150,N_4969,N_4574);
or U7151 (N_7151,N_4694,N_4620);
nand U7152 (N_7152,N_4562,N_3165);
or U7153 (N_7153,N_4733,N_5993);
xor U7154 (N_7154,N_3467,N_3508);
nor U7155 (N_7155,N_3385,N_4756);
or U7156 (N_7156,N_5650,N_3645);
or U7157 (N_7157,N_3888,N_5470);
or U7158 (N_7158,N_4030,N_3028);
nor U7159 (N_7159,N_4284,N_4964);
or U7160 (N_7160,N_5822,N_4439);
and U7161 (N_7161,N_3668,N_3247);
nor U7162 (N_7162,N_3166,N_5785);
nand U7163 (N_7163,N_4470,N_5774);
or U7164 (N_7164,N_4978,N_3161);
or U7165 (N_7165,N_4557,N_3827);
and U7166 (N_7166,N_3408,N_5647);
nor U7167 (N_7167,N_4457,N_3080);
and U7168 (N_7168,N_5407,N_4151);
nand U7169 (N_7169,N_3005,N_4928);
or U7170 (N_7170,N_5935,N_5295);
or U7171 (N_7171,N_4315,N_4155);
nand U7172 (N_7172,N_5626,N_3613);
nand U7173 (N_7173,N_5108,N_4583);
xnor U7174 (N_7174,N_5549,N_3040);
or U7175 (N_7175,N_5671,N_3732);
or U7176 (N_7176,N_4820,N_4328);
and U7177 (N_7177,N_3422,N_4540);
xnor U7178 (N_7178,N_5918,N_5123);
xor U7179 (N_7179,N_3347,N_4815);
nor U7180 (N_7180,N_4570,N_5186);
nor U7181 (N_7181,N_4011,N_3814);
nor U7182 (N_7182,N_4533,N_5577);
nand U7183 (N_7183,N_3634,N_5228);
and U7184 (N_7184,N_4480,N_4677);
nor U7185 (N_7185,N_5606,N_3264);
or U7186 (N_7186,N_5358,N_5181);
nor U7187 (N_7187,N_5432,N_5831);
and U7188 (N_7188,N_5554,N_5881);
nor U7189 (N_7189,N_4141,N_4176);
xnor U7190 (N_7190,N_4445,N_4430);
nor U7191 (N_7191,N_3940,N_4206);
and U7192 (N_7192,N_5552,N_5100);
xor U7193 (N_7193,N_5185,N_5919);
nor U7194 (N_7194,N_4438,N_5224);
and U7195 (N_7195,N_3160,N_4692);
and U7196 (N_7196,N_3871,N_4547);
nand U7197 (N_7197,N_4670,N_5976);
nor U7198 (N_7198,N_4374,N_3739);
and U7199 (N_7199,N_4877,N_3796);
or U7200 (N_7200,N_3954,N_4136);
nor U7201 (N_7201,N_4324,N_5294);
or U7202 (N_7202,N_5221,N_5686);
xor U7203 (N_7203,N_3078,N_5625);
or U7204 (N_7204,N_5392,N_3147);
or U7205 (N_7205,N_5561,N_3213);
nor U7206 (N_7206,N_3594,N_3767);
xor U7207 (N_7207,N_4882,N_5527);
nor U7208 (N_7208,N_5878,N_3286);
nor U7209 (N_7209,N_4595,N_4875);
nor U7210 (N_7210,N_5899,N_4375);
nand U7211 (N_7211,N_5078,N_3609);
and U7212 (N_7212,N_3901,N_5730);
nand U7213 (N_7213,N_4190,N_5442);
nor U7214 (N_7214,N_4391,N_3983);
xor U7215 (N_7215,N_4455,N_4124);
and U7216 (N_7216,N_4405,N_5525);
nand U7217 (N_7217,N_3199,N_5808);
or U7218 (N_7218,N_4936,N_4471);
or U7219 (N_7219,N_4512,N_3201);
nand U7220 (N_7220,N_4254,N_5032);
xor U7221 (N_7221,N_4053,N_4440);
nand U7222 (N_7222,N_3676,N_3791);
nor U7223 (N_7223,N_5337,N_4384);
nor U7224 (N_7224,N_3601,N_5350);
nand U7225 (N_7225,N_5811,N_3560);
xnor U7226 (N_7226,N_4223,N_4173);
nand U7227 (N_7227,N_4309,N_3320);
nor U7228 (N_7228,N_5418,N_5102);
xor U7229 (N_7229,N_4703,N_5466);
xor U7230 (N_7230,N_5867,N_4655);
xor U7231 (N_7231,N_4965,N_5933);
xor U7232 (N_7232,N_5997,N_4497);
xor U7233 (N_7233,N_3924,N_4752);
and U7234 (N_7234,N_4883,N_3938);
or U7235 (N_7235,N_5112,N_5323);
nand U7236 (N_7236,N_4437,N_5870);
or U7237 (N_7237,N_3094,N_5010);
and U7238 (N_7238,N_3790,N_3297);
nand U7239 (N_7239,N_5719,N_4252);
and U7240 (N_7240,N_5115,N_3276);
and U7241 (N_7241,N_3757,N_5202);
nand U7242 (N_7242,N_4584,N_4048);
nand U7243 (N_7243,N_3356,N_4539);
nand U7244 (N_7244,N_5464,N_4664);
and U7245 (N_7245,N_5038,N_3629);
nor U7246 (N_7246,N_4713,N_4074);
nand U7247 (N_7247,N_3638,N_4491);
nand U7248 (N_7248,N_3006,N_5786);
nor U7249 (N_7249,N_5370,N_4693);
and U7250 (N_7250,N_4095,N_3083);
xnor U7251 (N_7251,N_5941,N_4404);
and U7252 (N_7252,N_5439,N_4084);
or U7253 (N_7253,N_5622,N_3612);
nand U7254 (N_7254,N_5898,N_3495);
or U7255 (N_7255,N_5005,N_5217);
nor U7256 (N_7256,N_4394,N_5973);
and U7257 (N_7257,N_4975,N_5489);
xnor U7258 (N_7258,N_4698,N_3191);
and U7259 (N_7259,N_3642,N_5304);
or U7260 (N_7260,N_5128,N_4876);
or U7261 (N_7261,N_3801,N_4731);
or U7262 (N_7262,N_3132,N_4906);
nor U7263 (N_7263,N_3936,N_4886);
and U7264 (N_7264,N_4388,N_5261);
nor U7265 (N_7265,N_3208,N_5880);
or U7266 (N_7266,N_3665,N_5642);
nand U7267 (N_7267,N_3493,N_3643);
nor U7268 (N_7268,N_3125,N_3035);
xnor U7269 (N_7269,N_3460,N_4047);
and U7270 (N_7270,N_4410,N_4255);
nor U7271 (N_7271,N_4361,N_5306);
nand U7272 (N_7272,N_4369,N_5968);
nand U7273 (N_7273,N_5534,N_5320);
and U7274 (N_7274,N_5530,N_4063);
or U7275 (N_7275,N_4558,N_3443);
and U7276 (N_7276,N_4789,N_3046);
and U7277 (N_7277,N_3999,N_3666);
nor U7278 (N_7278,N_4643,N_3713);
xnor U7279 (N_7279,N_4096,N_5284);
and U7280 (N_7280,N_3374,N_5590);
nor U7281 (N_7281,N_4197,N_3939);
xor U7282 (N_7282,N_4646,N_3724);
nor U7283 (N_7283,N_5361,N_3736);
and U7284 (N_7284,N_5013,N_5168);
nand U7285 (N_7285,N_5317,N_5285);
or U7286 (N_7286,N_4496,N_3929);
and U7287 (N_7287,N_5007,N_4895);
and U7288 (N_7288,N_3428,N_5594);
and U7289 (N_7289,N_5036,N_5782);
nand U7290 (N_7290,N_5355,N_3253);
or U7291 (N_7291,N_4656,N_5875);
nand U7292 (N_7292,N_5451,N_5175);
nand U7293 (N_7293,N_3935,N_3673);
or U7294 (N_7294,N_4214,N_3391);
or U7295 (N_7295,N_3274,N_4434);
or U7296 (N_7296,N_4271,N_3621);
nand U7297 (N_7297,N_4231,N_5083);
and U7298 (N_7298,N_4941,N_5420);
nand U7299 (N_7299,N_4831,N_4519);
nand U7300 (N_7300,N_3386,N_3205);
nor U7301 (N_7301,N_4959,N_4077);
or U7302 (N_7302,N_3607,N_5396);
and U7303 (N_7303,N_5296,N_5923);
or U7304 (N_7304,N_3807,N_3776);
or U7305 (N_7305,N_3914,N_5540);
nand U7306 (N_7306,N_3159,N_3372);
nor U7307 (N_7307,N_3301,N_4660);
nand U7308 (N_7308,N_3307,N_5280);
and U7309 (N_7309,N_5131,N_5009);
or U7310 (N_7310,N_5619,N_5907);
and U7311 (N_7311,N_4407,N_3298);
and U7312 (N_7312,N_4399,N_4640);
nand U7313 (N_7313,N_5299,N_5251);
nor U7314 (N_7314,N_3218,N_5772);
nor U7315 (N_7315,N_4241,N_3027);
or U7316 (N_7316,N_3239,N_3916);
nand U7317 (N_7317,N_5999,N_5110);
or U7318 (N_7318,N_4226,N_5954);
and U7319 (N_7319,N_4800,N_5257);
or U7320 (N_7320,N_3998,N_4996);
nor U7321 (N_7321,N_5609,N_5826);
or U7322 (N_7322,N_5725,N_3967);
or U7323 (N_7323,N_4428,N_5050);
or U7324 (N_7324,N_5329,N_3395);
nand U7325 (N_7325,N_4180,N_4543);
xnor U7326 (N_7326,N_5474,N_3392);
and U7327 (N_7327,N_5071,N_5177);
and U7328 (N_7328,N_3488,N_5289);
or U7329 (N_7329,N_5243,N_4759);
nor U7330 (N_7330,N_3902,N_3928);
nand U7331 (N_7331,N_5885,N_3380);
nand U7332 (N_7332,N_5937,N_4307);
and U7333 (N_7333,N_4572,N_3137);
and U7334 (N_7334,N_5500,N_3326);
xnor U7335 (N_7335,N_3294,N_4395);
and U7336 (N_7336,N_5427,N_3344);
xor U7337 (N_7337,N_4299,N_3765);
or U7338 (N_7338,N_3619,N_4121);
nor U7339 (N_7339,N_5853,N_5928);
nor U7340 (N_7340,N_5824,N_4348);
nand U7341 (N_7341,N_5536,N_5176);
nand U7342 (N_7342,N_4599,N_4627);
nor U7343 (N_7343,N_5378,N_5001);
nand U7344 (N_7344,N_4653,N_4750);
nor U7345 (N_7345,N_4148,N_4010);
xnor U7346 (N_7346,N_5978,N_4306);
nor U7347 (N_7347,N_4177,N_5136);
and U7348 (N_7348,N_3635,N_3152);
nand U7349 (N_7349,N_5344,N_5193);
nand U7350 (N_7350,N_4087,N_5610);
xor U7351 (N_7351,N_3707,N_5290);
nor U7352 (N_7352,N_4500,N_4942);
and U7353 (N_7353,N_3819,N_5030);
nand U7354 (N_7354,N_3285,N_5640);
and U7355 (N_7355,N_3196,N_5127);
and U7356 (N_7356,N_4041,N_4224);
nand U7357 (N_7357,N_5070,N_3341);
and U7358 (N_7358,N_4730,N_3184);
or U7359 (N_7359,N_3188,N_4592);
nor U7360 (N_7360,N_5643,N_4037);
or U7361 (N_7361,N_5424,N_4839);
xnor U7362 (N_7362,N_3857,N_3641);
nand U7363 (N_7363,N_5528,N_5501);
nand U7364 (N_7364,N_3845,N_3332);
and U7365 (N_7365,N_4379,N_5906);
and U7366 (N_7366,N_3423,N_5117);
nand U7367 (N_7367,N_3965,N_5776);
xnor U7368 (N_7368,N_3511,N_3660);
and U7369 (N_7369,N_5792,N_3506);
or U7370 (N_7370,N_5375,N_3803);
nand U7371 (N_7371,N_4161,N_5668);
xnor U7372 (N_7372,N_3664,N_4747);
nor U7373 (N_7373,N_5029,N_3590);
or U7374 (N_7374,N_3763,N_5118);
and U7375 (N_7375,N_3782,N_5207);
nand U7376 (N_7376,N_5487,N_5376);
nor U7377 (N_7377,N_5092,N_5480);
nand U7378 (N_7378,N_3896,N_3748);
nand U7379 (N_7379,N_3774,N_4844);
or U7380 (N_7380,N_3357,N_3384);
nand U7381 (N_7381,N_4210,N_3413);
xnor U7382 (N_7382,N_4899,N_4779);
nand U7383 (N_7383,N_5547,N_4166);
nand U7384 (N_7384,N_4249,N_5618);
and U7385 (N_7385,N_4986,N_3472);
and U7386 (N_7386,N_5646,N_5002);
and U7387 (N_7387,N_3022,N_5889);
xor U7388 (N_7388,N_4795,N_4762);
and U7389 (N_7389,N_5137,N_5584);
and U7390 (N_7390,N_5938,N_3365);
nand U7391 (N_7391,N_3882,N_5960);
and U7392 (N_7392,N_4422,N_4257);
and U7393 (N_7393,N_4983,N_5122);
nor U7394 (N_7394,N_3490,N_3259);
and U7395 (N_7395,N_3140,N_5454);
nor U7396 (N_7396,N_5068,N_4336);
and U7397 (N_7397,N_4753,N_3572);
nor U7398 (N_7398,N_5860,N_4409);
and U7399 (N_7399,N_4536,N_3931);
and U7400 (N_7400,N_3785,N_5060);
or U7401 (N_7401,N_3445,N_5096);
nand U7402 (N_7402,N_5673,N_5656);
and U7403 (N_7403,N_4447,N_4298);
and U7404 (N_7404,N_5106,N_4668);
nor U7405 (N_7405,N_3565,N_4567);
and U7406 (N_7406,N_5372,N_5249);
or U7407 (N_7407,N_4191,N_4884);
and U7408 (N_7408,N_3669,N_4596);
or U7409 (N_7409,N_5912,N_4264);
and U7410 (N_7410,N_3768,N_4460);
or U7411 (N_7411,N_3900,N_3381);
or U7412 (N_7412,N_5076,N_3095);
or U7413 (N_7413,N_5498,N_3266);
or U7414 (N_7414,N_5632,N_3947);
xor U7415 (N_7415,N_5678,N_4683);
nor U7416 (N_7416,N_5612,N_3114);
or U7417 (N_7417,N_5301,N_4209);
xor U7418 (N_7418,N_5253,N_3730);
and U7419 (N_7419,N_4322,N_3415);
or U7420 (N_7420,N_4390,N_3306);
xnor U7421 (N_7421,N_4023,N_4981);
and U7422 (N_7422,N_3788,N_5797);
nor U7423 (N_7423,N_5756,N_3489);
nor U7424 (N_7424,N_5738,N_5963);
and U7425 (N_7425,N_3593,N_4424);
nor U7426 (N_7426,N_5287,N_5259);
nor U7427 (N_7427,N_5230,N_3265);
or U7428 (N_7428,N_5872,N_5864);
nand U7429 (N_7429,N_3661,N_5235);
and U7430 (N_7430,N_4024,N_3655);
nor U7431 (N_7431,N_3275,N_4463);
and U7432 (N_7432,N_5593,N_4458);
xnor U7433 (N_7433,N_4459,N_5769);
nand U7434 (N_7434,N_3671,N_4930);
nand U7435 (N_7435,N_3831,N_4349);
nor U7436 (N_7436,N_5598,N_3280);
and U7437 (N_7437,N_3877,N_3627);
nor U7438 (N_7438,N_4172,N_3727);
nand U7439 (N_7439,N_5753,N_5616);
nand U7440 (N_7440,N_5247,N_5596);
or U7441 (N_7441,N_5955,N_5795);
nand U7442 (N_7442,N_5801,N_4020);
or U7443 (N_7443,N_5021,N_4901);
nand U7444 (N_7444,N_3054,N_4685);
nor U7445 (N_7445,N_4442,N_3179);
nand U7446 (N_7446,N_5948,N_3705);
and U7447 (N_7447,N_5194,N_4647);
nand U7448 (N_7448,N_4732,N_4565);
nor U7449 (N_7449,N_3960,N_4666);
nand U7450 (N_7450,N_3077,N_5094);
nand U7451 (N_7451,N_4933,N_3451);
nor U7452 (N_7452,N_4426,N_4993);
or U7453 (N_7453,N_3501,N_4707);
or U7454 (N_7454,N_5755,N_3829);
nand U7455 (N_7455,N_4829,N_4712);
nor U7456 (N_7456,N_4598,N_3695);
xor U7457 (N_7457,N_5761,N_4111);
or U7458 (N_7458,N_4862,N_5158);
and U7459 (N_7459,N_5183,N_4436);
or U7460 (N_7460,N_3248,N_4865);
and U7461 (N_7461,N_4090,N_4566);
nor U7462 (N_7462,N_3798,N_4612);
and U7463 (N_7463,N_3543,N_4027);
and U7464 (N_7464,N_5841,N_4775);
xnor U7465 (N_7465,N_4597,N_4552);
or U7466 (N_7466,N_4393,N_4808);
nand U7467 (N_7467,N_4408,N_5660);
nor U7468 (N_7468,N_5048,N_3211);
nand U7469 (N_7469,N_3835,N_4832);
and U7470 (N_7470,N_5802,N_5838);
or U7471 (N_7471,N_3373,N_4979);
nand U7472 (N_7472,N_3299,N_5157);
and U7473 (N_7473,N_4380,N_4973);
nor U7474 (N_7474,N_3331,N_5515);
and U7475 (N_7475,N_3781,N_5861);
nand U7476 (N_7476,N_4984,N_4156);
nand U7477 (N_7477,N_3361,N_4345);
nor U7478 (N_7478,N_5482,N_4891);
nand U7479 (N_7479,N_4236,N_4974);
xnor U7480 (N_7480,N_4413,N_4267);
nand U7481 (N_7481,N_5958,N_4937);
and U7482 (N_7482,N_5508,N_4946);
and U7483 (N_7483,N_4319,N_4591);
nor U7484 (N_7484,N_5876,N_4652);
and U7485 (N_7485,N_4330,N_4067);
or U7486 (N_7486,N_5718,N_3000);
or U7487 (N_7487,N_4094,N_4398);
and U7488 (N_7488,N_3431,N_5644);
and U7489 (N_7489,N_5226,N_5099);
or U7490 (N_7490,N_4276,N_4128);
and U7491 (N_7491,N_5608,N_5319);
or U7492 (N_7492,N_5199,N_3795);
nor U7493 (N_7493,N_3561,N_4587);
xnor U7494 (N_7494,N_5807,N_5636);
or U7495 (N_7495,N_5810,N_5269);
or U7496 (N_7496,N_4687,N_4711);
or U7497 (N_7497,N_3047,N_5426);
nand U7498 (N_7498,N_3295,N_3865);
nor U7499 (N_7499,N_5930,N_3930);
or U7500 (N_7500,N_3693,N_3952);
nor U7501 (N_7501,N_5497,N_4142);
nand U7502 (N_7502,N_5681,N_4087);
nor U7503 (N_7503,N_4849,N_5600);
nor U7504 (N_7504,N_4499,N_3832);
nor U7505 (N_7505,N_5232,N_5009);
nand U7506 (N_7506,N_5451,N_5629);
xor U7507 (N_7507,N_4941,N_4733);
nand U7508 (N_7508,N_4030,N_3375);
and U7509 (N_7509,N_3686,N_3113);
or U7510 (N_7510,N_5680,N_5655);
xor U7511 (N_7511,N_4231,N_4193);
and U7512 (N_7512,N_3968,N_5741);
nand U7513 (N_7513,N_5030,N_5387);
or U7514 (N_7514,N_4791,N_4104);
and U7515 (N_7515,N_4401,N_5520);
nand U7516 (N_7516,N_3522,N_4827);
or U7517 (N_7517,N_5788,N_5998);
xor U7518 (N_7518,N_5261,N_3631);
or U7519 (N_7519,N_3461,N_3534);
or U7520 (N_7520,N_4008,N_3505);
and U7521 (N_7521,N_5226,N_4956);
nand U7522 (N_7522,N_5748,N_3119);
xnor U7523 (N_7523,N_3995,N_5116);
and U7524 (N_7524,N_5225,N_3001);
xnor U7525 (N_7525,N_5034,N_5231);
and U7526 (N_7526,N_5069,N_4243);
xor U7527 (N_7527,N_4384,N_4993);
and U7528 (N_7528,N_4993,N_3546);
nor U7529 (N_7529,N_4069,N_3490);
or U7530 (N_7530,N_3717,N_3741);
or U7531 (N_7531,N_3070,N_4361);
and U7532 (N_7532,N_5640,N_5072);
nand U7533 (N_7533,N_3457,N_4180);
nand U7534 (N_7534,N_4152,N_5159);
and U7535 (N_7535,N_3264,N_3129);
nor U7536 (N_7536,N_3666,N_4305);
and U7537 (N_7537,N_4645,N_5772);
nand U7538 (N_7538,N_5916,N_3362);
nor U7539 (N_7539,N_4455,N_3807);
and U7540 (N_7540,N_3319,N_5221);
nor U7541 (N_7541,N_4636,N_4200);
and U7542 (N_7542,N_4637,N_4207);
and U7543 (N_7543,N_5319,N_4868);
and U7544 (N_7544,N_5020,N_5597);
xor U7545 (N_7545,N_4700,N_4456);
or U7546 (N_7546,N_4064,N_5173);
and U7547 (N_7547,N_4893,N_4522);
or U7548 (N_7548,N_5892,N_4393);
nor U7549 (N_7549,N_3324,N_4018);
and U7550 (N_7550,N_4284,N_3769);
nand U7551 (N_7551,N_3448,N_3333);
nand U7552 (N_7552,N_5518,N_3246);
xor U7553 (N_7553,N_5560,N_5808);
nand U7554 (N_7554,N_5891,N_5740);
or U7555 (N_7555,N_5450,N_3186);
xor U7556 (N_7556,N_3424,N_4829);
nand U7557 (N_7557,N_4636,N_3551);
nand U7558 (N_7558,N_4490,N_5381);
and U7559 (N_7559,N_4086,N_5364);
and U7560 (N_7560,N_3457,N_4986);
nor U7561 (N_7561,N_5470,N_4664);
nor U7562 (N_7562,N_3089,N_3535);
nand U7563 (N_7563,N_3354,N_4360);
or U7564 (N_7564,N_5820,N_3095);
or U7565 (N_7565,N_5323,N_4560);
or U7566 (N_7566,N_4026,N_5717);
nor U7567 (N_7567,N_4366,N_3772);
nor U7568 (N_7568,N_4028,N_4258);
nor U7569 (N_7569,N_5812,N_3642);
nor U7570 (N_7570,N_5069,N_3188);
and U7571 (N_7571,N_5432,N_5794);
and U7572 (N_7572,N_3194,N_4461);
nor U7573 (N_7573,N_4406,N_5306);
nand U7574 (N_7574,N_3631,N_5537);
and U7575 (N_7575,N_5768,N_3000);
nand U7576 (N_7576,N_4479,N_5031);
nor U7577 (N_7577,N_3486,N_3805);
or U7578 (N_7578,N_3305,N_4345);
and U7579 (N_7579,N_4625,N_5425);
and U7580 (N_7580,N_4937,N_4115);
or U7581 (N_7581,N_5057,N_5957);
or U7582 (N_7582,N_4979,N_4653);
or U7583 (N_7583,N_5494,N_4551);
nor U7584 (N_7584,N_3479,N_4957);
or U7585 (N_7585,N_3348,N_3847);
nand U7586 (N_7586,N_3245,N_3014);
or U7587 (N_7587,N_4966,N_4487);
nor U7588 (N_7588,N_3797,N_5680);
or U7589 (N_7589,N_4794,N_3835);
nor U7590 (N_7590,N_4235,N_3592);
and U7591 (N_7591,N_5805,N_3344);
nor U7592 (N_7592,N_4875,N_4798);
and U7593 (N_7593,N_5406,N_4913);
and U7594 (N_7594,N_4869,N_3597);
nor U7595 (N_7595,N_5985,N_4541);
and U7596 (N_7596,N_4381,N_4480);
and U7597 (N_7597,N_4903,N_5038);
and U7598 (N_7598,N_5602,N_5068);
nand U7599 (N_7599,N_5346,N_3918);
and U7600 (N_7600,N_3117,N_3693);
or U7601 (N_7601,N_3667,N_5364);
and U7602 (N_7602,N_5126,N_5696);
nand U7603 (N_7603,N_5378,N_3711);
and U7604 (N_7604,N_3357,N_3510);
or U7605 (N_7605,N_5949,N_3700);
or U7606 (N_7606,N_4456,N_3718);
nand U7607 (N_7607,N_4400,N_3078);
nand U7608 (N_7608,N_5738,N_3503);
nor U7609 (N_7609,N_5445,N_3987);
nor U7610 (N_7610,N_4449,N_4000);
nor U7611 (N_7611,N_5383,N_5216);
nand U7612 (N_7612,N_3162,N_3568);
and U7613 (N_7613,N_3375,N_4555);
and U7614 (N_7614,N_5648,N_4239);
and U7615 (N_7615,N_3039,N_4385);
or U7616 (N_7616,N_4888,N_4927);
nor U7617 (N_7617,N_5688,N_3827);
and U7618 (N_7618,N_3465,N_4729);
nand U7619 (N_7619,N_3754,N_5852);
nor U7620 (N_7620,N_5620,N_3034);
nand U7621 (N_7621,N_3093,N_3734);
and U7622 (N_7622,N_5088,N_3447);
nand U7623 (N_7623,N_4284,N_5468);
nor U7624 (N_7624,N_5776,N_3178);
or U7625 (N_7625,N_5128,N_3618);
nor U7626 (N_7626,N_5204,N_3420);
nand U7627 (N_7627,N_4779,N_4183);
xnor U7628 (N_7628,N_4226,N_5155);
nor U7629 (N_7629,N_4550,N_3170);
or U7630 (N_7630,N_3302,N_4018);
and U7631 (N_7631,N_3960,N_4743);
and U7632 (N_7632,N_4459,N_3292);
or U7633 (N_7633,N_4305,N_5254);
nor U7634 (N_7634,N_4824,N_3777);
nor U7635 (N_7635,N_3355,N_5719);
nor U7636 (N_7636,N_5554,N_4402);
nand U7637 (N_7637,N_5562,N_5281);
xor U7638 (N_7638,N_3615,N_3097);
xnor U7639 (N_7639,N_4175,N_5183);
and U7640 (N_7640,N_5509,N_3426);
xor U7641 (N_7641,N_5328,N_4290);
or U7642 (N_7642,N_5457,N_4723);
nand U7643 (N_7643,N_3626,N_3620);
nor U7644 (N_7644,N_3821,N_5373);
xnor U7645 (N_7645,N_3497,N_5140);
nor U7646 (N_7646,N_4720,N_4322);
xor U7647 (N_7647,N_5004,N_4832);
or U7648 (N_7648,N_5344,N_4988);
or U7649 (N_7649,N_3458,N_5561);
and U7650 (N_7650,N_5541,N_4117);
nand U7651 (N_7651,N_5522,N_5299);
nand U7652 (N_7652,N_4180,N_5987);
nor U7653 (N_7653,N_5792,N_4975);
xor U7654 (N_7654,N_4718,N_4830);
or U7655 (N_7655,N_3395,N_4291);
nand U7656 (N_7656,N_5122,N_4776);
nor U7657 (N_7657,N_5987,N_5030);
nor U7658 (N_7658,N_3663,N_3805);
and U7659 (N_7659,N_5617,N_3383);
or U7660 (N_7660,N_3498,N_4522);
or U7661 (N_7661,N_4729,N_3849);
nor U7662 (N_7662,N_3064,N_5600);
and U7663 (N_7663,N_5098,N_4464);
or U7664 (N_7664,N_3303,N_4059);
nand U7665 (N_7665,N_5888,N_5702);
or U7666 (N_7666,N_3584,N_5893);
nor U7667 (N_7667,N_3086,N_5381);
nor U7668 (N_7668,N_3551,N_5057);
and U7669 (N_7669,N_5948,N_4339);
or U7670 (N_7670,N_5949,N_3698);
nand U7671 (N_7671,N_5400,N_5770);
nand U7672 (N_7672,N_4403,N_4088);
or U7673 (N_7673,N_5374,N_5731);
nand U7674 (N_7674,N_3853,N_5696);
xnor U7675 (N_7675,N_4060,N_5028);
nor U7676 (N_7676,N_5489,N_4018);
nor U7677 (N_7677,N_5271,N_4817);
and U7678 (N_7678,N_5188,N_4717);
or U7679 (N_7679,N_4026,N_5828);
or U7680 (N_7680,N_3824,N_4306);
nor U7681 (N_7681,N_5594,N_4653);
or U7682 (N_7682,N_3721,N_3528);
and U7683 (N_7683,N_4892,N_4241);
or U7684 (N_7684,N_4363,N_5237);
nand U7685 (N_7685,N_4278,N_5058);
and U7686 (N_7686,N_4130,N_5637);
and U7687 (N_7687,N_4880,N_5269);
and U7688 (N_7688,N_4329,N_3622);
nand U7689 (N_7689,N_4149,N_3835);
xnor U7690 (N_7690,N_5263,N_3040);
or U7691 (N_7691,N_3160,N_3998);
nand U7692 (N_7692,N_5128,N_5539);
and U7693 (N_7693,N_4788,N_5117);
and U7694 (N_7694,N_4243,N_5542);
and U7695 (N_7695,N_4764,N_4107);
or U7696 (N_7696,N_4002,N_5534);
and U7697 (N_7697,N_3585,N_3872);
and U7698 (N_7698,N_4490,N_4619);
or U7699 (N_7699,N_4631,N_3825);
nand U7700 (N_7700,N_3763,N_5638);
and U7701 (N_7701,N_5692,N_3131);
nand U7702 (N_7702,N_5334,N_3402);
or U7703 (N_7703,N_4732,N_3274);
nor U7704 (N_7704,N_5960,N_5846);
and U7705 (N_7705,N_3197,N_3919);
nand U7706 (N_7706,N_3492,N_4862);
or U7707 (N_7707,N_4305,N_4799);
or U7708 (N_7708,N_4900,N_5367);
or U7709 (N_7709,N_5905,N_5030);
and U7710 (N_7710,N_5992,N_3655);
or U7711 (N_7711,N_5192,N_4246);
and U7712 (N_7712,N_5563,N_5071);
nor U7713 (N_7713,N_4860,N_3205);
and U7714 (N_7714,N_5177,N_4813);
nand U7715 (N_7715,N_3250,N_3618);
nor U7716 (N_7716,N_4881,N_3588);
and U7717 (N_7717,N_5023,N_4244);
or U7718 (N_7718,N_4835,N_3009);
or U7719 (N_7719,N_3942,N_3950);
nor U7720 (N_7720,N_3043,N_3773);
or U7721 (N_7721,N_4258,N_5979);
nand U7722 (N_7722,N_5501,N_3483);
nand U7723 (N_7723,N_3549,N_5455);
nor U7724 (N_7724,N_4294,N_4095);
nand U7725 (N_7725,N_5054,N_5915);
and U7726 (N_7726,N_4070,N_4533);
or U7727 (N_7727,N_5945,N_5582);
xor U7728 (N_7728,N_5562,N_5514);
xnor U7729 (N_7729,N_4495,N_5753);
nand U7730 (N_7730,N_4564,N_3569);
or U7731 (N_7731,N_5545,N_5305);
and U7732 (N_7732,N_5567,N_3825);
and U7733 (N_7733,N_5439,N_5841);
or U7734 (N_7734,N_4355,N_4390);
or U7735 (N_7735,N_4245,N_3769);
nor U7736 (N_7736,N_3737,N_5033);
and U7737 (N_7737,N_4932,N_4822);
nor U7738 (N_7738,N_5813,N_3528);
xnor U7739 (N_7739,N_5782,N_5552);
xor U7740 (N_7740,N_3444,N_3522);
nor U7741 (N_7741,N_4742,N_5445);
nand U7742 (N_7742,N_5873,N_4511);
and U7743 (N_7743,N_5511,N_4152);
and U7744 (N_7744,N_5832,N_4963);
nor U7745 (N_7745,N_4915,N_4689);
xnor U7746 (N_7746,N_3502,N_3762);
nand U7747 (N_7747,N_3358,N_5793);
nand U7748 (N_7748,N_3327,N_4759);
and U7749 (N_7749,N_4844,N_3034);
and U7750 (N_7750,N_4922,N_4285);
nor U7751 (N_7751,N_5532,N_5917);
or U7752 (N_7752,N_4178,N_5757);
nand U7753 (N_7753,N_3780,N_5508);
and U7754 (N_7754,N_4979,N_4699);
nand U7755 (N_7755,N_3683,N_5395);
nor U7756 (N_7756,N_3335,N_4226);
nor U7757 (N_7757,N_4056,N_5188);
and U7758 (N_7758,N_5110,N_3014);
or U7759 (N_7759,N_4178,N_3443);
xor U7760 (N_7760,N_3966,N_4070);
or U7761 (N_7761,N_4993,N_3853);
nand U7762 (N_7762,N_5599,N_4574);
and U7763 (N_7763,N_4749,N_5043);
or U7764 (N_7764,N_4619,N_4626);
xor U7765 (N_7765,N_3695,N_4670);
and U7766 (N_7766,N_3061,N_3122);
and U7767 (N_7767,N_5546,N_4234);
nand U7768 (N_7768,N_3711,N_3355);
nand U7769 (N_7769,N_3112,N_4112);
nor U7770 (N_7770,N_5553,N_5717);
xor U7771 (N_7771,N_5142,N_5999);
or U7772 (N_7772,N_4215,N_3187);
nor U7773 (N_7773,N_3871,N_3881);
or U7774 (N_7774,N_5457,N_3351);
or U7775 (N_7775,N_4371,N_5533);
nor U7776 (N_7776,N_5980,N_3943);
or U7777 (N_7777,N_4597,N_5448);
and U7778 (N_7778,N_4833,N_5102);
xor U7779 (N_7779,N_4243,N_5525);
and U7780 (N_7780,N_4408,N_4349);
and U7781 (N_7781,N_5621,N_4635);
nand U7782 (N_7782,N_3717,N_4161);
or U7783 (N_7783,N_5503,N_4775);
nor U7784 (N_7784,N_4333,N_3761);
xor U7785 (N_7785,N_4435,N_3171);
nand U7786 (N_7786,N_5012,N_4033);
xnor U7787 (N_7787,N_3742,N_5265);
or U7788 (N_7788,N_4711,N_4587);
or U7789 (N_7789,N_5678,N_3654);
nor U7790 (N_7790,N_5962,N_3910);
and U7791 (N_7791,N_4701,N_5339);
nand U7792 (N_7792,N_5318,N_3712);
or U7793 (N_7793,N_3316,N_5070);
nand U7794 (N_7794,N_4347,N_4125);
nor U7795 (N_7795,N_3792,N_5484);
or U7796 (N_7796,N_3196,N_5878);
xor U7797 (N_7797,N_4909,N_5125);
nand U7798 (N_7798,N_4586,N_4851);
or U7799 (N_7799,N_3777,N_5264);
and U7800 (N_7800,N_4406,N_5994);
nand U7801 (N_7801,N_4407,N_5934);
and U7802 (N_7802,N_5755,N_4606);
nand U7803 (N_7803,N_5559,N_3745);
nand U7804 (N_7804,N_5274,N_4851);
nand U7805 (N_7805,N_4681,N_4020);
nand U7806 (N_7806,N_4588,N_5863);
or U7807 (N_7807,N_3377,N_3072);
nor U7808 (N_7808,N_4415,N_3616);
nand U7809 (N_7809,N_3548,N_4173);
xnor U7810 (N_7810,N_3091,N_4923);
or U7811 (N_7811,N_4866,N_5456);
or U7812 (N_7812,N_3342,N_5564);
nor U7813 (N_7813,N_4911,N_4239);
and U7814 (N_7814,N_4123,N_3717);
or U7815 (N_7815,N_3099,N_5663);
nand U7816 (N_7816,N_4956,N_3651);
nor U7817 (N_7817,N_3216,N_3142);
and U7818 (N_7818,N_4118,N_5987);
or U7819 (N_7819,N_3385,N_4705);
nand U7820 (N_7820,N_3148,N_5208);
or U7821 (N_7821,N_4129,N_5597);
and U7822 (N_7822,N_3636,N_3851);
and U7823 (N_7823,N_5095,N_4368);
nor U7824 (N_7824,N_4494,N_3764);
nand U7825 (N_7825,N_5799,N_3008);
nand U7826 (N_7826,N_3506,N_5192);
or U7827 (N_7827,N_4086,N_5387);
nor U7828 (N_7828,N_3520,N_3868);
or U7829 (N_7829,N_3805,N_4503);
nor U7830 (N_7830,N_5707,N_4850);
and U7831 (N_7831,N_3344,N_3285);
xor U7832 (N_7832,N_4671,N_3021);
and U7833 (N_7833,N_3885,N_4472);
xor U7834 (N_7834,N_4334,N_3425);
nand U7835 (N_7835,N_5945,N_4513);
nand U7836 (N_7836,N_5384,N_4640);
nor U7837 (N_7837,N_5662,N_5387);
nor U7838 (N_7838,N_5592,N_5176);
or U7839 (N_7839,N_4534,N_5815);
or U7840 (N_7840,N_5634,N_5666);
nand U7841 (N_7841,N_3726,N_4425);
and U7842 (N_7842,N_4491,N_5399);
nor U7843 (N_7843,N_4213,N_5579);
nor U7844 (N_7844,N_4426,N_4150);
and U7845 (N_7845,N_5996,N_3777);
nand U7846 (N_7846,N_4892,N_3076);
nor U7847 (N_7847,N_4332,N_4315);
or U7848 (N_7848,N_4244,N_4938);
or U7849 (N_7849,N_4571,N_3677);
nor U7850 (N_7850,N_4282,N_5545);
xnor U7851 (N_7851,N_3070,N_3529);
nand U7852 (N_7852,N_3501,N_4802);
nor U7853 (N_7853,N_5114,N_4192);
nor U7854 (N_7854,N_3179,N_3228);
or U7855 (N_7855,N_5421,N_5850);
xor U7856 (N_7856,N_5127,N_4886);
nand U7857 (N_7857,N_4502,N_5934);
or U7858 (N_7858,N_4723,N_5638);
nor U7859 (N_7859,N_3989,N_4772);
xor U7860 (N_7860,N_4462,N_5545);
nor U7861 (N_7861,N_4484,N_5956);
nand U7862 (N_7862,N_3635,N_4352);
or U7863 (N_7863,N_5944,N_4260);
xor U7864 (N_7864,N_5689,N_4660);
nand U7865 (N_7865,N_3845,N_4646);
and U7866 (N_7866,N_4109,N_4141);
and U7867 (N_7867,N_4826,N_3667);
xor U7868 (N_7868,N_4705,N_3071);
and U7869 (N_7869,N_4585,N_4889);
and U7870 (N_7870,N_3106,N_4160);
nand U7871 (N_7871,N_3046,N_4604);
and U7872 (N_7872,N_5752,N_5753);
xnor U7873 (N_7873,N_5165,N_3332);
nand U7874 (N_7874,N_3083,N_3766);
nor U7875 (N_7875,N_4999,N_4249);
or U7876 (N_7876,N_5892,N_3584);
nor U7877 (N_7877,N_4073,N_5498);
nand U7878 (N_7878,N_3119,N_4173);
nand U7879 (N_7879,N_3405,N_4024);
and U7880 (N_7880,N_4676,N_4846);
nor U7881 (N_7881,N_4074,N_5479);
and U7882 (N_7882,N_3643,N_3978);
nand U7883 (N_7883,N_5073,N_3586);
and U7884 (N_7884,N_3678,N_3103);
xnor U7885 (N_7885,N_5622,N_5763);
nor U7886 (N_7886,N_5234,N_4617);
nor U7887 (N_7887,N_4882,N_5468);
nor U7888 (N_7888,N_5135,N_4203);
and U7889 (N_7889,N_3007,N_5029);
nor U7890 (N_7890,N_5971,N_4269);
and U7891 (N_7891,N_3093,N_5644);
and U7892 (N_7892,N_4264,N_4754);
nor U7893 (N_7893,N_5867,N_4869);
and U7894 (N_7894,N_5654,N_4230);
and U7895 (N_7895,N_4180,N_5937);
or U7896 (N_7896,N_4456,N_5257);
and U7897 (N_7897,N_5852,N_4009);
nor U7898 (N_7898,N_4569,N_4740);
nand U7899 (N_7899,N_5218,N_5700);
nor U7900 (N_7900,N_5424,N_5873);
or U7901 (N_7901,N_4957,N_4023);
nand U7902 (N_7902,N_4831,N_3594);
nand U7903 (N_7903,N_4907,N_5185);
nor U7904 (N_7904,N_5161,N_5159);
or U7905 (N_7905,N_5465,N_4480);
nor U7906 (N_7906,N_5588,N_4034);
and U7907 (N_7907,N_4683,N_4585);
or U7908 (N_7908,N_4255,N_4790);
nor U7909 (N_7909,N_4482,N_3670);
and U7910 (N_7910,N_5717,N_4584);
or U7911 (N_7911,N_4413,N_5546);
nand U7912 (N_7912,N_4038,N_5381);
nor U7913 (N_7913,N_4811,N_3464);
nor U7914 (N_7914,N_5173,N_4239);
and U7915 (N_7915,N_5332,N_5996);
nand U7916 (N_7916,N_5078,N_5189);
or U7917 (N_7917,N_5603,N_3415);
nand U7918 (N_7918,N_3946,N_3485);
and U7919 (N_7919,N_5905,N_5507);
nor U7920 (N_7920,N_4014,N_5033);
nor U7921 (N_7921,N_3509,N_4098);
nand U7922 (N_7922,N_3746,N_4321);
xnor U7923 (N_7923,N_5737,N_3959);
or U7924 (N_7924,N_3822,N_4007);
or U7925 (N_7925,N_4517,N_5428);
nand U7926 (N_7926,N_3924,N_4654);
or U7927 (N_7927,N_4170,N_5093);
nand U7928 (N_7928,N_5684,N_3059);
nand U7929 (N_7929,N_4084,N_5330);
and U7930 (N_7930,N_5337,N_3998);
and U7931 (N_7931,N_5934,N_4882);
nand U7932 (N_7932,N_5988,N_5221);
nand U7933 (N_7933,N_3401,N_3735);
nand U7934 (N_7934,N_5138,N_5031);
nand U7935 (N_7935,N_4857,N_3851);
and U7936 (N_7936,N_5651,N_5738);
nor U7937 (N_7937,N_3555,N_3496);
nor U7938 (N_7938,N_5902,N_5633);
nand U7939 (N_7939,N_5600,N_3219);
or U7940 (N_7940,N_3764,N_5607);
or U7941 (N_7941,N_4147,N_4970);
or U7942 (N_7942,N_4114,N_4088);
or U7943 (N_7943,N_4226,N_4950);
nor U7944 (N_7944,N_3660,N_3986);
nor U7945 (N_7945,N_5525,N_5286);
or U7946 (N_7946,N_4233,N_5692);
or U7947 (N_7947,N_3132,N_5597);
xnor U7948 (N_7948,N_5574,N_5160);
nand U7949 (N_7949,N_4214,N_5482);
or U7950 (N_7950,N_3692,N_4235);
or U7951 (N_7951,N_4775,N_5515);
nand U7952 (N_7952,N_3871,N_3326);
nand U7953 (N_7953,N_4317,N_4802);
nand U7954 (N_7954,N_5889,N_3763);
or U7955 (N_7955,N_3743,N_3543);
or U7956 (N_7956,N_5571,N_4895);
nand U7957 (N_7957,N_3254,N_4556);
and U7958 (N_7958,N_3060,N_4066);
nand U7959 (N_7959,N_4795,N_3992);
nor U7960 (N_7960,N_5046,N_5875);
or U7961 (N_7961,N_4047,N_5198);
nor U7962 (N_7962,N_3768,N_4160);
nor U7963 (N_7963,N_3957,N_5967);
nor U7964 (N_7964,N_3178,N_3181);
nand U7965 (N_7965,N_5013,N_3509);
nand U7966 (N_7966,N_5765,N_5066);
and U7967 (N_7967,N_3780,N_4369);
or U7968 (N_7968,N_5426,N_4291);
or U7969 (N_7969,N_5122,N_5094);
and U7970 (N_7970,N_3653,N_5739);
and U7971 (N_7971,N_5537,N_4555);
nor U7972 (N_7972,N_5763,N_4525);
nor U7973 (N_7973,N_5286,N_3352);
and U7974 (N_7974,N_5082,N_3671);
xnor U7975 (N_7975,N_5812,N_5660);
or U7976 (N_7976,N_3088,N_3852);
nand U7977 (N_7977,N_5319,N_5111);
nand U7978 (N_7978,N_3093,N_5136);
nor U7979 (N_7979,N_5473,N_5146);
and U7980 (N_7980,N_5968,N_5839);
or U7981 (N_7981,N_5005,N_3883);
and U7982 (N_7982,N_4561,N_5044);
nor U7983 (N_7983,N_4602,N_5507);
xor U7984 (N_7984,N_3402,N_3694);
nand U7985 (N_7985,N_3194,N_4612);
or U7986 (N_7986,N_4139,N_5979);
nand U7987 (N_7987,N_5664,N_3893);
or U7988 (N_7988,N_5244,N_5986);
or U7989 (N_7989,N_4536,N_3359);
nand U7990 (N_7990,N_4582,N_3183);
or U7991 (N_7991,N_3920,N_4086);
or U7992 (N_7992,N_4137,N_5667);
nand U7993 (N_7993,N_5123,N_5211);
and U7994 (N_7994,N_3887,N_5411);
nor U7995 (N_7995,N_4947,N_4626);
or U7996 (N_7996,N_5783,N_5807);
or U7997 (N_7997,N_5048,N_3023);
nand U7998 (N_7998,N_5809,N_4820);
nand U7999 (N_7999,N_3010,N_5144);
and U8000 (N_8000,N_5144,N_4365);
xor U8001 (N_8001,N_5759,N_3887);
nand U8002 (N_8002,N_4447,N_3289);
and U8003 (N_8003,N_3489,N_5181);
nand U8004 (N_8004,N_5807,N_4538);
nand U8005 (N_8005,N_4411,N_4129);
and U8006 (N_8006,N_3620,N_5821);
nor U8007 (N_8007,N_5969,N_3535);
nand U8008 (N_8008,N_5885,N_5744);
or U8009 (N_8009,N_5772,N_5103);
nand U8010 (N_8010,N_4604,N_3957);
or U8011 (N_8011,N_3704,N_4115);
and U8012 (N_8012,N_3431,N_5578);
nor U8013 (N_8013,N_5247,N_4677);
and U8014 (N_8014,N_5375,N_4520);
nor U8015 (N_8015,N_4932,N_4388);
or U8016 (N_8016,N_5329,N_5704);
nand U8017 (N_8017,N_4307,N_4223);
nand U8018 (N_8018,N_4786,N_4569);
nor U8019 (N_8019,N_4181,N_3963);
nand U8020 (N_8020,N_5629,N_4330);
or U8021 (N_8021,N_4631,N_4278);
or U8022 (N_8022,N_4919,N_5281);
nand U8023 (N_8023,N_4683,N_3079);
and U8024 (N_8024,N_3312,N_5729);
nand U8025 (N_8025,N_5701,N_5062);
nor U8026 (N_8026,N_5212,N_3599);
or U8027 (N_8027,N_4477,N_4676);
and U8028 (N_8028,N_5218,N_3733);
xor U8029 (N_8029,N_3187,N_5470);
and U8030 (N_8030,N_5897,N_3710);
or U8031 (N_8031,N_3724,N_4957);
nand U8032 (N_8032,N_4733,N_4375);
and U8033 (N_8033,N_5636,N_5644);
or U8034 (N_8034,N_5719,N_5312);
nand U8035 (N_8035,N_3444,N_5441);
or U8036 (N_8036,N_3915,N_4198);
and U8037 (N_8037,N_3344,N_4309);
nor U8038 (N_8038,N_4893,N_5292);
nor U8039 (N_8039,N_5813,N_5664);
nor U8040 (N_8040,N_5801,N_5494);
nand U8041 (N_8041,N_3759,N_3173);
and U8042 (N_8042,N_5119,N_4974);
nand U8043 (N_8043,N_3165,N_5680);
nor U8044 (N_8044,N_3617,N_5103);
and U8045 (N_8045,N_3034,N_5311);
nor U8046 (N_8046,N_4242,N_4832);
xor U8047 (N_8047,N_3163,N_5933);
xnor U8048 (N_8048,N_3603,N_3675);
or U8049 (N_8049,N_5560,N_3102);
or U8050 (N_8050,N_5387,N_3474);
nand U8051 (N_8051,N_5774,N_3641);
nor U8052 (N_8052,N_3699,N_3702);
or U8053 (N_8053,N_5864,N_4865);
and U8054 (N_8054,N_5046,N_5038);
and U8055 (N_8055,N_4768,N_5614);
nor U8056 (N_8056,N_3865,N_3326);
xnor U8057 (N_8057,N_5616,N_4294);
and U8058 (N_8058,N_5453,N_3581);
nand U8059 (N_8059,N_3441,N_3690);
nor U8060 (N_8060,N_3089,N_4089);
xor U8061 (N_8061,N_4668,N_4540);
nand U8062 (N_8062,N_5694,N_3467);
and U8063 (N_8063,N_3109,N_4876);
and U8064 (N_8064,N_5517,N_5429);
xor U8065 (N_8065,N_4290,N_5314);
nor U8066 (N_8066,N_3285,N_4639);
nor U8067 (N_8067,N_3417,N_3663);
nand U8068 (N_8068,N_3797,N_3115);
and U8069 (N_8069,N_4495,N_3388);
nor U8070 (N_8070,N_3770,N_5470);
nor U8071 (N_8071,N_4678,N_4281);
or U8072 (N_8072,N_3969,N_5814);
nand U8073 (N_8073,N_4887,N_3537);
nand U8074 (N_8074,N_5090,N_4428);
nand U8075 (N_8075,N_4140,N_3747);
nand U8076 (N_8076,N_4892,N_5365);
nor U8077 (N_8077,N_3470,N_3372);
nor U8078 (N_8078,N_5857,N_5393);
xnor U8079 (N_8079,N_4249,N_5652);
and U8080 (N_8080,N_5786,N_5704);
nor U8081 (N_8081,N_4958,N_4352);
nand U8082 (N_8082,N_5032,N_3549);
nor U8083 (N_8083,N_5163,N_5063);
and U8084 (N_8084,N_4311,N_3129);
or U8085 (N_8085,N_4075,N_5260);
or U8086 (N_8086,N_4217,N_5809);
or U8087 (N_8087,N_3236,N_3230);
nor U8088 (N_8088,N_3073,N_5695);
nand U8089 (N_8089,N_3734,N_4801);
nor U8090 (N_8090,N_3058,N_3702);
and U8091 (N_8091,N_3965,N_5564);
nor U8092 (N_8092,N_3731,N_4872);
nor U8093 (N_8093,N_5545,N_4593);
nand U8094 (N_8094,N_3777,N_4976);
xor U8095 (N_8095,N_4440,N_3427);
or U8096 (N_8096,N_5855,N_5297);
or U8097 (N_8097,N_4509,N_4546);
nor U8098 (N_8098,N_4054,N_3769);
nand U8099 (N_8099,N_5207,N_3275);
nand U8100 (N_8100,N_4004,N_4587);
and U8101 (N_8101,N_3553,N_4215);
xnor U8102 (N_8102,N_4687,N_5264);
and U8103 (N_8103,N_3397,N_4019);
nor U8104 (N_8104,N_4625,N_3234);
nand U8105 (N_8105,N_3167,N_3004);
or U8106 (N_8106,N_3827,N_3964);
or U8107 (N_8107,N_4300,N_5361);
and U8108 (N_8108,N_4107,N_4938);
and U8109 (N_8109,N_5167,N_5472);
nor U8110 (N_8110,N_5824,N_3344);
xor U8111 (N_8111,N_3959,N_5363);
xor U8112 (N_8112,N_5225,N_3342);
nand U8113 (N_8113,N_3458,N_5347);
nor U8114 (N_8114,N_4938,N_5558);
and U8115 (N_8115,N_3418,N_4434);
nand U8116 (N_8116,N_4553,N_3018);
nor U8117 (N_8117,N_5327,N_3214);
xnor U8118 (N_8118,N_3355,N_5995);
nor U8119 (N_8119,N_3495,N_4842);
nor U8120 (N_8120,N_5504,N_3035);
nor U8121 (N_8121,N_3014,N_5956);
nor U8122 (N_8122,N_4787,N_5058);
nor U8123 (N_8123,N_5171,N_3228);
or U8124 (N_8124,N_4075,N_5493);
xnor U8125 (N_8125,N_4180,N_5835);
or U8126 (N_8126,N_4263,N_4232);
or U8127 (N_8127,N_4591,N_5651);
xor U8128 (N_8128,N_4877,N_5945);
nand U8129 (N_8129,N_3428,N_4728);
and U8130 (N_8130,N_5092,N_4883);
xor U8131 (N_8131,N_4769,N_4590);
or U8132 (N_8132,N_3392,N_4503);
or U8133 (N_8133,N_4376,N_4382);
nor U8134 (N_8134,N_4154,N_4766);
and U8135 (N_8135,N_5206,N_5004);
nand U8136 (N_8136,N_4899,N_4135);
or U8137 (N_8137,N_5807,N_5713);
and U8138 (N_8138,N_3539,N_4988);
nor U8139 (N_8139,N_3688,N_4052);
or U8140 (N_8140,N_3533,N_4505);
nor U8141 (N_8141,N_4511,N_4289);
or U8142 (N_8142,N_5968,N_4722);
nand U8143 (N_8143,N_4899,N_3253);
or U8144 (N_8144,N_4817,N_3201);
nand U8145 (N_8145,N_5712,N_5297);
or U8146 (N_8146,N_4295,N_3171);
nor U8147 (N_8147,N_5390,N_5238);
xor U8148 (N_8148,N_4377,N_4831);
nor U8149 (N_8149,N_4283,N_5991);
xnor U8150 (N_8150,N_4332,N_5467);
xnor U8151 (N_8151,N_5459,N_5951);
nor U8152 (N_8152,N_4065,N_5994);
or U8153 (N_8153,N_5588,N_3059);
or U8154 (N_8154,N_4401,N_3572);
and U8155 (N_8155,N_4296,N_4872);
and U8156 (N_8156,N_5810,N_4549);
and U8157 (N_8157,N_5531,N_3639);
or U8158 (N_8158,N_4814,N_5317);
nor U8159 (N_8159,N_3684,N_5294);
xor U8160 (N_8160,N_5433,N_4290);
and U8161 (N_8161,N_4602,N_4095);
and U8162 (N_8162,N_4585,N_4078);
or U8163 (N_8163,N_3285,N_5729);
nand U8164 (N_8164,N_5896,N_3665);
nor U8165 (N_8165,N_3362,N_3496);
nor U8166 (N_8166,N_3751,N_3387);
or U8167 (N_8167,N_5392,N_5477);
or U8168 (N_8168,N_5318,N_4407);
nand U8169 (N_8169,N_4519,N_3746);
and U8170 (N_8170,N_5626,N_4952);
nand U8171 (N_8171,N_4091,N_4000);
xor U8172 (N_8172,N_5155,N_5230);
and U8173 (N_8173,N_5785,N_4422);
nand U8174 (N_8174,N_3269,N_5195);
and U8175 (N_8175,N_5726,N_5929);
or U8176 (N_8176,N_4306,N_5282);
or U8177 (N_8177,N_4787,N_5305);
xnor U8178 (N_8178,N_4391,N_3132);
nand U8179 (N_8179,N_4040,N_4697);
or U8180 (N_8180,N_3629,N_5016);
nand U8181 (N_8181,N_5055,N_3972);
nand U8182 (N_8182,N_5975,N_5688);
and U8183 (N_8183,N_4981,N_4290);
and U8184 (N_8184,N_4417,N_4824);
and U8185 (N_8185,N_5694,N_3516);
and U8186 (N_8186,N_4914,N_5246);
nor U8187 (N_8187,N_4034,N_5093);
xor U8188 (N_8188,N_3764,N_5557);
nand U8189 (N_8189,N_4942,N_5535);
xor U8190 (N_8190,N_3844,N_4813);
nand U8191 (N_8191,N_3428,N_3383);
or U8192 (N_8192,N_4835,N_5038);
and U8193 (N_8193,N_4673,N_5812);
and U8194 (N_8194,N_4917,N_4903);
and U8195 (N_8195,N_3345,N_4545);
nand U8196 (N_8196,N_5329,N_3070);
nand U8197 (N_8197,N_3972,N_3892);
nor U8198 (N_8198,N_3045,N_5242);
and U8199 (N_8199,N_5972,N_3423);
and U8200 (N_8200,N_3036,N_5183);
nor U8201 (N_8201,N_4788,N_4393);
or U8202 (N_8202,N_4698,N_4684);
nor U8203 (N_8203,N_3523,N_4060);
nor U8204 (N_8204,N_4761,N_3203);
nor U8205 (N_8205,N_4882,N_5816);
and U8206 (N_8206,N_5998,N_5371);
or U8207 (N_8207,N_4473,N_3399);
nand U8208 (N_8208,N_3586,N_4603);
nor U8209 (N_8209,N_3603,N_4811);
nor U8210 (N_8210,N_3079,N_5249);
and U8211 (N_8211,N_5719,N_5045);
nand U8212 (N_8212,N_5847,N_4016);
and U8213 (N_8213,N_3087,N_3576);
nor U8214 (N_8214,N_5375,N_3687);
and U8215 (N_8215,N_5255,N_5625);
and U8216 (N_8216,N_4518,N_5961);
and U8217 (N_8217,N_5315,N_4751);
or U8218 (N_8218,N_5564,N_4389);
xor U8219 (N_8219,N_4490,N_5435);
or U8220 (N_8220,N_4099,N_4741);
and U8221 (N_8221,N_4767,N_3224);
and U8222 (N_8222,N_4588,N_3936);
nor U8223 (N_8223,N_4296,N_5147);
nor U8224 (N_8224,N_5741,N_4771);
or U8225 (N_8225,N_4056,N_5441);
nor U8226 (N_8226,N_5830,N_5191);
xnor U8227 (N_8227,N_3915,N_5620);
and U8228 (N_8228,N_4895,N_5869);
nand U8229 (N_8229,N_3346,N_3254);
nor U8230 (N_8230,N_4650,N_4249);
and U8231 (N_8231,N_3932,N_4752);
and U8232 (N_8232,N_4533,N_5793);
nand U8233 (N_8233,N_3577,N_5557);
xor U8234 (N_8234,N_3694,N_4130);
and U8235 (N_8235,N_5713,N_3919);
and U8236 (N_8236,N_5148,N_3935);
nand U8237 (N_8237,N_4145,N_5940);
xor U8238 (N_8238,N_3090,N_4652);
and U8239 (N_8239,N_3448,N_5993);
nand U8240 (N_8240,N_4475,N_4739);
nor U8241 (N_8241,N_4856,N_3718);
and U8242 (N_8242,N_5766,N_4199);
or U8243 (N_8243,N_3997,N_3628);
or U8244 (N_8244,N_5092,N_3588);
and U8245 (N_8245,N_4718,N_4623);
and U8246 (N_8246,N_4447,N_5777);
and U8247 (N_8247,N_4496,N_5949);
nand U8248 (N_8248,N_4884,N_4854);
and U8249 (N_8249,N_5419,N_5290);
and U8250 (N_8250,N_3000,N_4477);
nor U8251 (N_8251,N_3567,N_4968);
and U8252 (N_8252,N_3509,N_3985);
nor U8253 (N_8253,N_5503,N_4919);
nor U8254 (N_8254,N_4229,N_5202);
nor U8255 (N_8255,N_5066,N_3602);
nor U8256 (N_8256,N_5908,N_4937);
or U8257 (N_8257,N_5183,N_5675);
nand U8258 (N_8258,N_3545,N_3524);
nor U8259 (N_8259,N_4150,N_4398);
nor U8260 (N_8260,N_5551,N_5539);
nand U8261 (N_8261,N_4047,N_4377);
or U8262 (N_8262,N_5644,N_3843);
and U8263 (N_8263,N_3440,N_5083);
or U8264 (N_8264,N_5770,N_5989);
and U8265 (N_8265,N_4324,N_3242);
nand U8266 (N_8266,N_3575,N_5200);
nand U8267 (N_8267,N_3466,N_3386);
nand U8268 (N_8268,N_4205,N_4400);
nand U8269 (N_8269,N_4490,N_3829);
and U8270 (N_8270,N_4883,N_3343);
nand U8271 (N_8271,N_5278,N_5588);
or U8272 (N_8272,N_4739,N_4978);
nor U8273 (N_8273,N_5088,N_3356);
or U8274 (N_8274,N_4871,N_3357);
and U8275 (N_8275,N_4694,N_5870);
or U8276 (N_8276,N_3988,N_4904);
nor U8277 (N_8277,N_3487,N_3854);
xor U8278 (N_8278,N_3306,N_4936);
and U8279 (N_8279,N_5858,N_5456);
xor U8280 (N_8280,N_4617,N_5606);
or U8281 (N_8281,N_4151,N_4690);
or U8282 (N_8282,N_5569,N_5062);
xor U8283 (N_8283,N_5058,N_5050);
and U8284 (N_8284,N_3239,N_4980);
nor U8285 (N_8285,N_3828,N_5486);
or U8286 (N_8286,N_5685,N_3218);
nor U8287 (N_8287,N_5021,N_4598);
nand U8288 (N_8288,N_5487,N_3855);
or U8289 (N_8289,N_5672,N_3039);
nand U8290 (N_8290,N_5855,N_5607);
or U8291 (N_8291,N_4084,N_5466);
nand U8292 (N_8292,N_5193,N_3260);
nor U8293 (N_8293,N_4578,N_3390);
and U8294 (N_8294,N_5477,N_4167);
nand U8295 (N_8295,N_3626,N_4096);
nor U8296 (N_8296,N_5430,N_5483);
and U8297 (N_8297,N_5637,N_3338);
nor U8298 (N_8298,N_4205,N_3465);
and U8299 (N_8299,N_5425,N_4378);
nor U8300 (N_8300,N_4664,N_5322);
and U8301 (N_8301,N_4178,N_4961);
and U8302 (N_8302,N_3726,N_5742);
and U8303 (N_8303,N_5819,N_4346);
nand U8304 (N_8304,N_3360,N_4149);
and U8305 (N_8305,N_4073,N_5422);
nand U8306 (N_8306,N_3796,N_3890);
nor U8307 (N_8307,N_5109,N_3968);
or U8308 (N_8308,N_4743,N_4583);
or U8309 (N_8309,N_5418,N_3329);
or U8310 (N_8310,N_5083,N_3615);
nor U8311 (N_8311,N_3332,N_5453);
and U8312 (N_8312,N_5845,N_4183);
and U8313 (N_8313,N_4351,N_5418);
or U8314 (N_8314,N_4012,N_3186);
nand U8315 (N_8315,N_5162,N_4172);
or U8316 (N_8316,N_4579,N_3307);
nand U8317 (N_8317,N_3418,N_4757);
nor U8318 (N_8318,N_4664,N_3133);
and U8319 (N_8319,N_4819,N_4943);
or U8320 (N_8320,N_4807,N_5912);
nor U8321 (N_8321,N_3675,N_3084);
or U8322 (N_8322,N_4842,N_4498);
and U8323 (N_8323,N_5109,N_3929);
nor U8324 (N_8324,N_5291,N_3878);
nand U8325 (N_8325,N_3644,N_4645);
or U8326 (N_8326,N_5730,N_4210);
and U8327 (N_8327,N_5370,N_3838);
nor U8328 (N_8328,N_4759,N_5841);
nor U8329 (N_8329,N_5264,N_4277);
nand U8330 (N_8330,N_3428,N_3768);
nor U8331 (N_8331,N_4292,N_3819);
and U8332 (N_8332,N_3170,N_4615);
nand U8333 (N_8333,N_4668,N_4649);
and U8334 (N_8334,N_3983,N_3933);
and U8335 (N_8335,N_4606,N_4453);
and U8336 (N_8336,N_4992,N_3453);
or U8337 (N_8337,N_3920,N_5207);
xor U8338 (N_8338,N_4031,N_3081);
or U8339 (N_8339,N_3554,N_3056);
or U8340 (N_8340,N_3580,N_4440);
xor U8341 (N_8341,N_3718,N_3389);
or U8342 (N_8342,N_3244,N_3521);
or U8343 (N_8343,N_5468,N_5854);
and U8344 (N_8344,N_5730,N_5374);
and U8345 (N_8345,N_5193,N_5217);
and U8346 (N_8346,N_4445,N_5264);
xor U8347 (N_8347,N_4005,N_3941);
xor U8348 (N_8348,N_4543,N_5793);
nand U8349 (N_8349,N_3654,N_5473);
and U8350 (N_8350,N_5530,N_5131);
or U8351 (N_8351,N_3323,N_5137);
nand U8352 (N_8352,N_4231,N_4759);
nor U8353 (N_8353,N_5283,N_4093);
and U8354 (N_8354,N_4952,N_5986);
and U8355 (N_8355,N_3478,N_5543);
and U8356 (N_8356,N_5442,N_5311);
xor U8357 (N_8357,N_4817,N_3300);
and U8358 (N_8358,N_4773,N_5469);
xor U8359 (N_8359,N_4792,N_4162);
xnor U8360 (N_8360,N_5641,N_4459);
or U8361 (N_8361,N_4727,N_3415);
and U8362 (N_8362,N_3632,N_5237);
and U8363 (N_8363,N_5344,N_3910);
and U8364 (N_8364,N_5678,N_3929);
or U8365 (N_8365,N_4544,N_5268);
xor U8366 (N_8366,N_4154,N_5060);
or U8367 (N_8367,N_5869,N_3979);
or U8368 (N_8368,N_5640,N_5028);
nand U8369 (N_8369,N_4081,N_5644);
nor U8370 (N_8370,N_5638,N_4617);
and U8371 (N_8371,N_5491,N_3009);
nand U8372 (N_8372,N_5311,N_5372);
or U8373 (N_8373,N_4976,N_5125);
or U8374 (N_8374,N_3043,N_5837);
or U8375 (N_8375,N_3711,N_3558);
or U8376 (N_8376,N_4556,N_3689);
or U8377 (N_8377,N_4226,N_5758);
nand U8378 (N_8378,N_5550,N_4553);
and U8379 (N_8379,N_3619,N_5610);
or U8380 (N_8380,N_4453,N_5561);
nand U8381 (N_8381,N_4587,N_3448);
xor U8382 (N_8382,N_4585,N_3124);
or U8383 (N_8383,N_3683,N_5477);
xor U8384 (N_8384,N_3893,N_5785);
or U8385 (N_8385,N_5463,N_4620);
nor U8386 (N_8386,N_3441,N_5133);
nand U8387 (N_8387,N_4074,N_5733);
and U8388 (N_8388,N_5630,N_4643);
and U8389 (N_8389,N_3568,N_4083);
nand U8390 (N_8390,N_3385,N_5108);
nor U8391 (N_8391,N_5539,N_3957);
nand U8392 (N_8392,N_5151,N_3136);
nand U8393 (N_8393,N_4324,N_4132);
nor U8394 (N_8394,N_3071,N_4075);
or U8395 (N_8395,N_4457,N_5297);
nand U8396 (N_8396,N_4070,N_4613);
nor U8397 (N_8397,N_3361,N_5695);
and U8398 (N_8398,N_5959,N_5853);
nor U8399 (N_8399,N_5374,N_3105);
and U8400 (N_8400,N_4826,N_5318);
xnor U8401 (N_8401,N_5246,N_5774);
or U8402 (N_8402,N_3043,N_4699);
nor U8403 (N_8403,N_3867,N_3144);
xnor U8404 (N_8404,N_3253,N_4304);
or U8405 (N_8405,N_5728,N_3408);
and U8406 (N_8406,N_5811,N_4468);
xor U8407 (N_8407,N_5940,N_4359);
or U8408 (N_8408,N_5447,N_5293);
nand U8409 (N_8409,N_4058,N_5434);
and U8410 (N_8410,N_3210,N_4262);
xor U8411 (N_8411,N_5508,N_3490);
and U8412 (N_8412,N_3933,N_3885);
or U8413 (N_8413,N_3512,N_5712);
xor U8414 (N_8414,N_3157,N_3564);
and U8415 (N_8415,N_5457,N_4659);
and U8416 (N_8416,N_5174,N_5336);
nand U8417 (N_8417,N_5654,N_3166);
nor U8418 (N_8418,N_4531,N_3164);
or U8419 (N_8419,N_4929,N_3743);
or U8420 (N_8420,N_4815,N_4896);
and U8421 (N_8421,N_4134,N_4561);
nand U8422 (N_8422,N_5194,N_4444);
nor U8423 (N_8423,N_3899,N_5635);
or U8424 (N_8424,N_3378,N_3374);
nand U8425 (N_8425,N_5596,N_3388);
or U8426 (N_8426,N_3258,N_5002);
or U8427 (N_8427,N_4406,N_5707);
nor U8428 (N_8428,N_4149,N_3108);
or U8429 (N_8429,N_3218,N_3614);
or U8430 (N_8430,N_3069,N_5425);
and U8431 (N_8431,N_3867,N_4373);
or U8432 (N_8432,N_3623,N_3854);
and U8433 (N_8433,N_5048,N_4802);
and U8434 (N_8434,N_5548,N_3425);
or U8435 (N_8435,N_4608,N_3601);
nor U8436 (N_8436,N_4509,N_4323);
and U8437 (N_8437,N_5860,N_4421);
or U8438 (N_8438,N_3211,N_3892);
nor U8439 (N_8439,N_3399,N_3409);
xor U8440 (N_8440,N_3848,N_3046);
xnor U8441 (N_8441,N_5812,N_4602);
and U8442 (N_8442,N_5227,N_3181);
nand U8443 (N_8443,N_3144,N_4978);
and U8444 (N_8444,N_3169,N_5730);
and U8445 (N_8445,N_3830,N_4921);
nor U8446 (N_8446,N_3252,N_4567);
nor U8447 (N_8447,N_5255,N_4390);
nor U8448 (N_8448,N_5754,N_5974);
and U8449 (N_8449,N_3292,N_3068);
nand U8450 (N_8450,N_4170,N_5213);
or U8451 (N_8451,N_3535,N_3364);
nand U8452 (N_8452,N_3585,N_3897);
nor U8453 (N_8453,N_3679,N_5862);
xor U8454 (N_8454,N_4175,N_3569);
and U8455 (N_8455,N_3950,N_3330);
nand U8456 (N_8456,N_3409,N_4599);
and U8457 (N_8457,N_3998,N_3891);
nand U8458 (N_8458,N_4893,N_5058);
or U8459 (N_8459,N_4270,N_4767);
and U8460 (N_8460,N_3697,N_5193);
xor U8461 (N_8461,N_4109,N_4933);
and U8462 (N_8462,N_3480,N_4066);
nor U8463 (N_8463,N_3073,N_3521);
nor U8464 (N_8464,N_3521,N_4540);
and U8465 (N_8465,N_5675,N_3565);
nand U8466 (N_8466,N_3084,N_3615);
nand U8467 (N_8467,N_3907,N_5117);
nand U8468 (N_8468,N_4443,N_5421);
or U8469 (N_8469,N_4824,N_3373);
or U8470 (N_8470,N_5781,N_3888);
nor U8471 (N_8471,N_3022,N_3433);
nand U8472 (N_8472,N_4155,N_4262);
nand U8473 (N_8473,N_4378,N_3590);
nand U8474 (N_8474,N_5123,N_4091);
nand U8475 (N_8475,N_3743,N_3381);
or U8476 (N_8476,N_5857,N_4958);
or U8477 (N_8477,N_4029,N_5567);
xnor U8478 (N_8478,N_5862,N_4521);
nand U8479 (N_8479,N_3902,N_3603);
nor U8480 (N_8480,N_3102,N_4392);
nand U8481 (N_8481,N_5579,N_3476);
nand U8482 (N_8482,N_5010,N_3770);
or U8483 (N_8483,N_3172,N_4699);
nor U8484 (N_8484,N_3667,N_5367);
and U8485 (N_8485,N_4352,N_4603);
or U8486 (N_8486,N_3585,N_4774);
and U8487 (N_8487,N_5561,N_3050);
or U8488 (N_8488,N_5887,N_3011);
or U8489 (N_8489,N_4217,N_4042);
nand U8490 (N_8490,N_5433,N_5507);
and U8491 (N_8491,N_4399,N_4620);
or U8492 (N_8492,N_4898,N_4644);
or U8493 (N_8493,N_4134,N_4495);
nand U8494 (N_8494,N_4829,N_4389);
and U8495 (N_8495,N_3956,N_3494);
or U8496 (N_8496,N_5587,N_3089);
nor U8497 (N_8497,N_4731,N_3803);
xor U8498 (N_8498,N_5695,N_3656);
nand U8499 (N_8499,N_5555,N_5937);
nand U8500 (N_8500,N_5154,N_4836);
and U8501 (N_8501,N_3303,N_5662);
nand U8502 (N_8502,N_5619,N_5686);
nor U8503 (N_8503,N_4261,N_4476);
and U8504 (N_8504,N_5383,N_4568);
or U8505 (N_8505,N_4807,N_3061);
or U8506 (N_8506,N_5346,N_4479);
and U8507 (N_8507,N_5515,N_5320);
xor U8508 (N_8508,N_3024,N_3014);
or U8509 (N_8509,N_3147,N_5977);
or U8510 (N_8510,N_4514,N_5377);
xor U8511 (N_8511,N_3439,N_3672);
nand U8512 (N_8512,N_4975,N_3174);
or U8513 (N_8513,N_4758,N_4211);
xnor U8514 (N_8514,N_3712,N_4919);
nand U8515 (N_8515,N_5846,N_5336);
nor U8516 (N_8516,N_4016,N_5733);
nand U8517 (N_8517,N_3598,N_5807);
and U8518 (N_8518,N_4309,N_3162);
and U8519 (N_8519,N_5333,N_3083);
or U8520 (N_8520,N_5053,N_4215);
nor U8521 (N_8521,N_5731,N_4514);
nand U8522 (N_8522,N_4358,N_3749);
nor U8523 (N_8523,N_5137,N_3027);
xnor U8524 (N_8524,N_4775,N_3032);
or U8525 (N_8525,N_5566,N_5912);
nor U8526 (N_8526,N_3320,N_3431);
nor U8527 (N_8527,N_3174,N_4011);
and U8528 (N_8528,N_5608,N_5915);
nand U8529 (N_8529,N_5329,N_4556);
nand U8530 (N_8530,N_5736,N_3651);
nand U8531 (N_8531,N_3606,N_5954);
and U8532 (N_8532,N_4462,N_5592);
and U8533 (N_8533,N_3650,N_5476);
and U8534 (N_8534,N_3773,N_5873);
and U8535 (N_8535,N_5264,N_5661);
nand U8536 (N_8536,N_3203,N_3299);
and U8537 (N_8537,N_3257,N_4722);
nand U8538 (N_8538,N_5767,N_3991);
nand U8539 (N_8539,N_3672,N_5360);
nor U8540 (N_8540,N_3888,N_3279);
nor U8541 (N_8541,N_5793,N_5049);
or U8542 (N_8542,N_5430,N_5787);
xnor U8543 (N_8543,N_4673,N_4688);
or U8544 (N_8544,N_5714,N_5762);
or U8545 (N_8545,N_3558,N_5371);
and U8546 (N_8546,N_3599,N_5943);
or U8547 (N_8547,N_3586,N_3610);
nor U8548 (N_8548,N_4038,N_3964);
or U8549 (N_8549,N_5505,N_4852);
nand U8550 (N_8550,N_3796,N_4095);
nor U8551 (N_8551,N_3496,N_5621);
or U8552 (N_8552,N_4309,N_3219);
and U8553 (N_8553,N_4135,N_3131);
and U8554 (N_8554,N_5301,N_4270);
or U8555 (N_8555,N_5521,N_3286);
and U8556 (N_8556,N_5360,N_3341);
nor U8557 (N_8557,N_3619,N_5327);
nor U8558 (N_8558,N_5615,N_3157);
or U8559 (N_8559,N_4451,N_3220);
nor U8560 (N_8560,N_3630,N_5419);
xnor U8561 (N_8561,N_4188,N_3142);
xnor U8562 (N_8562,N_5761,N_5039);
and U8563 (N_8563,N_3004,N_3635);
xnor U8564 (N_8564,N_4442,N_3096);
nor U8565 (N_8565,N_5478,N_4465);
nor U8566 (N_8566,N_5584,N_3158);
nor U8567 (N_8567,N_5630,N_5953);
nor U8568 (N_8568,N_4316,N_4203);
nor U8569 (N_8569,N_4177,N_3823);
xnor U8570 (N_8570,N_3115,N_5600);
xor U8571 (N_8571,N_3388,N_5060);
nor U8572 (N_8572,N_3029,N_5335);
or U8573 (N_8573,N_4098,N_3913);
nand U8574 (N_8574,N_5400,N_3576);
xor U8575 (N_8575,N_3718,N_4311);
and U8576 (N_8576,N_3835,N_5176);
or U8577 (N_8577,N_5428,N_4128);
or U8578 (N_8578,N_4753,N_4736);
nand U8579 (N_8579,N_3777,N_3239);
xor U8580 (N_8580,N_4533,N_3072);
nand U8581 (N_8581,N_5631,N_3212);
and U8582 (N_8582,N_4809,N_4231);
and U8583 (N_8583,N_5412,N_4608);
nor U8584 (N_8584,N_4029,N_5825);
and U8585 (N_8585,N_5732,N_3780);
and U8586 (N_8586,N_4224,N_5544);
and U8587 (N_8587,N_4758,N_3207);
and U8588 (N_8588,N_5702,N_3752);
or U8589 (N_8589,N_4224,N_4510);
or U8590 (N_8590,N_3366,N_5415);
nand U8591 (N_8591,N_4980,N_4589);
nor U8592 (N_8592,N_4242,N_4605);
and U8593 (N_8593,N_3104,N_5417);
xor U8594 (N_8594,N_3116,N_4497);
and U8595 (N_8595,N_5317,N_5566);
nand U8596 (N_8596,N_4046,N_4432);
nor U8597 (N_8597,N_5007,N_3570);
nand U8598 (N_8598,N_5372,N_4969);
and U8599 (N_8599,N_5699,N_3059);
nand U8600 (N_8600,N_3924,N_3936);
nor U8601 (N_8601,N_3658,N_5130);
nor U8602 (N_8602,N_5288,N_4130);
or U8603 (N_8603,N_5862,N_5556);
nor U8604 (N_8604,N_4176,N_5741);
nand U8605 (N_8605,N_3684,N_5995);
nand U8606 (N_8606,N_4010,N_4438);
or U8607 (N_8607,N_5254,N_5813);
or U8608 (N_8608,N_3772,N_4096);
nor U8609 (N_8609,N_5887,N_4772);
and U8610 (N_8610,N_3877,N_4820);
or U8611 (N_8611,N_5746,N_5933);
nor U8612 (N_8612,N_3001,N_5067);
xor U8613 (N_8613,N_3348,N_5029);
and U8614 (N_8614,N_5806,N_3891);
and U8615 (N_8615,N_4407,N_5127);
nor U8616 (N_8616,N_3338,N_4584);
nand U8617 (N_8617,N_5893,N_4778);
or U8618 (N_8618,N_3872,N_3709);
or U8619 (N_8619,N_3516,N_4054);
and U8620 (N_8620,N_4071,N_4363);
and U8621 (N_8621,N_4681,N_5089);
nor U8622 (N_8622,N_4977,N_3023);
nand U8623 (N_8623,N_3403,N_4486);
nor U8624 (N_8624,N_4094,N_3401);
and U8625 (N_8625,N_5787,N_5445);
nand U8626 (N_8626,N_5786,N_3905);
nand U8627 (N_8627,N_4677,N_4997);
or U8628 (N_8628,N_5380,N_3457);
or U8629 (N_8629,N_3760,N_4443);
xnor U8630 (N_8630,N_5156,N_4474);
nand U8631 (N_8631,N_3752,N_3600);
or U8632 (N_8632,N_5851,N_3741);
or U8633 (N_8633,N_4986,N_5181);
nand U8634 (N_8634,N_5672,N_5850);
nor U8635 (N_8635,N_3971,N_5558);
or U8636 (N_8636,N_3102,N_3492);
and U8637 (N_8637,N_3812,N_3312);
nand U8638 (N_8638,N_5615,N_3878);
nand U8639 (N_8639,N_5804,N_4443);
or U8640 (N_8640,N_3782,N_5146);
and U8641 (N_8641,N_4189,N_3488);
or U8642 (N_8642,N_4075,N_4170);
xor U8643 (N_8643,N_5610,N_5757);
and U8644 (N_8644,N_4612,N_3242);
xor U8645 (N_8645,N_3661,N_3963);
and U8646 (N_8646,N_5113,N_4074);
and U8647 (N_8647,N_4387,N_4069);
nor U8648 (N_8648,N_4403,N_5306);
nor U8649 (N_8649,N_4197,N_4517);
nand U8650 (N_8650,N_4672,N_4687);
nand U8651 (N_8651,N_3438,N_4802);
nor U8652 (N_8652,N_4975,N_3091);
nor U8653 (N_8653,N_4177,N_3542);
nor U8654 (N_8654,N_3730,N_4211);
nand U8655 (N_8655,N_5949,N_3445);
nand U8656 (N_8656,N_4769,N_3966);
nand U8657 (N_8657,N_4727,N_4992);
and U8658 (N_8658,N_4204,N_4937);
nor U8659 (N_8659,N_5013,N_5545);
and U8660 (N_8660,N_3472,N_4717);
or U8661 (N_8661,N_4671,N_4936);
and U8662 (N_8662,N_4062,N_4042);
or U8663 (N_8663,N_5100,N_3974);
xor U8664 (N_8664,N_3819,N_5500);
or U8665 (N_8665,N_4905,N_4891);
and U8666 (N_8666,N_3576,N_4378);
or U8667 (N_8667,N_4155,N_3311);
nor U8668 (N_8668,N_4837,N_3013);
nand U8669 (N_8669,N_5482,N_5450);
nand U8670 (N_8670,N_4622,N_4252);
and U8671 (N_8671,N_3258,N_4575);
and U8672 (N_8672,N_5239,N_3466);
nor U8673 (N_8673,N_4393,N_4632);
and U8674 (N_8674,N_3270,N_5188);
nor U8675 (N_8675,N_5252,N_3166);
or U8676 (N_8676,N_5683,N_3746);
nand U8677 (N_8677,N_5770,N_5516);
or U8678 (N_8678,N_3790,N_4052);
or U8679 (N_8679,N_4647,N_3518);
nand U8680 (N_8680,N_5875,N_3797);
or U8681 (N_8681,N_4348,N_3673);
nor U8682 (N_8682,N_5872,N_5360);
nor U8683 (N_8683,N_3440,N_4241);
or U8684 (N_8684,N_4796,N_5326);
nor U8685 (N_8685,N_3144,N_5268);
nor U8686 (N_8686,N_4725,N_3992);
nand U8687 (N_8687,N_4119,N_3241);
nor U8688 (N_8688,N_3107,N_3575);
and U8689 (N_8689,N_3729,N_4304);
nor U8690 (N_8690,N_5512,N_5890);
and U8691 (N_8691,N_4052,N_4671);
nand U8692 (N_8692,N_3882,N_5875);
or U8693 (N_8693,N_4237,N_4716);
and U8694 (N_8694,N_3483,N_4017);
nor U8695 (N_8695,N_3601,N_5660);
or U8696 (N_8696,N_4017,N_4692);
nor U8697 (N_8697,N_3945,N_4855);
nand U8698 (N_8698,N_4739,N_3010);
nand U8699 (N_8699,N_5467,N_5393);
nor U8700 (N_8700,N_5399,N_4271);
and U8701 (N_8701,N_3864,N_5020);
or U8702 (N_8702,N_4095,N_3292);
nor U8703 (N_8703,N_5757,N_5043);
nand U8704 (N_8704,N_3487,N_5351);
or U8705 (N_8705,N_3181,N_5475);
or U8706 (N_8706,N_3147,N_5765);
and U8707 (N_8707,N_4778,N_3084);
and U8708 (N_8708,N_3067,N_3785);
nor U8709 (N_8709,N_4259,N_5901);
nor U8710 (N_8710,N_3315,N_5340);
nand U8711 (N_8711,N_4149,N_4079);
and U8712 (N_8712,N_3841,N_5954);
nand U8713 (N_8713,N_3657,N_3138);
xnor U8714 (N_8714,N_4647,N_3116);
and U8715 (N_8715,N_4747,N_5482);
nand U8716 (N_8716,N_3919,N_5674);
and U8717 (N_8717,N_3448,N_3676);
nor U8718 (N_8718,N_5695,N_5462);
or U8719 (N_8719,N_5398,N_3053);
and U8720 (N_8720,N_4741,N_3333);
nand U8721 (N_8721,N_4669,N_4744);
and U8722 (N_8722,N_5762,N_5241);
or U8723 (N_8723,N_3616,N_5537);
and U8724 (N_8724,N_5020,N_3279);
nand U8725 (N_8725,N_4194,N_3850);
or U8726 (N_8726,N_4514,N_5817);
nor U8727 (N_8727,N_3030,N_5346);
nor U8728 (N_8728,N_4956,N_4868);
xnor U8729 (N_8729,N_4260,N_5875);
nand U8730 (N_8730,N_5307,N_3255);
or U8731 (N_8731,N_5829,N_4358);
or U8732 (N_8732,N_4697,N_3155);
nand U8733 (N_8733,N_3866,N_5470);
nand U8734 (N_8734,N_5176,N_4418);
and U8735 (N_8735,N_4277,N_3650);
or U8736 (N_8736,N_3919,N_4491);
xor U8737 (N_8737,N_3570,N_3988);
and U8738 (N_8738,N_5033,N_4182);
nand U8739 (N_8739,N_5421,N_3253);
and U8740 (N_8740,N_4409,N_5733);
or U8741 (N_8741,N_3586,N_3969);
nor U8742 (N_8742,N_4422,N_5866);
nor U8743 (N_8743,N_4174,N_5742);
nor U8744 (N_8744,N_4291,N_4397);
or U8745 (N_8745,N_5749,N_3958);
xor U8746 (N_8746,N_3172,N_4906);
nand U8747 (N_8747,N_4374,N_3698);
xnor U8748 (N_8748,N_3479,N_3481);
and U8749 (N_8749,N_5179,N_4968);
or U8750 (N_8750,N_4027,N_3244);
nor U8751 (N_8751,N_4795,N_5808);
or U8752 (N_8752,N_5725,N_5526);
and U8753 (N_8753,N_5184,N_3369);
nor U8754 (N_8754,N_3893,N_4652);
nor U8755 (N_8755,N_5928,N_4563);
nand U8756 (N_8756,N_4349,N_3469);
and U8757 (N_8757,N_5078,N_4748);
and U8758 (N_8758,N_4868,N_5167);
or U8759 (N_8759,N_3640,N_3979);
or U8760 (N_8760,N_3146,N_3728);
nor U8761 (N_8761,N_3696,N_3104);
and U8762 (N_8762,N_4691,N_4764);
nand U8763 (N_8763,N_4428,N_4203);
or U8764 (N_8764,N_4996,N_3402);
or U8765 (N_8765,N_5917,N_3434);
nand U8766 (N_8766,N_5048,N_4331);
and U8767 (N_8767,N_3650,N_5159);
nor U8768 (N_8768,N_3736,N_5707);
nand U8769 (N_8769,N_4726,N_3820);
nor U8770 (N_8770,N_3946,N_4209);
and U8771 (N_8771,N_4320,N_5838);
nor U8772 (N_8772,N_4148,N_4516);
or U8773 (N_8773,N_4691,N_5348);
nor U8774 (N_8774,N_5477,N_4109);
nor U8775 (N_8775,N_4854,N_5121);
nor U8776 (N_8776,N_5100,N_4911);
nand U8777 (N_8777,N_5440,N_4012);
nand U8778 (N_8778,N_5528,N_5880);
nand U8779 (N_8779,N_4024,N_4789);
and U8780 (N_8780,N_5642,N_4573);
nand U8781 (N_8781,N_4870,N_5673);
and U8782 (N_8782,N_3276,N_5716);
and U8783 (N_8783,N_5923,N_4173);
nor U8784 (N_8784,N_4815,N_5327);
and U8785 (N_8785,N_5171,N_4293);
nand U8786 (N_8786,N_4394,N_4730);
nor U8787 (N_8787,N_5533,N_4879);
nor U8788 (N_8788,N_5027,N_4323);
nand U8789 (N_8789,N_5364,N_5848);
nor U8790 (N_8790,N_4624,N_4528);
or U8791 (N_8791,N_3390,N_3620);
and U8792 (N_8792,N_5033,N_3712);
or U8793 (N_8793,N_3052,N_3383);
or U8794 (N_8794,N_5478,N_4100);
xnor U8795 (N_8795,N_3653,N_3853);
and U8796 (N_8796,N_3459,N_5913);
xnor U8797 (N_8797,N_3583,N_5976);
or U8798 (N_8798,N_5964,N_5728);
nand U8799 (N_8799,N_4123,N_5135);
nand U8800 (N_8800,N_4260,N_4738);
and U8801 (N_8801,N_3122,N_3685);
nand U8802 (N_8802,N_3725,N_4628);
or U8803 (N_8803,N_4954,N_5552);
xnor U8804 (N_8804,N_3508,N_5966);
and U8805 (N_8805,N_5060,N_5020);
or U8806 (N_8806,N_3263,N_3431);
nand U8807 (N_8807,N_4811,N_4963);
or U8808 (N_8808,N_3015,N_4549);
and U8809 (N_8809,N_4798,N_4720);
nand U8810 (N_8810,N_5203,N_4151);
nand U8811 (N_8811,N_3014,N_5506);
nor U8812 (N_8812,N_4580,N_4538);
and U8813 (N_8813,N_4227,N_4912);
and U8814 (N_8814,N_5766,N_4342);
or U8815 (N_8815,N_3844,N_3512);
or U8816 (N_8816,N_4743,N_4911);
nor U8817 (N_8817,N_3887,N_3628);
xor U8818 (N_8818,N_3725,N_4094);
and U8819 (N_8819,N_3251,N_5781);
nor U8820 (N_8820,N_5573,N_3292);
nand U8821 (N_8821,N_5324,N_4598);
or U8822 (N_8822,N_5712,N_5783);
nand U8823 (N_8823,N_5105,N_4910);
and U8824 (N_8824,N_5494,N_5683);
or U8825 (N_8825,N_4508,N_4393);
nor U8826 (N_8826,N_3783,N_4694);
nand U8827 (N_8827,N_4380,N_3993);
and U8828 (N_8828,N_5146,N_3956);
nor U8829 (N_8829,N_4959,N_4471);
nor U8830 (N_8830,N_4202,N_3124);
and U8831 (N_8831,N_4995,N_4720);
nand U8832 (N_8832,N_5701,N_3708);
and U8833 (N_8833,N_4597,N_5841);
and U8834 (N_8834,N_4384,N_3022);
nand U8835 (N_8835,N_4546,N_5717);
and U8836 (N_8836,N_4476,N_5940);
and U8837 (N_8837,N_4933,N_4704);
nand U8838 (N_8838,N_3750,N_4594);
and U8839 (N_8839,N_5778,N_5119);
or U8840 (N_8840,N_5901,N_3999);
nor U8841 (N_8841,N_3164,N_3008);
or U8842 (N_8842,N_5714,N_5802);
and U8843 (N_8843,N_3637,N_4774);
or U8844 (N_8844,N_3353,N_4003);
nand U8845 (N_8845,N_3914,N_4591);
or U8846 (N_8846,N_5322,N_4728);
and U8847 (N_8847,N_5929,N_3874);
and U8848 (N_8848,N_4738,N_5806);
nand U8849 (N_8849,N_3380,N_5423);
nand U8850 (N_8850,N_4562,N_3201);
nand U8851 (N_8851,N_4834,N_5421);
and U8852 (N_8852,N_5713,N_4086);
or U8853 (N_8853,N_4310,N_3323);
xor U8854 (N_8854,N_4234,N_3285);
or U8855 (N_8855,N_4196,N_5587);
or U8856 (N_8856,N_5728,N_3005);
or U8857 (N_8857,N_3386,N_5976);
nand U8858 (N_8858,N_3206,N_4033);
or U8859 (N_8859,N_4491,N_4374);
or U8860 (N_8860,N_3414,N_4529);
nand U8861 (N_8861,N_4365,N_4306);
nand U8862 (N_8862,N_5009,N_5065);
and U8863 (N_8863,N_5743,N_4711);
nand U8864 (N_8864,N_3756,N_3930);
or U8865 (N_8865,N_3573,N_4766);
nand U8866 (N_8866,N_3490,N_5015);
xor U8867 (N_8867,N_4448,N_5554);
nor U8868 (N_8868,N_4792,N_5268);
xor U8869 (N_8869,N_3428,N_3328);
and U8870 (N_8870,N_4026,N_5288);
nand U8871 (N_8871,N_5638,N_5149);
xnor U8872 (N_8872,N_3686,N_4262);
nand U8873 (N_8873,N_5302,N_3701);
nand U8874 (N_8874,N_4229,N_5818);
nand U8875 (N_8875,N_3606,N_4728);
and U8876 (N_8876,N_4538,N_4240);
or U8877 (N_8877,N_4986,N_5314);
nor U8878 (N_8878,N_5080,N_4557);
nand U8879 (N_8879,N_5910,N_4594);
nand U8880 (N_8880,N_4079,N_5417);
or U8881 (N_8881,N_3818,N_4830);
nor U8882 (N_8882,N_3612,N_4043);
nor U8883 (N_8883,N_5074,N_3639);
nand U8884 (N_8884,N_4710,N_5626);
and U8885 (N_8885,N_5488,N_3640);
or U8886 (N_8886,N_5379,N_4952);
nor U8887 (N_8887,N_5657,N_5034);
and U8888 (N_8888,N_3628,N_4700);
and U8889 (N_8889,N_5036,N_4749);
and U8890 (N_8890,N_4371,N_4896);
nor U8891 (N_8891,N_3083,N_5068);
nand U8892 (N_8892,N_4617,N_4656);
and U8893 (N_8893,N_3559,N_3834);
nor U8894 (N_8894,N_3520,N_5039);
or U8895 (N_8895,N_5671,N_5409);
nor U8896 (N_8896,N_3986,N_3541);
nand U8897 (N_8897,N_4650,N_4931);
xor U8898 (N_8898,N_4848,N_5044);
nor U8899 (N_8899,N_4142,N_5985);
nand U8900 (N_8900,N_4477,N_3545);
nor U8901 (N_8901,N_5015,N_4034);
or U8902 (N_8902,N_5914,N_5245);
or U8903 (N_8903,N_4185,N_5251);
and U8904 (N_8904,N_4925,N_3751);
or U8905 (N_8905,N_3950,N_5875);
or U8906 (N_8906,N_5296,N_3142);
and U8907 (N_8907,N_5725,N_3162);
or U8908 (N_8908,N_5540,N_3592);
xnor U8909 (N_8909,N_4962,N_4622);
or U8910 (N_8910,N_5384,N_3201);
nor U8911 (N_8911,N_4322,N_3293);
or U8912 (N_8912,N_3584,N_4279);
and U8913 (N_8913,N_3329,N_4208);
nand U8914 (N_8914,N_4959,N_4816);
xor U8915 (N_8915,N_5037,N_4720);
or U8916 (N_8916,N_5531,N_5871);
nand U8917 (N_8917,N_4144,N_4109);
or U8918 (N_8918,N_4414,N_3942);
and U8919 (N_8919,N_4623,N_3600);
xor U8920 (N_8920,N_4479,N_5271);
nor U8921 (N_8921,N_5779,N_5270);
and U8922 (N_8922,N_5294,N_4905);
or U8923 (N_8923,N_5107,N_5948);
nand U8924 (N_8924,N_3326,N_5986);
nand U8925 (N_8925,N_3450,N_4096);
xnor U8926 (N_8926,N_3507,N_5617);
nand U8927 (N_8927,N_4029,N_5497);
nand U8928 (N_8928,N_3676,N_3507);
and U8929 (N_8929,N_5803,N_3278);
and U8930 (N_8930,N_4407,N_5532);
or U8931 (N_8931,N_4575,N_3504);
nor U8932 (N_8932,N_4080,N_5509);
or U8933 (N_8933,N_4940,N_3096);
and U8934 (N_8934,N_3760,N_4940);
and U8935 (N_8935,N_3852,N_4142);
and U8936 (N_8936,N_4499,N_4753);
xor U8937 (N_8937,N_5452,N_3891);
or U8938 (N_8938,N_4286,N_5566);
nor U8939 (N_8939,N_4327,N_4531);
or U8940 (N_8940,N_4538,N_5747);
and U8941 (N_8941,N_3854,N_3031);
nand U8942 (N_8942,N_3575,N_3416);
and U8943 (N_8943,N_5606,N_3431);
nor U8944 (N_8944,N_3163,N_5057);
nor U8945 (N_8945,N_3951,N_3477);
or U8946 (N_8946,N_5847,N_4722);
or U8947 (N_8947,N_5879,N_4674);
nor U8948 (N_8948,N_4261,N_4759);
and U8949 (N_8949,N_3036,N_3694);
nor U8950 (N_8950,N_4242,N_5123);
and U8951 (N_8951,N_5905,N_4888);
and U8952 (N_8952,N_5557,N_5636);
and U8953 (N_8953,N_5033,N_5702);
or U8954 (N_8954,N_3502,N_3131);
or U8955 (N_8955,N_3987,N_4590);
xnor U8956 (N_8956,N_4485,N_4172);
and U8957 (N_8957,N_4647,N_3636);
and U8958 (N_8958,N_3853,N_5401);
and U8959 (N_8959,N_5818,N_5700);
nand U8960 (N_8960,N_3746,N_5665);
nor U8961 (N_8961,N_4145,N_4191);
or U8962 (N_8962,N_5366,N_5620);
nand U8963 (N_8963,N_5225,N_4120);
and U8964 (N_8964,N_4532,N_5557);
nor U8965 (N_8965,N_4648,N_5808);
xnor U8966 (N_8966,N_4452,N_4731);
or U8967 (N_8967,N_3531,N_5974);
nand U8968 (N_8968,N_4599,N_4335);
xnor U8969 (N_8969,N_3296,N_4944);
and U8970 (N_8970,N_4262,N_3464);
nor U8971 (N_8971,N_4389,N_3741);
nand U8972 (N_8972,N_4530,N_5530);
xor U8973 (N_8973,N_4248,N_5694);
nor U8974 (N_8974,N_3152,N_5923);
nor U8975 (N_8975,N_3855,N_4458);
xor U8976 (N_8976,N_3942,N_4174);
nor U8977 (N_8977,N_4169,N_3748);
nand U8978 (N_8978,N_5526,N_4636);
or U8979 (N_8979,N_3346,N_4953);
or U8980 (N_8980,N_4136,N_4037);
or U8981 (N_8981,N_3478,N_5777);
or U8982 (N_8982,N_3155,N_3907);
or U8983 (N_8983,N_4279,N_5203);
nand U8984 (N_8984,N_4044,N_5887);
and U8985 (N_8985,N_4923,N_3705);
and U8986 (N_8986,N_3101,N_4758);
nor U8987 (N_8987,N_3591,N_5283);
nor U8988 (N_8988,N_3562,N_4904);
and U8989 (N_8989,N_5280,N_4401);
nand U8990 (N_8990,N_5928,N_3771);
xor U8991 (N_8991,N_5803,N_3719);
nand U8992 (N_8992,N_3548,N_5107);
and U8993 (N_8993,N_4985,N_5043);
and U8994 (N_8994,N_5546,N_5269);
or U8995 (N_8995,N_4973,N_5698);
or U8996 (N_8996,N_3970,N_4886);
nor U8997 (N_8997,N_5883,N_4074);
or U8998 (N_8998,N_5167,N_3359);
nor U8999 (N_8999,N_3337,N_4402);
and U9000 (N_9000,N_7066,N_6337);
and U9001 (N_9001,N_6142,N_6499);
xnor U9002 (N_9002,N_7762,N_7420);
xnor U9003 (N_9003,N_8178,N_8203);
nand U9004 (N_9004,N_6920,N_8875);
or U9005 (N_9005,N_8416,N_7781);
nor U9006 (N_9006,N_7785,N_8516);
or U9007 (N_9007,N_7570,N_7324);
and U9008 (N_9008,N_7281,N_6533);
nand U9009 (N_9009,N_6619,N_8720);
nor U9010 (N_9010,N_6542,N_7597);
and U9011 (N_9011,N_8149,N_8774);
and U9012 (N_9012,N_6366,N_8307);
nand U9013 (N_9013,N_7106,N_6959);
or U9014 (N_9014,N_7512,N_7796);
nand U9015 (N_9015,N_6438,N_7942);
and U9016 (N_9016,N_6174,N_8739);
xnor U9017 (N_9017,N_8843,N_8487);
nor U9018 (N_9018,N_7121,N_6018);
nand U9019 (N_9019,N_8861,N_7059);
nand U9020 (N_9020,N_6097,N_8294);
and U9021 (N_9021,N_6595,N_6076);
nor U9022 (N_9022,N_6528,N_6033);
and U9023 (N_9023,N_8333,N_6613);
xnor U9024 (N_9024,N_6943,N_8039);
nor U9025 (N_9025,N_6351,N_8618);
nand U9026 (N_9026,N_6704,N_7409);
and U9027 (N_9027,N_6857,N_7936);
or U9028 (N_9028,N_6537,N_8023);
nor U9029 (N_9029,N_8250,N_6709);
nand U9030 (N_9030,N_7923,N_8556);
or U9031 (N_9031,N_6792,N_7323);
xor U9032 (N_9032,N_6056,N_7898);
nand U9033 (N_9033,N_8331,N_6338);
or U9034 (N_9034,N_7929,N_8763);
nand U9035 (N_9035,N_8276,N_6911);
or U9036 (N_9036,N_6095,N_7239);
or U9037 (N_9037,N_8120,N_8508);
and U9038 (N_9038,N_7246,N_7742);
nand U9039 (N_9039,N_6853,N_6517);
xnor U9040 (N_9040,N_7398,N_8346);
and U9041 (N_9041,N_6488,N_6482);
nand U9042 (N_9042,N_7958,N_8765);
or U9043 (N_9043,N_7410,N_8850);
and U9044 (N_9044,N_8075,N_7071);
and U9045 (N_9045,N_8891,N_6820);
nor U9046 (N_9046,N_7542,N_7452);
nor U9047 (N_9047,N_8472,N_8274);
or U9048 (N_9048,N_8478,N_8283);
nand U9049 (N_9049,N_8839,N_6627);
xor U9050 (N_9050,N_6070,N_6423);
nor U9051 (N_9051,N_8162,N_8696);
or U9052 (N_9052,N_8224,N_8725);
or U9053 (N_9053,N_8761,N_7481);
nand U9054 (N_9054,N_8738,N_8393);
or U9055 (N_9055,N_7435,N_7102);
nand U9056 (N_9056,N_6526,N_7661);
nor U9057 (N_9057,N_7638,N_8076);
nand U9058 (N_9058,N_7617,N_7747);
and U9059 (N_9059,N_8827,N_6226);
and U9060 (N_9060,N_6635,N_7471);
nand U9061 (N_9061,N_8954,N_7133);
nand U9062 (N_9062,N_6347,N_7558);
xnor U9063 (N_9063,N_7307,N_6220);
nand U9064 (N_9064,N_8981,N_8812);
or U9065 (N_9065,N_7244,N_8136);
nand U9066 (N_9066,N_8630,N_6117);
nor U9067 (N_9067,N_7562,N_6399);
or U9068 (N_9068,N_7088,N_7003);
or U9069 (N_9069,N_8833,N_8906);
nor U9070 (N_9070,N_6088,N_6433);
nor U9071 (N_9071,N_6082,N_6014);
nand U9072 (N_9072,N_6730,N_6872);
nor U9073 (N_9073,N_7596,N_7778);
nand U9074 (N_9074,N_7705,N_8522);
or U9075 (N_9075,N_8364,N_7317);
xor U9076 (N_9076,N_7684,N_8639);
nor U9077 (N_9077,N_6944,N_8375);
nor U9078 (N_9078,N_8986,N_6013);
or U9079 (N_9079,N_8080,N_7702);
nor U9080 (N_9080,N_6908,N_6600);
and U9081 (N_9081,N_7527,N_6910);
nor U9082 (N_9082,N_7026,N_7791);
nor U9083 (N_9083,N_8313,N_6825);
nand U9084 (N_9084,N_8649,N_8892);
nor U9085 (N_9085,N_8118,N_7127);
nand U9086 (N_9086,N_7884,N_7730);
or U9087 (N_9087,N_7557,N_6444);
nor U9088 (N_9088,N_8942,N_6673);
or U9089 (N_9089,N_6477,N_6991);
and U9090 (N_9090,N_7683,N_8612);
nor U9091 (N_9091,N_6929,N_8360);
and U9092 (N_9092,N_6674,N_8785);
or U9093 (N_9093,N_6880,N_7966);
nor U9094 (N_9094,N_6605,N_7708);
or U9095 (N_9095,N_6536,N_7342);
and U9096 (N_9096,N_8316,N_6415);
and U9097 (N_9097,N_7017,N_6064);
and U9098 (N_9098,N_8090,N_7011);
nand U9099 (N_9099,N_7192,N_8175);
nand U9100 (N_9100,N_6371,N_8025);
or U9101 (N_9101,N_7788,N_6222);
nor U9102 (N_9102,N_6522,N_6104);
nor U9103 (N_9103,N_6207,N_7369);
nor U9104 (N_9104,N_8383,N_6624);
nor U9105 (N_9105,N_6296,N_8820);
or U9106 (N_9106,N_6967,N_8066);
and U9107 (N_9107,N_6826,N_6471);
nor U9108 (N_9108,N_7439,N_7874);
nor U9109 (N_9109,N_8259,N_6119);
or U9110 (N_9110,N_6312,N_7326);
xnor U9111 (N_9111,N_8211,N_7228);
nand U9112 (N_9112,N_7852,N_7279);
nand U9113 (N_9113,N_8151,N_8251);
and U9114 (N_9114,N_8733,N_8400);
or U9115 (N_9115,N_6360,N_6722);
nand U9116 (N_9116,N_7673,N_7651);
and U9117 (N_9117,N_7338,N_7247);
and U9118 (N_9118,N_6954,N_6553);
nor U9119 (N_9119,N_6166,N_7816);
nand U9120 (N_9120,N_7120,N_7010);
nand U9121 (N_9121,N_8356,N_7212);
or U9122 (N_9122,N_7496,N_8239);
or U9123 (N_9123,N_8964,N_7081);
or U9124 (N_9124,N_6282,N_8409);
nor U9125 (N_9125,N_8226,N_7767);
or U9126 (N_9126,N_8079,N_6968);
or U9127 (N_9127,N_7207,N_7187);
nand U9128 (N_9128,N_6003,N_8081);
nand U9129 (N_9129,N_7652,N_6241);
and U9130 (N_9130,N_7349,N_7196);
nor U9131 (N_9131,N_7610,N_7018);
or U9132 (N_9132,N_7225,N_7206);
or U9133 (N_9133,N_7209,N_6496);
nor U9134 (N_9134,N_6218,N_7887);
nor U9135 (N_9135,N_6210,N_7714);
xor U9136 (N_9136,N_6414,N_6974);
or U9137 (N_9137,N_6020,N_8880);
nor U9138 (N_9138,N_6180,N_8626);
and U9139 (N_9139,N_7448,N_8576);
xnor U9140 (N_9140,N_6294,N_7387);
and U9141 (N_9141,N_8474,N_8061);
or U9142 (N_9142,N_7182,N_8663);
or U9143 (N_9143,N_8143,N_6118);
and U9144 (N_9144,N_8886,N_8037);
nor U9145 (N_9145,N_7311,N_7715);
or U9146 (N_9146,N_7843,N_8811);
nand U9147 (N_9147,N_7735,N_6669);
xor U9148 (N_9148,N_7532,N_8575);
nand U9149 (N_9149,N_8742,N_7365);
nand U9150 (N_9150,N_8834,N_6592);
or U9151 (N_9151,N_8732,N_6171);
xnor U9152 (N_9152,N_6390,N_7722);
nor U9153 (N_9153,N_8193,N_6301);
or U9154 (N_9154,N_7539,N_8927);
or U9155 (N_9155,N_6325,N_8545);
nand U9156 (N_9156,N_6846,N_8538);
or U9157 (N_9157,N_7918,N_8008);
or U9158 (N_9158,N_8321,N_6632);
nor U9159 (N_9159,N_8229,N_6672);
xnor U9160 (N_9160,N_7129,N_7613);
or U9161 (N_9161,N_8623,N_6176);
or U9162 (N_9162,N_8172,N_6128);
nor U9163 (N_9163,N_7441,N_7998);
nor U9164 (N_9164,N_6755,N_8152);
and U9165 (N_9165,N_7477,N_7497);
xnor U9166 (N_9166,N_6870,N_7516);
nand U9167 (N_9167,N_8897,N_6563);
xor U9168 (N_9168,N_6330,N_6614);
and U9169 (N_9169,N_8507,N_8985);
nor U9170 (N_9170,N_7343,N_7175);
or U9171 (N_9171,N_7486,N_7056);
and U9172 (N_9172,N_6668,N_7748);
or U9173 (N_9173,N_8314,N_8987);
or U9174 (N_9174,N_8493,N_8913);
xnor U9175 (N_9175,N_8481,N_7725);
xnor U9176 (N_9176,N_8320,N_6456);
nand U9177 (N_9177,N_6594,N_6903);
or U9178 (N_9178,N_7992,N_6052);
or U9179 (N_9179,N_6250,N_6469);
nand U9180 (N_9180,N_7803,N_8371);
nand U9181 (N_9181,N_7085,N_6584);
or U9182 (N_9182,N_6894,N_8931);
or U9183 (N_9183,N_7920,N_7857);
nand U9184 (N_9184,N_7689,N_8134);
or U9185 (N_9185,N_6935,N_8971);
or U9186 (N_9186,N_6050,N_8595);
and U9187 (N_9187,N_8990,N_6113);
nand U9188 (N_9188,N_7181,N_8504);
and U9189 (N_9189,N_6208,N_8367);
nand U9190 (N_9190,N_6623,N_6815);
nor U9191 (N_9191,N_8145,N_7216);
and U9192 (N_9192,N_6646,N_7863);
and U9193 (N_9193,N_7197,N_8675);
nor U9194 (N_9194,N_8455,N_6086);
and U9195 (N_9195,N_8597,N_7541);
nor U9196 (N_9196,N_8216,N_7663);
and U9197 (N_9197,N_8022,N_6487);
nor U9198 (N_9198,N_8072,N_6251);
nand U9199 (N_9199,N_6108,N_8632);
and U9200 (N_9200,N_8670,N_8949);
nand U9201 (N_9201,N_7022,N_8298);
nand U9202 (N_9202,N_8074,N_7814);
and U9203 (N_9203,N_6998,N_7960);
or U9204 (N_9204,N_6655,N_7728);
nor U9205 (N_9205,N_7895,N_7798);
nor U9206 (N_9206,N_6689,N_6648);
and U9207 (N_9207,N_8108,N_8401);
nor U9208 (N_9208,N_6562,N_6112);
xnor U9209 (N_9209,N_8608,N_8713);
nor U9210 (N_9210,N_6643,N_6365);
xor U9211 (N_9211,N_6634,N_6694);
nand U9212 (N_9212,N_7480,N_6239);
xor U9213 (N_9213,N_7238,N_6859);
nand U9214 (N_9214,N_6856,N_8857);
nand U9215 (N_9215,N_7147,N_7520);
nand U9216 (N_9216,N_8621,N_7930);
nor U9217 (N_9217,N_8984,N_6083);
nand U9218 (N_9218,N_6626,N_6593);
or U9219 (N_9219,N_6551,N_8132);
and U9220 (N_9220,N_6742,N_6280);
nor U9221 (N_9221,N_8727,N_7912);
nor U9222 (N_9222,N_8315,N_7425);
or U9223 (N_9223,N_8104,N_6111);
and U9224 (N_9224,N_8633,N_6025);
or U9225 (N_9225,N_7716,N_8362);
nand U9226 (N_9226,N_7686,N_7283);
nand U9227 (N_9227,N_8106,N_6193);
and U9228 (N_9228,N_7602,N_7176);
and U9229 (N_9229,N_8789,N_7350);
or U9230 (N_9230,N_7633,N_7125);
nand U9231 (N_9231,N_6890,N_8484);
xnor U9232 (N_9232,N_7894,N_6383);
nor U9233 (N_9233,N_8323,N_7867);
and U9234 (N_9234,N_8438,N_8164);
nor U9235 (N_9235,N_8688,N_6028);
nand U9236 (N_9236,N_6687,N_7556);
nor U9237 (N_9237,N_7351,N_6568);
xor U9238 (N_9238,N_7935,N_8920);
xor U9239 (N_9239,N_6952,N_7959);
nor U9240 (N_9240,N_6402,N_8397);
and U9241 (N_9241,N_6152,N_8835);
and U9242 (N_9242,N_7380,N_6115);
or U9243 (N_9243,N_6934,N_6369);
or U9244 (N_9244,N_8405,N_6363);
or U9245 (N_9245,N_7063,N_8267);
or U9246 (N_9246,N_8404,N_8135);
nand U9247 (N_9247,N_8205,N_7759);
xor U9248 (N_9248,N_6726,N_8643);
or U9249 (N_9249,N_6212,N_6631);
xor U9250 (N_9250,N_7161,N_8542);
xor U9251 (N_9251,N_8710,N_8050);
or U9252 (N_9252,N_7726,N_8183);
or U9253 (N_9253,N_6746,N_6322);
nand U9254 (N_9254,N_8836,N_6247);
xnor U9255 (N_9255,N_7620,N_8559);
nor U9256 (N_9256,N_7094,N_8144);
xor U9257 (N_9257,N_8728,N_7679);
nand U9258 (N_9258,N_7939,N_7891);
xor U9259 (N_9259,N_8589,N_6573);
nor U9260 (N_9260,N_7103,N_6607);
xnor U9261 (N_9261,N_6127,N_6449);
nand U9262 (N_9262,N_6513,N_8345);
nor U9263 (N_9263,N_8754,N_7772);
nand U9264 (N_9264,N_6201,N_6610);
nor U9265 (N_9265,N_6472,N_8529);
nand U9266 (N_9266,N_6510,N_8411);
or U9267 (N_9267,N_6670,N_8204);
nand U9268 (N_9268,N_8432,N_8815);
or U9269 (N_9269,N_7653,N_7255);
or U9270 (N_9270,N_6440,N_8924);
or U9271 (N_9271,N_8454,N_6860);
and U9272 (N_9272,N_7347,N_7944);
nand U9273 (N_9273,N_8282,N_6413);
xnor U9274 (N_9274,N_8809,N_7348);
nand U9275 (N_9275,N_6447,N_7404);
nand U9276 (N_9276,N_6838,N_6574);
nor U9277 (N_9277,N_7148,N_7509);
nor U9278 (N_9278,N_7447,N_6649);
nand U9279 (N_9279,N_6179,N_8846);
nor U9280 (N_9280,N_8067,N_6340);
nand U9281 (N_9281,N_8552,N_8723);
nand U9282 (N_9282,N_6286,N_7254);
and U9283 (N_9283,N_7158,N_6063);
or U9284 (N_9284,N_6266,N_7925);
or U9285 (N_9285,N_7240,N_7336);
nand U9286 (N_9286,N_7752,N_8297);
and U9287 (N_9287,N_6979,N_7185);
nor U9288 (N_9288,N_7657,N_8300);
or U9289 (N_9289,N_7205,N_7799);
nand U9290 (N_9290,N_7450,N_8369);
xnor U9291 (N_9291,N_6540,N_6389);
nor U9292 (N_9292,N_7988,N_7099);
nand U9293 (N_9293,N_6891,N_7737);
xor U9294 (N_9294,N_8157,N_6348);
nand U9295 (N_9295,N_6804,N_7353);
and U9296 (N_9296,N_8035,N_8122);
or U9297 (N_9297,N_6992,N_7828);
and U9298 (N_9298,N_6039,N_6831);
xnor U9299 (N_9299,N_6552,N_8430);
or U9300 (N_9300,N_7849,N_7897);
nor U9301 (N_9301,N_8755,N_6711);
nand U9302 (N_9302,N_6803,N_8690);
nor U9303 (N_9303,N_8534,N_8165);
nor U9304 (N_9304,N_8693,N_7036);
nand U9305 (N_9305,N_6502,N_7286);
xor U9306 (N_9306,N_6256,N_6021);
nor U9307 (N_9307,N_8860,N_7972);
nand U9308 (N_9308,N_8709,N_7515);
or U9309 (N_9309,N_8977,N_8002);
or U9310 (N_9310,N_7294,N_6651);
nor U9311 (N_9311,N_8588,N_8995);
and U9312 (N_9312,N_8909,N_8309);
and U9313 (N_9313,N_7717,N_6221);
or U9314 (N_9314,N_7491,N_7669);
and U9315 (N_9315,N_8856,N_7007);
nand U9316 (N_9316,N_6942,N_7917);
nor U9317 (N_9317,N_8457,N_7789);
xnor U9318 (N_9318,N_7124,N_7068);
and U9319 (N_9319,N_7974,N_8392);
or U9320 (N_9320,N_6147,N_8291);
nor U9321 (N_9321,N_6524,N_8653);
or U9322 (N_9322,N_6625,N_6227);
nor U9323 (N_9323,N_6566,N_7523);
nor U9324 (N_9324,N_7522,N_7694);
nand U9325 (N_9325,N_8989,N_8547);
nand U9326 (N_9326,N_6008,N_6145);
nor U9327 (N_9327,N_8398,N_6955);
nor U9328 (N_9328,N_8441,N_6802);
xor U9329 (N_9329,N_7779,N_8168);
nor U9330 (N_9330,N_7070,N_7979);
nor U9331 (N_9331,N_7401,N_8791);
or U9332 (N_9332,N_8933,N_8792);
nand U9333 (N_9333,N_6421,N_6044);
xnor U9334 (N_9334,N_8661,N_7832);
nor U9335 (N_9335,N_7528,N_6267);
and U9336 (N_9336,N_6791,N_7329);
and U9337 (N_9337,N_6662,N_6367);
or U9338 (N_9338,N_6609,N_6769);
nor U9339 (N_9339,N_8156,N_6011);
or U9340 (N_9340,N_7659,N_7553);
xnor U9341 (N_9341,N_8444,N_8744);
nand U9342 (N_9342,N_7418,N_7634);
or U9343 (N_9343,N_7640,N_8794);
nand U9344 (N_9344,N_6597,N_7322);
and U9345 (N_9345,N_7400,N_6426);
or U9346 (N_9346,N_7984,N_7868);
nand U9347 (N_9347,N_7215,N_6437);
nor U9348 (N_9348,N_7731,N_6724);
xor U9349 (N_9349,N_6130,N_7589);
or U9350 (N_9350,N_8182,N_7015);
nand U9351 (N_9351,N_6906,N_7519);
nor U9352 (N_9352,N_6985,N_8396);
nor U9353 (N_9353,N_8296,N_6938);
nor U9354 (N_9354,N_7882,N_8112);
nand U9355 (N_9355,N_7275,N_8519);
or U9356 (N_9356,N_7630,N_6777);
nand U9357 (N_9357,N_8098,N_7821);
nand U9358 (N_9358,N_6110,N_6637);
nor U9359 (N_9359,N_8213,N_6315);
and U9360 (N_9360,N_7855,N_6589);
nand U9361 (N_9361,N_8940,N_8569);
and U9362 (N_9362,N_7628,N_6292);
and U9363 (N_9363,N_8530,N_8553);
or U9364 (N_9364,N_8466,N_8221);
nor U9365 (N_9365,N_7755,N_8206);
nor U9366 (N_9366,N_6381,N_8852);
and U9367 (N_9367,N_8718,N_6124);
xor U9368 (N_9368,N_8459,N_8359);
nor U9369 (N_9369,N_8303,N_8353);
nand U9370 (N_9370,N_6022,N_8272);
and U9371 (N_9371,N_8434,N_8721);
or U9372 (N_9372,N_7381,N_8795);
nor U9373 (N_9373,N_6969,N_6768);
and U9374 (N_9374,N_7318,N_6029);
and U9375 (N_9375,N_8853,N_7529);
nand U9376 (N_9376,N_8439,N_7262);
nor U9377 (N_9377,N_7222,N_6745);
and U9378 (N_9378,N_7211,N_7325);
and U9379 (N_9379,N_8844,N_7954);
or U9380 (N_9380,N_8919,N_8573);
or U9381 (N_9381,N_7267,N_8338);
nand U9382 (N_9382,N_8113,N_8972);
xnor U9383 (N_9383,N_8230,N_7438);
nor U9384 (N_9384,N_6065,N_8572);
or U9385 (N_9385,N_6773,N_8053);
and U9386 (N_9386,N_6936,N_7965);
nor U9387 (N_9387,N_6590,N_6658);
xnor U9388 (N_9388,N_6284,N_7858);
nand U9389 (N_9389,N_6930,N_7670);
nor U9390 (N_9390,N_6408,N_6972);
xnor U9391 (N_9391,N_7793,N_6343);
nand U9392 (N_9392,N_7727,N_7290);
xor U9393 (N_9393,N_6149,N_7665);
nor U9394 (N_9394,N_7047,N_6904);
and U9395 (N_9395,N_6059,N_6303);
xor U9396 (N_9396,N_8443,N_7810);
and U9397 (N_9397,N_8288,N_8306);
nor U9398 (N_9398,N_6706,N_8277);
or U9399 (N_9399,N_8190,N_7574);
or U9400 (N_9400,N_7004,N_6578);
or U9401 (N_9401,N_7546,N_8918);
or U9402 (N_9402,N_8257,N_6475);
or U9403 (N_9403,N_7055,N_6228);
or U9404 (N_9404,N_7943,N_6754);
nand U9405 (N_9405,N_6956,N_6692);
or U9406 (N_9406,N_7741,N_8528);
and U9407 (N_9407,N_7335,N_6454);
nand U9408 (N_9408,N_6547,N_7449);
nor U9409 (N_9409,N_8505,N_6764);
and U9410 (N_9410,N_6009,N_6479);
and U9411 (N_9411,N_6231,N_6883);
nand U9412 (N_9412,N_7846,N_7534);
nor U9413 (N_9413,N_8117,N_7345);
nor U9414 (N_9414,N_6630,N_6380);
or U9415 (N_9415,N_7252,N_6283);
and U9416 (N_9416,N_6265,N_8100);
or U9417 (N_9417,N_7388,N_7896);
and U9418 (N_9418,N_8776,N_7700);
or U9419 (N_9419,N_7355,N_7698);
nor U9420 (N_9420,N_7417,N_8818);
or U9421 (N_9421,N_6154,N_8352);
nand U9422 (N_9422,N_7560,N_6306);
nor U9423 (N_9423,N_7406,N_8268);
nand U9424 (N_9424,N_6081,N_8593);
nand U9425 (N_9425,N_7079,N_7879);
xnor U9426 (N_9426,N_8249,N_8305);
or U9427 (N_9427,N_6721,N_8446);
and U9428 (N_9428,N_7889,N_8677);
nand U9429 (N_9429,N_7565,N_7552);
and U9430 (N_9430,N_6144,N_8148);
or U9431 (N_9431,N_8415,N_6480);
or U9432 (N_9432,N_6539,N_8581);
or U9433 (N_9433,N_8908,N_7189);
or U9434 (N_9434,N_6734,N_8683);
or U9435 (N_9435,N_8520,N_8837);
nand U9436 (N_9436,N_7809,N_6506);
nand U9437 (N_9437,N_6258,N_6780);
or U9438 (N_9438,N_8021,N_6527);
nand U9439 (N_9439,N_6202,N_6173);
nor U9440 (N_9440,N_7744,N_6917);
and U9441 (N_9441,N_7263,N_7921);
or U9442 (N_9442,N_8917,N_8563);
and U9443 (N_9443,N_6928,N_8662);
or U9444 (N_9444,N_8408,N_7834);
or U9445 (N_9445,N_7680,N_6765);
and U9446 (N_9446,N_8094,N_7397);
or U9447 (N_9447,N_8043,N_8322);
and U9448 (N_9448,N_6782,N_8379);
nand U9449 (N_9449,N_8800,N_7976);
and U9450 (N_9450,N_8627,N_7871);
nor U9451 (N_9451,N_7819,N_8475);
or U9452 (N_9452,N_6786,N_8819);
or U9453 (N_9453,N_7764,N_8914);
or U9454 (N_9454,N_6854,N_8109);
nor U9455 (N_9455,N_7945,N_6277);
and U9456 (N_9456,N_6901,N_7152);
nor U9457 (N_9457,N_7374,N_7547);
or U9458 (N_9458,N_8708,N_7822);
nor U9459 (N_9459,N_6778,N_7877);
or U9460 (N_9460,N_7373,N_8807);
nand U9461 (N_9461,N_7854,N_7636);
nor U9462 (N_9462,N_7902,N_7616);
nand U9463 (N_9463,N_7352,N_6983);
or U9464 (N_9464,N_8731,N_6733);
nor U9465 (N_9465,N_7501,N_7464);
nand U9466 (N_9466,N_8026,N_7375);
nor U9467 (N_9467,N_7853,N_8361);
and U9468 (N_9468,N_8937,N_6183);
and U9469 (N_9469,N_6404,N_6159);
nor U9470 (N_9470,N_8802,N_7469);
nand U9471 (N_9471,N_8966,N_8453);
and U9472 (N_9472,N_8712,N_6523);
nand U9473 (N_9473,N_8565,N_8616);
nor U9474 (N_9474,N_7316,N_7763);
nor U9475 (N_9475,N_8804,N_6571);
nand U9476 (N_9476,N_6185,N_7399);
and U9477 (N_9477,N_6123,N_7130);
nand U9478 (N_9478,N_6187,N_8052);
nor U9479 (N_9479,N_7622,N_7376);
nor U9480 (N_9480,N_6581,N_7223);
nand U9481 (N_9481,N_6428,N_6680);
and U9482 (N_9482,N_8749,N_6849);
or U9483 (N_9483,N_7746,N_6165);
and U9484 (N_9484,N_7037,N_7339);
and U9485 (N_9485,N_8884,N_8953);
or U9486 (N_9486,N_8236,N_6761);
nor U9487 (N_9487,N_8746,N_7947);
xnor U9488 (N_9488,N_8289,N_7555);
and U9489 (N_9489,N_8228,N_6355);
nand U9490 (N_9490,N_7572,N_8851);
and U9491 (N_9491,N_8261,N_7297);
nand U9492 (N_9492,N_6896,N_7384);
nand U9493 (N_9493,N_7985,N_6155);
and U9494 (N_9494,N_8063,N_7140);
and U9495 (N_9495,N_7493,N_7199);
or U9496 (N_9496,N_6871,N_8491);
nor U9497 (N_9497,N_7467,N_6401);
and U9498 (N_9498,N_8978,N_7485);
nor U9499 (N_9499,N_8996,N_7364);
nand U9500 (N_9500,N_7549,N_8730);
and U9501 (N_9501,N_6806,N_6823);
or U9502 (N_9502,N_7430,N_8264);
or U9503 (N_9503,N_8770,N_7824);
and U9504 (N_9504,N_7289,N_8604);
and U9505 (N_9505,N_7259,N_8059);
nand U9506 (N_9506,N_6394,N_7051);
or U9507 (N_9507,N_8017,N_8904);
nand U9508 (N_9508,N_8872,N_6652);
or U9509 (N_9509,N_6771,N_8780);
nor U9510 (N_9510,N_8704,N_8412);
nor U9511 (N_9511,N_7790,N_8901);
and U9512 (N_9512,N_7386,N_6981);
or U9513 (N_9513,N_7039,N_8467);
nor U9514 (N_9514,N_6750,N_6398);
xnor U9515 (N_9515,N_8018,N_7359);
or U9516 (N_9516,N_7331,N_8970);
and U9517 (N_9517,N_6462,N_7975);
or U9518 (N_9518,N_7993,N_8011);
nand U9519 (N_9519,N_6912,N_7413);
nand U9520 (N_9520,N_6078,N_8231);
or U9521 (N_9521,N_7787,N_8005);
or U9522 (N_9522,N_7682,N_8195);
or U9523 (N_9523,N_7455,N_8429);
or U9524 (N_9524,N_8636,N_6388);
xnor U9525 (N_9525,N_8372,N_7113);
nand U9526 (N_9526,N_8512,N_7458);
and U9527 (N_9527,N_7110,N_8447);
and U9528 (N_9528,N_7710,N_7378);
and U9529 (N_9529,N_8994,N_7724);
or U9530 (N_9530,N_7554,N_7649);
nand U9531 (N_9531,N_6068,N_6298);
nor U9532 (N_9532,N_8155,N_8170);
nor U9533 (N_9533,N_8934,N_7642);
nor U9534 (N_9534,N_6217,N_7507);
nor U9535 (N_9535,N_8969,N_7531);
or U9536 (N_9536,N_8496,N_7606);
or U9537 (N_9537,N_6817,N_6837);
nand U9538 (N_9538,N_8262,N_7027);
nor U9539 (N_9539,N_7414,N_7083);
or U9540 (N_9540,N_8344,N_7321);
nand U9541 (N_9541,N_8130,N_6580);
and U9542 (N_9542,N_7118,N_8847);
nand U9543 (N_9543,N_6374,N_7862);
and U9544 (N_9544,N_8480,N_8406);
nand U9545 (N_9545,N_7478,N_6727);
or U9546 (N_9546,N_6720,N_8854);
nand U9547 (N_9547,N_6372,N_7237);
or U9548 (N_9548,N_8606,N_7666);
or U9549 (N_9549,N_6425,N_7548);
or U9550 (N_9550,N_6191,N_7733);
nand U9551 (N_9551,N_8982,N_6946);
or U9552 (N_9552,N_8062,N_7431);
or U9553 (N_9553,N_6342,N_8896);
nand U9554 (N_9554,N_7214,N_8773);
and U9555 (N_9555,N_6478,N_6335);
or U9556 (N_9556,N_7170,N_8237);
or U9557 (N_9557,N_6719,N_6010);
nor U9558 (N_9558,N_6881,N_6172);
nand U9559 (N_9559,N_8388,N_7002);
and U9560 (N_9560,N_8357,N_7905);
nand U9561 (N_9561,N_6121,N_6075);
or U9562 (N_9562,N_6424,N_8285);
xnor U9563 (N_9563,N_7500,N_7899);
or U9564 (N_9564,N_6816,N_8787);
or U9565 (N_9565,N_8330,N_7179);
or U9566 (N_9566,N_7440,N_6723);
and U9567 (N_9567,N_6705,N_7208);
nor U9568 (N_9568,N_8308,N_8925);
or U9569 (N_9569,N_7220,N_8500);
or U9570 (N_9570,N_6302,N_8568);
nor U9571 (N_9571,N_6798,N_8105);
nor U9572 (N_9572,N_6924,N_6461);
nand U9573 (N_9573,N_6840,N_6189);
or U9574 (N_9574,N_6120,N_8290);
xor U9575 (N_9575,N_8110,N_8596);
or U9576 (N_9576,N_8139,N_8567);
nor U9577 (N_9577,N_7804,N_6148);
and U9578 (N_9578,N_7258,N_6975);
or U9579 (N_9579,N_7136,N_7720);
and U9580 (N_9580,N_6074,N_7860);
and U9581 (N_9581,N_6834,N_8238);
nand U9582 (N_9582,N_6876,N_6358);
or U9583 (N_9583,N_8784,N_6067);
nor U9584 (N_9584,N_8351,N_8952);
xor U9585 (N_9585,N_6060,N_7122);
nor U9586 (N_9586,N_7568,N_6957);
nor U9587 (N_9587,N_6184,N_7062);
nor U9588 (N_9588,N_8463,N_6026);
nor U9589 (N_9589,N_7719,N_7241);
nand U9590 (N_9590,N_6162,N_6178);
nor U9591 (N_9591,N_7607,N_6485);
or U9592 (N_9592,N_8209,N_7437);
xor U9593 (N_9593,N_8647,N_7692);
nor U9594 (N_9594,N_8778,N_8796);
and U9595 (N_9595,N_8701,N_6707);
xor U9596 (N_9596,N_6055,N_8826);
and U9597 (N_9597,N_6511,N_8049);
nand U9598 (N_9598,N_6084,N_6457);
or U9599 (N_9599,N_6695,N_6040);
or U9600 (N_9600,N_7598,N_7487);
nor U9601 (N_9601,N_7505,N_6601);
nand U9602 (N_9602,N_6560,N_7138);
or U9603 (N_9603,N_8210,N_7341);
nor U9604 (N_9604,N_7233,N_6268);
nor U9605 (N_9605,N_7457,N_6776);
nor U9606 (N_9606,N_7382,N_8325);
xor U9607 (N_9607,N_8509,N_7550);
and U9608 (N_9608,N_7770,N_8585);
nor U9609 (N_9609,N_7981,N_7173);
nand U9610 (N_9610,N_7032,N_7451);
nor U9611 (N_9611,N_6422,N_8876);
nand U9612 (N_9612,N_7713,N_6855);
or U9613 (N_9613,N_8115,N_6261);
nand U9614 (N_9614,N_7693,N_7075);
and U9615 (N_9615,N_7490,N_6257);
nor U9616 (N_9616,N_8564,N_8085);
or U9617 (N_9617,N_7699,N_8214);
or U9618 (N_9618,N_8980,N_7315);
or U9619 (N_9619,N_8417,N_6346);
or U9620 (N_9620,N_6644,N_8863);
nand U9621 (N_9621,N_6445,N_7583);
nor U9622 (N_9622,N_8032,N_6557);
and U9623 (N_9623,N_7096,N_7842);
nor U9624 (N_9624,N_8497,N_6681);
and U9625 (N_9625,N_8384,N_8460);
or U9626 (N_9626,N_8867,N_6314);
or U9627 (N_9627,N_8657,N_8410);
nor U9628 (N_9628,N_7775,N_8560);
nand U9629 (N_9629,N_8768,N_6384);
xnor U9630 (N_9630,N_8674,N_6588);
and U9631 (N_9631,N_6240,N_6464);
nor U9632 (N_9632,N_6213,N_8137);
and U9633 (N_9633,N_6710,N_6490);
xor U9634 (N_9634,N_8327,N_8341);
and U9635 (N_9635,N_7656,N_7569);
and U9636 (N_9636,N_8879,N_6103);
or U9637 (N_9637,N_6435,N_8997);
nor U9638 (N_9638,N_6933,N_7543);
nand U9639 (N_9639,N_6168,N_7685);
nand U9640 (N_9640,N_7517,N_6535);
and U9641 (N_9641,N_8407,N_8620);
nand U9642 (N_9642,N_6679,N_6085);
nand U9643 (N_9643,N_8012,N_8855);
nand U9644 (N_9644,N_8788,N_6125);
xnor U9645 (N_9645,N_8328,N_6715);
or U9646 (N_9646,N_7119,N_6285);
or U9647 (N_9647,N_6945,N_7276);
and U9648 (N_9648,N_6843,N_6555);
nor U9649 (N_9649,N_8946,N_6886);
nand U9650 (N_9650,N_7098,N_6518);
nor U9651 (N_9651,N_7866,N_8207);
or U9652 (N_9652,N_8006,N_7436);
or U9653 (N_9653,N_6309,N_6970);
and U9654 (N_9654,N_7908,N_6001);
nor U9655 (N_9655,N_6885,N_8199);
nand U9656 (N_9656,N_7890,N_6829);
nor U9657 (N_9657,N_7328,N_8034);
and U9658 (N_9658,N_6543,N_7116);
nor U9659 (N_9659,N_6129,N_8234);
or U9660 (N_9660,N_8571,N_6199);
xnor U9661 (N_9661,N_7495,N_6332);
or U9662 (N_9662,N_8471,N_8227);
nor U9663 (N_9663,N_8087,N_8686);
nand U9664 (N_9664,N_8699,N_8260);
xnor U9665 (N_9665,N_6749,N_7463);
nor U9666 (N_9666,N_6153,N_8698);
nor U9667 (N_9667,N_6450,N_8584);
and U9668 (N_9668,N_8324,N_8965);
and U9669 (N_9669,N_8885,N_6950);
nand U9670 (N_9670,N_8993,N_8889);
nand U9671 (N_9671,N_8051,N_7107);
and U9672 (N_9672,N_8842,N_6140);
nor U9673 (N_9673,N_7780,N_7601);
nor U9674 (N_9674,N_8869,N_7971);
or U9675 (N_9675,N_6532,N_7260);
or U9676 (N_9676,N_8158,N_6851);
or U9677 (N_9677,N_6019,N_6216);
nand U9678 (N_9678,N_7644,N_8629);
xor U9679 (N_9679,N_7551,N_6832);
nor U9680 (N_9680,N_8511,N_8935);
and U9681 (N_9681,N_7864,N_6913);
and U9682 (N_9682,N_6598,N_6385);
and U9683 (N_9683,N_6416,N_6441);
nor U9684 (N_9684,N_7014,N_6156);
nand U9685 (N_9685,N_7291,N_7978);
or U9686 (N_9686,N_6747,N_7732);
nand U9687 (N_9687,N_7844,N_7023);
nor U9688 (N_9688,N_8114,N_7080);
or U9689 (N_9689,N_6549,N_7266);
nand U9690 (N_9690,N_7219,N_6544);
nand U9691 (N_9691,N_7900,N_7149);
and U9692 (N_9692,N_8941,N_6807);
xnor U9693 (N_9693,N_7801,N_7403);
and U9694 (N_9694,N_8814,N_6693);
nand U9695 (N_9695,N_7180,N_6494);
or U9696 (N_9696,N_7021,N_8923);
or U9697 (N_9697,N_8001,N_6182);
and U9698 (N_9698,N_6708,N_8271);
or U9699 (N_9699,N_7020,N_6486);
and U9700 (N_9700,N_8808,N_6038);
nand U9701 (N_9701,N_7061,N_6386);
nand U9702 (N_9702,N_8829,N_7545);
nand U9703 (N_9703,N_6034,N_8273);
and U9704 (N_9704,N_8561,N_7671);
nor U9705 (N_9705,N_7786,N_8577);
nand U9706 (N_9706,N_7906,N_8968);
nand U9707 (N_9707,N_7766,N_7655);
nand U9708 (N_9708,N_8777,N_6575);
or U9709 (N_9709,N_6654,N_8579);
or U9710 (N_9710,N_8930,N_7242);
nor U9711 (N_9711,N_7200,N_8929);
nor U9712 (N_9712,N_7295,N_6525);
and U9713 (N_9713,N_7870,N_8166);
nor U9714 (N_9714,N_6107,N_7327);
nand U9715 (N_9715,N_8583,N_7980);
nor U9716 (N_9716,N_8945,N_7177);
nor U9717 (N_9717,N_7035,N_6516);
nor U9718 (N_9718,N_8461,N_6900);
nand U9719 (N_9719,N_6203,N_6259);
nand U9720 (N_9720,N_7218,N_6146);
or U9721 (N_9721,N_6281,N_7285);
or U9722 (N_9722,N_7624,N_7028);
xnor U9723 (N_9723,N_6501,N_6387);
and U9724 (N_9724,N_8449,N_8082);
xor U9725 (N_9725,N_7104,N_7594);
nand U9726 (N_9726,N_6550,N_8350);
or U9727 (N_9727,N_6509,N_7544);
nor U9728 (N_9728,N_6275,N_7802);
and U9729 (N_9729,N_7604,N_8926);
and U9730 (N_9730,N_8269,N_7082);
nand U9731 (N_9731,N_8526,N_6219);
and U9732 (N_9732,N_6205,N_6775);
and U9733 (N_9733,N_8592,N_6043);
nand U9734 (N_9734,N_7030,N_6599);
nor U9735 (N_9735,N_7184,N_8963);
xor U9736 (N_9736,N_8436,N_6994);
nor U9737 (N_9737,N_8533,N_6729);
xor U9738 (N_9738,N_8655,N_8707);
nand U9739 (N_9739,N_8672,N_8890);
xnor U9740 (N_9740,N_6801,N_6864);
xnor U9741 (N_9741,N_6812,N_6683);
xnor U9742 (N_9742,N_8380,N_8423);
nand U9743 (N_9743,N_6430,N_6396);
and U9744 (N_9744,N_6045,N_8735);
or U9745 (N_9745,N_7421,N_6379);
nor U9746 (N_9746,N_8724,N_7314);
nand U9747 (N_9747,N_7191,N_8562);
nand U9748 (N_9748,N_8223,N_8241);
nor U9749 (N_9749,N_6737,N_8456);
and U9750 (N_9750,N_8295,N_7818);
or U9751 (N_9751,N_7888,N_7797);
nand U9752 (N_9752,N_7836,N_8091);
nand U9753 (N_9753,N_7639,N_7703);
or U9754 (N_9754,N_8343,N_7579);
nor U9755 (N_9755,N_7114,N_8821);
nand U9756 (N_9756,N_7052,N_6211);
nor U9757 (N_9757,N_6287,N_8745);
nor U9758 (N_9758,N_6080,N_8126);
or U9759 (N_9759,N_7193,N_6743);
or U9760 (N_9760,N_8376,N_7695);
and U9761 (N_9761,N_7615,N_6465);
or U9762 (N_9762,N_8402,N_7337);
or U9763 (N_9763,N_8046,N_6640);
xnor U9764 (N_9764,N_8816,N_8270);
nor U9765 (N_9765,N_6079,N_7243);
and U9766 (N_9766,N_8607,N_6419);
or U9767 (N_9767,N_8582,N_6554);
nor U9768 (N_9768,N_8342,N_6666);
or U9769 (N_9769,N_6731,N_7646);
nand U9770 (N_9770,N_8525,N_6352);
nand U9771 (N_9771,N_8898,N_8775);
nand U9772 (N_9772,N_7812,N_7932);
nor U9773 (N_9773,N_8883,N_7511);
and U9774 (N_9774,N_7091,N_8557);
nand U9775 (N_9775,N_6628,N_7995);
nand U9776 (N_9776,N_6645,N_6090);
and U9777 (N_9777,N_8753,N_8611);
and U9778 (N_9778,N_7648,N_6126);
xnor U9779 (N_9779,N_6307,N_8452);
and U9780 (N_9780,N_6783,N_8121);
nand U9781 (N_9781,N_7629,N_8888);
nor U9782 (N_9782,N_8830,N_7643);
nor U9783 (N_9783,N_6446,N_8275);
nand U9784 (N_9784,N_7234,N_8358);
nor U9785 (N_9785,N_6997,N_7881);
or U9786 (N_9786,N_8813,N_6617);
nor U9787 (N_9787,N_8244,N_6098);
xnor U9788 (N_9788,N_8403,N_8658);
nor U9789 (N_9789,N_8133,N_8640);
or U9790 (N_9790,N_7174,N_6135);
xor U9791 (N_9791,N_6253,N_8541);
nor U9792 (N_9792,N_6263,N_8385);
xnor U9793 (N_9793,N_7603,N_7142);
xor U9794 (N_9794,N_6236,N_6685);
nand U9795 (N_9795,N_7001,N_6561);
or U9796 (N_9796,N_7827,N_8233);
nand U9797 (N_9797,N_6299,N_6223);
nand U9798 (N_9798,N_8422,N_8973);
nor U9799 (N_9799,N_7293,N_6844);
xor U9800 (N_9800,N_7996,N_6295);
nand U9801 (N_9801,N_7696,N_6888);
xor U9802 (N_9802,N_8609,N_6861);
and U9803 (N_9803,N_8279,N_7672);
nor U9804 (N_9804,N_7753,N_8428);
nand U9805 (N_9805,N_8740,N_7090);
nand U9806 (N_9806,N_7751,N_6473);
or U9807 (N_9807,N_6741,N_8469);
nand U9808 (N_9808,N_7296,N_8060);
and U9809 (N_9809,N_6538,N_7272);
nor U9810 (N_9810,N_7600,N_7235);
or U9811 (N_9811,N_8549,N_6684);
nor U9812 (N_9812,N_6072,N_6922);
and U9813 (N_9813,N_6862,N_8651);
or U9814 (N_9814,N_6006,N_8181);
xor U9815 (N_9815,N_8377,N_7904);
nand U9816 (N_9816,N_6254,N_6865);
nand U9817 (N_9817,N_7278,N_7134);
nand U9818 (N_9818,N_8550,N_6940);
and U9819 (N_9819,N_6897,N_7911);
or U9820 (N_9820,N_8286,N_8660);
and U9821 (N_9821,N_6377,N_8786);
or U9822 (N_9822,N_6827,N_7280);
xnor U9823 (N_9823,N_8603,N_7588);
or U9824 (N_9824,N_6905,N_7195);
or U9825 (N_9825,N_7422,N_6558);
xnor U9826 (N_9826,N_8347,N_7424);
and U9827 (N_9827,N_7169,N_7587);
and U9828 (N_9828,N_7577,N_7277);
nand U9829 (N_9829,N_6873,N_8769);
or U9830 (N_9830,N_8858,N_6805);
and U9831 (N_9831,N_6845,N_8326);
xor U9832 (N_9832,N_7584,N_8910);
nor U9833 (N_9833,N_8645,N_8058);
or U9834 (N_9834,N_8705,N_8492);
and U9835 (N_9835,N_6937,N_8427);
and U9836 (N_9836,N_7883,N_7371);
nand U9837 (N_9837,N_6238,N_6272);
or U9838 (N_9838,N_7483,N_7955);
nand U9839 (N_9839,N_6368,N_7590);
nor U9840 (N_9840,N_6839,N_8679);
nand U9841 (N_9841,N_6418,N_8695);
and U9842 (N_9842,N_8605,N_7303);
nor U9843 (N_9843,N_7711,N_8319);
nand U9844 (N_9844,N_8840,N_7361);
or U9845 (N_9845,N_8697,N_8479);
nand U9846 (N_9846,N_7249,N_7390);
nand U9847 (N_9847,N_6887,N_6869);
or U9848 (N_9848,N_8865,N_6740);
or U9849 (N_9849,N_7078,N_8691);
xnor U9850 (N_9850,N_8414,N_6448);
xnor U9851 (N_9851,N_7474,N_7922);
and U9852 (N_9852,N_8766,N_6691);
nand U9853 (N_9853,N_6493,N_7396);
nand U9854 (N_9854,N_8225,N_6818);
nand U9855 (N_9855,N_8922,N_8154);
or U9856 (N_9856,N_6252,N_6925);
nand U9857 (N_9857,N_7627,N_8532);
or U9858 (N_9858,N_6546,N_6042);
xor U9859 (N_9859,N_8668,N_6249);
nand U9860 (N_9860,N_8825,N_6797);
and U9861 (N_9861,N_8450,N_6565);
or U9862 (N_9862,N_8998,N_8988);
nand U9863 (N_9863,N_6977,N_6116);
and U9864 (N_9864,N_7203,N_8128);
nor U9865 (N_9865,N_7563,N_8395);
xnor U9866 (N_9866,N_7054,N_7982);
or U9867 (N_9867,N_7907,N_6569);
nand U9868 (N_9868,N_7566,N_7006);
or U9869 (N_9869,N_6023,N_7823);
or U9870 (N_9870,N_7518,N_7538);
and U9871 (N_9871,N_6293,N_6432);
or U9872 (N_9872,N_8413,N_7647);
nand U9873 (N_9873,N_7952,N_6770);
or U9874 (N_9874,N_8458,N_8235);
and U9875 (N_9875,N_6996,N_6066);
nor U9876 (N_9876,N_8488,N_6353);
nor U9877 (N_9877,N_6143,N_6093);
nand U9878 (N_9878,N_8041,N_6759);
xor U9879 (N_9879,N_8646,N_7513);
nor U9880 (N_9880,N_6406,N_8348);
nor U9881 (N_9881,N_6200,N_8332);
nor U9882 (N_9882,N_6393,N_7132);
or U9883 (N_9883,N_6429,N_8084);
or U9884 (N_9884,N_7878,N_6138);
and U9885 (N_9885,N_8881,N_8150);
and U9886 (N_9886,N_6586,N_7928);
or U9887 (N_9887,N_8031,N_6463);
and U9888 (N_9888,N_8514,N_6427);
and U9889 (N_9889,N_7060,N_6987);
nor U9890 (N_9890,N_8044,N_6460);
or U9891 (N_9891,N_7826,N_6712);
nor U9892 (N_9892,N_7997,N_6304);
and U9893 (N_9893,N_6622,N_8900);
and U9894 (N_9894,N_6545,N_7926);
and U9895 (N_9895,N_8748,N_6736);
and U9896 (N_9896,N_6504,N_7739);
and U9897 (N_9897,N_6874,N_6245);
and U9898 (N_9898,N_7412,N_8517);
nand U9899 (N_9899,N_6273,N_6382);
and U9900 (N_9900,N_7991,N_6169);
and U9901 (N_9901,N_8464,N_6452);
or U9902 (N_9902,N_8702,N_6647);
nand U9903 (N_9903,N_7383,N_8020);
xor U9904 (N_9904,N_7757,N_8979);
and U9905 (N_9905,N_8793,N_7137);
nand U9906 (N_9906,N_6246,N_7968);
nand U9907 (N_9907,N_7363,N_8722);
and U9908 (N_9908,N_6373,N_7178);
nor U9909 (N_9909,N_7740,N_7476);
or U9910 (N_9910,N_7334,N_7101);
and U9911 (N_9911,N_7442,N_6122);
and U9912 (N_9912,N_6319,N_7210);
nand U9913 (N_9913,N_6868,N_7167);
or U9914 (N_9914,N_6051,N_6015);
nand U9915 (N_9915,N_6787,N_7631);
nor U9916 (N_9916,N_7662,N_8714);
or U9917 (N_9917,N_6007,N_6999);
and U9918 (N_9918,N_8038,N_7619);
nor U9919 (N_9919,N_8760,N_6030);
or U9920 (N_9920,N_8681,N_6262);
nor U9921 (N_9921,N_6682,N_8329);
or U9922 (N_9922,N_8266,N_8916);
or U9923 (N_9923,N_8127,N_7154);
and U9924 (N_9924,N_8200,N_8667);
and U9925 (N_9925,N_7284,N_8280);
nand U9926 (N_9926,N_8246,N_6233);
nor U9927 (N_9927,N_8911,N_8893);
nand U9928 (N_9928,N_6134,N_8201);
or U9929 (N_9929,N_8167,N_8907);
or U9930 (N_9930,N_7248,N_7084);
and U9931 (N_9931,N_7813,N_7468);
and U9932 (N_9932,N_6615,N_8363);
or U9933 (N_9933,N_6037,N_8097);
nand U9934 (N_9934,N_6359,N_7432);
and U9935 (N_9935,N_6850,N_6579);
nor U9936 (N_9936,N_8539,N_7164);
or U9937 (N_9937,N_6559,N_6106);
or U9938 (N_9938,N_6320,N_7264);
or U9939 (N_9939,N_6830,N_8255);
and U9940 (N_9940,N_6809,N_7446);
nand U9941 (N_9941,N_6376,N_8111);
or U9942 (N_9942,N_6713,N_6902);
xnor U9943 (N_9943,N_8614,N_8253);
nand U9944 (N_9944,N_8684,N_8659);
nand U9945 (N_9945,N_6931,N_7183);
and U9946 (N_9946,N_8554,N_8921);
or U9947 (N_9947,N_8310,N_8381);
or U9948 (N_9948,N_7367,N_8064);
nor U9949 (N_9949,N_8171,N_8191);
or U9950 (N_9950,N_6650,N_6519);
or U9951 (N_9951,N_8426,N_6828);
or U9952 (N_9952,N_8102,N_6800);
nand U9953 (N_9953,N_7141,N_6327);
and U9954 (N_9954,N_8146,N_8445);
and U9955 (N_9955,N_7416,N_8197);
or U9956 (N_9956,N_7903,N_7479);
and U9957 (N_9957,N_7990,N_6529);
and U9958 (N_9958,N_6163,N_8502);
or U9959 (N_9959,N_6316,N_6431);
nand U9960 (N_9960,N_7658,N_7934);
nor U9961 (N_9961,N_7190,N_7144);
nand U9962 (N_9962,N_8706,N_7592);
nand U9963 (N_9963,N_7667,N_6069);
nor U9964 (N_9964,N_7226,N_6500);
and U9965 (N_9965,N_6161,N_8265);
and U9966 (N_9966,N_8418,N_7298);
nor U9967 (N_9967,N_7924,N_7963);
and U9968 (N_9968,N_6058,N_8700);
or U9969 (N_9969,N_7394,N_8240);
nor U9970 (N_9970,N_6244,N_7095);
nand U9971 (N_9971,N_6167,N_8368);
or U9972 (N_9972,N_7795,N_6339);
nor U9973 (N_9973,N_8510,N_7426);
nand U9974 (N_9974,N_8421,N_7815);
or U9975 (N_9975,N_7213,N_7330);
or U9976 (N_9976,N_8186,N_7768);
nor U9977 (N_9977,N_6671,N_6753);
or U9978 (N_9978,N_6714,N_7931);
nand U9979 (N_9979,N_6451,N_7150);
or U9980 (N_9980,N_8912,N_8024);
xnor U9981 (N_9981,N_7163,N_7808);
and U9982 (N_9982,N_8220,N_8215);
or U9983 (N_9983,N_6915,N_6716);
and U9984 (N_9984,N_8057,N_7654);
nor U9985 (N_9985,N_7777,N_7729);
nand U9986 (N_9986,N_7265,N_6760);
or U9987 (N_9987,N_8254,N_8386);
nand U9988 (N_9988,N_8635,N_7044);
or U9989 (N_9989,N_7034,N_6728);
nand U9990 (N_9990,N_7256,N_6214);
and U9991 (N_9991,N_7964,N_6795);
nor U9992 (N_9992,N_6949,N_7612);
nand U9993 (N_9993,N_6548,N_7157);
nor U9994 (N_9994,N_8587,N_6483);
nor U9995 (N_9995,N_8419,N_8599);
nor U9996 (N_9996,N_6114,N_8797);
nand U9997 (N_9997,N_7681,N_8304);
nor U9998 (N_9998,N_7301,N_6150);
and U9999 (N_9999,N_6961,N_6198);
or U10000 (N_10000,N_8174,N_6260);
nand U10001 (N_10001,N_6988,N_6923);
nor U10002 (N_10002,N_7675,N_7305);
nor U10003 (N_10003,N_6035,N_7475);
and U10004 (N_10004,N_6410,N_6206);
nor U10005 (N_10005,N_6274,N_7756);
nor U10006 (N_10006,N_7031,N_7876);
or U10007 (N_10007,N_8431,N_8093);
nand U10008 (N_10008,N_8956,N_7245);
nor U10009 (N_10009,N_6953,N_7428);
nand U10010 (N_10010,N_7230,N_8828);
nand U10011 (N_10011,N_7368,N_7346);
and U10012 (N_10012,N_6175,N_7835);
nor U10013 (N_10013,N_8991,N_6629);
or U10014 (N_10014,N_8301,N_7973);
nor U10015 (N_10015,N_8083,N_8619);
nand U10016 (N_10016,N_7792,N_6094);
nand U10017 (N_10017,N_7058,N_6596);
or U10018 (N_10018,N_7783,N_7395);
and U10019 (N_10019,N_8664,N_7046);
xnor U10020 (N_10020,N_7049,N_8382);
or U10021 (N_10021,N_8284,N_7126);
nand U10022 (N_10022,N_6781,N_8756);
or U10023 (N_10023,N_8184,N_8801);
or U10024 (N_10024,N_7856,N_6417);
nand U10025 (N_10025,N_8548,N_8866);
nor U10026 (N_10026,N_7434,N_7635);
nand U10027 (N_10027,N_8859,N_8951);
or U10028 (N_10028,N_8349,N_7970);
and U10029 (N_10029,N_7459,N_7847);
nor U10030 (N_10030,N_8877,N_8494);
nand U10031 (N_10031,N_7204,N_6892);
nor U10032 (N_10032,N_8506,N_6718);
and U10033 (N_10033,N_8437,N_7875);
nand U10034 (N_10034,N_8425,N_6092);
or U10035 (N_10035,N_7155,N_7489);
nor U10036 (N_10036,N_8943,N_8317);
and U10037 (N_10037,N_6311,N_8007);
and U10038 (N_10038,N_8641,N_7758);
and U10039 (N_10039,N_8870,N_8845);
or U10040 (N_10040,N_6884,N_7251);
or U10041 (N_10041,N_6841,N_7537);
or U10042 (N_10042,N_8955,N_6279);
and U10043 (N_10043,N_6875,N_6442);
or U10044 (N_10044,N_7618,N_7774);
and U10045 (N_10045,N_7503,N_8958);
and U10046 (N_10046,N_7227,N_8232);
or U10047 (N_10047,N_7029,N_7077);
or U10048 (N_10048,N_7938,N_8355);
nand U10049 (N_10049,N_8101,N_7776);
and U10050 (N_10050,N_6895,N_7313);
and U10051 (N_10051,N_7462,N_6602);
nand U10052 (N_10052,N_8540,N_6842);
or U10053 (N_10053,N_8600,N_7839);
nand U10054 (N_10054,N_7865,N_8936);
or U10055 (N_10055,N_8365,N_7829);
and U10056 (N_10056,N_7609,N_7344);
and U10057 (N_10057,N_7989,N_7626);
nor U10058 (N_10058,N_7358,N_7625);
xor U10059 (N_10059,N_8462,N_8389);
nor U10060 (N_10060,N_6349,N_8019);
nand U10061 (N_10061,N_7166,N_8518);
nor U10062 (N_10062,N_7872,N_7535);
nor U10063 (N_10063,N_6434,N_7461);
or U10064 (N_10064,N_7806,N_6392);
nand U10065 (N_10065,N_8281,N_6909);
and U10066 (N_10066,N_6725,N_8805);
and U10067 (N_10067,N_6164,N_7038);
nor U10068 (N_10068,N_8095,N_7040);
nand U10069 (N_10069,N_8823,N_8903);
xor U10070 (N_10070,N_8747,N_6197);
xnor U10071 (N_10071,N_6919,N_7377);
nand U10072 (N_10072,N_7953,N_7749);
nor U10073 (N_10073,N_7043,N_8928);
nand U10074 (N_10074,N_8374,N_8194);
or U10075 (N_10075,N_7445,N_7292);
or U10076 (N_10076,N_7009,N_7482);
nor U10077 (N_10077,N_8803,N_8451);
and U10078 (N_10078,N_8424,N_7309);
or U10079 (N_10079,N_7525,N_6639);
and U10080 (N_10080,N_6514,N_8003);
nor U10081 (N_10081,N_7608,N_8198);
or U10082 (N_10082,N_8521,N_7151);
and U10083 (N_10083,N_8864,N_7453);
nor U10084 (N_10084,N_8715,N_6836);
nor U10085 (N_10085,N_6735,N_8687);
nor U10086 (N_10086,N_8782,N_8124);
and U10087 (N_10087,N_8337,N_6621);
nor U10088 (N_10088,N_8065,N_6893);
or U10089 (N_10089,N_8680,N_8524);
nand U10090 (N_10090,N_7194,N_7961);
xnor U10091 (N_10091,N_8694,N_6530);
or U10092 (N_10092,N_7019,N_6484);
xnor U10093 (N_10093,N_6420,N_7354);
and U10094 (N_10094,N_8515,N_7074);
nor U10095 (N_10095,N_8887,N_7392);
and U10096 (N_10096,N_8399,N_6512);
or U10097 (N_10097,N_7250,N_6324);
nand U10098 (N_10098,N_8366,N_8831);
nand U10099 (N_10099,N_6758,N_8141);
nor U10100 (N_10100,N_7357,N_7372);
xnor U10101 (N_10101,N_8947,N_7162);
nand U10102 (N_10102,N_6591,N_8513);
and U10103 (N_10103,N_6660,N_7611);
nor U10104 (N_10104,N_6196,N_7969);
nor U10105 (N_10105,N_7736,N_8440);
nand U10106 (N_10106,N_8495,N_7614);
or U10107 (N_10107,N_7087,N_6364);
and U10108 (N_10108,N_8692,N_8486);
xor U10109 (N_10109,N_8726,N_6289);
and U10110 (N_10110,N_7811,N_8116);
nand U10111 (N_10111,N_8088,N_8586);
nor U10112 (N_10112,N_6192,N_6047);
and U10113 (N_10113,N_7721,N_8523);
xor U10114 (N_10114,N_7319,N_8033);
nand U10115 (N_10115,N_8817,N_7738);
and U10116 (N_10116,N_8666,N_6046);
and U10117 (N_10117,N_8179,N_6515);
and U10118 (N_10118,N_7273,N_8652);
and U10119 (N_10119,N_6772,N_7300);
nand U10120 (N_10120,N_7402,N_8711);
nor U10121 (N_10121,N_6481,N_6474);
xnor U10122 (N_10122,N_8783,N_8737);
and U10123 (N_10123,N_6012,N_7419);
and U10124 (N_10124,N_6766,N_8055);
xnor U10125 (N_10125,N_8189,N_7946);
xnor U10126 (N_10126,N_7465,N_8070);
or U10127 (N_10127,N_8476,N_8196);
and U10128 (N_10128,N_8716,N_6467);
and U10129 (N_10129,N_8799,N_7706);
nand U10130 (N_10130,N_6752,N_8676);
nor U10131 (N_10131,N_8634,N_7712);
or U10132 (N_10132,N_8734,N_7366);
nand U10133 (N_10133,N_8040,N_7072);
or U10134 (N_10134,N_8242,N_6459);
xor U10135 (N_10135,N_7701,N_8160);
or U10136 (N_10136,N_7820,N_8669);
or U10137 (N_10137,N_6087,N_6748);
nand U10138 (N_10138,N_8477,N_7573);
or U10139 (N_10139,N_7000,N_6099);
nand U10140 (N_10140,N_7585,N_6336);
nor U10141 (N_10141,N_6497,N_6697);
or U10142 (N_10142,N_6224,N_8762);
or U10143 (N_10143,N_8391,N_8483);
or U10144 (N_10144,N_7723,N_8278);
xnor U10145 (N_10145,N_7108,N_8119);
xnor U10146 (N_10146,N_7645,N_7914);
and U10147 (N_10147,N_8771,N_8222);
or U10148 (N_10148,N_7005,N_7521);
nor U10149 (N_10149,N_7510,N_8047);
or U10150 (N_10150,N_6852,N_6255);
nand U10151 (N_10151,N_6799,N_8590);
and U10152 (N_10152,N_8535,N_8570);
and U10153 (N_10153,N_8263,N_8107);
nor U10154 (N_10154,N_8976,N_6344);
or U10155 (N_10155,N_8613,N_7718);
nand U10156 (N_10156,N_6264,N_6405);
and U10157 (N_10157,N_7269,N_6833);
and U10158 (N_10158,N_7578,N_8899);
nand U10159 (N_10159,N_6305,N_7745);
nor U10160 (N_10160,N_7885,N_7582);
nor U10161 (N_10161,N_7253,N_7909);
nor U10162 (N_10162,N_8610,N_7869);
nand U10163 (N_10163,N_6785,N_8673);
nor U10164 (N_10164,N_6661,N_7041);
xor U10165 (N_10165,N_8959,N_6779);
nand U10166 (N_10166,N_6326,N_7837);
nor U10167 (N_10167,N_7707,N_6071);
and U10168 (N_10168,N_6470,N_6916);
or U10169 (N_10169,N_6989,N_7229);
nand U10170 (N_10170,N_8781,N_8628);
nor U10171 (N_10171,N_8950,N_6411);
or U10172 (N_10172,N_6498,N_6102);
nor U10173 (N_10173,N_6941,N_6698);
or U10174 (N_10174,N_7427,N_6636);
or U10175 (N_10175,N_7687,N_7506);
and U10176 (N_10176,N_8779,N_7128);
xor U10177 (N_10177,N_6822,N_7595);
and U10178 (N_10178,N_8339,N_8873);
xnor U10179 (N_10179,N_6101,N_6520);
nor U10180 (N_10180,N_6412,N_8717);
xor U10181 (N_10181,N_8465,N_6848);
nand U10182 (N_10182,N_7910,N_8536);
and U10183 (N_10183,N_7013,N_6700);
nand U10184 (N_10184,N_7533,N_7580);
nor U10185 (N_10185,N_7977,N_7025);
or U10186 (N_10186,N_7957,N_8537);
xnor U10187 (N_10187,N_6603,N_6907);
or U10188 (N_10188,N_6986,N_6248);
nor U10189 (N_10189,N_8642,N_8054);
nor U10190 (N_10190,N_8252,N_7299);
and U10191 (N_10191,N_8482,N_8566);
or U10192 (N_10192,N_6717,N_7073);
nor U10193 (N_10193,N_6939,N_6756);
nand U10194 (N_10194,N_7873,N_6328);
xnor U10195 (N_10195,N_6541,N_6229);
nor U10196 (N_10196,N_8125,N_8665);
nand U10197 (N_10197,N_7389,N_6204);
and U10198 (N_10198,N_6141,N_7678);
and U10199 (N_10199,N_6951,N_7575);
nand U10200 (N_10200,N_7567,N_7466);
nor U10201 (N_10201,N_8293,N_6814);
nor U10202 (N_10202,N_6170,N_7008);
nand U10203 (N_10203,N_6331,N_7494);
xnor U10204 (N_10204,N_6409,N_6604);
and U10205 (N_10205,N_8615,N_6215);
xnor U10206 (N_10206,N_8824,N_8948);
nor U10207 (N_10207,N_6918,N_6136);
nand U10208 (N_10208,N_6276,N_7526);
and U10209 (N_10209,N_6503,N_7217);
and U10210 (N_10210,N_7850,N_6195);
and U10211 (N_10211,N_7743,N_6638);
and U10212 (N_10212,N_7840,N_6663);
and U10213 (N_10213,N_8131,N_7800);
and U10214 (N_10214,N_7188,N_6002);
nand U10215 (N_10215,N_8009,N_7817);
or U10216 (N_10216,N_6190,N_6863);
nor U10217 (N_10217,N_7288,N_7605);
and U10218 (N_10218,N_8173,N_7391);
or U10219 (N_10219,N_6774,N_6158);
or U10220 (N_10220,N_6354,N_6308);
nor U10221 (N_10221,N_8299,N_7473);
and U10222 (N_10222,N_7664,N_7621);
nand U10223 (N_10223,N_7704,N_7236);
and U10224 (N_10224,N_8624,N_6947);
nor U10225 (N_10225,N_7760,N_7880);
nand U10226 (N_10226,N_7105,N_7650);
nand U10227 (N_10227,N_7825,N_8433);
and U10228 (N_10228,N_6278,N_7202);
and U10229 (N_10229,N_6921,N_8638);
or U10230 (N_10230,N_8163,N_7057);
xnor U10231 (N_10231,N_7861,N_7660);
and U10232 (N_10232,N_8967,N_7232);
or U10233 (N_10233,N_6867,N_7139);
and U10234 (N_10234,N_7224,N_8882);
and U10235 (N_10235,N_8849,N_8622);
nor U10236 (N_10236,N_8123,N_8485);
nand U10237 (N_10237,N_6024,N_6813);
or U10238 (N_10238,N_6318,N_7937);
or U10239 (N_10239,N_8336,N_8719);
nor U10240 (N_10240,N_7076,N_6960);
nand U10241 (N_10241,N_8752,N_6958);
nor U10242 (N_10242,N_7257,N_7986);
or U10243 (N_10243,N_6824,N_7949);
or U10244 (N_10244,N_6109,N_8180);
and U10245 (N_10245,N_8961,N_7362);
or U10246 (N_10246,N_7201,N_7131);
and U10247 (N_10247,N_7593,N_6847);
or U10248 (N_10248,N_7159,N_6225);
and U10249 (N_10249,N_8378,N_6054);
nor U10250 (N_10250,N_6209,N_7123);
or U10251 (N_10251,N_8312,N_7393);
xor U10252 (N_10252,N_6567,N_7045);
xor U10253 (N_10253,N_7287,N_7143);
and U10254 (N_10254,N_6585,N_7423);
or U10255 (N_10255,N_6675,N_8140);
nor U10256 (N_10256,N_8772,N_8069);
xor U10257 (N_10257,N_8758,N_6665);
and U10258 (N_10258,N_7145,N_6443);
xor U10259 (N_10259,N_6131,N_7093);
or U10260 (N_10260,N_8256,N_7050);
or U10261 (N_10261,N_6310,N_7411);
or U10262 (N_10262,N_8617,N_6317);
xnor U10263 (N_10263,N_6041,N_8689);
nand U10264 (N_10264,N_8015,N_7271);
nor U10265 (N_10265,N_7064,N_6990);
and U10266 (N_10266,N_8340,N_7112);
nor U10267 (N_10267,N_7012,N_8531);
and U10268 (N_10268,N_6703,N_7146);
and U10269 (N_10269,N_7165,N_7933);
xor U10270 (N_10270,N_7771,N_6468);
and U10271 (N_10271,N_6300,N_6188);
or U10272 (N_10272,N_7916,N_7690);
and U10273 (N_10273,N_8503,N_7408);
or U10274 (N_10274,N_6100,N_8177);
nor U10275 (N_10275,N_8601,N_8648);
nand U10276 (N_10276,N_8501,N_7951);
nor U10277 (N_10277,N_6962,N_6132);
nand U10278 (N_10278,N_8318,N_8678);
or U10279 (N_10279,N_7308,N_7499);
and U10280 (N_10280,N_6608,N_6105);
and U10281 (N_10281,N_7892,N_7559);
nor U10282 (N_10282,N_7488,N_7320);
or U10283 (N_10283,N_8962,N_6879);
nand U10284 (N_10284,N_8580,N_6403);
nor U10285 (N_10285,N_6091,N_7310);
xor U10286 (N_10286,N_6089,N_8878);
nand U10287 (N_10287,N_7508,N_6329);
nor U10288 (N_10288,N_8045,N_6032);
or U10289 (N_10289,N_6570,N_6980);
and U10290 (N_10290,N_7765,N_7987);
xnor U10291 (N_10291,N_6971,N_6641);
nand U10292 (N_10292,N_7231,N_8644);
nor U10293 (N_10293,N_6948,N_6656);
and U10294 (N_10294,N_6521,N_6507);
and U10295 (N_10295,N_7172,N_7794);
nor U10296 (N_10296,N_7668,N_6739);
or U10297 (N_10297,N_8243,N_6965);
nor U10298 (N_10298,N_8435,N_7641);
or U10299 (N_10299,N_7999,N_8089);
nor U10300 (N_10300,N_7379,N_8473);
and U10301 (N_10301,N_7198,N_7333);
or U10302 (N_10302,N_6194,N_6362);
and U10303 (N_10303,N_7067,N_6036);
xor U10304 (N_10304,N_8868,N_7913);
xnor U10305 (N_10305,N_6606,N_8370);
or U10306 (N_10306,N_8999,N_7919);
or U10307 (N_10307,N_8161,N_8671);
nor U10308 (N_10308,N_6508,N_7429);
and U10309 (N_10309,N_8311,N_7576);
nand U10310 (N_10310,N_8185,N_7282);
nand U10311 (N_10311,N_8068,N_7370);
nand U10312 (N_10312,N_6690,N_8757);
nor U10313 (N_10313,N_6794,N_6341);
nand U10314 (N_10314,N_6096,N_6288);
and U10315 (N_10315,N_6978,N_8932);
xor U10316 (N_10316,N_6004,N_7688);
nor U10317 (N_10317,N_7433,N_8292);
nor U10318 (N_10318,N_6757,N_8468);
and U10319 (N_10319,N_7599,N_6407);
nand U10320 (N_10320,N_8974,N_8656);
or U10321 (N_10321,N_6572,N_8874);
nor U10322 (N_10322,N_8138,N_8142);
nor U10323 (N_10323,N_8208,N_8848);
xnor U10324 (N_10324,N_7117,N_8056);
nor U10325 (N_10325,N_8806,N_8598);
nand U10326 (N_10326,N_8014,N_8741);
or U10327 (N_10327,N_8004,N_6618);
nand U10328 (N_10328,N_8096,N_7274);
or U10329 (N_10329,N_8759,N_7385);
or U10330 (N_10330,N_8092,N_8751);
nor U10331 (N_10331,N_6914,N_7940);
or U10332 (N_10332,N_6858,N_6732);
nand U10333 (N_10333,N_6375,N_7586);
and U10334 (N_10334,N_6458,N_8767);
nor U10335 (N_10335,N_8373,N_8498);
nor U10336 (N_10336,N_6620,N_8387);
xnor U10337 (N_10337,N_6878,N_7312);
xor U10338 (N_10338,N_6061,N_8822);
nand U10339 (N_10339,N_8578,N_8558);
or U10340 (N_10340,N_6230,N_6899);
nor U10341 (N_10341,N_6611,N_8245);
nand U10342 (N_10342,N_6476,N_6657);
xnor U10343 (N_10343,N_7530,N_6321);
or U10344 (N_10344,N_6653,N_6232);
nand U10345 (N_10345,N_6234,N_8938);
and U10346 (N_10346,N_8028,N_7472);
or U10347 (N_10347,N_6889,N_6927);
and U10348 (N_10348,N_6489,N_8187);
or U10349 (N_10349,N_6243,N_7571);
xor U10350 (N_10350,N_6031,N_7927);
xor U10351 (N_10351,N_7053,N_6993);
nor U10352 (N_10352,N_8915,N_6378);
and U10353 (N_10353,N_6391,N_8071);
and U10354 (N_10354,N_6017,N_6077);
nor U10355 (N_10355,N_8129,N_7581);
nand U10356 (N_10356,N_6701,N_7065);
and U10357 (N_10357,N_7086,N_8871);
or U10358 (N_10358,N_7270,N_7983);
and U10359 (N_10359,N_6984,N_8489);
nor U10360 (N_10360,N_6439,N_8810);
or U10361 (N_10361,N_8099,N_7268);
or U10362 (N_10362,N_8902,N_6790);
nand U10363 (N_10363,N_7100,N_8750);
nand U10364 (N_10364,N_7492,N_6767);
nand U10365 (N_10365,N_6808,N_8077);
nor U10366 (N_10366,N_6395,N_7097);
nand U10367 (N_10367,N_7186,N_6676);
and U10368 (N_10368,N_6898,N_7691);
and U10369 (N_10369,N_7676,N_8010);
or U10370 (N_10370,N_8048,N_8992);
or U10371 (N_10371,N_6702,N_6696);
or U10372 (N_10372,N_7845,N_7750);
xor U10373 (N_10373,N_7504,N_6576);
and U10374 (N_10374,N_7153,N_7261);
xnor U10375 (N_10375,N_8442,N_7536);
nor U10376 (N_10376,N_6291,N_8448);
nor U10377 (N_10377,N_8176,N_6583);
and U10378 (N_10378,N_7697,N_7470);
and U10379 (N_10379,N_7859,N_6738);
nand U10380 (N_10380,N_7805,N_7340);
nand U10381 (N_10381,N_8302,N_6397);
nand U10382 (N_10382,N_6290,N_8470);
and U10383 (N_10383,N_6789,N_6505);
or U10384 (N_10384,N_8029,N_8905);
or U10385 (N_10385,N_7561,N_8591);
nand U10386 (N_10386,N_6062,N_8192);
or U10387 (N_10387,N_6133,N_6361);
or U10388 (N_10388,N_8217,N_6835);
nor U10389 (N_10389,N_6556,N_6139);
nand U10390 (N_10390,N_7502,N_8939);
or U10391 (N_10391,N_7841,N_7456);
nor U10392 (N_10392,N_8335,N_6577);
nor U10393 (N_10393,N_7734,N_7024);
and U10394 (N_10394,N_6271,N_6177);
nand U10395 (N_10395,N_8247,N_6982);
nand U10396 (N_10396,N_8650,N_7838);
nor U10397 (N_10397,N_6667,N_8832);
or U10398 (N_10398,N_7674,N_6762);
nor U10399 (N_10399,N_6453,N_8895);
nor U10400 (N_10400,N_6882,N_8703);
or U10401 (N_10401,N_6877,N_7901);
nor U10402 (N_10402,N_7994,N_8894);
and U10403 (N_10403,N_6491,N_6821);
and U10404 (N_10404,N_6313,N_8390);
nand U10405 (N_10405,N_6564,N_7135);
and U10406 (N_10406,N_7115,N_7893);
nor U10407 (N_10407,N_8016,N_7941);
or U10408 (N_10408,N_7851,N_6323);
nand U10409 (N_10409,N_8574,N_6976);
xor U10410 (N_10410,N_8169,N_8073);
nand U10411 (N_10411,N_6664,N_6612);
and U10412 (N_10412,N_6181,N_7033);
nand U10413 (N_10413,N_8736,N_7069);
or U10414 (N_10414,N_6582,N_6995);
nand U10415 (N_10415,N_8287,N_7089);
nand U10416 (N_10416,N_6926,N_8602);
and U10417 (N_10417,N_6297,N_8212);
nand U10418 (N_10418,N_8159,N_8147);
nor U10419 (N_10419,N_7356,N_6151);
and U10420 (N_10420,N_8798,N_6370);
or U10421 (N_10421,N_8258,N_7831);
or U10422 (N_10422,N_6964,N_6053);
nor U10423 (N_10423,N_7048,N_6400);
and U10424 (N_10424,N_7109,N_7848);
nand U10425 (N_10425,N_8086,N_8637);
and U10426 (N_10426,N_6796,N_8790);
or U10427 (N_10427,N_7160,N_6793);
or U10428 (N_10428,N_7360,N_7304);
xnor U10429 (N_10429,N_7460,N_8354);
nor U10430 (N_10430,N_7092,N_6237);
and U10431 (N_10431,N_6973,N_8499);
nor U10432 (N_10432,N_7405,N_7498);
or U10433 (N_10433,N_6350,N_8682);
and U10434 (N_10434,N_8654,N_7807);
and U10435 (N_10435,N_6966,N_8983);
xor U10436 (N_10436,N_7956,N_6810);
or U10437 (N_10437,N_6678,N_6659);
and U10438 (N_10438,N_8000,N_7111);
nor U10439 (N_10439,N_8013,N_7677);
or U10440 (N_10440,N_8960,N_6531);
nor U10441 (N_10441,N_8218,N_8036);
and U10442 (N_10442,N_6633,N_6357);
nor U10443 (N_10443,N_7306,N_7833);
nand U10444 (N_10444,N_7830,N_7886);
nand U10445 (N_10445,N_6027,N_6642);
and U10446 (N_10446,N_6049,N_6016);
or U10447 (N_10447,N_8103,N_8202);
xor U10448 (N_10448,N_6819,N_7454);
nor U10449 (N_10449,N_8543,N_6186);
or U10450 (N_10450,N_8394,N_6932);
and U10451 (N_10451,N_7415,N_8027);
and U10452 (N_10452,N_7754,N_7156);
nand U10453 (N_10453,N_8975,N_8420);
nand U10454 (N_10454,N_6334,N_8078);
nand U10455 (N_10455,N_6866,N_7524);
nand U10456 (N_10456,N_6495,N_8546);
and U10457 (N_10457,N_6466,N_6763);
and U10458 (N_10458,N_6811,N_6270);
and U10459 (N_10459,N_8248,N_7540);
and U10460 (N_10460,N_8841,N_6356);
or U10461 (N_10461,N_6436,N_8544);
or U10462 (N_10462,N_7042,N_6688);
or U10463 (N_10463,N_6534,N_8527);
xor U10464 (N_10464,N_8743,N_6242);
and U10465 (N_10465,N_7709,N_7962);
and U10466 (N_10466,N_6333,N_6000);
or U10467 (N_10467,N_7948,N_6269);
nand U10468 (N_10468,N_7407,N_6587);
nand U10469 (N_10469,N_8944,N_6157);
and U10470 (N_10470,N_6751,N_6345);
nand U10471 (N_10471,N_6963,N_7514);
nand U10472 (N_10472,N_7761,N_7773);
nand U10473 (N_10473,N_6057,N_7564);
xor U10474 (N_10474,N_8219,N_8555);
nor U10475 (N_10475,N_8188,N_8594);
and U10476 (N_10476,N_7784,N_7168);
nor U10477 (N_10477,N_8862,N_7591);
or U10478 (N_10478,N_7221,N_6455);
or U10479 (N_10479,N_6048,N_6744);
nor U10480 (N_10480,N_8764,N_8490);
nand U10481 (N_10481,N_6073,N_7637);
nor U10482 (N_10482,N_7332,N_8729);
nor U10483 (N_10483,N_7443,N_7769);
or U10484 (N_10484,N_7623,N_8030);
nor U10485 (N_10485,N_7915,N_8625);
nand U10486 (N_10486,N_6788,N_8334);
nand U10487 (N_10487,N_7302,N_7484);
xor U10488 (N_10488,N_6492,N_6005);
nand U10489 (N_10489,N_7967,N_7171);
nand U10490 (N_10490,N_6699,N_7950);
or U10491 (N_10491,N_6784,N_7016);
xnor U10492 (N_10492,N_8685,N_6677);
or U10493 (N_10493,N_8631,N_6235);
xnor U10494 (N_10494,N_6686,N_8153);
or U10495 (N_10495,N_6160,N_8551);
or U10496 (N_10496,N_6616,N_7782);
nor U10497 (N_10497,N_8838,N_7632);
or U10498 (N_10498,N_8957,N_7444);
or U10499 (N_10499,N_6137,N_8042);
nor U10500 (N_10500,N_7190,N_8649);
or U10501 (N_10501,N_8630,N_6986);
nor U10502 (N_10502,N_6246,N_6156);
nand U10503 (N_10503,N_8632,N_6408);
nor U10504 (N_10504,N_7707,N_8960);
nand U10505 (N_10505,N_8181,N_8067);
nor U10506 (N_10506,N_8396,N_7018);
nor U10507 (N_10507,N_6218,N_6994);
or U10508 (N_10508,N_6644,N_8654);
nand U10509 (N_10509,N_7799,N_7200);
nor U10510 (N_10510,N_6920,N_8736);
and U10511 (N_10511,N_7363,N_7256);
and U10512 (N_10512,N_8269,N_7344);
nor U10513 (N_10513,N_7700,N_8374);
nand U10514 (N_10514,N_7799,N_8470);
xor U10515 (N_10515,N_7562,N_8823);
or U10516 (N_10516,N_7906,N_6939);
nand U10517 (N_10517,N_8837,N_7902);
nor U10518 (N_10518,N_7171,N_7094);
or U10519 (N_10519,N_8856,N_6945);
or U10520 (N_10520,N_8156,N_6855);
or U10521 (N_10521,N_8805,N_8948);
and U10522 (N_10522,N_6021,N_8315);
or U10523 (N_10523,N_8039,N_7008);
and U10524 (N_10524,N_7811,N_7970);
nor U10525 (N_10525,N_8178,N_8353);
xor U10526 (N_10526,N_8088,N_7623);
nor U10527 (N_10527,N_6907,N_7762);
or U10528 (N_10528,N_8649,N_6935);
nand U10529 (N_10529,N_8564,N_8593);
nor U10530 (N_10530,N_7755,N_7156);
nor U10531 (N_10531,N_8978,N_8015);
or U10532 (N_10532,N_7216,N_7836);
and U10533 (N_10533,N_6245,N_6018);
nor U10534 (N_10534,N_8392,N_8792);
nor U10535 (N_10535,N_6570,N_8735);
or U10536 (N_10536,N_7533,N_7866);
or U10537 (N_10537,N_8670,N_8052);
nand U10538 (N_10538,N_8067,N_8426);
or U10539 (N_10539,N_7695,N_6467);
or U10540 (N_10540,N_8499,N_7469);
and U10541 (N_10541,N_7549,N_8499);
and U10542 (N_10542,N_7164,N_6407);
nand U10543 (N_10543,N_7794,N_6072);
or U10544 (N_10544,N_8487,N_6996);
xnor U10545 (N_10545,N_8478,N_7570);
nor U10546 (N_10546,N_6973,N_8960);
nand U10547 (N_10547,N_6355,N_7294);
nand U10548 (N_10548,N_7171,N_8852);
nor U10549 (N_10549,N_6134,N_7973);
nor U10550 (N_10550,N_8595,N_6268);
nand U10551 (N_10551,N_6213,N_6576);
nand U10552 (N_10552,N_6282,N_8704);
xor U10553 (N_10553,N_7687,N_6690);
nor U10554 (N_10554,N_6382,N_6338);
nand U10555 (N_10555,N_8362,N_7721);
or U10556 (N_10556,N_8011,N_6684);
nand U10557 (N_10557,N_7941,N_8115);
xnor U10558 (N_10558,N_6416,N_8202);
or U10559 (N_10559,N_7937,N_7712);
or U10560 (N_10560,N_8832,N_8670);
nand U10561 (N_10561,N_6687,N_7825);
and U10562 (N_10562,N_7355,N_8420);
xor U10563 (N_10563,N_8642,N_7304);
and U10564 (N_10564,N_7678,N_6515);
or U10565 (N_10565,N_8142,N_6536);
nand U10566 (N_10566,N_7652,N_6133);
nor U10567 (N_10567,N_6842,N_8718);
and U10568 (N_10568,N_7058,N_8611);
nand U10569 (N_10569,N_8948,N_8832);
nand U10570 (N_10570,N_8154,N_7974);
and U10571 (N_10571,N_6213,N_8993);
nor U10572 (N_10572,N_6164,N_8359);
nand U10573 (N_10573,N_6888,N_6055);
and U10574 (N_10574,N_7906,N_7571);
nor U10575 (N_10575,N_8293,N_7689);
or U10576 (N_10576,N_6055,N_7555);
nand U10577 (N_10577,N_7374,N_8485);
and U10578 (N_10578,N_6091,N_8937);
and U10579 (N_10579,N_7269,N_7923);
xor U10580 (N_10580,N_7314,N_8261);
xnor U10581 (N_10581,N_6103,N_7538);
nor U10582 (N_10582,N_6730,N_7474);
nand U10583 (N_10583,N_7672,N_8191);
or U10584 (N_10584,N_8756,N_7061);
or U10585 (N_10585,N_8314,N_6275);
nor U10586 (N_10586,N_6565,N_6993);
and U10587 (N_10587,N_6900,N_6269);
or U10588 (N_10588,N_6770,N_7682);
xor U10589 (N_10589,N_7081,N_6527);
nand U10590 (N_10590,N_8918,N_7861);
nand U10591 (N_10591,N_8953,N_8676);
nand U10592 (N_10592,N_7255,N_8125);
and U10593 (N_10593,N_8593,N_8866);
nor U10594 (N_10594,N_6515,N_6981);
or U10595 (N_10595,N_8774,N_6606);
xor U10596 (N_10596,N_7044,N_6059);
or U10597 (N_10597,N_6014,N_8102);
nor U10598 (N_10598,N_7030,N_7697);
nor U10599 (N_10599,N_7683,N_8202);
and U10600 (N_10600,N_8018,N_6351);
and U10601 (N_10601,N_6203,N_8410);
xnor U10602 (N_10602,N_7200,N_6373);
and U10603 (N_10603,N_6885,N_8004);
nand U10604 (N_10604,N_7183,N_8990);
and U10605 (N_10605,N_7994,N_8254);
or U10606 (N_10606,N_8528,N_7394);
nor U10607 (N_10607,N_8852,N_6396);
or U10608 (N_10608,N_8142,N_7662);
or U10609 (N_10609,N_8848,N_6091);
and U10610 (N_10610,N_8208,N_8658);
or U10611 (N_10611,N_7926,N_7211);
nand U10612 (N_10612,N_6302,N_7477);
nor U10613 (N_10613,N_6095,N_8895);
or U10614 (N_10614,N_6254,N_7418);
and U10615 (N_10615,N_7062,N_8465);
xor U10616 (N_10616,N_7858,N_6561);
nor U10617 (N_10617,N_6143,N_8380);
xor U10618 (N_10618,N_6284,N_8570);
nor U10619 (N_10619,N_8891,N_6473);
or U10620 (N_10620,N_8005,N_7371);
and U10621 (N_10621,N_6718,N_8190);
nor U10622 (N_10622,N_8547,N_7752);
or U10623 (N_10623,N_7944,N_8636);
and U10624 (N_10624,N_7086,N_7439);
nand U10625 (N_10625,N_8565,N_7491);
nor U10626 (N_10626,N_8579,N_6272);
or U10627 (N_10627,N_6091,N_6431);
or U10628 (N_10628,N_8106,N_6086);
or U10629 (N_10629,N_7417,N_7316);
xor U10630 (N_10630,N_7615,N_6846);
nand U10631 (N_10631,N_7782,N_7102);
and U10632 (N_10632,N_6553,N_7162);
and U10633 (N_10633,N_7796,N_8553);
and U10634 (N_10634,N_6981,N_7351);
nor U10635 (N_10635,N_8903,N_6586);
and U10636 (N_10636,N_8227,N_7987);
or U10637 (N_10637,N_6207,N_6777);
xor U10638 (N_10638,N_7110,N_8251);
or U10639 (N_10639,N_7136,N_6299);
nand U10640 (N_10640,N_7955,N_6952);
or U10641 (N_10641,N_8252,N_7388);
or U10642 (N_10642,N_7609,N_6921);
nand U10643 (N_10643,N_8063,N_6172);
xor U10644 (N_10644,N_7356,N_7515);
xnor U10645 (N_10645,N_7407,N_7680);
nor U10646 (N_10646,N_6429,N_7014);
nor U10647 (N_10647,N_6286,N_7878);
and U10648 (N_10648,N_8522,N_6880);
nand U10649 (N_10649,N_7739,N_7240);
nand U10650 (N_10650,N_8534,N_7544);
nor U10651 (N_10651,N_6968,N_6756);
xor U10652 (N_10652,N_7346,N_7269);
nor U10653 (N_10653,N_7894,N_6805);
or U10654 (N_10654,N_8466,N_6220);
or U10655 (N_10655,N_8060,N_8062);
nand U10656 (N_10656,N_6640,N_8658);
and U10657 (N_10657,N_6661,N_7951);
and U10658 (N_10658,N_8439,N_6958);
xor U10659 (N_10659,N_8656,N_6315);
and U10660 (N_10660,N_8714,N_8790);
nor U10661 (N_10661,N_7131,N_7619);
and U10662 (N_10662,N_8559,N_7624);
nand U10663 (N_10663,N_7116,N_8210);
nand U10664 (N_10664,N_6850,N_8492);
and U10665 (N_10665,N_6113,N_6453);
or U10666 (N_10666,N_8228,N_6981);
or U10667 (N_10667,N_7945,N_6947);
nor U10668 (N_10668,N_7546,N_7118);
or U10669 (N_10669,N_6920,N_6400);
and U10670 (N_10670,N_6420,N_7463);
xnor U10671 (N_10671,N_8158,N_8840);
xnor U10672 (N_10672,N_7163,N_7433);
and U10673 (N_10673,N_7263,N_8855);
xor U10674 (N_10674,N_6285,N_8588);
nand U10675 (N_10675,N_6018,N_8495);
nor U10676 (N_10676,N_7362,N_6664);
or U10677 (N_10677,N_8915,N_6287);
or U10678 (N_10678,N_7252,N_6196);
nor U10679 (N_10679,N_8343,N_7334);
nor U10680 (N_10680,N_7456,N_7911);
xnor U10681 (N_10681,N_7251,N_6072);
and U10682 (N_10682,N_6473,N_7881);
or U10683 (N_10683,N_6654,N_7106);
and U10684 (N_10684,N_8835,N_7880);
nand U10685 (N_10685,N_6312,N_8314);
nand U10686 (N_10686,N_8430,N_8729);
and U10687 (N_10687,N_6033,N_7989);
or U10688 (N_10688,N_8602,N_7168);
and U10689 (N_10689,N_6363,N_8018);
and U10690 (N_10690,N_7890,N_8231);
or U10691 (N_10691,N_7626,N_6157);
xor U10692 (N_10692,N_8606,N_6071);
nor U10693 (N_10693,N_8088,N_6356);
nor U10694 (N_10694,N_7536,N_8636);
xnor U10695 (N_10695,N_6002,N_8405);
nand U10696 (N_10696,N_8817,N_7050);
and U10697 (N_10697,N_6913,N_7403);
xnor U10698 (N_10698,N_7345,N_6424);
and U10699 (N_10699,N_6079,N_8685);
or U10700 (N_10700,N_8242,N_6324);
nor U10701 (N_10701,N_6174,N_6076);
nand U10702 (N_10702,N_7165,N_7511);
xnor U10703 (N_10703,N_8170,N_8100);
nand U10704 (N_10704,N_7424,N_7969);
and U10705 (N_10705,N_8770,N_6346);
nand U10706 (N_10706,N_7560,N_8473);
or U10707 (N_10707,N_8112,N_8902);
xnor U10708 (N_10708,N_8560,N_7526);
xnor U10709 (N_10709,N_6652,N_8343);
and U10710 (N_10710,N_7761,N_8668);
or U10711 (N_10711,N_6978,N_8027);
and U10712 (N_10712,N_8086,N_7557);
nand U10713 (N_10713,N_8803,N_8916);
nor U10714 (N_10714,N_7968,N_8014);
nand U10715 (N_10715,N_6464,N_7818);
nor U10716 (N_10716,N_7003,N_6383);
nand U10717 (N_10717,N_6402,N_8911);
or U10718 (N_10718,N_8400,N_8743);
nand U10719 (N_10719,N_8418,N_8525);
nor U10720 (N_10720,N_6817,N_7631);
xor U10721 (N_10721,N_6045,N_8129);
nor U10722 (N_10722,N_8760,N_6345);
and U10723 (N_10723,N_7803,N_7307);
nand U10724 (N_10724,N_7912,N_7994);
or U10725 (N_10725,N_8960,N_8170);
and U10726 (N_10726,N_7025,N_6046);
nand U10727 (N_10727,N_6534,N_7213);
and U10728 (N_10728,N_7884,N_6895);
nand U10729 (N_10729,N_7667,N_8337);
nor U10730 (N_10730,N_8456,N_6387);
nor U10731 (N_10731,N_6322,N_8636);
nand U10732 (N_10732,N_7585,N_8926);
and U10733 (N_10733,N_7633,N_8307);
nor U10734 (N_10734,N_8129,N_8580);
or U10735 (N_10735,N_8934,N_8142);
and U10736 (N_10736,N_8358,N_8481);
and U10737 (N_10737,N_7561,N_8974);
and U10738 (N_10738,N_6731,N_8185);
nor U10739 (N_10739,N_7180,N_8785);
nor U10740 (N_10740,N_6802,N_6804);
or U10741 (N_10741,N_7154,N_6963);
nand U10742 (N_10742,N_7565,N_7991);
xor U10743 (N_10743,N_8298,N_7428);
nand U10744 (N_10744,N_8953,N_6102);
and U10745 (N_10745,N_8399,N_8362);
and U10746 (N_10746,N_6566,N_6045);
and U10747 (N_10747,N_7695,N_6905);
nand U10748 (N_10748,N_6217,N_6811);
nand U10749 (N_10749,N_6141,N_6170);
and U10750 (N_10750,N_7131,N_7292);
xnor U10751 (N_10751,N_6851,N_6795);
or U10752 (N_10752,N_7942,N_6092);
xor U10753 (N_10753,N_8611,N_8680);
nand U10754 (N_10754,N_6496,N_8380);
or U10755 (N_10755,N_7232,N_6924);
nor U10756 (N_10756,N_7580,N_7175);
nor U10757 (N_10757,N_6232,N_8304);
or U10758 (N_10758,N_8559,N_7153);
or U10759 (N_10759,N_6240,N_6803);
nand U10760 (N_10760,N_6885,N_6797);
or U10761 (N_10761,N_7595,N_7824);
nor U10762 (N_10762,N_8689,N_7553);
nor U10763 (N_10763,N_7372,N_7300);
nor U10764 (N_10764,N_7036,N_7288);
or U10765 (N_10765,N_6524,N_8402);
and U10766 (N_10766,N_8346,N_7722);
nor U10767 (N_10767,N_7028,N_6866);
xnor U10768 (N_10768,N_7740,N_6425);
nor U10769 (N_10769,N_6847,N_6265);
and U10770 (N_10770,N_8855,N_7442);
xnor U10771 (N_10771,N_7019,N_6066);
and U10772 (N_10772,N_8085,N_6448);
or U10773 (N_10773,N_7858,N_7562);
and U10774 (N_10774,N_6966,N_8953);
nand U10775 (N_10775,N_6711,N_8124);
nor U10776 (N_10776,N_8583,N_6206);
and U10777 (N_10777,N_8689,N_6680);
xor U10778 (N_10778,N_6681,N_7446);
and U10779 (N_10779,N_6137,N_7395);
nand U10780 (N_10780,N_8974,N_8743);
xnor U10781 (N_10781,N_8136,N_6885);
or U10782 (N_10782,N_8548,N_6360);
nand U10783 (N_10783,N_8976,N_8746);
and U10784 (N_10784,N_7287,N_8809);
nand U10785 (N_10785,N_6206,N_8754);
and U10786 (N_10786,N_8094,N_6219);
nand U10787 (N_10787,N_7856,N_7947);
nand U10788 (N_10788,N_6472,N_6839);
and U10789 (N_10789,N_8916,N_6924);
xnor U10790 (N_10790,N_6034,N_8789);
nand U10791 (N_10791,N_7292,N_7441);
or U10792 (N_10792,N_7023,N_8768);
and U10793 (N_10793,N_8913,N_6154);
nand U10794 (N_10794,N_8009,N_6348);
nor U10795 (N_10795,N_6539,N_8584);
nand U10796 (N_10796,N_6574,N_7835);
nor U10797 (N_10797,N_6902,N_7490);
and U10798 (N_10798,N_6096,N_6710);
nand U10799 (N_10799,N_6745,N_7269);
or U10800 (N_10800,N_8768,N_6069);
and U10801 (N_10801,N_7656,N_7993);
nor U10802 (N_10802,N_6809,N_7734);
or U10803 (N_10803,N_8295,N_6691);
and U10804 (N_10804,N_7919,N_6293);
nand U10805 (N_10805,N_8500,N_7724);
or U10806 (N_10806,N_6226,N_6425);
nand U10807 (N_10807,N_7034,N_6159);
xnor U10808 (N_10808,N_7443,N_8504);
or U10809 (N_10809,N_7008,N_6424);
and U10810 (N_10810,N_7362,N_7540);
or U10811 (N_10811,N_8716,N_8926);
or U10812 (N_10812,N_7642,N_6331);
xnor U10813 (N_10813,N_8089,N_7632);
nand U10814 (N_10814,N_6021,N_6088);
nor U10815 (N_10815,N_8299,N_6917);
nand U10816 (N_10816,N_7015,N_8782);
and U10817 (N_10817,N_7851,N_6382);
nor U10818 (N_10818,N_8812,N_6206);
nand U10819 (N_10819,N_6503,N_6624);
or U10820 (N_10820,N_6867,N_7123);
or U10821 (N_10821,N_7746,N_7416);
and U10822 (N_10822,N_8086,N_6176);
or U10823 (N_10823,N_7156,N_6108);
and U10824 (N_10824,N_6443,N_8262);
xor U10825 (N_10825,N_6302,N_8290);
nand U10826 (N_10826,N_6640,N_7500);
nand U10827 (N_10827,N_6629,N_8167);
nor U10828 (N_10828,N_8921,N_6706);
nand U10829 (N_10829,N_6118,N_8975);
xnor U10830 (N_10830,N_7652,N_8948);
and U10831 (N_10831,N_6205,N_6846);
nor U10832 (N_10832,N_6373,N_6005);
nand U10833 (N_10833,N_7232,N_6124);
xnor U10834 (N_10834,N_7557,N_6737);
xnor U10835 (N_10835,N_7911,N_8174);
nor U10836 (N_10836,N_8381,N_6590);
or U10837 (N_10837,N_8743,N_7179);
nand U10838 (N_10838,N_8204,N_8928);
or U10839 (N_10839,N_6000,N_8038);
and U10840 (N_10840,N_7757,N_6817);
nand U10841 (N_10841,N_6334,N_7111);
nor U10842 (N_10842,N_7914,N_8051);
xor U10843 (N_10843,N_8781,N_7097);
and U10844 (N_10844,N_7685,N_7565);
and U10845 (N_10845,N_6898,N_7668);
nand U10846 (N_10846,N_6372,N_7626);
nor U10847 (N_10847,N_8316,N_8396);
nand U10848 (N_10848,N_7897,N_8601);
nand U10849 (N_10849,N_8233,N_8248);
and U10850 (N_10850,N_8751,N_6974);
and U10851 (N_10851,N_6219,N_6235);
nand U10852 (N_10852,N_8520,N_6736);
and U10853 (N_10853,N_8881,N_8817);
nand U10854 (N_10854,N_7551,N_8760);
and U10855 (N_10855,N_7627,N_6691);
nor U10856 (N_10856,N_6930,N_8737);
or U10857 (N_10857,N_6266,N_6880);
nand U10858 (N_10858,N_6962,N_8795);
and U10859 (N_10859,N_6564,N_8598);
nand U10860 (N_10860,N_7649,N_8476);
or U10861 (N_10861,N_7861,N_7195);
nand U10862 (N_10862,N_6646,N_6589);
nand U10863 (N_10863,N_6911,N_6045);
nand U10864 (N_10864,N_8669,N_8331);
and U10865 (N_10865,N_6261,N_6756);
and U10866 (N_10866,N_6556,N_8193);
or U10867 (N_10867,N_8243,N_7843);
nand U10868 (N_10868,N_6206,N_6081);
or U10869 (N_10869,N_6610,N_8702);
and U10870 (N_10870,N_6294,N_7268);
nor U10871 (N_10871,N_7590,N_6107);
nor U10872 (N_10872,N_7520,N_7286);
and U10873 (N_10873,N_6153,N_7956);
xnor U10874 (N_10874,N_6206,N_6990);
nand U10875 (N_10875,N_6425,N_8883);
xnor U10876 (N_10876,N_8181,N_8745);
or U10877 (N_10877,N_7011,N_7910);
and U10878 (N_10878,N_6512,N_6933);
and U10879 (N_10879,N_8085,N_7474);
and U10880 (N_10880,N_6853,N_8069);
nor U10881 (N_10881,N_6018,N_7246);
and U10882 (N_10882,N_7565,N_8679);
or U10883 (N_10883,N_7545,N_8271);
nor U10884 (N_10884,N_6382,N_7940);
or U10885 (N_10885,N_8569,N_6407);
and U10886 (N_10886,N_6834,N_6600);
nor U10887 (N_10887,N_6524,N_7742);
or U10888 (N_10888,N_6067,N_8039);
nand U10889 (N_10889,N_7714,N_6757);
and U10890 (N_10890,N_7486,N_7835);
and U10891 (N_10891,N_8217,N_6997);
nand U10892 (N_10892,N_6378,N_6930);
and U10893 (N_10893,N_6043,N_8895);
xor U10894 (N_10894,N_8028,N_7316);
nand U10895 (N_10895,N_6941,N_8036);
nor U10896 (N_10896,N_7838,N_6511);
xor U10897 (N_10897,N_6747,N_8009);
and U10898 (N_10898,N_6954,N_8911);
xor U10899 (N_10899,N_6093,N_8739);
or U10900 (N_10900,N_8810,N_6079);
and U10901 (N_10901,N_8682,N_7134);
nand U10902 (N_10902,N_8569,N_7626);
or U10903 (N_10903,N_6899,N_6033);
xnor U10904 (N_10904,N_8930,N_6941);
or U10905 (N_10905,N_7152,N_6498);
or U10906 (N_10906,N_8477,N_6071);
or U10907 (N_10907,N_8002,N_8965);
or U10908 (N_10908,N_7438,N_6835);
and U10909 (N_10909,N_8162,N_7012);
nand U10910 (N_10910,N_6580,N_8396);
nor U10911 (N_10911,N_7645,N_7526);
or U10912 (N_10912,N_8972,N_7383);
nand U10913 (N_10913,N_7537,N_8571);
or U10914 (N_10914,N_7217,N_7621);
nand U10915 (N_10915,N_6759,N_6444);
and U10916 (N_10916,N_8412,N_8859);
nor U10917 (N_10917,N_8202,N_6875);
nand U10918 (N_10918,N_6265,N_8197);
xnor U10919 (N_10919,N_8072,N_7056);
and U10920 (N_10920,N_6806,N_8134);
xnor U10921 (N_10921,N_7674,N_7827);
and U10922 (N_10922,N_7561,N_6969);
xnor U10923 (N_10923,N_6713,N_8159);
nand U10924 (N_10924,N_7167,N_7457);
nand U10925 (N_10925,N_8594,N_8664);
or U10926 (N_10926,N_8896,N_6379);
and U10927 (N_10927,N_6751,N_7717);
and U10928 (N_10928,N_6342,N_6157);
nor U10929 (N_10929,N_6172,N_6664);
or U10930 (N_10930,N_8614,N_7200);
or U10931 (N_10931,N_8268,N_8661);
xor U10932 (N_10932,N_7324,N_7284);
nand U10933 (N_10933,N_6132,N_7858);
or U10934 (N_10934,N_8006,N_6712);
nand U10935 (N_10935,N_7693,N_8918);
nand U10936 (N_10936,N_6240,N_6666);
or U10937 (N_10937,N_8612,N_8128);
nor U10938 (N_10938,N_8255,N_6495);
or U10939 (N_10939,N_6827,N_8804);
nor U10940 (N_10940,N_7684,N_7171);
and U10941 (N_10941,N_6947,N_8178);
nor U10942 (N_10942,N_8203,N_6967);
xnor U10943 (N_10943,N_7225,N_6634);
or U10944 (N_10944,N_6203,N_8535);
xor U10945 (N_10945,N_8519,N_7278);
and U10946 (N_10946,N_6479,N_7338);
and U10947 (N_10947,N_7112,N_6537);
nand U10948 (N_10948,N_6228,N_7028);
and U10949 (N_10949,N_8423,N_7754);
or U10950 (N_10950,N_6507,N_6056);
nand U10951 (N_10951,N_6959,N_7555);
or U10952 (N_10952,N_7649,N_7765);
nand U10953 (N_10953,N_6700,N_6113);
or U10954 (N_10954,N_6723,N_8032);
xor U10955 (N_10955,N_7970,N_8269);
nor U10956 (N_10956,N_8910,N_7063);
nor U10957 (N_10957,N_7482,N_8705);
xor U10958 (N_10958,N_6387,N_7496);
nand U10959 (N_10959,N_7008,N_6793);
and U10960 (N_10960,N_8929,N_6615);
xor U10961 (N_10961,N_6960,N_8710);
or U10962 (N_10962,N_7881,N_6620);
nor U10963 (N_10963,N_8145,N_6603);
and U10964 (N_10964,N_7327,N_7144);
or U10965 (N_10965,N_6053,N_8892);
or U10966 (N_10966,N_6187,N_7284);
nand U10967 (N_10967,N_6591,N_6316);
and U10968 (N_10968,N_6604,N_6805);
nand U10969 (N_10969,N_7565,N_6812);
and U10970 (N_10970,N_8614,N_8841);
nand U10971 (N_10971,N_8258,N_7179);
nand U10972 (N_10972,N_6920,N_6251);
and U10973 (N_10973,N_7075,N_7184);
or U10974 (N_10974,N_7775,N_8795);
nor U10975 (N_10975,N_7134,N_7852);
nand U10976 (N_10976,N_6169,N_8313);
or U10977 (N_10977,N_8072,N_8408);
or U10978 (N_10978,N_8491,N_7201);
and U10979 (N_10979,N_6699,N_8969);
nand U10980 (N_10980,N_7972,N_7683);
or U10981 (N_10981,N_8736,N_6311);
nor U10982 (N_10982,N_8693,N_7309);
nand U10983 (N_10983,N_6054,N_8423);
or U10984 (N_10984,N_6457,N_8750);
nand U10985 (N_10985,N_8372,N_7027);
or U10986 (N_10986,N_7649,N_8247);
nand U10987 (N_10987,N_6741,N_8230);
nand U10988 (N_10988,N_7959,N_8293);
xnor U10989 (N_10989,N_6901,N_7653);
xnor U10990 (N_10990,N_8531,N_8749);
or U10991 (N_10991,N_8362,N_7072);
or U10992 (N_10992,N_7588,N_6754);
xor U10993 (N_10993,N_7622,N_7681);
nand U10994 (N_10994,N_8987,N_8830);
xnor U10995 (N_10995,N_8110,N_8682);
or U10996 (N_10996,N_7706,N_7400);
and U10997 (N_10997,N_6903,N_6984);
nor U10998 (N_10998,N_8524,N_6939);
nor U10999 (N_10999,N_7608,N_7049);
nand U11000 (N_11000,N_8334,N_6041);
and U11001 (N_11001,N_7432,N_6779);
nand U11002 (N_11002,N_6222,N_6975);
nor U11003 (N_11003,N_7386,N_8638);
and U11004 (N_11004,N_6538,N_7323);
nand U11005 (N_11005,N_7549,N_8140);
and U11006 (N_11006,N_7766,N_6942);
and U11007 (N_11007,N_6384,N_7231);
and U11008 (N_11008,N_6747,N_6680);
xnor U11009 (N_11009,N_6585,N_6142);
and U11010 (N_11010,N_7645,N_6310);
nor U11011 (N_11011,N_8779,N_8325);
nor U11012 (N_11012,N_7197,N_6728);
nand U11013 (N_11013,N_8840,N_7701);
nand U11014 (N_11014,N_7383,N_6362);
nand U11015 (N_11015,N_6875,N_7585);
or U11016 (N_11016,N_6142,N_8940);
or U11017 (N_11017,N_7671,N_7972);
or U11018 (N_11018,N_8413,N_8220);
nor U11019 (N_11019,N_7850,N_7151);
nand U11020 (N_11020,N_7940,N_8697);
or U11021 (N_11021,N_6843,N_8653);
xor U11022 (N_11022,N_8125,N_8435);
or U11023 (N_11023,N_6002,N_6531);
nor U11024 (N_11024,N_8693,N_8471);
xnor U11025 (N_11025,N_6283,N_7376);
nand U11026 (N_11026,N_6962,N_7705);
or U11027 (N_11027,N_8222,N_6838);
and U11028 (N_11028,N_8803,N_7881);
or U11029 (N_11029,N_6762,N_8216);
nor U11030 (N_11030,N_8313,N_6380);
and U11031 (N_11031,N_6892,N_8840);
nor U11032 (N_11032,N_8909,N_7831);
xnor U11033 (N_11033,N_7570,N_8858);
nand U11034 (N_11034,N_8654,N_8684);
and U11035 (N_11035,N_6941,N_7402);
nor U11036 (N_11036,N_8936,N_8468);
or U11037 (N_11037,N_8825,N_7418);
or U11038 (N_11038,N_6497,N_8468);
nor U11039 (N_11039,N_7546,N_8155);
and U11040 (N_11040,N_7159,N_6728);
nor U11041 (N_11041,N_8675,N_7252);
xor U11042 (N_11042,N_7267,N_8298);
or U11043 (N_11043,N_8721,N_8425);
nand U11044 (N_11044,N_7561,N_8556);
or U11045 (N_11045,N_6628,N_6040);
nand U11046 (N_11046,N_7695,N_6334);
xor U11047 (N_11047,N_6902,N_8152);
or U11048 (N_11048,N_6034,N_6429);
and U11049 (N_11049,N_7363,N_7860);
nor U11050 (N_11050,N_7492,N_6257);
or U11051 (N_11051,N_8169,N_8156);
or U11052 (N_11052,N_7349,N_7319);
nor U11053 (N_11053,N_6365,N_7210);
and U11054 (N_11054,N_7730,N_7558);
nand U11055 (N_11055,N_6869,N_8446);
xnor U11056 (N_11056,N_8524,N_7248);
or U11057 (N_11057,N_8096,N_7394);
nor U11058 (N_11058,N_7188,N_7042);
nand U11059 (N_11059,N_7948,N_6876);
nor U11060 (N_11060,N_6147,N_6732);
xor U11061 (N_11061,N_6406,N_6924);
nor U11062 (N_11062,N_6946,N_8748);
or U11063 (N_11063,N_6218,N_6616);
and U11064 (N_11064,N_6561,N_6698);
or U11065 (N_11065,N_8164,N_7718);
xnor U11066 (N_11066,N_6983,N_7194);
nand U11067 (N_11067,N_8232,N_7499);
and U11068 (N_11068,N_8405,N_6953);
nand U11069 (N_11069,N_7676,N_7650);
and U11070 (N_11070,N_7263,N_6207);
nand U11071 (N_11071,N_6616,N_6630);
or U11072 (N_11072,N_7043,N_6372);
nand U11073 (N_11073,N_8445,N_7547);
and U11074 (N_11074,N_7248,N_8523);
nand U11075 (N_11075,N_8856,N_6185);
nor U11076 (N_11076,N_6936,N_6327);
xnor U11077 (N_11077,N_8942,N_7204);
or U11078 (N_11078,N_8740,N_8647);
xor U11079 (N_11079,N_8796,N_6438);
and U11080 (N_11080,N_7535,N_8704);
or U11081 (N_11081,N_8220,N_6826);
nand U11082 (N_11082,N_7957,N_6664);
nand U11083 (N_11083,N_7353,N_6718);
nor U11084 (N_11084,N_6758,N_7011);
nor U11085 (N_11085,N_8455,N_8637);
nand U11086 (N_11086,N_8790,N_6599);
nand U11087 (N_11087,N_6244,N_6100);
and U11088 (N_11088,N_6805,N_8443);
and U11089 (N_11089,N_8387,N_8514);
nand U11090 (N_11090,N_8600,N_7683);
or U11091 (N_11091,N_8638,N_8937);
or U11092 (N_11092,N_7844,N_8826);
nor U11093 (N_11093,N_8964,N_7160);
and U11094 (N_11094,N_6406,N_6733);
xnor U11095 (N_11095,N_8579,N_7212);
and U11096 (N_11096,N_8118,N_8797);
and U11097 (N_11097,N_8335,N_7350);
or U11098 (N_11098,N_8129,N_8893);
nand U11099 (N_11099,N_6482,N_6274);
xnor U11100 (N_11100,N_6640,N_6077);
nor U11101 (N_11101,N_6572,N_8447);
nand U11102 (N_11102,N_6954,N_7045);
nand U11103 (N_11103,N_6347,N_6446);
or U11104 (N_11104,N_7180,N_7624);
xor U11105 (N_11105,N_7973,N_6280);
or U11106 (N_11106,N_8384,N_6986);
nor U11107 (N_11107,N_6056,N_6525);
nor U11108 (N_11108,N_8498,N_6212);
or U11109 (N_11109,N_6343,N_8402);
and U11110 (N_11110,N_7965,N_6591);
and U11111 (N_11111,N_7595,N_6925);
xor U11112 (N_11112,N_8095,N_8993);
nor U11113 (N_11113,N_8417,N_6502);
and U11114 (N_11114,N_8829,N_7515);
xnor U11115 (N_11115,N_7613,N_8390);
nor U11116 (N_11116,N_6582,N_6423);
nand U11117 (N_11117,N_6642,N_6678);
or U11118 (N_11118,N_8120,N_7989);
or U11119 (N_11119,N_6494,N_7243);
and U11120 (N_11120,N_8126,N_7614);
and U11121 (N_11121,N_6665,N_6447);
nand U11122 (N_11122,N_8063,N_8579);
xnor U11123 (N_11123,N_6721,N_6510);
nand U11124 (N_11124,N_7088,N_7239);
or U11125 (N_11125,N_8012,N_6189);
nand U11126 (N_11126,N_8758,N_6131);
nand U11127 (N_11127,N_7547,N_7666);
and U11128 (N_11128,N_7053,N_6787);
nand U11129 (N_11129,N_8008,N_8868);
nand U11130 (N_11130,N_6193,N_7147);
nand U11131 (N_11131,N_7301,N_7683);
and U11132 (N_11132,N_8006,N_8934);
nand U11133 (N_11133,N_8909,N_6620);
or U11134 (N_11134,N_7231,N_8474);
and U11135 (N_11135,N_7003,N_7632);
nor U11136 (N_11136,N_8187,N_8370);
nand U11137 (N_11137,N_6027,N_8102);
nor U11138 (N_11138,N_6564,N_8305);
nand U11139 (N_11139,N_6523,N_8338);
nand U11140 (N_11140,N_6930,N_7093);
and U11141 (N_11141,N_6125,N_7336);
nor U11142 (N_11142,N_8661,N_6542);
and U11143 (N_11143,N_8869,N_7432);
and U11144 (N_11144,N_7246,N_8108);
nor U11145 (N_11145,N_8522,N_7432);
xnor U11146 (N_11146,N_8818,N_6167);
nand U11147 (N_11147,N_7755,N_6361);
nor U11148 (N_11148,N_6865,N_8291);
nand U11149 (N_11149,N_8929,N_6108);
and U11150 (N_11150,N_8582,N_7260);
nor U11151 (N_11151,N_6049,N_8176);
nand U11152 (N_11152,N_7061,N_8754);
nand U11153 (N_11153,N_7615,N_8982);
nor U11154 (N_11154,N_6709,N_6416);
nor U11155 (N_11155,N_6465,N_8656);
and U11156 (N_11156,N_7024,N_8600);
xnor U11157 (N_11157,N_6916,N_6815);
and U11158 (N_11158,N_7229,N_6393);
nand U11159 (N_11159,N_8797,N_6468);
nor U11160 (N_11160,N_7874,N_7512);
nand U11161 (N_11161,N_6121,N_8112);
xnor U11162 (N_11162,N_7237,N_8960);
or U11163 (N_11163,N_8678,N_6874);
or U11164 (N_11164,N_8100,N_7259);
xor U11165 (N_11165,N_7327,N_8267);
nand U11166 (N_11166,N_6990,N_8707);
nand U11167 (N_11167,N_8931,N_8884);
xor U11168 (N_11168,N_8032,N_6885);
nand U11169 (N_11169,N_8744,N_8003);
xor U11170 (N_11170,N_7079,N_7395);
and U11171 (N_11171,N_7770,N_8775);
and U11172 (N_11172,N_8688,N_8622);
nand U11173 (N_11173,N_8490,N_6706);
nand U11174 (N_11174,N_8581,N_7527);
and U11175 (N_11175,N_8189,N_7676);
or U11176 (N_11176,N_7298,N_7255);
nor U11177 (N_11177,N_8514,N_7269);
nand U11178 (N_11178,N_6793,N_8576);
and U11179 (N_11179,N_6860,N_8654);
nor U11180 (N_11180,N_7199,N_8202);
or U11181 (N_11181,N_7751,N_8202);
nor U11182 (N_11182,N_6248,N_7228);
nand U11183 (N_11183,N_6514,N_8134);
xor U11184 (N_11184,N_6217,N_8623);
xnor U11185 (N_11185,N_8026,N_8278);
or U11186 (N_11186,N_8306,N_7753);
and U11187 (N_11187,N_7983,N_6787);
nand U11188 (N_11188,N_8240,N_6318);
nor U11189 (N_11189,N_7121,N_8247);
nor U11190 (N_11190,N_7133,N_7103);
nor U11191 (N_11191,N_7078,N_6441);
and U11192 (N_11192,N_8809,N_7335);
and U11193 (N_11193,N_7010,N_7829);
and U11194 (N_11194,N_8853,N_8158);
xnor U11195 (N_11195,N_6522,N_8550);
and U11196 (N_11196,N_8928,N_7461);
and U11197 (N_11197,N_8322,N_7725);
or U11198 (N_11198,N_6621,N_8173);
and U11199 (N_11199,N_6836,N_8441);
or U11200 (N_11200,N_7665,N_7233);
nor U11201 (N_11201,N_7983,N_7281);
or U11202 (N_11202,N_6100,N_8670);
nand U11203 (N_11203,N_7270,N_6188);
nor U11204 (N_11204,N_6877,N_7592);
nor U11205 (N_11205,N_6246,N_6477);
or U11206 (N_11206,N_6228,N_6560);
or U11207 (N_11207,N_7629,N_7011);
and U11208 (N_11208,N_8549,N_6901);
and U11209 (N_11209,N_8159,N_7770);
nand U11210 (N_11210,N_7874,N_8997);
or U11211 (N_11211,N_7158,N_7668);
and U11212 (N_11212,N_7571,N_8074);
and U11213 (N_11213,N_8643,N_8883);
or U11214 (N_11214,N_8291,N_7397);
or U11215 (N_11215,N_6163,N_6801);
nand U11216 (N_11216,N_7114,N_7489);
nand U11217 (N_11217,N_8073,N_8957);
nand U11218 (N_11218,N_6399,N_7219);
nor U11219 (N_11219,N_8250,N_8802);
nand U11220 (N_11220,N_6040,N_6112);
and U11221 (N_11221,N_7419,N_7093);
and U11222 (N_11222,N_8576,N_7699);
nor U11223 (N_11223,N_6287,N_8102);
nand U11224 (N_11224,N_8425,N_7684);
and U11225 (N_11225,N_7680,N_7717);
nand U11226 (N_11226,N_8578,N_7198);
or U11227 (N_11227,N_7001,N_7499);
nand U11228 (N_11228,N_8905,N_7229);
nor U11229 (N_11229,N_6975,N_7547);
nand U11230 (N_11230,N_8444,N_7296);
and U11231 (N_11231,N_8917,N_6431);
or U11232 (N_11232,N_6078,N_8186);
nor U11233 (N_11233,N_7258,N_6728);
or U11234 (N_11234,N_7546,N_6001);
nor U11235 (N_11235,N_6601,N_6094);
and U11236 (N_11236,N_8096,N_6016);
nor U11237 (N_11237,N_6775,N_6810);
or U11238 (N_11238,N_6819,N_8080);
and U11239 (N_11239,N_7823,N_6238);
and U11240 (N_11240,N_6086,N_6746);
nand U11241 (N_11241,N_6228,N_8825);
nand U11242 (N_11242,N_7398,N_8125);
and U11243 (N_11243,N_8731,N_8578);
or U11244 (N_11244,N_7845,N_7019);
xnor U11245 (N_11245,N_8440,N_6103);
and U11246 (N_11246,N_6444,N_7013);
nor U11247 (N_11247,N_8795,N_7481);
nand U11248 (N_11248,N_8603,N_7365);
nand U11249 (N_11249,N_7655,N_7187);
and U11250 (N_11250,N_6874,N_6404);
nand U11251 (N_11251,N_8497,N_7932);
or U11252 (N_11252,N_6487,N_8073);
and U11253 (N_11253,N_7344,N_7223);
or U11254 (N_11254,N_7738,N_8686);
or U11255 (N_11255,N_7408,N_6557);
or U11256 (N_11256,N_6169,N_6694);
or U11257 (N_11257,N_6872,N_8964);
and U11258 (N_11258,N_8988,N_8877);
nand U11259 (N_11259,N_7326,N_6918);
and U11260 (N_11260,N_6435,N_8346);
nor U11261 (N_11261,N_7573,N_8244);
xor U11262 (N_11262,N_8163,N_6963);
or U11263 (N_11263,N_6554,N_6037);
or U11264 (N_11264,N_8319,N_6274);
nor U11265 (N_11265,N_6542,N_6954);
nor U11266 (N_11266,N_7323,N_8725);
nor U11267 (N_11267,N_8863,N_6991);
nand U11268 (N_11268,N_8141,N_7353);
nor U11269 (N_11269,N_8320,N_8098);
nand U11270 (N_11270,N_7996,N_7089);
and U11271 (N_11271,N_8466,N_8387);
and U11272 (N_11272,N_6574,N_7866);
nor U11273 (N_11273,N_7089,N_8766);
and U11274 (N_11274,N_6601,N_6494);
nor U11275 (N_11275,N_7392,N_6839);
and U11276 (N_11276,N_8070,N_6188);
nor U11277 (N_11277,N_6707,N_6173);
nor U11278 (N_11278,N_6926,N_8984);
and U11279 (N_11279,N_6600,N_7652);
nand U11280 (N_11280,N_6261,N_7710);
and U11281 (N_11281,N_7072,N_8872);
nand U11282 (N_11282,N_7419,N_8087);
or U11283 (N_11283,N_6870,N_7155);
nand U11284 (N_11284,N_8585,N_8780);
nor U11285 (N_11285,N_7152,N_6775);
nand U11286 (N_11286,N_6018,N_6835);
nand U11287 (N_11287,N_6144,N_6558);
xor U11288 (N_11288,N_6095,N_7421);
or U11289 (N_11289,N_6040,N_7546);
nand U11290 (N_11290,N_7869,N_8814);
nor U11291 (N_11291,N_6988,N_6394);
and U11292 (N_11292,N_8101,N_7286);
and U11293 (N_11293,N_7996,N_7330);
nand U11294 (N_11294,N_6929,N_8798);
nand U11295 (N_11295,N_7889,N_6255);
nor U11296 (N_11296,N_7122,N_6131);
nand U11297 (N_11297,N_7225,N_8971);
xnor U11298 (N_11298,N_6411,N_8795);
or U11299 (N_11299,N_8824,N_7963);
or U11300 (N_11300,N_6802,N_8240);
nand U11301 (N_11301,N_7528,N_6996);
nor U11302 (N_11302,N_6430,N_7956);
xor U11303 (N_11303,N_8057,N_7109);
nand U11304 (N_11304,N_8404,N_6686);
and U11305 (N_11305,N_8049,N_8504);
and U11306 (N_11306,N_7966,N_8068);
and U11307 (N_11307,N_7025,N_6606);
or U11308 (N_11308,N_8923,N_8817);
or U11309 (N_11309,N_7844,N_7242);
nor U11310 (N_11310,N_8049,N_8832);
nor U11311 (N_11311,N_8290,N_8722);
nand U11312 (N_11312,N_7780,N_7087);
nor U11313 (N_11313,N_8032,N_8869);
or U11314 (N_11314,N_7824,N_6724);
and U11315 (N_11315,N_6159,N_6709);
or U11316 (N_11316,N_6392,N_8173);
and U11317 (N_11317,N_6603,N_6277);
or U11318 (N_11318,N_6807,N_6341);
and U11319 (N_11319,N_6907,N_7200);
or U11320 (N_11320,N_6685,N_7403);
nor U11321 (N_11321,N_8352,N_7691);
nand U11322 (N_11322,N_6720,N_7580);
nor U11323 (N_11323,N_8875,N_7999);
and U11324 (N_11324,N_7334,N_6798);
nor U11325 (N_11325,N_6669,N_6781);
and U11326 (N_11326,N_6063,N_8746);
nor U11327 (N_11327,N_7097,N_7685);
nand U11328 (N_11328,N_6407,N_6572);
and U11329 (N_11329,N_8891,N_6662);
and U11330 (N_11330,N_6417,N_8214);
and U11331 (N_11331,N_8247,N_8457);
nand U11332 (N_11332,N_8241,N_8148);
or U11333 (N_11333,N_8648,N_8767);
nand U11334 (N_11334,N_6986,N_6879);
and U11335 (N_11335,N_6088,N_8651);
nor U11336 (N_11336,N_8996,N_6641);
xnor U11337 (N_11337,N_7604,N_8141);
xnor U11338 (N_11338,N_8106,N_6974);
nand U11339 (N_11339,N_7716,N_6219);
xnor U11340 (N_11340,N_8456,N_6211);
xnor U11341 (N_11341,N_8784,N_8168);
or U11342 (N_11342,N_7310,N_6338);
nor U11343 (N_11343,N_7563,N_7189);
and U11344 (N_11344,N_6289,N_6445);
and U11345 (N_11345,N_7186,N_6667);
nor U11346 (N_11346,N_6545,N_8124);
and U11347 (N_11347,N_7018,N_8087);
nor U11348 (N_11348,N_7759,N_8794);
nand U11349 (N_11349,N_8007,N_7394);
nor U11350 (N_11350,N_6379,N_7087);
and U11351 (N_11351,N_6743,N_8160);
xor U11352 (N_11352,N_8377,N_7677);
nand U11353 (N_11353,N_7513,N_6909);
nand U11354 (N_11354,N_6013,N_6247);
or U11355 (N_11355,N_7839,N_8314);
and U11356 (N_11356,N_6528,N_6920);
nand U11357 (N_11357,N_8566,N_7638);
nor U11358 (N_11358,N_8261,N_6029);
xnor U11359 (N_11359,N_8254,N_6719);
nor U11360 (N_11360,N_7825,N_7892);
nor U11361 (N_11361,N_6682,N_8013);
and U11362 (N_11362,N_7496,N_6214);
nor U11363 (N_11363,N_6496,N_8503);
nand U11364 (N_11364,N_7457,N_8531);
nand U11365 (N_11365,N_8860,N_7893);
nand U11366 (N_11366,N_8668,N_6809);
nor U11367 (N_11367,N_7007,N_8588);
and U11368 (N_11368,N_7086,N_7451);
or U11369 (N_11369,N_7240,N_6717);
or U11370 (N_11370,N_6556,N_7890);
or U11371 (N_11371,N_6776,N_7537);
or U11372 (N_11372,N_8887,N_7697);
xor U11373 (N_11373,N_6416,N_6701);
and U11374 (N_11374,N_6876,N_8221);
nor U11375 (N_11375,N_8559,N_6843);
xor U11376 (N_11376,N_6031,N_6491);
and U11377 (N_11377,N_8775,N_7519);
or U11378 (N_11378,N_6653,N_8502);
and U11379 (N_11379,N_8896,N_6250);
and U11380 (N_11380,N_8728,N_7236);
nand U11381 (N_11381,N_6367,N_8682);
and U11382 (N_11382,N_7227,N_6115);
xor U11383 (N_11383,N_7783,N_7048);
nand U11384 (N_11384,N_6699,N_8072);
and U11385 (N_11385,N_6098,N_6664);
and U11386 (N_11386,N_6121,N_7164);
or U11387 (N_11387,N_7542,N_8604);
or U11388 (N_11388,N_7861,N_8802);
and U11389 (N_11389,N_8999,N_7991);
nand U11390 (N_11390,N_7839,N_8988);
or U11391 (N_11391,N_8697,N_7231);
and U11392 (N_11392,N_6665,N_7274);
and U11393 (N_11393,N_8090,N_6984);
or U11394 (N_11394,N_7789,N_6269);
nand U11395 (N_11395,N_7707,N_7934);
or U11396 (N_11396,N_8505,N_6824);
nand U11397 (N_11397,N_7391,N_6735);
or U11398 (N_11398,N_6850,N_6072);
and U11399 (N_11399,N_7466,N_8112);
or U11400 (N_11400,N_8124,N_8434);
nor U11401 (N_11401,N_8494,N_7392);
nand U11402 (N_11402,N_7130,N_7502);
nand U11403 (N_11403,N_7913,N_6954);
nand U11404 (N_11404,N_6386,N_6791);
nand U11405 (N_11405,N_8540,N_7479);
nand U11406 (N_11406,N_6242,N_7635);
or U11407 (N_11407,N_7021,N_7720);
and U11408 (N_11408,N_6082,N_7689);
nor U11409 (N_11409,N_8140,N_7734);
or U11410 (N_11410,N_8411,N_7587);
nand U11411 (N_11411,N_6399,N_8424);
nor U11412 (N_11412,N_7522,N_8360);
or U11413 (N_11413,N_7535,N_8898);
and U11414 (N_11414,N_7946,N_7617);
and U11415 (N_11415,N_6903,N_8565);
nand U11416 (N_11416,N_6568,N_8950);
xnor U11417 (N_11417,N_6811,N_6588);
nor U11418 (N_11418,N_8679,N_8618);
or U11419 (N_11419,N_7712,N_8470);
and U11420 (N_11420,N_7080,N_8255);
or U11421 (N_11421,N_8656,N_6529);
nor U11422 (N_11422,N_6554,N_8087);
xnor U11423 (N_11423,N_7992,N_6506);
and U11424 (N_11424,N_8453,N_7931);
or U11425 (N_11425,N_8450,N_7000);
and U11426 (N_11426,N_6519,N_7169);
xor U11427 (N_11427,N_7085,N_8786);
and U11428 (N_11428,N_8937,N_6139);
and U11429 (N_11429,N_6239,N_7328);
and U11430 (N_11430,N_8679,N_7991);
or U11431 (N_11431,N_8767,N_6597);
nand U11432 (N_11432,N_7160,N_8280);
xnor U11433 (N_11433,N_8647,N_7849);
nand U11434 (N_11434,N_7426,N_7507);
and U11435 (N_11435,N_8871,N_8638);
nand U11436 (N_11436,N_8149,N_6375);
xnor U11437 (N_11437,N_8083,N_8805);
nor U11438 (N_11438,N_6361,N_8611);
or U11439 (N_11439,N_7532,N_8199);
and U11440 (N_11440,N_7620,N_6258);
or U11441 (N_11441,N_6805,N_8836);
or U11442 (N_11442,N_6431,N_7389);
nand U11443 (N_11443,N_8070,N_6348);
and U11444 (N_11444,N_6481,N_7379);
or U11445 (N_11445,N_8305,N_6388);
and U11446 (N_11446,N_6902,N_8316);
or U11447 (N_11447,N_6682,N_7094);
or U11448 (N_11448,N_6446,N_6890);
and U11449 (N_11449,N_8812,N_7804);
xor U11450 (N_11450,N_6669,N_8521);
nor U11451 (N_11451,N_6653,N_6152);
nor U11452 (N_11452,N_8778,N_8883);
and U11453 (N_11453,N_7946,N_7805);
nor U11454 (N_11454,N_8620,N_8129);
xor U11455 (N_11455,N_7955,N_8909);
nor U11456 (N_11456,N_6086,N_8186);
nand U11457 (N_11457,N_6579,N_6955);
and U11458 (N_11458,N_8096,N_6623);
nand U11459 (N_11459,N_7239,N_8631);
nor U11460 (N_11460,N_6965,N_8799);
nand U11461 (N_11461,N_6823,N_7144);
or U11462 (N_11462,N_7648,N_8825);
or U11463 (N_11463,N_8148,N_8431);
nor U11464 (N_11464,N_6603,N_7407);
nor U11465 (N_11465,N_8821,N_7132);
or U11466 (N_11466,N_7527,N_6116);
nand U11467 (N_11467,N_8491,N_6723);
nor U11468 (N_11468,N_8221,N_6029);
and U11469 (N_11469,N_7754,N_6737);
and U11470 (N_11470,N_8802,N_8565);
or U11471 (N_11471,N_7508,N_6312);
and U11472 (N_11472,N_6501,N_7957);
nand U11473 (N_11473,N_7912,N_6260);
or U11474 (N_11474,N_7279,N_8945);
and U11475 (N_11475,N_6959,N_7409);
nand U11476 (N_11476,N_8822,N_6123);
xnor U11477 (N_11477,N_6973,N_8238);
or U11478 (N_11478,N_6474,N_6779);
nor U11479 (N_11479,N_8520,N_8549);
and U11480 (N_11480,N_6799,N_6780);
nand U11481 (N_11481,N_8725,N_7136);
nand U11482 (N_11482,N_8344,N_6368);
nor U11483 (N_11483,N_6762,N_6913);
nand U11484 (N_11484,N_8161,N_7910);
nor U11485 (N_11485,N_7061,N_6455);
or U11486 (N_11486,N_7940,N_7634);
xnor U11487 (N_11487,N_8839,N_7237);
and U11488 (N_11488,N_7468,N_7815);
nor U11489 (N_11489,N_6092,N_7335);
nand U11490 (N_11490,N_7170,N_6636);
nor U11491 (N_11491,N_7916,N_8145);
and U11492 (N_11492,N_6650,N_7307);
and U11493 (N_11493,N_6689,N_8249);
and U11494 (N_11494,N_8908,N_6381);
nor U11495 (N_11495,N_6839,N_6451);
nor U11496 (N_11496,N_6697,N_8772);
nand U11497 (N_11497,N_8839,N_6730);
and U11498 (N_11498,N_8666,N_7162);
nand U11499 (N_11499,N_8346,N_7199);
nand U11500 (N_11500,N_6357,N_8323);
or U11501 (N_11501,N_8252,N_6574);
xor U11502 (N_11502,N_7435,N_6954);
nor U11503 (N_11503,N_8891,N_8340);
nor U11504 (N_11504,N_8009,N_7482);
and U11505 (N_11505,N_6324,N_6288);
nor U11506 (N_11506,N_8795,N_7735);
xor U11507 (N_11507,N_7171,N_7524);
nand U11508 (N_11508,N_8750,N_7992);
and U11509 (N_11509,N_8103,N_8800);
and U11510 (N_11510,N_8338,N_6325);
or U11511 (N_11511,N_8496,N_6379);
xnor U11512 (N_11512,N_7738,N_6305);
or U11513 (N_11513,N_6903,N_6988);
xnor U11514 (N_11514,N_6618,N_6961);
nor U11515 (N_11515,N_7409,N_6949);
or U11516 (N_11516,N_7008,N_6534);
and U11517 (N_11517,N_6686,N_7711);
nor U11518 (N_11518,N_6815,N_7325);
nor U11519 (N_11519,N_7615,N_7107);
or U11520 (N_11520,N_7666,N_7746);
or U11521 (N_11521,N_6446,N_6709);
and U11522 (N_11522,N_6362,N_8903);
and U11523 (N_11523,N_6671,N_8263);
or U11524 (N_11524,N_7478,N_6923);
nand U11525 (N_11525,N_8060,N_8348);
or U11526 (N_11526,N_6458,N_6428);
nor U11527 (N_11527,N_6790,N_8048);
nand U11528 (N_11528,N_6391,N_6311);
nor U11529 (N_11529,N_8417,N_7195);
and U11530 (N_11530,N_6748,N_6975);
nor U11531 (N_11531,N_7935,N_7271);
and U11532 (N_11532,N_6184,N_8220);
and U11533 (N_11533,N_7792,N_6690);
and U11534 (N_11534,N_6212,N_7911);
nor U11535 (N_11535,N_8295,N_8181);
and U11536 (N_11536,N_8252,N_6514);
and U11537 (N_11537,N_8387,N_8177);
nand U11538 (N_11538,N_8721,N_8799);
xnor U11539 (N_11539,N_8261,N_7348);
nand U11540 (N_11540,N_7389,N_6421);
or U11541 (N_11541,N_6811,N_7182);
or U11542 (N_11542,N_7919,N_7469);
and U11543 (N_11543,N_7686,N_8212);
and U11544 (N_11544,N_8226,N_7418);
and U11545 (N_11545,N_8846,N_7728);
and U11546 (N_11546,N_7326,N_7919);
or U11547 (N_11547,N_6351,N_7716);
nor U11548 (N_11548,N_8570,N_8996);
nand U11549 (N_11549,N_7415,N_6875);
or U11550 (N_11550,N_6343,N_7430);
nand U11551 (N_11551,N_8120,N_8938);
nand U11552 (N_11552,N_8943,N_7629);
nand U11553 (N_11553,N_6527,N_7579);
nand U11554 (N_11554,N_6867,N_7942);
and U11555 (N_11555,N_6991,N_7122);
nand U11556 (N_11556,N_8109,N_7588);
and U11557 (N_11557,N_6553,N_7694);
and U11558 (N_11558,N_6369,N_8874);
nor U11559 (N_11559,N_7869,N_8575);
or U11560 (N_11560,N_8581,N_6414);
or U11561 (N_11561,N_8375,N_6126);
or U11562 (N_11562,N_8470,N_8800);
or U11563 (N_11563,N_7728,N_8644);
nand U11564 (N_11564,N_7694,N_6488);
and U11565 (N_11565,N_7519,N_7151);
nor U11566 (N_11566,N_8149,N_8339);
nand U11567 (N_11567,N_6923,N_7346);
or U11568 (N_11568,N_8793,N_6066);
nor U11569 (N_11569,N_8226,N_8316);
nand U11570 (N_11570,N_6616,N_8329);
and U11571 (N_11571,N_6202,N_7424);
nor U11572 (N_11572,N_6700,N_6018);
nor U11573 (N_11573,N_7755,N_8135);
xor U11574 (N_11574,N_7183,N_6908);
and U11575 (N_11575,N_6066,N_7416);
nor U11576 (N_11576,N_6765,N_8568);
or U11577 (N_11577,N_6689,N_7760);
nand U11578 (N_11578,N_8398,N_7413);
xnor U11579 (N_11579,N_7884,N_7744);
nand U11580 (N_11580,N_8701,N_6798);
and U11581 (N_11581,N_8584,N_8357);
and U11582 (N_11582,N_8410,N_6861);
or U11583 (N_11583,N_7422,N_6650);
and U11584 (N_11584,N_8694,N_7060);
or U11585 (N_11585,N_7278,N_7058);
or U11586 (N_11586,N_7816,N_8410);
nor U11587 (N_11587,N_7549,N_6510);
and U11588 (N_11588,N_7181,N_8801);
xnor U11589 (N_11589,N_6171,N_6805);
and U11590 (N_11590,N_8432,N_6236);
nor U11591 (N_11591,N_8503,N_8474);
nor U11592 (N_11592,N_8708,N_7081);
or U11593 (N_11593,N_6369,N_8326);
nor U11594 (N_11594,N_8149,N_8089);
and U11595 (N_11595,N_6606,N_6863);
and U11596 (N_11596,N_6677,N_6086);
or U11597 (N_11597,N_6134,N_6657);
nor U11598 (N_11598,N_7080,N_6800);
and U11599 (N_11599,N_6045,N_8888);
or U11600 (N_11600,N_7547,N_6892);
or U11601 (N_11601,N_6135,N_7725);
nor U11602 (N_11602,N_7146,N_7086);
xnor U11603 (N_11603,N_8583,N_7284);
nor U11604 (N_11604,N_8032,N_6287);
and U11605 (N_11605,N_7717,N_6086);
nand U11606 (N_11606,N_8430,N_6405);
nor U11607 (N_11607,N_8151,N_6224);
and U11608 (N_11608,N_8393,N_7888);
nor U11609 (N_11609,N_6050,N_7642);
and U11610 (N_11610,N_8447,N_8089);
nor U11611 (N_11611,N_6104,N_7345);
or U11612 (N_11612,N_7699,N_7776);
nand U11613 (N_11613,N_8297,N_7111);
and U11614 (N_11614,N_6622,N_8189);
or U11615 (N_11615,N_6818,N_8347);
and U11616 (N_11616,N_6535,N_7618);
or U11617 (N_11617,N_8438,N_6105);
and U11618 (N_11618,N_6518,N_7458);
or U11619 (N_11619,N_8000,N_7876);
or U11620 (N_11620,N_6286,N_6507);
nand U11621 (N_11621,N_7875,N_8354);
and U11622 (N_11622,N_6878,N_7049);
nand U11623 (N_11623,N_8127,N_6886);
xnor U11624 (N_11624,N_8017,N_6770);
and U11625 (N_11625,N_8608,N_6425);
nor U11626 (N_11626,N_8122,N_6571);
and U11627 (N_11627,N_7324,N_6170);
nand U11628 (N_11628,N_8293,N_7124);
nand U11629 (N_11629,N_7242,N_8280);
or U11630 (N_11630,N_6774,N_7123);
and U11631 (N_11631,N_8232,N_7984);
nand U11632 (N_11632,N_7141,N_7900);
nand U11633 (N_11633,N_8070,N_6277);
and U11634 (N_11634,N_7988,N_7639);
and U11635 (N_11635,N_6869,N_7778);
xor U11636 (N_11636,N_6434,N_7672);
or U11637 (N_11637,N_6596,N_7268);
or U11638 (N_11638,N_6042,N_6512);
nor U11639 (N_11639,N_6898,N_7020);
nor U11640 (N_11640,N_6740,N_8234);
nor U11641 (N_11641,N_6617,N_8708);
and U11642 (N_11642,N_7859,N_7112);
or U11643 (N_11643,N_8549,N_8668);
nor U11644 (N_11644,N_7168,N_8148);
and U11645 (N_11645,N_7130,N_7880);
or U11646 (N_11646,N_7788,N_8442);
nand U11647 (N_11647,N_6065,N_7006);
and U11648 (N_11648,N_7617,N_7293);
or U11649 (N_11649,N_8729,N_8401);
or U11650 (N_11650,N_8582,N_6451);
or U11651 (N_11651,N_8948,N_8908);
and U11652 (N_11652,N_8967,N_7506);
nand U11653 (N_11653,N_8011,N_6502);
nand U11654 (N_11654,N_7118,N_7513);
nor U11655 (N_11655,N_8361,N_8926);
nand U11656 (N_11656,N_6736,N_8778);
nor U11657 (N_11657,N_8428,N_8305);
nor U11658 (N_11658,N_7308,N_7741);
nor U11659 (N_11659,N_8597,N_6723);
nand U11660 (N_11660,N_7448,N_6188);
and U11661 (N_11661,N_7010,N_6913);
nor U11662 (N_11662,N_7077,N_8885);
or U11663 (N_11663,N_7115,N_7362);
nor U11664 (N_11664,N_6897,N_7640);
nor U11665 (N_11665,N_6615,N_7211);
and U11666 (N_11666,N_8093,N_7568);
xnor U11667 (N_11667,N_8753,N_8703);
nand U11668 (N_11668,N_8380,N_6190);
nor U11669 (N_11669,N_8935,N_8271);
xor U11670 (N_11670,N_6901,N_6044);
or U11671 (N_11671,N_6213,N_8805);
nor U11672 (N_11672,N_6036,N_7737);
and U11673 (N_11673,N_6908,N_8680);
nand U11674 (N_11674,N_8577,N_6884);
nand U11675 (N_11675,N_8702,N_6851);
and U11676 (N_11676,N_6354,N_8756);
nor U11677 (N_11677,N_8487,N_8353);
nor U11678 (N_11678,N_8154,N_7126);
or U11679 (N_11679,N_6931,N_8585);
and U11680 (N_11680,N_6114,N_7535);
or U11681 (N_11681,N_8293,N_7139);
or U11682 (N_11682,N_8308,N_6839);
and U11683 (N_11683,N_7128,N_8108);
nand U11684 (N_11684,N_8573,N_7122);
nand U11685 (N_11685,N_6411,N_6888);
and U11686 (N_11686,N_6125,N_8278);
nand U11687 (N_11687,N_8293,N_6071);
nor U11688 (N_11688,N_6410,N_7946);
nor U11689 (N_11689,N_8357,N_8647);
and U11690 (N_11690,N_6803,N_8224);
nand U11691 (N_11691,N_8510,N_6919);
or U11692 (N_11692,N_6502,N_6030);
or U11693 (N_11693,N_8548,N_7082);
and U11694 (N_11694,N_7432,N_7422);
and U11695 (N_11695,N_6508,N_8057);
nand U11696 (N_11696,N_7965,N_6755);
or U11697 (N_11697,N_7036,N_8141);
nand U11698 (N_11698,N_8311,N_6179);
and U11699 (N_11699,N_6284,N_6461);
xnor U11700 (N_11700,N_6225,N_7681);
or U11701 (N_11701,N_7383,N_8408);
and U11702 (N_11702,N_7835,N_8853);
nand U11703 (N_11703,N_8405,N_7329);
and U11704 (N_11704,N_7716,N_8655);
and U11705 (N_11705,N_8936,N_8372);
nor U11706 (N_11706,N_8135,N_7484);
and U11707 (N_11707,N_8631,N_7416);
nand U11708 (N_11708,N_7752,N_6072);
nor U11709 (N_11709,N_8683,N_6908);
and U11710 (N_11710,N_8539,N_7667);
nand U11711 (N_11711,N_6120,N_8348);
nor U11712 (N_11712,N_6991,N_7420);
nor U11713 (N_11713,N_6440,N_6523);
xor U11714 (N_11714,N_8009,N_6693);
and U11715 (N_11715,N_8015,N_6984);
nor U11716 (N_11716,N_8331,N_7809);
nor U11717 (N_11717,N_6289,N_8344);
or U11718 (N_11718,N_7421,N_8438);
nand U11719 (N_11719,N_6168,N_6437);
nor U11720 (N_11720,N_7358,N_6178);
and U11721 (N_11721,N_7448,N_8995);
xor U11722 (N_11722,N_6020,N_7046);
or U11723 (N_11723,N_7295,N_7728);
xor U11724 (N_11724,N_7142,N_7023);
nor U11725 (N_11725,N_6058,N_8828);
or U11726 (N_11726,N_7277,N_7495);
nor U11727 (N_11727,N_6201,N_8242);
or U11728 (N_11728,N_8714,N_6694);
nor U11729 (N_11729,N_7154,N_7844);
nor U11730 (N_11730,N_6616,N_8488);
nor U11731 (N_11731,N_6952,N_8865);
nor U11732 (N_11732,N_8191,N_6863);
or U11733 (N_11733,N_6911,N_6727);
or U11734 (N_11734,N_7802,N_8147);
and U11735 (N_11735,N_7736,N_6683);
xor U11736 (N_11736,N_7891,N_8350);
nand U11737 (N_11737,N_7302,N_8856);
nand U11738 (N_11738,N_8877,N_8050);
nand U11739 (N_11739,N_6211,N_7165);
nor U11740 (N_11740,N_6652,N_7805);
nor U11741 (N_11741,N_7947,N_7621);
nor U11742 (N_11742,N_8603,N_7534);
nor U11743 (N_11743,N_7091,N_6653);
and U11744 (N_11744,N_6274,N_8676);
xnor U11745 (N_11745,N_7526,N_8168);
nor U11746 (N_11746,N_8317,N_7014);
and U11747 (N_11747,N_8102,N_6116);
or U11748 (N_11748,N_8254,N_8238);
nand U11749 (N_11749,N_6089,N_8658);
nand U11750 (N_11750,N_6752,N_6341);
nand U11751 (N_11751,N_7668,N_6422);
nand U11752 (N_11752,N_7576,N_7829);
nor U11753 (N_11753,N_6111,N_6889);
nand U11754 (N_11754,N_8942,N_6719);
or U11755 (N_11755,N_8294,N_6840);
xnor U11756 (N_11756,N_6543,N_7864);
nor U11757 (N_11757,N_7641,N_6402);
nand U11758 (N_11758,N_6479,N_7004);
nor U11759 (N_11759,N_7532,N_7583);
xnor U11760 (N_11760,N_6015,N_8865);
and U11761 (N_11761,N_7052,N_6507);
or U11762 (N_11762,N_6435,N_8334);
nor U11763 (N_11763,N_8229,N_8705);
or U11764 (N_11764,N_6117,N_7664);
or U11765 (N_11765,N_7963,N_7398);
nand U11766 (N_11766,N_6864,N_7969);
nor U11767 (N_11767,N_8244,N_7940);
nand U11768 (N_11768,N_8652,N_6474);
nor U11769 (N_11769,N_6760,N_6654);
nor U11770 (N_11770,N_7212,N_6137);
nand U11771 (N_11771,N_7802,N_6390);
nor U11772 (N_11772,N_7126,N_7799);
or U11773 (N_11773,N_6479,N_7407);
nor U11774 (N_11774,N_6071,N_6914);
or U11775 (N_11775,N_8305,N_7952);
or U11776 (N_11776,N_7889,N_8131);
and U11777 (N_11777,N_7257,N_6082);
or U11778 (N_11778,N_7189,N_6847);
and U11779 (N_11779,N_6019,N_8527);
nand U11780 (N_11780,N_7794,N_6265);
nand U11781 (N_11781,N_6156,N_6081);
and U11782 (N_11782,N_6016,N_7507);
and U11783 (N_11783,N_8728,N_8624);
nor U11784 (N_11784,N_7317,N_6450);
and U11785 (N_11785,N_7223,N_8664);
and U11786 (N_11786,N_6066,N_6542);
nand U11787 (N_11787,N_7151,N_8921);
nor U11788 (N_11788,N_6545,N_8343);
and U11789 (N_11789,N_6504,N_7561);
nor U11790 (N_11790,N_6278,N_6119);
nand U11791 (N_11791,N_6997,N_7550);
and U11792 (N_11792,N_7119,N_8886);
or U11793 (N_11793,N_8237,N_6227);
nand U11794 (N_11794,N_7657,N_7199);
xor U11795 (N_11795,N_8678,N_6138);
nor U11796 (N_11796,N_7195,N_6011);
nand U11797 (N_11797,N_8146,N_6374);
and U11798 (N_11798,N_7316,N_6089);
or U11799 (N_11799,N_7754,N_6480);
or U11800 (N_11800,N_7771,N_7109);
nor U11801 (N_11801,N_8870,N_7683);
nand U11802 (N_11802,N_6305,N_8141);
xnor U11803 (N_11803,N_7475,N_7176);
or U11804 (N_11804,N_7194,N_6277);
and U11805 (N_11805,N_8307,N_6434);
and U11806 (N_11806,N_6716,N_6474);
and U11807 (N_11807,N_7526,N_6782);
and U11808 (N_11808,N_7687,N_8332);
or U11809 (N_11809,N_8373,N_8283);
nor U11810 (N_11810,N_7215,N_8857);
nand U11811 (N_11811,N_6081,N_7893);
or U11812 (N_11812,N_6251,N_8556);
xnor U11813 (N_11813,N_6711,N_7339);
nor U11814 (N_11814,N_6212,N_8993);
and U11815 (N_11815,N_8721,N_8942);
nand U11816 (N_11816,N_6722,N_6784);
or U11817 (N_11817,N_8475,N_6906);
nand U11818 (N_11818,N_7485,N_7291);
nor U11819 (N_11819,N_6187,N_7306);
or U11820 (N_11820,N_8208,N_6730);
nor U11821 (N_11821,N_7924,N_7826);
nor U11822 (N_11822,N_6397,N_8564);
nand U11823 (N_11823,N_6016,N_8913);
nor U11824 (N_11824,N_8168,N_6656);
nand U11825 (N_11825,N_6263,N_8702);
or U11826 (N_11826,N_6940,N_7626);
or U11827 (N_11827,N_6396,N_6747);
nand U11828 (N_11828,N_8924,N_8100);
or U11829 (N_11829,N_6497,N_7721);
xnor U11830 (N_11830,N_6883,N_6375);
nor U11831 (N_11831,N_6051,N_7186);
nor U11832 (N_11832,N_7643,N_7450);
and U11833 (N_11833,N_8944,N_7101);
nor U11834 (N_11834,N_6999,N_8000);
or U11835 (N_11835,N_8028,N_7817);
nor U11836 (N_11836,N_7048,N_7895);
or U11837 (N_11837,N_7023,N_8800);
nor U11838 (N_11838,N_6258,N_7175);
nand U11839 (N_11839,N_8064,N_8367);
or U11840 (N_11840,N_6543,N_7778);
or U11841 (N_11841,N_7734,N_6253);
xnor U11842 (N_11842,N_8598,N_8122);
and U11843 (N_11843,N_8977,N_7772);
nand U11844 (N_11844,N_6077,N_7539);
nor U11845 (N_11845,N_8177,N_7332);
or U11846 (N_11846,N_8814,N_6320);
nor U11847 (N_11847,N_6021,N_6460);
and U11848 (N_11848,N_8280,N_6732);
xnor U11849 (N_11849,N_7262,N_6253);
nand U11850 (N_11850,N_8944,N_7613);
and U11851 (N_11851,N_7302,N_6790);
nor U11852 (N_11852,N_7254,N_8240);
nor U11853 (N_11853,N_6304,N_8120);
and U11854 (N_11854,N_7857,N_7401);
nor U11855 (N_11855,N_6163,N_7073);
nor U11856 (N_11856,N_8601,N_6352);
nand U11857 (N_11857,N_8676,N_7164);
and U11858 (N_11858,N_8121,N_6182);
nand U11859 (N_11859,N_8565,N_8443);
or U11860 (N_11860,N_8245,N_6933);
nand U11861 (N_11861,N_6360,N_8664);
and U11862 (N_11862,N_7971,N_7684);
and U11863 (N_11863,N_7707,N_6722);
or U11864 (N_11864,N_6491,N_8213);
and U11865 (N_11865,N_6490,N_8226);
and U11866 (N_11866,N_6706,N_8412);
xor U11867 (N_11867,N_8990,N_7746);
and U11868 (N_11868,N_8350,N_8074);
and U11869 (N_11869,N_6174,N_6185);
and U11870 (N_11870,N_7677,N_6940);
nand U11871 (N_11871,N_7312,N_6352);
nand U11872 (N_11872,N_7994,N_6384);
nor U11873 (N_11873,N_8494,N_7450);
or U11874 (N_11874,N_8696,N_7270);
or U11875 (N_11875,N_8091,N_6160);
nor U11876 (N_11876,N_8647,N_6272);
nor U11877 (N_11877,N_6818,N_7747);
xor U11878 (N_11878,N_8995,N_7758);
nand U11879 (N_11879,N_6015,N_8401);
nand U11880 (N_11880,N_8186,N_8351);
xnor U11881 (N_11881,N_8762,N_6808);
nor U11882 (N_11882,N_6947,N_6818);
xor U11883 (N_11883,N_8211,N_8791);
and U11884 (N_11884,N_8434,N_7227);
or U11885 (N_11885,N_8617,N_6057);
or U11886 (N_11886,N_6933,N_7842);
and U11887 (N_11887,N_7148,N_7726);
and U11888 (N_11888,N_7717,N_6364);
and U11889 (N_11889,N_7025,N_6841);
nand U11890 (N_11890,N_8680,N_7707);
nand U11891 (N_11891,N_6430,N_7788);
nand U11892 (N_11892,N_6025,N_7843);
nand U11893 (N_11893,N_7328,N_7197);
nand U11894 (N_11894,N_6775,N_6308);
xor U11895 (N_11895,N_8396,N_6096);
or U11896 (N_11896,N_7101,N_6372);
nand U11897 (N_11897,N_8784,N_8628);
or U11898 (N_11898,N_8251,N_7612);
nand U11899 (N_11899,N_7040,N_6417);
nand U11900 (N_11900,N_7435,N_6723);
and U11901 (N_11901,N_6321,N_6005);
nor U11902 (N_11902,N_6875,N_7623);
and U11903 (N_11903,N_8884,N_6176);
nor U11904 (N_11904,N_6035,N_8522);
or U11905 (N_11905,N_6213,N_7819);
nand U11906 (N_11906,N_8679,N_8759);
or U11907 (N_11907,N_6831,N_6386);
xor U11908 (N_11908,N_7607,N_6498);
or U11909 (N_11909,N_7620,N_8004);
and U11910 (N_11910,N_7164,N_8621);
nand U11911 (N_11911,N_7858,N_6250);
nand U11912 (N_11912,N_8805,N_7169);
and U11913 (N_11913,N_8975,N_6347);
nand U11914 (N_11914,N_7118,N_8160);
or U11915 (N_11915,N_7022,N_7929);
xor U11916 (N_11916,N_6053,N_6841);
nor U11917 (N_11917,N_6080,N_8558);
xnor U11918 (N_11918,N_6951,N_7547);
nor U11919 (N_11919,N_7362,N_6681);
or U11920 (N_11920,N_8327,N_6838);
and U11921 (N_11921,N_7179,N_6926);
nor U11922 (N_11922,N_7139,N_8157);
nor U11923 (N_11923,N_7397,N_8487);
and U11924 (N_11924,N_6288,N_8159);
nor U11925 (N_11925,N_8502,N_6326);
nor U11926 (N_11926,N_8380,N_7553);
xor U11927 (N_11927,N_8348,N_7951);
or U11928 (N_11928,N_7825,N_7283);
and U11929 (N_11929,N_7338,N_7783);
and U11930 (N_11930,N_8922,N_6192);
or U11931 (N_11931,N_6266,N_7012);
nand U11932 (N_11932,N_6646,N_8709);
nand U11933 (N_11933,N_7874,N_8338);
and U11934 (N_11934,N_7896,N_6666);
nor U11935 (N_11935,N_8021,N_6642);
nor U11936 (N_11936,N_6749,N_6970);
xor U11937 (N_11937,N_6895,N_8418);
nand U11938 (N_11938,N_8401,N_8842);
or U11939 (N_11939,N_8148,N_6435);
xnor U11940 (N_11940,N_7297,N_7897);
nor U11941 (N_11941,N_6312,N_7631);
nand U11942 (N_11942,N_6077,N_8330);
nand U11943 (N_11943,N_7804,N_7475);
or U11944 (N_11944,N_7991,N_6129);
nor U11945 (N_11945,N_7874,N_6585);
nand U11946 (N_11946,N_6200,N_6776);
nor U11947 (N_11947,N_7247,N_8593);
nor U11948 (N_11948,N_6919,N_6345);
or U11949 (N_11949,N_7775,N_7509);
nand U11950 (N_11950,N_7043,N_7741);
or U11951 (N_11951,N_6549,N_8791);
or U11952 (N_11952,N_8235,N_7047);
nand U11953 (N_11953,N_8964,N_7483);
nor U11954 (N_11954,N_8884,N_8978);
nand U11955 (N_11955,N_6943,N_8599);
and U11956 (N_11956,N_8674,N_8198);
xnor U11957 (N_11957,N_8006,N_8167);
nor U11958 (N_11958,N_6659,N_8914);
nand U11959 (N_11959,N_7605,N_6026);
and U11960 (N_11960,N_6264,N_6134);
or U11961 (N_11961,N_8152,N_7613);
nor U11962 (N_11962,N_8009,N_8264);
or U11963 (N_11963,N_8586,N_6023);
and U11964 (N_11964,N_8089,N_7136);
or U11965 (N_11965,N_8984,N_6215);
nand U11966 (N_11966,N_8671,N_6684);
and U11967 (N_11967,N_7148,N_8856);
nand U11968 (N_11968,N_7657,N_6509);
xnor U11969 (N_11969,N_7154,N_6134);
nand U11970 (N_11970,N_8800,N_8108);
and U11971 (N_11971,N_7077,N_8345);
xor U11972 (N_11972,N_6416,N_7562);
and U11973 (N_11973,N_6541,N_6677);
and U11974 (N_11974,N_6361,N_8699);
or U11975 (N_11975,N_8395,N_8513);
nor U11976 (N_11976,N_7835,N_8031);
nor U11977 (N_11977,N_7286,N_8812);
nand U11978 (N_11978,N_8354,N_6814);
nand U11979 (N_11979,N_8174,N_7821);
and U11980 (N_11980,N_6882,N_6513);
or U11981 (N_11981,N_8639,N_6957);
and U11982 (N_11982,N_7052,N_7897);
or U11983 (N_11983,N_8783,N_7264);
or U11984 (N_11984,N_7592,N_6912);
nor U11985 (N_11985,N_6694,N_7621);
or U11986 (N_11986,N_7901,N_8612);
nor U11987 (N_11987,N_8349,N_6398);
and U11988 (N_11988,N_7924,N_7020);
nor U11989 (N_11989,N_7257,N_8204);
xnor U11990 (N_11990,N_7418,N_6648);
nor U11991 (N_11991,N_6121,N_7244);
xor U11992 (N_11992,N_7707,N_7219);
nor U11993 (N_11993,N_6303,N_6402);
nor U11994 (N_11994,N_6628,N_7584);
or U11995 (N_11995,N_8549,N_8685);
and U11996 (N_11996,N_8625,N_6861);
and U11997 (N_11997,N_6198,N_8735);
nand U11998 (N_11998,N_8267,N_7762);
nor U11999 (N_11999,N_6661,N_7388);
or U12000 (N_12000,N_10357,N_9790);
and U12001 (N_12001,N_10282,N_11645);
or U12002 (N_12002,N_11707,N_11202);
or U12003 (N_12003,N_9518,N_11460);
and U12004 (N_12004,N_11459,N_9531);
or U12005 (N_12005,N_10973,N_9835);
nor U12006 (N_12006,N_10052,N_9774);
and U12007 (N_12007,N_9442,N_9168);
and U12008 (N_12008,N_11930,N_9973);
nor U12009 (N_12009,N_9077,N_9002);
nor U12010 (N_12010,N_9311,N_10695);
nand U12011 (N_12011,N_10903,N_10868);
or U12012 (N_12012,N_9356,N_10270);
and U12013 (N_12013,N_11754,N_9722);
xnor U12014 (N_12014,N_11805,N_11725);
nand U12015 (N_12015,N_10978,N_10960);
or U12016 (N_12016,N_11906,N_9213);
or U12017 (N_12017,N_11745,N_10897);
nand U12018 (N_12018,N_11405,N_9252);
nand U12019 (N_12019,N_10110,N_11799);
nand U12020 (N_12020,N_9841,N_10666);
or U12021 (N_12021,N_11087,N_10992);
or U12022 (N_12022,N_9096,N_11187);
nor U12023 (N_12023,N_11137,N_9146);
nor U12024 (N_12024,N_10882,N_10100);
xnor U12025 (N_12025,N_10125,N_10640);
nand U12026 (N_12026,N_9102,N_11017);
xor U12027 (N_12027,N_10917,N_11908);
or U12028 (N_12028,N_10124,N_9831);
or U12029 (N_12029,N_9454,N_9052);
and U12030 (N_12030,N_9475,N_11368);
or U12031 (N_12031,N_9093,N_9240);
nor U12032 (N_12032,N_9085,N_10624);
or U12033 (N_12033,N_9009,N_10271);
xnor U12034 (N_12034,N_11406,N_9760);
and U12035 (N_12035,N_9643,N_11741);
or U12036 (N_12036,N_11516,N_9840);
nor U12037 (N_12037,N_10998,N_10557);
and U12038 (N_12038,N_9290,N_11367);
and U12039 (N_12039,N_11461,N_9821);
or U12040 (N_12040,N_11288,N_9349);
nand U12041 (N_12041,N_9169,N_11131);
or U12042 (N_12042,N_9268,N_11861);
nand U12043 (N_12043,N_9108,N_9269);
nand U12044 (N_12044,N_11918,N_10250);
or U12045 (N_12045,N_11657,N_10525);
or U12046 (N_12046,N_11231,N_9890);
xor U12047 (N_12047,N_10537,N_10795);
nand U12048 (N_12048,N_9471,N_9872);
and U12049 (N_12049,N_9985,N_10989);
and U12050 (N_12050,N_9786,N_9981);
nand U12051 (N_12051,N_10389,N_10018);
nor U12052 (N_12052,N_11124,N_10997);
or U12053 (N_12053,N_10353,N_11129);
nor U12054 (N_12054,N_10546,N_9119);
or U12055 (N_12055,N_10059,N_10149);
nor U12056 (N_12056,N_10941,N_10912);
nand U12057 (N_12057,N_9614,N_9669);
nand U12058 (N_12058,N_10962,N_9181);
or U12059 (N_12059,N_11032,N_9881);
xnor U12060 (N_12060,N_10220,N_11715);
nor U12061 (N_12061,N_9803,N_9113);
nor U12062 (N_12062,N_10435,N_9399);
and U12063 (N_12063,N_9978,N_11012);
and U12064 (N_12064,N_10735,N_9036);
nor U12065 (N_12065,N_9325,N_11445);
xnor U12066 (N_12066,N_9548,N_10055);
nand U12067 (N_12067,N_10115,N_9069);
nor U12068 (N_12068,N_11652,N_10713);
nor U12069 (N_12069,N_11259,N_9289);
xor U12070 (N_12070,N_9633,N_9051);
xnor U12071 (N_12071,N_10551,N_11230);
and U12072 (N_12072,N_10488,N_9745);
nand U12073 (N_12073,N_9467,N_9435);
xnor U12074 (N_12074,N_11197,N_9566);
xor U12075 (N_12075,N_9788,N_9083);
and U12076 (N_12076,N_10225,N_10456);
and U12077 (N_12077,N_10919,N_11214);
and U12078 (N_12078,N_10970,N_9323);
or U12079 (N_12079,N_9486,N_9006);
and U12080 (N_12080,N_10050,N_11082);
nand U12081 (N_12081,N_10610,N_11569);
or U12082 (N_12082,N_11661,N_11552);
or U12083 (N_12083,N_9133,N_9228);
nor U12084 (N_12084,N_9709,N_11207);
nor U12085 (N_12085,N_9142,N_10209);
nand U12086 (N_12086,N_10684,N_11440);
nor U12087 (N_12087,N_10049,N_9933);
and U12088 (N_12088,N_10300,N_9297);
nor U12089 (N_12089,N_11026,N_11083);
and U12090 (N_12090,N_9880,N_10460);
nand U12091 (N_12091,N_10676,N_11609);
and U12092 (N_12092,N_9087,N_9075);
nor U12093 (N_12093,N_11956,N_9209);
xnor U12094 (N_12094,N_9928,N_9470);
nand U12095 (N_12095,N_10630,N_11967);
nand U12096 (N_12096,N_10237,N_10378);
or U12097 (N_12097,N_10348,N_10333);
and U12098 (N_12098,N_10368,N_9971);
nand U12099 (N_12099,N_9613,N_10665);
or U12100 (N_12100,N_11226,N_9128);
nor U12101 (N_12101,N_9538,N_10858);
nor U12102 (N_12102,N_11040,N_11785);
or U12103 (N_12103,N_11765,N_10890);
nor U12104 (N_12104,N_10079,N_9187);
nand U12105 (N_12105,N_10185,N_9752);
and U12106 (N_12106,N_11423,N_11344);
or U12107 (N_12107,N_10545,N_11162);
nand U12108 (N_12108,N_9299,N_9092);
nand U12109 (N_12109,N_11984,N_11727);
nor U12110 (N_12110,N_9529,N_10136);
nand U12111 (N_12111,N_9173,N_9911);
xnor U12112 (N_12112,N_10518,N_11734);
nor U12113 (N_12113,N_10806,N_9878);
nand U12114 (N_12114,N_10345,N_11695);
or U12115 (N_12115,N_9528,N_9089);
and U12116 (N_12116,N_11110,N_9353);
nor U12117 (N_12117,N_11605,N_11009);
nand U12118 (N_12118,N_11262,N_11993);
and U12119 (N_12119,N_10672,N_10755);
or U12120 (N_12120,N_9319,N_10527);
and U12121 (N_12121,N_10264,N_11890);
or U12122 (N_12122,N_11400,N_10422);
or U12123 (N_12123,N_11211,N_10823);
nor U12124 (N_12124,N_11052,N_11146);
nor U12125 (N_12125,N_11870,N_10490);
nor U12126 (N_12126,N_9152,N_11311);
nor U12127 (N_12127,N_10967,N_9065);
nand U12128 (N_12128,N_9879,N_11468);
nand U12129 (N_12129,N_11261,N_9818);
or U12130 (N_12130,N_9759,N_10238);
or U12131 (N_12131,N_10524,N_10671);
nor U12132 (N_12132,N_9592,N_11486);
or U12133 (N_12133,N_11008,N_10257);
nand U12134 (N_12134,N_10338,N_9479);
or U12135 (N_12135,N_10475,N_9585);
and U12136 (N_12136,N_9666,N_11023);
nand U12137 (N_12137,N_9233,N_10776);
nor U12138 (N_12138,N_9622,N_10117);
nand U12139 (N_12139,N_11410,N_11517);
nor U12140 (N_12140,N_9720,N_9569);
nand U12141 (N_12141,N_9799,N_10246);
and U12142 (N_12142,N_10476,N_9648);
or U12143 (N_12143,N_9322,N_10639);
or U12144 (N_12144,N_9428,N_11381);
and U12145 (N_12145,N_11104,N_11560);
nand U12146 (N_12146,N_10213,N_10285);
or U12147 (N_12147,N_11491,N_10090);
nand U12148 (N_12148,N_9285,N_9673);
nand U12149 (N_12149,N_10299,N_10797);
or U12150 (N_12150,N_10060,N_9210);
and U12151 (N_12151,N_9452,N_10714);
nand U12152 (N_12152,N_11498,N_9870);
nand U12153 (N_12153,N_10502,N_9656);
and U12154 (N_12154,N_10116,N_10195);
nor U12155 (N_12155,N_9256,N_9789);
and U12156 (N_12156,N_11228,N_11896);
or U12157 (N_12157,N_10219,N_10884);
and U12158 (N_12158,N_11313,N_10278);
or U12159 (N_12159,N_11921,N_10581);
nand U12160 (N_12160,N_10170,N_10226);
nor U12161 (N_12161,N_11597,N_10556);
or U12162 (N_12162,N_9387,N_10274);
nand U12163 (N_12163,N_10145,N_11111);
and U12164 (N_12164,N_10153,N_9743);
nor U12165 (N_12165,N_10076,N_10986);
nor U12166 (N_12166,N_9432,N_11522);
xnor U12167 (N_12167,N_9557,N_11308);
and U12168 (N_12168,N_10382,N_9603);
nor U12169 (N_12169,N_10984,N_9834);
and U12170 (N_12170,N_10608,N_11565);
nor U12171 (N_12171,N_10341,N_10501);
and U12172 (N_12172,N_10114,N_11169);
xor U12173 (N_12173,N_10730,N_11135);
nor U12174 (N_12174,N_10854,N_11603);
nand U12175 (N_12175,N_9849,N_10315);
and U12176 (N_12176,N_10165,N_11935);
nor U12177 (N_12177,N_11443,N_9282);
nand U12178 (N_12178,N_10003,N_9016);
or U12179 (N_12179,N_11800,N_11458);
nor U12180 (N_12180,N_11359,N_9386);
nor U12181 (N_12181,N_9175,N_11672);
nor U12182 (N_12182,N_10011,N_11441);
xor U12183 (N_12183,N_9868,N_11816);
nand U12184 (N_12184,N_10982,N_9650);
and U12185 (N_12185,N_9995,N_9559);
or U12186 (N_12186,N_10470,N_11966);
and U12187 (N_12187,N_9207,N_10664);
or U12188 (N_12188,N_11619,N_9645);
and U12189 (N_12189,N_10739,N_10439);
or U12190 (N_12190,N_9655,N_10363);
nor U12191 (N_12191,N_10881,N_11212);
nand U12192 (N_12192,N_11171,N_11824);
nor U12193 (N_12193,N_10016,N_11648);
nand U12194 (N_12194,N_11225,N_10214);
nor U12195 (N_12195,N_11769,N_9511);
or U12196 (N_12196,N_11549,N_11699);
and U12197 (N_12197,N_10134,N_9057);
nor U12198 (N_12198,N_10221,N_10373);
nor U12199 (N_12199,N_9573,N_11398);
and U12200 (N_12200,N_9136,N_9354);
or U12201 (N_12201,N_9130,N_10971);
or U12202 (N_12202,N_10930,N_11404);
nand U12203 (N_12203,N_9012,N_10876);
or U12204 (N_12204,N_9010,N_9658);
nand U12205 (N_12205,N_9318,N_11312);
and U12206 (N_12206,N_10494,N_9484);
nor U12207 (N_12207,N_11036,N_10308);
or U12208 (N_12208,N_9338,N_9632);
and U12209 (N_12209,N_10179,N_11938);
or U12210 (N_12210,N_9994,N_11991);
and U12211 (N_12211,N_11088,N_11886);
nand U12212 (N_12212,N_10482,N_10148);
nand U12213 (N_12213,N_11815,N_10601);
nand U12214 (N_12214,N_9558,N_11842);
nand U12215 (N_12215,N_11422,N_9215);
or U12216 (N_12216,N_10168,N_11182);
or U12217 (N_12217,N_11823,N_11901);
nand U12218 (N_12218,N_10491,N_10269);
xnor U12219 (N_12219,N_9616,N_10392);
or U12220 (N_12220,N_9764,N_10463);
nand U12221 (N_12221,N_9114,N_9198);
nor U12222 (N_12222,N_10385,N_10994);
nor U12223 (N_12223,N_9575,N_11188);
nor U12224 (N_12224,N_9015,N_10505);
xor U12225 (N_12225,N_11485,N_11252);
nor U12226 (N_12226,N_10289,N_11833);
and U12227 (N_12227,N_9698,N_9716);
nand U12228 (N_12228,N_11393,N_11616);
nor U12229 (N_12229,N_9327,N_10840);
or U12230 (N_12230,N_9466,N_10945);
or U12231 (N_12231,N_9577,N_9986);
nor U12232 (N_12232,N_11472,N_10774);
nor U12233 (N_12233,N_9823,N_10745);
or U12234 (N_12234,N_11857,N_10754);
and U12235 (N_12235,N_9007,N_11513);
nor U12236 (N_12236,N_11607,N_11810);
or U12237 (N_12237,N_9062,N_9811);
and U12238 (N_12238,N_10925,N_11253);
nor U12239 (N_12239,N_10584,N_10592);
nor U12240 (N_12240,N_9064,N_11949);
nor U12241 (N_12241,N_10779,N_10874);
or U12242 (N_12242,N_10659,N_10885);
xnor U12243 (N_12243,N_11469,N_10056);
or U12244 (N_12244,N_10102,N_11594);
nand U12245 (N_12245,N_10020,N_9920);
xnor U12246 (N_12246,N_11903,N_11487);
or U12247 (N_12247,N_10705,N_10983);
nor U12248 (N_12248,N_10094,N_10586);
or U12249 (N_12249,N_9974,N_11470);
and U12250 (N_12250,N_9508,N_11412);
and U12251 (N_12251,N_9004,N_11070);
nor U12252 (N_12252,N_9433,N_9249);
nor U12253 (N_12253,N_9226,N_9121);
nand U12254 (N_12254,N_10837,N_11974);
or U12255 (N_12255,N_11771,N_11576);
xor U12256 (N_12256,N_10523,N_10273);
nor U12257 (N_12257,N_10403,N_11527);
nor U12258 (N_12258,N_9101,N_10267);
or U12259 (N_12259,N_11478,N_10820);
nor U12260 (N_12260,N_9443,N_10051);
nand U12261 (N_12261,N_9839,N_11455);
or U12262 (N_12262,N_9343,N_9138);
nor U12263 (N_12263,N_11978,N_10555);
xnor U12264 (N_12264,N_11326,N_10542);
nand U12265 (N_12265,N_9397,N_11747);
or U12266 (N_12266,N_11170,N_9251);
or U12267 (N_12267,N_9731,N_9150);
nor U12268 (N_12268,N_11858,N_9234);
and U12269 (N_12269,N_11025,N_9693);
xor U12270 (N_12270,N_9229,N_11150);
or U12271 (N_12271,N_10072,N_10048);
and U12272 (N_12272,N_11389,N_10550);
or U12273 (N_12273,N_11743,N_11094);
or U12274 (N_12274,N_10182,N_10126);
and U12275 (N_12275,N_11219,N_9676);
nand U12276 (N_12276,N_10272,N_11977);
and U12277 (N_12277,N_10139,N_10559);
nor U12278 (N_12278,N_10914,N_11065);
or U12279 (N_12279,N_10744,N_9188);
xnor U12280 (N_12280,N_11397,N_9339);
nor U12281 (N_12281,N_11489,N_11245);
nand U12282 (N_12282,N_11531,N_11911);
and U12283 (N_12283,N_9125,N_10040);
and U12284 (N_12284,N_9286,N_10748);
and U12285 (N_12285,N_10395,N_9407);
and U12286 (N_12286,N_10216,N_11375);
and U12287 (N_12287,N_10570,N_11760);
xor U12288 (N_12288,N_9785,N_10192);
nor U12289 (N_12289,N_9374,N_10256);
and U12290 (N_12290,N_11946,N_10266);
or U12291 (N_12291,N_9491,N_9337);
nand U12292 (N_12292,N_10162,N_11784);
nand U12293 (N_12293,N_9111,N_9259);
and U12294 (N_12294,N_10397,N_10762);
or U12295 (N_12295,N_10813,N_9347);
nand U12296 (N_12296,N_11347,N_10449);
xnor U12297 (N_12297,N_10263,N_11377);
nor U12298 (N_12298,N_11637,N_11889);
nor U12299 (N_12299,N_11315,N_10712);
nor U12300 (N_12300,N_9706,N_11192);
and U12301 (N_12301,N_11421,N_11562);
and U12302 (N_12302,N_9024,N_9663);
and U12303 (N_12303,N_11394,N_10576);
xnor U12304 (N_12304,N_11872,N_9516);
nand U12305 (N_12305,N_10109,N_11456);
and U12306 (N_12306,N_9043,N_9419);
nand U12307 (N_12307,N_10694,N_11763);
nor U12308 (N_12308,N_11692,N_10954);
and U12309 (N_12309,N_9238,N_11073);
nand U12310 (N_12310,N_9812,N_9448);
nor U12311 (N_12311,N_11586,N_9266);
nand U12312 (N_12312,N_11767,N_10222);
nor U12313 (N_12313,N_11762,N_11797);
and U12314 (N_12314,N_11439,N_11418);
xor U12315 (N_12315,N_10894,N_11272);
and U12316 (N_12316,N_10690,N_9157);
nor U12317 (N_12317,N_11650,N_11305);
or U12318 (N_12318,N_9357,N_10901);
or U12319 (N_12319,N_9710,N_10807);
nand U12320 (N_12320,N_9951,N_11257);
and U12321 (N_12321,N_11484,N_10122);
or U12322 (N_12322,N_11668,N_9615);
nand U12323 (N_12323,N_10727,N_10471);
and U12324 (N_12324,N_10859,N_10822);
nor U12325 (N_12325,N_11866,N_9711);
nor U12326 (N_12326,N_11595,N_11343);
nand U12327 (N_12327,N_9179,N_10260);
nor U12328 (N_12328,N_11399,N_10497);
nand U12329 (N_12329,N_10321,N_10204);
nand U12330 (N_12330,N_9915,N_10438);
nor U12331 (N_12331,N_9131,N_11233);
nor U12332 (N_12332,N_11497,N_10996);
and U12333 (N_12333,N_9684,N_10635);
and U12334 (N_12334,N_11270,N_11107);
nor U12335 (N_12335,N_9017,N_11604);
nand U12336 (N_12336,N_11689,N_11499);
nor U12337 (N_12337,N_11798,N_9312);
nand U12338 (N_12338,N_9984,N_10087);
nand U12339 (N_12339,N_11566,N_11708);
nor U12340 (N_12340,N_9996,N_11772);
and U12341 (N_12341,N_9802,N_9081);
nor U12342 (N_12342,N_10814,N_10207);
or U12343 (N_12343,N_9330,N_11425);
or U12344 (N_12344,N_11213,N_10801);
nand U12345 (N_12345,N_10987,N_9851);
or U12346 (N_12346,N_10371,N_11812);
and U12347 (N_12347,N_10193,N_11471);
and U12348 (N_12348,N_9739,N_9172);
nand U12349 (N_12349,N_11931,N_11869);
nor U12350 (N_12350,N_9235,N_11995);
nand U12351 (N_12351,N_9298,N_11783);
or U12352 (N_12352,N_9916,N_9944);
xnor U12353 (N_12353,N_10606,N_11337);
and U12354 (N_12354,N_9754,N_10855);
xor U12355 (N_12355,N_11782,N_11356);
nand U12356 (N_12356,N_9814,N_11300);
or U12357 (N_12357,N_9847,N_9143);
or U12358 (N_12358,N_9830,N_11284);
nand U12359 (N_12359,N_11388,N_10787);
and U12360 (N_12360,N_9336,N_10492);
and U12361 (N_12361,N_11507,N_10878);
nor U12362 (N_12362,N_10759,N_11736);
and U12363 (N_12363,N_9401,N_10361);
or U12364 (N_12364,N_10377,N_10458);
nor U12365 (N_12365,N_10099,N_10831);
nor U12366 (N_12366,N_10623,N_9551);
or U12367 (N_12367,N_10086,N_11766);
nand U12368 (N_12368,N_11618,N_9091);
nand U12369 (N_12369,N_11593,N_9753);
and U12370 (N_12370,N_9171,N_9961);
xnor U12371 (N_12371,N_10811,N_11855);
nand U12372 (N_12372,N_10850,N_9713);
or U12373 (N_12373,N_9927,N_9054);
nand U12374 (N_12374,N_9744,N_9254);
and U12375 (N_12375,N_9857,N_11626);
or U12376 (N_12376,N_10303,N_10964);
xnor U12377 (N_12377,N_11319,N_11572);
xor U12378 (N_12378,N_11464,N_9140);
xor U12379 (N_12379,N_11492,N_11501);
nor U12380 (N_12380,N_10297,N_9977);
nor U12381 (N_12381,N_11140,N_9273);
nand U12382 (N_12382,N_10426,N_11899);
and U12383 (N_12383,N_9550,N_10547);
or U12384 (N_12384,N_9050,N_11295);
and U12385 (N_12385,N_10660,N_11427);
or U12386 (N_12386,N_10066,N_9261);
nor U12387 (N_12387,N_9560,N_11078);
nor U12388 (N_12388,N_9197,N_10612);
nand U12389 (N_12389,N_11885,N_11514);
or U12390 (N_12390,N_10766,N_9366);
xor U12391 (N_12391,N_11686,N_10414);
and U12392 (N_12392,N_10150,N_11058);
nand U12393 (N_12393,N_11003,N_10320);
nand U12394 (N_12394,N_10319,N_10186);
or U12395 (N_12395,N_11988,N_9141);
or U12396 (N_12396,N_10477,N_11072);
xor U12397 (N_12397,N_9598,N_10360);
nor U12398 (N_12398,N_9232,N_10138);
and U12399 (N_12399,N_11181,N_11742);
or U12400 (N_12400,N_9571,N_10942);
nor U12401 (N_12401,N_9733,N_11413);
nor U12402 (N_12402,N_10092,N_10008);
nor U12403 (N_12403,N_9084,N_9924);
nand U12404 (N_12404,N_11592,N_9301);
nor U12405 (N_12405,N_11675,N_11482);
nor U12406 (N_12406,N_9833,N_11887);
nor U12407 (N_12407,N_10835,N_11582);
and U12408 (N_12408,N_9523,N_11660);
or U12409 (N_12409,N_9378,N_9122);
nor U12410 (N_12410,N_10275,N_11221);
nor U12411 (N_12411,N_11787,N_9302);
or U12412 (N_12412,N_9646,N_10334);
nand U12413 (N_12413,N_10792,N_9183);
and U12414 (N_12414,N_9826,N_9599);
nand U12415 (N_12415,N_10541,N_11323);
nor U12416 (N_12416,N_10856,N_9061);
xor U12417 (N_12417,N_9923,N_11133);
and U12418 (N_12418,N_10956,N_11696);
nor U12419 (N_12419,N_11060,N_9783);
and U12420 (N_12420,N_9078,N_10733);
nand U12421 (N_12421,N_10832,N_10356);
or U12422 (N_12422,N_9132,N_10793);
nand U12423 (N_12423,N_10326,N_10317);
nand U12424 (N_12424,N_10808,N_9206);
or U12425 (N_12425,N_10722,N_10985);
or U12426 (N_12426,N_10327,N_9869);
nand U12427 (N_12427,N_9664,N_11051);
or U12428 (N_12428,N_10074,N_9100);
or U12429 (N_12429,N_11276,N_10844);
and U12430 (N_12430,N_9473,N_10388);
nor U12431 (N_12431,N_9605,N_9817);
and U12432 (N_12432,N_11307,N_9377);
nor U12433 (N_12433,N_10252,N_11704);
or U12434 (N_12434,N_10817,N_10924);
or U12435 (N_12435,N_11854,N_9824);
xor U12436 (N_12436,N_10863,N_11465);
xor U12437 (N_12437,N_9522,N_11969);
xnor U12438 (N_12438,N_10661,N_9705);
or U12439 (N_12439,N_9219,N_11524);
nor U12440 (N_12440,N_10654,N_10734);
and U12441 (N_12441,N_10819,N_9581);
and U12442 (N_12442,N_10104,N_10829);
or U12443 (N_12443,N_10773,N_9773);
xor U12444 (N_12444,N_11953,N_9192);
and U12445 (N_12445,N_10014,N_9647);
nor U12446 (N_12446,N_9549,N_11283);
or U12447 (N_12447,N_9341,N_10268);
nand U12448 (N_12448,N_11932,N_11098);
nor U12449 (N_12449,N_9056,N_11066);
nand U12450 (N_12450,N_9221,N_10702);
nor U12451 (N_12451,N_10340,N_11678);
nor U12452 (N_12452,N_11035,N_9193);
nor U12453 (N_12453,N_10459,N_11850);
xor U12454 (N_12454,N_11385,N_9820);
nand U12455 (N_12455,N_9950,N_10408);
or U12456 (N_12456,N_11010,N_11888);
nor U12457 (N_12457,N_10803,N_11613);
nor U12458 (N_12458,N_10228,N_11044);
or U12459 (N_12459,N_10129,N_9779);
or U12460 (N_12460,N_9941,N_9212);
and U12461 (N_12461,N_10335,N_9359);
nor U12462 (N_12462,N_9935,N_9604);
or U12463 (N_12463,N_10313,N_9342);
nor U12464 (N_12464,N_10633,N_9189);
and U12465 (N_12465,N_10331,N_9416);
and U12466 (N_12466,N_11334,N_10288);
nor U12467 (N_12467,N_10098,N_9991);
nand U12468 (N_12468,N_9253,N_9685);
nand U12469 (N_12469,N_9702,N_10637);
nor U12470 (N_12470,N_11860,N_10804);
nand U12471 (N_12471,N_10188,N_11673);
or U12472 (N_12472,N_10253,N_11021);
xnor U12473 (N_12473,N_11435,N_9149);
nand U12474 (N_12474,N_9524,N_11963);
xnor U12475 (N_12475,N_10693,N_9053);
or U12476 (N_12476,N_9761,N_11105);
nor U12477 (N_12477,N_9422,N_9757);
and U12478 (N_12478,N_9129,N_10151);
nor U12479 (N_12479,N_9842,N_11687);
nand U12480 (N_12480,N_10616,N_9853);
nor U12481 (N_12481,N_11155,N_9572);
or U12482 (N_12482,N_10425,N_11166);
xor U12483 (N_12483,N_10386,N_11744);
xor U12484 (N_12484,N_10034,N_11067);
xnor U12485 (N_12485,N_9939,N_10939);
and U12486 (N_12486,N_11683,N_9034);
and U12487 (N_12487,N_11955,N_11139);
nand U12488 (N_12488,N_11209,N_11480);
or U12489 (N_12489,N_9654,N_9597);
nor U12490 (N_12490,N_10668,N_9520);
or U12491 (N_12491,N_9690,N_10680);
nand U12492 (N_12492,N_11001,N_9909);
or U12493 (N_12493,N_10706,N_9202);
xor U12494 (N_12494,N_9222,N_11998);
or U12495 (N_12495,N_9208,N_11301);
nand U12496 (N_12496,N_10526,N_10108);
and U12497 (N_12497,N_10351,N_9782);
and U12498 (N_12498,N_11075,N_11016);
and U12499 (N_12499,N_11152,N_10775);
nand U12500 (N_12500,N_9037,N_11241);
nand U12501 (N_12501,N_10381,N_10375);
nor U12502 (N_12502,N_11898,N_9328);
nor U12503 (N_12503,N_11024,N_11416);
and U12504 (N_12504,N_11753,N_9430);
and U12505 (N_12505,N_9864,N_9755);
or U12506 (N_12506,N_10171,N_11014);
nor U12507 (N_12507,N_10558,N_10513);
and U12508 (N_12508,N_9126,N_10223);
and U12509 (N_12509,N_11851,N_9063);
nand U12510 (N_12510,N_10577,N_9892);
nand U12511 (N_12511,N_11680,N_11157);
nand U12512 (N_12512,N_10594,N_10405);
xnor U12513 (N_12513,N_9032,N_10133);
or U12514 (N_12514,N_10763,N_9746);
and U12515 (N_12515,N_10352,N_10084);
nor U12516 (N_12516,N_11488,N_11353);
or U12517 (N_12517,N_11142,N_9107);
and U12518 (N_12518,N_10609,N_9611);
nor U12519 (N_12519,N_11837,N_10590);
and U12520 (N_12520,N_11937,N_9079);
nand U12521 (N_12521,N_11018,N_9642);
nand U12522 (N_12522,N_11970,N_9271);
nor U12523 (N_12523,N_11322,N_10295);
and U12524 (N_12524,N_9947,N_11999);
and U12525 (N_12525,N_11390,N_10758);
nor U12526 (N_12526,N_11965,N_11362);
or U12527 (N_12527,N_9822,N_10589);
or U12528 (N_12528,N_11554,N_11190);
nand U12529 (N_12529,N_11145,N_9066);
nor U12530 (N_12530,N_11496,N_9035);
and U12531 (N_12531,N_10948,N_10215);
or U12532 (N_12532,N_11373,N_9934);
and U12533 (N_12533,N_11034,N_9242);
nor U12534 (N_12534,N_10009,N_11540);
nor U12535 (N_12535,N_10161,N_10652);
nor U12536 (N_12536,N_10017,N_10540);
or U12537 (N_12537,N_9768,N_11002);
or U12538 (N_12538,N_10281,N_11781);
nand U12539 (N_12539,N_11159,N_9871);
nor U12540 (N_12540,N_10958,N_10004);
xor U12541 (N_12541,N_11320,N_10398);
nor U12542 (N_12542,N_10444,N_10365);
nand U12543 (N_12543,N_10747,N_11710);
nand U12544 (N_12544,N_10071,N_9191);
or U12545 (N_12545,N_10199,N_11165);
and U12546 (N_12546,N_10889,N_11746);
or U12547 (N_12547,N_9556,N_11843);
nor U12548 (N_12548,N_10258,N_10484);
nor U12549 (N_12549,N_9696,N_11684);
or U12550 (N_12550,N_9778,N_11382);
or U12551 (N_12551,N_10111,N_11047);
nor U12552 (N_12552,N_11260,N_10175);
nand U12553 (N_12553,N_9792,N_11542);
nand U12554 (N_12554,N_10533,N_11574);
or U12555 (N_12555,N_10486,N_11895);
nor U12556 (N_12556,N_10241,N_9483);
xor U12557 (N_12557,N_10157,N_10140);
nand U12558 (N_12558,N_9413,N_10548);
nand U12559 (N_12559,N_10574,N_9772);
or U12560 (N_12560,N_11556,N_11844);
nor U12561 (N_12561,N_10479,N_10886);
nand U12562 (N_12562,N_10027,N_10614);
nand U12563 (N_12563,N_9636,N_10703);
nand U12564 (N_12564,N_11327,N_11128);
and U12565 (N_12565,N_11841,N_9026);
nor U12566 (N_12566,N_9660,N_11801);
and U12567 (N_12567,N_11666,N_9699);
nand U12568 (N_12568,N_10922,N_9588);
nand U12569 (N_12569,N_9608,N_9158);
and U12570 (N_12570,N_9068,N_10767);
and U12571 (N_12571,N_9809,N_9682);
nand U12572 (N_12572,N_10845,N_11519);
or U12573 (N_12573,N_9040,N_10154);
nor U12574 (N_12574,N_10362,N_9515);
and U12575 (N_12575,N_10218,N_11175);
or U12576 (N_12576,N_9177,N_10753);
nand U12577 (N_12577,N_11653,N_10167);
nand U12578 (N_12578,N_11467,N_11624);
nand U12579 (N_12579,N_9715,N_11822);
or U12580 (N_12580,N_9607,N_10196);
or U12581 (N_12581,N_10561,N_9384);
nor U12582 (N_12582,N_11280,N_10952);
nand U12583 (N_12583,N_11509,N_11185);
nor U12584 (N_12584,N_9888,N_9670);
and U12585 (N_12585,N_10909,N_9513);
nor U12586 (N_12586,N_11206,N_9963);
and U12587 (N_12587,N_10908,N_11396);
xnor U12588 (N_12588,N_10451,N_10674);
nor U12589 (N_12589,N_11452,N_10447);
and U12590 (N_12590,N_10217,N_9620);
nand U12591 (N_12591,N_9504,N_11013);
or U12592 (N_12592,N_9780,N_9895);
nand U12593 (N_12593,N_10708,N_11194);
xor U12594 (N_12594,N_9987,N_10880);
and U12595 (N_12595,N_11265,N_11109);
xnor U12596 (N_12596,N_11339,N_11050);
nand U12597 (N_12597,N_9553,N_9332);
and U12598 (N_12598,N_10756,N_10311);
nand U12599 (N_12599,N_11019,N_10254);
nor U12600 (N_12600,N_11670,N_11864);
nand U12601 (N_12601,N_9844,N_9031);
nand U12602 (N_12602,N_10239,N_9241);
nand U12603 (N_12603,N_11987,N_9310);
nand U12604 (N_12604,N_11877,N_9224);
xnor U12605 (N_12605,N_10532,N_11287);
or U12606 (N_12606,N_10716,N_10597);
nor U12607 (N_12607,N_9494,N_11697);
and U12608 (N_12608,N_11317,N_10453);
nor U12609 (N_12609,N_11525,N_11902);
or U12610 (N_12610,N_11596,N_11968);
and U12611 (N_12611,N_11957,N_11808);
and U12612 (N_12612,N_9949,N_10450);
or U12613 (N_12613,N_11701,N_11447);
xnor U12614 (N_12614,N_10077,N_11705);
nand U12615 (N_12615,N_9776,N_9153);
nand U12616 (N_12616,N_9546,N_11453);
nand U12617 (N_12617,N_10206,N_9184);
xnor U12618 (N_12618,N_10243,N_10409);
nor U12619 (N_12619,N_11273,N_10563);
or U12620 (N_12620,N_9567,N_9363);
and U12621 (N_12621,N_10857,N_11623);
xnor U12622 (N_12622,N_11982,N_11871);
nand U12623 (N_12623,N_11553,N_9362);
and U12624 (N_12624,N_11358,N_11494);
nand U12625 (N_12625,N_11638,N_11832);
nand U12626 (N_12626,N_9534,N_9369);
and U12627 (N_12627,N_11942,N_9703);
or U12628 (N_12628,N_9926,N_9431);
and U12629 (N_12629,N_10701,N_10043);
xor U12630 (N_12630,N_9852,N_11346);
and U12631 (N_12631,N_10743,N_9848);
or U12632 (N_12632,N_11395,N_11639);
or U12633 (N_12633,N_11933,N_11581);
and U12634 (N_12634,N_11493,N_9072);
nor U12635 (N_12635,N_10067,N_9270);
or U12636 (N_12636,N_10827,N_11417);
or U12637 (N_12637,N_10571,N_11118);
and U12638 (N_12638,N_9662,N_11384);
and U12639 (N_12639,N_10000,N_10015);
xor U12640 (N_12640,N_10106,N_9791);
nand U12641 (N_12641,N_9258,N_11309);
or U12642 (N_12642,N_10191,N_10805);
xor U12643 (N_12643,N_9794,N_11838);
or U12644 (N_12644,N_11759,N_11883);
nor U12645 (N_12645,N_9574,N_10957);
nor U12646 (N_12646,N_9729,N_11726);
nor U12647 (N_12647,N_10354,N_9738);
or U12648 (N_12648,N_10342,N_10499);
and U12649 (N_12649,N_11939,N_11442);
and U12650 (N_12650,N_9005,N_11299);
nor U12651 (N_12651,N_11239,N_11246);
nand U12652 (N_12652,N_11037,N_9919);
nor U12653 (N_12653,N_9306,N_11981);
nand U12654 (N_12654,N_10791,N_10057);
nor U12655 (N_12655,N_9815,N_11821);
nor U12656 (N_12656,N_9260,N_10189);
xnor U12657 (N_12657,N_10069,N_11476);
or U12658 (N_12658,N_11502,N_11789);
or U12659 (N_12659,N_10187,N_11224);
nand U12660 (N_12660,N_9589,N_11925);
or U12661 (N_12661,N_10893,N_9797);
nand U12662 (N_12662,N_9231,N_10596);
and U12663 (N_12663,N_10902,N_9583);
or U12664 (N_12664,N_11015,N_11649);
and U12665 (N_12665,N_9176,N_9810);
nand U12666 (N_12666,N_9813,N_11324);
and U12667 (N_12667,N_11117,N_9217);
and U12668 (N_12668,N_9292,N_9402);
or U12669 (N_12669,N_11829,N_9908);
nor U12670 (N_12670,N_11278,N_9281);
and U12671 (N_12671,N_11779,N_10132);
or U12672 (N_12672,N_9398,N_11229);
xor U12673 (N_12673,N_11281,N_9925);
and U12674 (N_12674,N_11430,N_9412);
and U12675 (N_12675,N_10224,N_10146);
and U12676 (N_12676,N_11160,N_11271);
xor U12677 (N_12677,N_10039,N_10585);
or U12678 (N_12678,N_10107,N_10830);
nor U12679 (N_12679,N_10294,N_10921);
xnor U12680 (N_12680,N_9340,N_10740);
xor U12681 (N_12681,N_10261,N_9859);
nor U12682 (N_12682,N_11371,N_9781);
nor U12683 (N_12683,N_10349,N_11457);
and U12684 (N_12684,N_9501,N_10166);
and U12685 (N_12685,N_10028,N_9400);
nand U12686 (N_12686,N_9250,N_10464);
nand U12687 (N_12687,N_9094,N_11227);
or U12688 (N_12688,N_11223,N_11845);
nor U12689 (N_12689,N_10042,N_11056);
xor U12690 (N_12690,N_9936,N_10276);
nand U12691 (N_12691,N_11602,N_11882);
and U12692 (N_12692,N_10742,N_11583);
or U12693 (N_12693,N_9059,N_9681);
and U12694 (N_12694,N_9204,N_9246);
nand U12695 (N_12695,N_9602,N_10875);
xnor U12696 (N_12696,N_10516,N_9041);
or U12697 (N_12697,N_9316,N_9262);
nor U12698 (N_12698,N_9736,N_9379);
nor U12699 (N_12699,N_9687,N_11092);
or U12700 (N_12700,N_10279,N_10828);
and U12701 (N_12701,N_10416,N_9194);
and U12702 (N_12702,N_10235,N_9364);
nand U12703 (N_12703,N_10259,N_11392);
or U12704 (N_12704,N_9450,N_10152);
and U12705 (N_12705,N_9784,N_11636);
nor U12706 (N_12706,N_9652,N_11512);
or U12707 (N_12707,N_10976,N_9203);
xnor U12708 (N_12708,N_11215,N_10907);
nor U12709 (N_12709,N_10205,N_10343);
nand U12710 (N_12710,N_11959,N_10434);
or U12711 (N_12711,N_9628,N_9495);
and U12712 (N_12712,N_9825,N_10862);
or U12713 (N_12713,N_11510,N_9904);
and U12714 (N_12714,N_9661,N_9544);
or U12715 (N_12715,N_11709,N_9634);
or U12716 (N_12716,N_9019,N_11080);
nand U12717 (N_12717,N_9727,N_10675);
or U12718 (N_12718,N_10302,N_9885);
nor U12719 (N_12719,N_9457,N_11729);
or U12720 (N_12720,N_11068,N_11136);
nand U12721 (N_12721,N_11409,N_10977);
and U12722 (N_12722,N_9686,N_10836);
and U12723 (N_12723,N_9943,N_10424);
nor U12724 (N_12724,N_9988,N_11504);
nand U12725 (N_12725,N_11929,N_9082);
or U12726 (N_12726,N_9510,N_11123);
nor U12727 (N_12727,N_11748,N_10815);
and U12728 (N_12728,N_9308,N_9361);
or U12729 (N_12729,N_11640,N_9594);
nand U12730 (N_12730,N_9671,N_10142);
nor U12731 (N_12731,N_11119,N_10053);
nor U12732 (N_12732,N_9900,N_11533);
nand U12733 (N_12733,N_9247,N_9721);
nand U12734 (N_12734,N_10044,N_9201);
xor U12735 (N_12735,N_11919,N_10529);
xnor U12736 (N_12736,N_10656,N_9547);
nor U12737 (N_12737,N_11536,N_9899);
and U12738 (N_12738,N_9955,N_9464);
nand U12739 (N_12739,N_9389,N_9893);
nand U12740 (N_12740,N_9953,N_9324);
or U12741 (N_12741,N_10515,N_11218);
xor U12742 (N_12742,N_10078,N_9463);
xor U12743 (N_12743,N_10565,N_10696);
nand U12744 (N_12744,N_9502,N_10975);
and U12745 (N_12745,N_11617,N_10641);
or U12746 (N_12746,N_11598,N_9816);
nand U12747 (N_12747,N_10887,N_9116);
and U12748 (N_12748,N_11149,N_11506);
or U12749 (N_12749,N_11986,N_9139);
or U12750 (N_12750,N_11242,N_9022);
nor U12751 (N_12751,N_11366,N_10201);
nand U12752 (N_12752,N_9071,N_10777);
and U12753 (N_12753,N_9856,N_11446);
nand U12754 (N_12754,N_11130,N_11330);
nand U12755 (N_12755,N_11293,N_10846);
nand U12756 (N_12756,N_11268,N_9537);
nor U12757 (N_12757,N_11076,N_9866);
xor U12758 (N_12758,N_9683,N_9708);
and U12759 (N_12759,N_9942,N_10915);
nor U12760 (N_12760,N_9403,N_9980);
nand U12761 (N_12761,N_11786,N_11818);
nand U12762 (N_12762,N_11756,N_11739);
xnor U12763 (N_12763,N_9156,N_11263);
or U12764 (N_12764,N_10121,N_11809);
and U12765 (N_12765,N_9545,N_11676);
nor U12766 (N_12766,N_11164,N_11546);
nor U12767 (N_12767,N_11755,N_11796);
or U12768 (N_12768,N_11625,N_11269);
and U12769 (N_12769,N_10741,N_11612);
and U12770 (N_12770,N_11345,N_11084);
and U12771 (N_12771,N_11958,N_9623);
or U12772 (N_12772,N_9758,N_11690);
nor U12773 (N_12773,N_10190,N_9329);
and U12774 (N_12774,N_10913,N_9627);
nand U12775 (N_12775,N_9901,N_10575);
and U12776 (N_12776,N_9771,N_9678);
nor U12777 (N_12777,N_11907,N_11718);
and U12778 (N_12778,N_9563,N_10323);
xnor U12779 (N_12779,N_10544,N_9320);
nand U12780 (N_12780,N_10782,N_9039);
and U12781 (N_12781,N_11940,N_11916);
and U12782 (N_12782,N_9346,N_10485);
nand U12783 (N_12783,N_10865,N_11057);
nor U12784 (N_12784,N_11302,N_9144);
nand U12785 (N_12785,N_10493,N_10026);
and U12786 (N_12786,N_10749,N_9962);
nand U12787 (N_12787,N_11862,N_11481);
or U12788 (N_12788,N_11189,N_10686);
or U12789 (N_12789,N_10657,N_10155);
xor U12790 (N_12790,N_11372,N_10093);
nand U12791 (N_12791,N_10920,N_11795);
or U12792 (N_12792,N_10006,N_9481);
or U12793 (N_12793,N_9489,N_11884);
or U12794 (N_12794,N_10041,N_10183);
nor U12795 (N_12795,N_10200,N_9373);
and U12796 (N_12796,N_11049,N_11575);
and U12797 (N_12797,N_10643,N_10536);
and U12798 (N_12798,N_11401,N_9801);
xnor U12799 (N_12799,N_9060,N_10322);
xor U12800 (N_12800,N_10135,N_11631);
nor U12801 (N_12801,N_11122,N_10265);
nand U12802 (N_12802,N_9874,N_9747);
nand U12803 (N_12803,N_11238,N_9110);
nor U12804 (N_12804,N_11768,N_11601);
or U12805 (N_12805,N_9088,N_11462);
nand U12806 (N_12806,N_11275,N_10440);
xnor U12807 (N_12807,N_10520,N_10174);
and U12808 (N_12808,N_10843,N_10130);
or U12809 (N_12809,N_9641,N_11731);
xnor U12810 (N_12810,N_10234,N_10158);
nor U12811 (N_12811,N_9960,N_10949);
nand U12812 (N_12812,N_11033,N_10979);
nand U12813 (N_12813,N_10923,N_9178);
and U12814 (N_12814,N_9283,N_9497);
xor U12815 (N_12815,N_9717,N_11632);
nor U12816 (N_12816,N_11232,N_10293);
nor U12817 (N_12817,N_11737,N_10128);
and U12818 (N_12818,N_11454,N_9411);
nor U12819 (N_12819,N_11848,N_9048);
or U12820 (N_12820,N_11538,N_9414);
and U12821 (N_12821,N_10812,N_10768);
or U12822 (N_12822,N_10173,N_11579);
or U12823 (N_12823,N_10113,N_11985);
or U12824 (N_12824,N_11839,N_10512);
xnor U12825 (N_12825,N_9601,N_11081);
or U12826 (N_12826,N_9498,N_9640);
or U12827 (N_12827,N_9503,N_9719);
nand U12828 (N_12828,N_10852,N_10968);
and U12829 (N_12829,N_9657,N_9982);
nor U12830 (N_12830,N_11924,N_11703);
xnor U12831 (N_12831,N_9993,N_9305);
and U12832 (N_12832,N_9458,N_11644);
and U12833 (N_12833,N_10534,N_10469);
and U12834 (N_12834,N_9959,N_10429);
nand U12835 (N_12835,N_10236,N_11904);
nand U12836 (N_12836,N_9418,N_9700);
nand U12837 (N_12837,N_11286,N_10172);
nor U12838 (N_12838,N_11589,N_9750);
or U12839 (N_12839,N_10798,N_11306);
or U12840 (N_12840,N_11148,N_11250);
and U12841 (N_12841,N_11174,N_10095);
and U12842 (N_12842,N_9263,N_10519);
nand U12843 (N_12843,N_10599,N_11584);
nor U12844 (N_12844,N_9855,N_10951);
xor U12845 (N_12845,N_11240,N_9367);
and U12846 (N_12846,N_9619,N_9630);
or U12847 (N_12847,N_11521,N_11134);
or U12848 (N_12848,N_11316,N_9304);
and U12849 (N_12849,N_11934,N_10232);
nand U12850 (N_12850,N_10514,N_10993);
and U12851 (N_12851,N_9562,N_11941);
xor U12852 (N_12852,N_11713,N_11975);
nor U12853 (N_12853,N_11217,N_10013);
nand U12854 (N_12854,N_9380,N_9287);
nand U12855 (N_12855,N_9166,N_9420);
and U12856 (N_12856,N_10507,N_9964);
nand U12857 (N_12857,N_11168,N_9417);
xor U12858 (N_12858,N_9104,N_11633);
nand U12859 (N_12859,N_9726,N_10420);
or U12860 (N_12860,N_11570,N_10929);
or U12861 (N_12861,N_10869,N_10202);
nor U12862 (N_12862,N_9679,N_9843);
nor U12863 (N_12863,N_11331,N_11115);
and U12864 (N_12864,N_10943,N_10277);
nand U12865 (N_12865,N_9930,N_11220);
nor U12866 (N_12866,N_9106,N_11659);
and U12867 (N_12867,N_11191,N_11951);
nand U12868 (N_12868,N_11061,N_9033);
nand U12869 (N_12869,N_11437,N_9368);
or U12870 (N_12870,N_11518,N_10802);
nand U12871 (N_12871,N_11585,N_11853);
or U12872 (N_12872,N_10963,N_10933);
and U12873 (N_12873,N_10001,N_10770);
and U12874 (N_12874,N_11794,N_10932);
nand U12875 (N_12875,N_10560,N_9164);
xnor U12876 (N_12876,N_11103,N_10649);
or U12877 (N_12877,N_11424,N_11622);
and U12878 (N_12878,N_10487,N_10936);
or U12879 (N_12879,N_11490,N_10950);
nand U12880 (N_12880,N_9526,N_10579);
xnor U12881 (N_12881,N_10437,N_11567);
nand U12882 (N_12882,N_11325,N_9109);
nor U12883 (N_12883,N_10396,N_11950);
nor U12884 (N_12884,N_10877,N_9462);
or U12885 (N_12885,N_10764,N_10461);
nor U12886 (N_12886,N_11528,N_10669);
nor U12887 (N_12887,N_9291,N_11151);
or U12888 (N_12888,N_11167,N_9968);
or U12889 (N_12889,N_9334,N_11062);
and U12890 (N_12890,N_9894,N_9421);
and U12891 (N_12891,N_9637,N_10771);
nand U12892 (N_12892,N_10628,N_10251);
nor U12893 (N_12893,N_11776,N_10685);
nand U12894 (N_12894,N_9393,N_10411);
nand U12895 (N_12895,N_9767,N_11006);
nor U12896 (N_12896,N_10626,N_11428);
or U12897 (N_12897,N_10417,N_10816);
or U12898 (N_12898,N_10022,N_10446);
and U12899 (N_12899,N_9046,N_9552);
nand U12900 (N_12900,N_10650,N_10953);
and U12901 (N_12901,N_9200,N_11545);
nor U12902 (N_12902,N_11420,N_9514);
nor U12903 (N_12903,N_11923,N_11629);
or U12904 (N_12904,N_9590,N_11335);
and U12905 (N_12905,N_11700,N_9989);
nor U12906 (N_12906,N_9023,N_10393);
nand U12907 (N_12907,N_9913,N_11063);
or U12908 (N_12908,N_11859,N_11717);
and U12909 (N_12909,N_11716,N_11780);
and U12910 (N_12910,N_10648,N_10483);
nand U12911 (N_12911,N_11577,N_10717);
or U12912 (N_12912,N_10306,N_10210);
xnor U12913 (N_12913,N_10032,N_10974);
or U12914 (N_12914,N_10367,N_11007);
nor U12915 (N_12915,N_11255,N_11720);
or U12916 (N_12916,N_9969,N_10242);
xor U12917 (N_12917,N_10012,N_9667);
nand U12918 (N_12918,N_11694,N_11750);
nor U12919 (N_12919,N_11203,N_9118);
and U12920 (N_12920,N_11928,N_11093);
nor U12921 (N_12921,N_11097,N_9769);
nor U12922 (N_12922,N_10070,N_10089);
and U12923 (N_12923,N_11178,N_9586);
nor U12924 (N_12924,N_9474,N_11927);
xor U12925 (N_12925,N_11282,N_11591);
nand U12926 (N_12926,N_10310,N_10298);
or U12927 (N_12927,N_10247,N_9692);
or U12928 (N_12928,N_10731,N_11376);
or U12929 (N_12929,N_9385,N_10081);
nand U12930 (N_12930,N_9554,N_10704);
nor U12931 (N_12931,N_10899,N_10045);
or U12932 (N_12932,N_9907,N_10620);
or U12933 (N_12933,N_9846,N_11945);
nor U12934 (N_12934,N_10062,N_9294);
and U12935 (N_12935,N_10412,N_11236);
nand U12936 (N_12936,N_9244,N_9718);
nand U12937 (N_12937,N_10587,N_11791);
and U12938 (N_12938,N_11059,N_10605);
nand U12939 (N_12939,N_11086,N_9272);
and U12940 (N_12940,N_10097,N_9438);
nor U12941 (N_12941,N_10181,N_10905);
and U12942 (N_12942,N_9858,N_10075);
or U12943 (N_12943,N_11728,N_9220);
or U12944 (N_12944,N_11354,N_11867);
and U12945 (N_12945,N_11407,N_11101);
and U12946 (N_12946,N_10384,N_9725);
or U12947 (N_12947,N_9940,N_11112);
and U12948 (N_12948,N_9929,N_9539);
nor U12949 (N_12949,N_10569,N_9030);
nand U12950 (N_12950,N_9530,N_11847);
nand U12951 (N_12951,N_9453,N_9321);
or U12952 (N_12952,N_11370,N_9997);
and U12953 (N_12953,N_11342,N_10796);
and U12954 (N_12954,N_10723,N_10752);
nor U12955 (N_12955,N_10988,N_11020);
nor U12956 (N_12956,N_11402,N_11761);
nand U12957 (N_12957,N_10245,N_10355);
and U12958 (N_12958,N_11436,N_11495);
xor U12959 (N_12959,N_10718,N_11106);
nor U12960 (N_12960,N_9808,N_11802);
xnor U12961 (N_12961,N_10799,N_9160);
nand U12962 (N_12962,N_11475,N_10506);
xor U12963 (N_12963,N_9127,N_9218);
nand U12964 (N_12964,N_10337,N_10866);
and U12965 (N_12965,N_9629,N_11827);
and U12966 (N_12966,N_10180,N_11500);
xor U12967 (N_12967,N_11749,N_9049);
nor U12968 (N_12968,N_11290,N_11874);
nand U12969 (N_12969,N_10602,N_9624);
or U12970 (N_12970,N_11677,N_9796);
nor U12971 (N_12971,N_9424,N_10208);
xor U12972 (N_12972,N_10593,N_10582);
and U12973 (N_12973,N_10318,N_10372);
nor U12974 (N_12974,N_9120,N_9360);
and U12975 (N_12975,N_9370,N_9979);
nand U12976 (N_12976,N_10631,N_9351);
nor U12977 (N_12977,N_9447,N_9074);
or U12978 (N_12978,N_10663,N_10123);
nor U12979 (N_12979,N_11364,N_9485);
nor U12980 (N_12980,N_9540,N_11688);
nor U12981 (N_12981,N_11873,N_11154);
nor U12982 (N_12982,N_11834,N_9689);
nand U12983 (N_12983,N_10480,N_9365);
xnor U12984 (N_12984,N_9519,N_9097);
or U12985 (N_12985,N_9013,N_11329);
and U12986 (N_12986,N_9000,N_9135);
nand U12987 (N_12987,N_11222,N_11674);
nand U12988 (N_12988,N_11962,N_9970);
nor U12989 (N_12989,N_10473,N_10679);
nand U12990 (N_12990,N_10019,N_9958);
or U12991 (N_12991,N_9429,N_10636);
nor U12992 (N_12992,N_9440,N_9196);
nand U12993 (N_12993,N_11156,N_10496);
nor U12994 (N_12994,N_9415,N_9806);
and U12995 (N_12995,N_11298,N_10838);
nand U12996 (N_12996,N_11089,N_9536);
and U12997 (N_12997,N_9492,N_10178);
nand U12998 (N_12998,N_10955,N_9090);
or U12999 (N_12999,N_10304,N_9257);
and U13000 (N_13000,N_10096,N_9649);
nor U13001 (N_13001,N_10143,N_10503);
nor U13002 (N_13002,N_9541,N_10233);
or U13003 (N_13003,N_11011,N_9606);
or U13004 (N_13004,N_9195,N_9735);
nand U13005 (N_13005,N_11195,N_9174);
nor U13006 (N_13006,N_10244,N_10410);
and U13007 (N_13007,N_11651,N_9564);
and U13008 (N_13008,N_11451,N_11947);
nor U13009 (N_13009,N_9891,N_9621);
or U13010 (N_13010,N_9478,N_11360);
xnor U13011 (N_13011,N_10644,N_10465);
and U13012 (N_13012,N_9288,N_9300);
and U13013 (N_13013,N_10364,N_11996);
nand U13014 (N_13014,N_9333,N_10010);
nand U13015 (N_13015,N_9922,N_9712);
nand U13016 (N_13016,N_9348,N_10699);
or U13017 (N_13017,N_10719,N_9375);
nor U13018 (N_13018,N_9570,N_9449);
nor U13019 (N_13019,N_9595,N_10634);
nand U13020 (N_13020,N_9468,N_9651);
and U13021 (N_13021,N_11773,N_10700);
and U13022 (N_13022,N_10212,N_9381);
nor U13023 (N_13023,N_11646,N_10961);
or U13024 (N_13024,N_11943,N_9954);
nand U13025 (N_13025,N_10495,N_10332);
xor U13026 (N_13026,N_10567,N_11944);
and U13027 (N_13027,N_11234,N_9600);
xnor U13028 (N_13028,N_9905,N_10578);
nand U13029 (N_13029,N_11172,N_10790);
xnor U13030 (N_13030,N_11635,N_9405);
nor U13031 (N_13031,N_11764,N_9832);
or U13032 (N_13032,N_11208,N_11658);
or U13033 (N_13033,N_11913,N_11551);
xnor U13034 (N_13034,N_11216,N_11863);
and U13035 (N_13035,N_11819,N_11264);
nand U13036 (N_13036,N_9395,N_9490);
nor U13037 (N_13037,N_10786,N_9838);
and U13038 (N_13038,N_9828,N_9532);
nand U13039 (N_13039,N_11095,N_10729);
nor U13040 (N_13040,N_10916,N_9055);
or U13041 (N_13041,N_11909,N_9798);
and U13042 (N_13042,N_11578,N_9728);
and U13043 (N_13043,N_9394,N_9274);
nor U13044 (N_13044,N_11643,N_11198);
and U13045 (N_13045,N_11813,N_9455);
or U13046 (N_13046,N_10478,N_11477);
and U13047 (N_13047,N_11807,N_9021);
nand U13048 (N_13048,N_10682,N_11332);
or U13049 (N_13049,N_9326,N_11127);
nor U13050 (N_13050,N_11997,N_10061);
or U13051 (N_13051,N_11350,N_11614);
nor U13052 (N_13052,N_9280,N_9555);
nand U13053 (N_13053,N_11917,N_11158);
nor U13054 (N_13054,N_9151,N_9639);
or U13055 (N_13055,N_9527,N_10725);
or U13056 (N_13056,N_10230,N_9578);
or U13057 (N_13057,N_10651,N_10966);
nand U13058 (N_13058,N_11900,N_11667);
nand U13059 (N_13059,N_11177,N_9423);
xnor U13060 (N_13060,N_11279,N_10248);
nor U13061 (N_13061,N_10427,N_9408);
and U13062 (N_13062,N_11757,N_11102);
or U13063 (N_13063,N_10662,N_10255);
nand U13064 (N_13064,N_11091,N_10583);
xor U13065 (N_13065,N_10508,N_10229);
nor U13066 (N_13066,N_10617,N_10607);
nor U13067 (N_13067,N_10504,N_9948);
nand U13068 (N_13068,N_9190,N_10772);
and U13069 (N_13069,N_11204,N_10572);
nand U13070 (N_13070,N_9499,N_10176);
nand U13071 (N_13071,N_10383,N_10860);
and U13072 (N_13072,N_9465,N_9344);
and U13073 (N_13073,N_9444,N_10091);
nor U13074 (N_13074,N_11983,N_11730);
nand U13075 (N_13075,N_9787,N_11778);
or U13076 (N_13076,N_11627,N_11735);
and U13077 (N_13077,N_10604,N_10387);
and U13078 (N_13078,N_10645,N_10600);
and U13079 (N_13079,N_11048,N_10455);
nor U13080 (N_13080,N_11587,N_9112);
nor U13081 (N_13081,N_10312,N_11074);
nor U13082 (N_13082,N_11125,N_10240);
nand U13083 (N_13083,N_9014,N_9827);
nand U13084 (N_13084,N_10284,N_9186);
nand U13085 (N_13085,N_9439,N_9284);
nand U13086 (N_13086,N_9314,N_10879);
and U13087 (N_13087,N_11630,N_10738);
and U13088 (N_13088,N_10911,N_11415);
or U13089 (N_13089,N_10436,N_11176);
and U13090 (N_13090,N_10359,N_10673);
or U13091 (N_13091,N_11806,N_9865);
nor U13092 (N_13092,N_9331,N_10746);
and U13093 (N_13093,N_9867,N_10737);
or U13094 (N_13094,N_10872,N_10562);
or U13095 (N_13095,N_9533,N_10934);
nor U13096 (N_13096,N_10035,N_11875);
or U13097 (N_13097,N_10280,N_9972);
nor U13098 (N_13098,N_11665,N_9741);
xnor U13099 (N_13099,N_11055,N_9999);
xor U13100 (N_13100,N_11248,N_10972);
xnor U13101 (N_13101,N_11647,N_11247);
and U13102 (N_13102,N_10689,N_9278);
nor U13103 (N_13103,N_9459,N_10670);
or U13104 (N_13104,N_10441,N_10751);
nand U13105 (N_13105,N_11143,N_9058);
or U13106 (N_13106,N_10419,N_10658);
xnor U13107 (N_13107,N_11153,N_9659);
nand U13108 (N_13108,N_11600,N_10033);
nand U13109 (N_13109,N_9469,N_11336);
and U13110 (N_13110,N_9618,N_11449);
nand U13111 (N_13111,N_9239,N_10543);
and U13112 (N_13112,N_11274,N_10023);
nor U13113 (N_13113,N_10144,N_9862);
or U13114 (N_13114,N_9044,N_11790);
nor U13115 (N_13115,N_11972,N_11314);
or U13116 (N_13116,N_11529,N_10653);
xor U13117 (N_13117,N_11429,N_10809);
nand U13118 (N_13118,N_10613,N_10231);
nand U13119 (N_13119,N_9296,N_11340);
and U13120 (N_13120,N_11912,N_10083);
and U13121 (N_13121,N_9680,N_11077);
and U13122 (N_13122,N_9313,N_11414);
or U13123 (N_13123,N_10105,N_9147);
xnor U13124 (N_13124,N_11291,N_11803);
nor U13125 (N_13125,N_9205,N_10370);
nor U13126 (N_13126,N_10709,N_9535);
nor U13127 (N_13127,N_10873,N_10037);
and U13128 (N_13128,N_9992,N_10517);
and U13129 (N_13129,N_11310,N_10646);
or U13130 (N_13130,N_10472,N_10394);
nand U13131 (N_13131,N_10141,N_11535);
or U13132 (N_13132,N_10927,N_9576);
and U13133 (N_13133,N_11479,N_10677);
nor U13134 (N_13134,N_10169,N_9267);
nand U13135 (N_13135,N_11555,N_11205);
or U13136 (N_13136,N_11508,N_10697);
and U13137 (N_13137,N_11722,N_11365);
and U13138 (N_13138,N_10788,N_10824);
nand U13139 (N_13139,N_11004,N_10910);
or U13140 (N_13140,N_10687,N_11920);
and U13141 (N_13141,N_10990,N_9376);
xor U13142 (N_13142,N_10007,N_9303);
nor U13143 (N_13143,N_10937,N_11113);
nor U13144 (N_13144,N_11539,N_11041);
xnor U13145 (N_13145,N_11723,N_10892);
xnor U13146 (N_13146,N_11355,N_9917);
or U13147 (N_13147,N_10421,N_9076);
nand U13148 (N_13148,N_11568,N_11053);
nand U13149 (N_13149,N_11180,N_11434);
nand U13150 (N_13150,N_9593,N_11881);
or U13151 (N_13151,N_9568,N_11321);
nand U13152 (N_13152,N_11523,N_11432);
and U13153 (N_13153,N_9170,N_9227);
and U13154 (N_13154,N_9243,N_9937);
or U13155 (N_13155,N_10826,N_9070);
xor U13156 (N_13156,N_9854,N_11254);
xnor U13157 (N_13157,N_11054,N_11561);
nand U13158 (N_13158,N_11893,N_10292);
and U13159 (N_13159,N_10969,N_10184);
or U13160 (N_13160,N_9625,N_9445);
nand U13161 (N_13161,N_9638,N_10522);
or U13162 (N_13162,N_11971,N_11530);
and U13163 (N_13163,N_11990,N_10851);
nand U13164 (N_13164,N_10430,N_10350);
or U13165 (N_13165,N_9446,N_9371);
or U13166 (N_13166,N_10871,N_11201);
or U13167 (N_13167,N_11711,N_9045);
nor U13168 (N_13168,N_10407,N_11046);
or U13169 (N_13169,N_11792,N_11865);
and U13170 (N_13170,N_11277,N_9350);
nand U13171 (N_13171,N_10789,N_11256);
nor U13172 (N_13172,N_11681,N_9612);
or U13173 (N_13173,N_9561,N_9461);
and U13174 (N_13174,N_11258,N_10400);
nand U13175 (N_13175,N_11936,N_11655);
nand U13176 (N_13176,N_9276,N_11615);
or U13177 (N_13177,N_11029,N_9001);
or U13178 (N_13178,N_9837,N_11431);
nor U13179 (N_13179,N_10466,N_10211);
or U13180 (N_13180,N_9793,N_10535);
or U13181 (N_13181,N_11770,N_10784);
nand U13182 (N_13182,N_10867,N_11285);
and U13183 (N_13183,N_11879,N_9688);
xor U13184 (N_13184,N_9740,N_11856);
nor U13185 (N_13185,N_11266,N_10065);
and U13186 (N_13186,N_11608,N_9277);
nand U13187 (N_13187,N_10005,N_10418);
and U13188 (N_13188,N_9123,N_10655);
or U13189 (N_13189,N_9884,N_9182);
or U13190 (N_13190,N_11071,N_11814);
and U13191 (N_13191,N_10286,N_9211);
nand U13192 (N_13192,N_10568,N_10728);
nor U13193 (N_13193,N_9580,N_10433);
xor U13194 (N_13194,N_11114,N_11548);
nand U13195 (N_13195,N_9584,N_11811);
xnor U13196 (N_13196,N_10765,N_11244);
or U13197 (N_13197,N_10842,N_10794);
or U13198 (N_13198,N_10564,N_9482);
nand U13199 (N_13199,N_11825,N_11419);
and U13200 (N_13200,N_9441,N_11922);
and U13201 (N_13201,N_10991,N_9742);
or U13202 (N_13202,N_11606,N_10539);
and U13203 (N_13203,N_9358,N_11173);
nand U13204 (N_13204,N_10301,N_11588);
and U13205 (N_13205,N_11199,N_9434);
nand U13206 (N_13206,N_10030,N_9161);
nand U13207 (N_13207,N_10642,N_9863);
nor U13208 (N_13208,N_9248,N_9777);
and U13209 (N_13209,N_9159,N_9237);
and U13210 (N_13210,N_11804,N_9695);
and U13211 (N_13211,N_9966,N_11369);
nor U13212 (N_13212,N_10980,N_11926);
and U13213 (N_13213,N_11503,N_11994);
xor U13214 (N_13214,N_11620,N_10940);
and U13215 (N_13215,N_9476,N_9011);
and U13216 (N_13216,N_9775,N_10119);
nor U13217 (N_13217,N_9099,N_11894);
nand U13218 (N_13218,N_11030,N_11777);
or U13219 (N_13219,N_11557,N_11463);
or U13220 (N_13220,N_9103,N_10625);
and U13221 (N_13221,N_10127,N_9472);
nand U13222 (N_13222,N_9488,N_10137);
nor U13223 (N_13223,N_9587,N_10521);
or U13224 (N_13224,N_11698,N_11835);
and U13225 (N_13225,N_11380,N_10549);
nand U13226 (N_13226,N_9807,N_11210);
nand U13227 (N_13227,N_11520,N_11836);
and U13228 (N_13228,N_11714,N_10888);
nor U13229 (N_13229,N_11656,N_11685);
xor U13230 (N_13230,N_11992,N_10330);
or U13231 (N_13231,N_11979,N_11438);
and U13232 (N_13232,N_10847,N_9644);
nand U13233 (N_13233,N_10667,N_11200);
nand U13234 (N_13234,N_9505,N_10432);
or U13235 (N_13235,N_9829,N_10316);
or U13236 (N_13236,N_11348,N_10336);
nand U13237 (N_13237,N_9406,N_11905);
xnor U13238 (N_13238,N_11628,N_9800);
and U13239 (N_13239,N_9749,N_10082);
nor U13240 (N_13240,N_10896,N_9542);
nand U13241 (N_13241,N_11544,N_11341);
and U13242 (N_13242,N_10580,N_9154);
and U13243 (N_13243,N_9025,N_11738);
and U13244 (N_13244,N_10720,N_11891);
xnor U13245 (N_13245,N_9990,N_10500);
nor U13246 (N_13246,N_10692,N_9819);
nor U13247 (N_13247,N_9672,N_11664);
xnor U13248 (N_13248,N_9889,N_10841);
and U13249 (N_13249,N_10757,N_9275);
or U13250 (N_13250,N_10198,N_10707);
and U13251 (N_13251,N_9734,N_10156);
nand U13252 (N_13252,N_9877,N_11817);
nor U13253 (N_13253,N_11186,N_11724);
and U13254 (N_13254,N_9902,N_9383);
or U13255 (N_13255,N_10938,N_11043);
xnor U13256 (N_13256,N_11914,N_10031);
nand U13257 (N_13257,N_10595,N_11547);
or U13258 (N_13258,N_9162,N_10413);
nand U13259 (N_13259,N_10538,N_9410);
nand U13260 (N_13260,N_10448,N_10622);
nor U13261 (N_13261,N_9042,N_9509);
nand U13262 (N_13262,N_9938,N_10112);
xor U13263 (N_13263,N_11184,N_9860);
xor U13264 (N_13264,N_11980,N_9883);
nand U13265 (N_13265,N_9279,N_10376);
nand U13266 (N_13266,N_10944,N_11915);
xor U13267 (N_13267,N_9255,N_10710);
nand U13268 (N_13268,N_11961,N_11251);
or U13269 (N_13269,N_10085,N_11774);
nand U13270 (N_13270,N_11752,N_10467);
nand U13271 (N_13271,N_10088,N_10678);
and U13272 (N_13272,N_10369,N_11138);
nand U13273 (N_13273,N_9098,N_11831);
or U13274 (N_13274,N_10629,N_11045);
nor U13275 (N_13275,N_11526,N_9456);
nand U13276 (N_13276,N_9425,N_10101);
or U13277 (N_13277,N_11642,N_9631);
and U13278 (N_13278,N_9437,N_9850);
nand U13279 (N_13279,N_9610,N_10783);
xor U13280 (N_13280,N_10839,N_11537);
and U13281 (N_13281,N_11541,N_10999);
and U13282 (N_13282,N_11391,N_11948);
or U13283 (N_13283,N_11039,N_9914);
and U13284 (N_13284,N_11712,N_9134);
and U13285 (N_13285,N_10415,N_11511);
nor U13286 (N_13286,N_9732,N_9500);
and U13287 (N_13287,N_10552,N_11662);
or U13288 (N_13288,N_11289,N_10995);
and U13289 (N_13289,N_9124,N_9665);
nor U13290 (N_13290,N_11363,N_9836);
nor U13291 (N_13291,N_10249,N_10891);
nand U13292 (N_13292,N_11543,N_9701);
nor U13293 (N_13293,N_11564,N_10926);
and U13294 (N_13294,N_10262,N_10864);
nand U13295 (N_13295,N_11196,N_11031);
nor U13296 (N_13296,N_10511,N_9897);
or U13297 (N_13297,N_10853,N_11294);
or U13298 (N_13298,N_11237,N_10760);
and U13299 (N_13299,N_10118,N_11559);
xnor U13300 (N_13300,N_10314,N_9117);
nor U13301 (N_13301,N_11296,N_11740);
nand U13302 (N_13302,N_11448,N_11849);
and U13303 (N_13303,N_9335,N_11590);
nand U13304 (N_13304,N_9512,N_9765);
and U13305 (N_13305,N_11027,N_11161);
nand U13306 (N_13306,N_9707,N_11304);
and U13307 (N_13307,N_10638,N_10931);
nand U13308 (N_13308,N_10147,N_9115);
and U13309 (N_13309,N_9264,N_9018);
xor U13310 (N_13310,N_9027,N_9436);
nand U13311 (N_13311,N_10825,N_10164);
nor U13312 (N_13312,N_10454,N_11534);
or U13313 (N_13313,N_11976,N_9861);
nand U13314 (N_13314,N_10848,N_11411);
nand U13315 (N_13315,N_11960,N_9770);
nand U13316 (N_13316,N_9038,N_10778);
and U13317 (N_13317,N_10870,N_10073);
and U13318 (N_13318,N_10615,N_10029);
or U13319 (N_13319,N_9579,N_10287);
or U13320 (N_13320,N_9845,N_10325);
nor U13321 (N_13321,N_10573,N_9898);
or U13322 (N_13322,N_10691,N_10025);
nand U13323 (N_13323,N_11163,N_9653);
nor U13324 (N_13324,N_9163,N_9691);
and U13325 (N_13325,N_9345,N_9525);
nand U13326 (N_13326,N_9976,N_10227);
or U13327 (N_13327,N_11550,N_11973);
nand U13328 (N_13328,N_11702,N_9675);
nand U13329 (N_13329,N_11147,N_11235);
nor U13330 (N_13330,N_9945,N_10928);
or U13331 (N_13331,N_9265,N_10366);
and U13332 (N_13332,N_10347,N_11641);
nor U13333 (N_13333,N_10619,N_11846);
nand U13334 (N_13334,N_9521,N_11910);
xor U13335 (N_13335,N_11179,N_11450);
nand U13336 (N_13336,N_11964,N_11338);
xor U13337 (N_13337,N_10688,N_11297);
nor U13338 (N_13338,N_11868,N_10390);
or U13339 (N_13339,N_10530,N_9427);
or U13340 (N_13340,N_10163,N_11571);
or U13341 (N_13341,N_9932,N_9047);
or U13342 (N_13342,N_10058,N_10800);
or U13343 (N_13343,N_9543,N_10598);
or U13344 (N_13344,N_10698,N_10468);
and U13345 (N_13345,N_10553,N_10197);
nand U13346 (N_13346,N_10721,N_9748);
nand U13347 (N_13347,N_11599,N_9008);
and U13348 (N_13348,N_10120,N_11876);
and U13349 (N_13349,N_10981,N_10324);
or U13350 (N_13350,N_10918,N_9426);
and U13351 (N_13351,N_11378,N_9493);
nor U13352 (N_13352,N_9496,N_11880);
nor U13353 (N_13353,N_11751,N_11108);
xor U13354 (N_13354,N_10724,N_10399);
and U13355 (N_13355,N_11669,N_10947);
nor U13356 (N_13356,N_10177,N_11663);
or U13357 (N_13357,N_9477,N_9596);
nor U13358 (N_13358,N_11679,N_9875);
or U13359 (N_13359,N_9668,N_11349);
nand U13360 (N_13360,N_10309,N_9697);
and U13361 (N_13361,N_11318,N_10785);
and U13362 (N_13362,N_10379,N_9236);
nand U13363 (N_13363,N_11144,N_10431);
nor U13364 (N_13364,N_9965,N_11249);
nand U13365 (N_13365,N_11611,N_11474);
or U13366 (N_13366,N_10965,N_11826);
nor U13367 (N_13367,N_9737,N_11085);
and U13368 (N_13368,N_9352,N_10732);
and U13369 (N_13369,N_10883,N_9714);
or U13370 (N_13370,N_11621,N_9095);
or U13371 (N_13371,N_11064,N_10194);
and U13372 (N_13372,N_10588,N_10358);
and U13373 (N_13373,N_11989,N_11038);
nand U13374 (N_13374,N_11952,N_9029);
xnor U13375 (N_13375,N_10603,N_9028);
nand U13376 (N_13376,N_10632,N_10510);
and U13377 (N_13377,N_9952,N_11120);
xor U13378 (N_13378,N_10959,N_11733);
and U13379 (N_13379,N_9921,N_9882);
nor U13380 (N_13380,N_9873,N_11473);
and U13381 (N_13381,N_10103,N_10591);
nor U13382 (N_13382,N_9694,N_10683);
and U13383 (N_13383,N_10404,N_9887);
nand U13384 (N_13384,N_10935,N_11193);
nor U13385 (N_13385,N_9382,N_11878);
or U13386 (N_13386,N_10566,N_10131);
and U13387 (N_13387,N_10328,N_9723);
and U13388 (N_13388,N_9309,N_11840);
and U13389 (N_13389,N_10736,N_10681);
and U13390 (N_13390,N_11580,N_10391);
xor U13391 (N_13391,N_10618,N_9295);
and U13392 (N_13392,N_10946,N_10861);
and U13393 (N_13393,N_11005,N_11426);
nand U13394 (N_13394,N_9591,N_10406);
and U13395 (N_13395,N_10428,N_9148);
xor U13396 (N_13396,N_10898,N_10481);
or U13397 (N_13397,N_9307,N_9372);
nor U13398 (N_13398,N_11361,N_9517);
and U13399 (N_13399,N_10457,N_11028);
nor U13400 (N_13400,N_9105,N_9635);
nand U13401 (N_13401,N_11022,N_10024);
nand U13402 (N_13402,N_11374,N_9315);
nand U13403 (N_13403,N_9626,N_11532);
nor U13404 (N_13404,N_9388,N_10818);
nor U13405 (N_13405,N_9216,N_9396);
nand U13406 (N_13406,N_9762,N_10346);
and U13407 (N_13407,N_9804,N_11721);
xnor U13408 (N_13408,N_9609,N_10442);
or U13409 (N_13409,N_10474,N_11141);
or U13410 (N_13410,N_9903,N_10750);
or U13411 (N_13411,N_11079,N_9391);
or U13412 (N_13412,N_10895,N_9763);
nand U13413 (N_13413,N_11132,N_10769);
and U13414 (N_13414,N_9912,N_11788);
or U13415 (N_13415,N_11267,N_10296);
or U13416 (N_13416,N_10904,N_10038);
and U13417 (N_13417,N_9565,N_10528);
and U13418 (N_13418,N_9230,N_10531);
nand U13419 (N_13419,N_11706,N_9392);
nor U13420 (N_13420,N_10900,N_9751);
and U13421 (N_13421,N_9674,N_11126);
nor U13422 (N_13422,N_10443,N_9223);
or U13423 (N_13423,N_11090,N_11610);
nor U13424 (N_13424,N_10380,N_10647);
nor U13425 (N_13425,N_11820,N_11828);
nand U13426 (N_13426,N_11775,N_11243);
nor U13427 (N_13427,N_9155,N_11379);
or U13428 (N_13428,N_11758,N_11852);
nor U13429 (N_13429,N_9225,N_10021);
xor U13430 (N_13430,N_9946,N_10068);
and U13431 (N_13431,N_10489,N_10283);
nor U13432 (N_13432,N_10402,N_10611);
or U13433 (N_13433,N_9983,N_9167);
and U13434 (N_13434,N_11682,N_9073);
nor U13435 (N_13435,N_10498,N_9180);
nand U13436 (N_13436,N_9487,N_9199);
or U13437 (N_13437,N_11351,N_11352);
nor U13438 (N_13438,N_9967,N_9931);
nor U13439 (N_13439,N_11096,N_11000);
and U13440 (N_13440,N_10290,N_11830);
xor U13441 (N_13441,N_9390,N_10849);
nand U13442 (N_13442,N_9355,N_10509);
and U13443 (N_13443,N_10160,N_11292);
nor U13444 (N_13444,N_9756,N_10833);
nand U13445 (N_13445,N_9165,N_10307);
nor U13446 (N_13446,N_9906,N_9086);
xor U13447 (N_13447,N_10462,N_11357);
and U13448 (N_13448,N_9730,N_11563);
nor U13449 (N_13449,N_9617,N_11328);
xor U13450 (N_13450,N_11383,N_9480);
and U13451 (N_13451,N_11483,N_9957);
and U13452 (N_13452,N_11433,N_9080);
nand U13453 (N_13453,N_11954,N_9293);
or U13454 (N_13454,N_9185,N_11671);
xnor U13455 (N_13455,N_10452,N_9214);
and U13456 (N_13456,N_10203,N_11897);
xnor U13457 (N_13457,N_10621,N_9975);
nand U13458 (N_13458,N_11515,N_11693);
nand U13459 (N_13459,N_9956,N_11116);
nand U13460 (N_13460,N_10374,N_10036);
and U13461 (N_13461,N_10834,N_11505);
xor U13462 (N_13462,N_9317,N_10159);
nor U13463 (N_13463,N_11303,N_9886);
or U13464 (N_13464,N_10554,N_10401);
nand U13465 (N_13465,N_9704,N_10080);
and U13466 (N_13466,N_9724,N_9460);
or U13467 (N_13467,N_9998,N_10329);
or U13468 (N_13468,N_9910,N_11121);
and U13469 (N_13469,N_9795,N_10821);
nand U13470 (N_13470,N_11444,N_9003);
or U13471 (N_13471,N_10063,N_11386);
or U13472 (N_13472,N_9677,N_9145);
or U13473 (N_13473,N_11719,N_11793);
nand U13474 (N_13474,N_9506,N_10810);
nor U13475 (N_13475,N_9245,N_10047);
or U13476 (N_13476,N_10780,N_9582);
nor U13477 (N_13477,N_11183,N_10339);
or U13478 (N_13478,N_9876,N_10445);
and U13479 (N_13479,N_11691,N_11558);
nand U13480 (N_13480,N_11732,N_11042);
xnor U13481 (N_13481,N_11466,N_9805);
and U13482 (N_13482,N_9766,N_9067);
or U13483 (N_13483,N_10054,N_11100);
nor U13484 (N_13484,N_9896,N_9507);
nor U13485 (N_13485,N_11408,N_9451);
nand U13486 (N_13486,N_11333,N_10715);
xnor U13487 (N_13487,N_11069,N_9137);
nor U13488 (N_13488,N_10726,N_11634);
nand U13489 (N_13489,N_11099,N_9404);
and U13490 (N_13490,N_11403,N_11892);
or U13491 (N_13491,N_11387,N_9020);
xor U13492 (N_13492,N_10906,N_10002);
nand U13493 (N_13493,N_10344,N_10627);
or U13494 (N_13494,N_10781,N_10711);
nor U13495 (N_13495,N_11573,N_10046);
and U13496 (N_13496,N_10761,N_10305);
nor U13497 (N_13497,N_9409,N_9918);
nor U13498 (N_13498,N_10423,N_10291);
and U13499 (N_13499,N_10064,N_11654);
nand U13500 (N_13500,N_11258,N_11288);
or U13501 (N_13501,N_9119,N_10534);
nand U13502 (N_13502,N_9102,N_9023);
nor U13503 (N_13503,N_9735,N_11687);
nand U13504 (N_13504,N_10357,N_11526);
or U13505 (N_13505,N_9284,N_11072);
and U13506 (N_13506,N_10379,N_11573);
or U13507 (N_13507,N_9140,N_11507);
nor U13508 (N_13508,N_11911,N_10574);
and U13509 (N_13509,N_11845,N_11556);
nor U13510 (N_13510,N_10639,N_11811);
nor U13511 (N_13511,N_9289,N_11244);
and U13512 (N_13512,N_11937,N_11827);
or U13513 (N_13513,N_10631,N_10714);
nand U13514 (N_13514,N_11696,N_9938);
and U13515 (N_13515,N_9921,N_11242);
or U13516 (N_13516,N_10278,N_11096);
nand U13517 (N_13517,N_10600,N_10474);
and U13518 (N_13518,N_11935,N_11500);
and U13519 (N_13519,N_10481,N_11234);
nand U13520 (N_13520,N_9128,N_10546);
and U13521 (N_13521,N_11875,N_10261);
nor U13522 (N_13522,N_11268,N_10262);
nand U13523 (N_13523,N_10290,N_11992);
or U13524 (N_13524,N_11782,N_11526);
nor U13525 (N_13525,N_11387,N_9919);
or U13526 (N_13526,N_9424,N_11099);
xor U13527 (N_13527,N_10321,N_9469);
and U13528 (N_13528,N_9647,N_11552);
and U13529 (N_13529,N_9325,N_10659);
nor U13530 (N_13530,N_10926,N_11465);
nand U13531 (N_13531,N_9665,N_11895);
or U13532 (N_13532,N_10695,N_9424);
or U13533 (N_13533,N_11775,N_10031);
and U13534 (N_13534,N_9700,N_11424);
and U13535 (N_13535,N_10057,N_9496);
or U13536 (N_13536,N_10126,N_10125);
and U13537 (N_13537,N_9651,N_10792);
nor U13538 (N_13538,N_11528,N_9851);
xnor U13539 (N_13539,N_11708,N_10297);
and U13540 (N_13540,N_10551,N_10786);
or U13541 (N_13541,N_10097,N_10480);
and U13542 (N_13542,N_11741,N_9012);
nand U13543 (N_13543,N_10713,N_10565);
nor U13544 (N_13544,N_11684,N_10022);
nand U13545 (N_13545,N_11835,N_9196);
xnor U13546 (N_13546,N_10758,N_11451);
or U13547 (N_13547,N_11988,N_9059);
xnor U13548 (N_13548,N_10724,N_9630);
or U13549 (N_13549,N_9213,N_9488);
or U13550 (N_13550,N_10794,N_9941);
nand U13551 (N_13551,N_9321,N_9388);
nand U13552 (N_13552,N_9260,N_11384);
nor U13553 (N_13553,N_9715,N_10494);
or U13554 (N_13554,N_10092,N_10726);
nor U13555 (N_13555,N_10780,N_9954);
nor U13556 (N_13556,N_11984,N_11448);
nor U13557 (N_13557,N_11347,N_9930);
nor U13558 (N_13558,N_11461,N_11886);
nand U13559 (N_13559,N_9527,N_10281);
or U13560 (N_13560,N_10894,N_9993);
and U13561 (N_13561,N_9032,N_9671);
and U13562 (N_13562,N_11306,N_10579);
nor U13563 (N_13563,N_11739,N_10855);
or U13564 (N_13564,N_11000,N_10913);
xnor U13565 (N_13565,N_10173,N_9731);
or U13566 (N_13566,N_9671,N_10523);
and U13567 (N_13567,N_9328,N_10334);
nor U13568 (N_13568,N_9830,N_9572);
nor U13569 (N_13569,N_9411,N_10421);
or U13570 (N_13570,N_11446,N_11337);
and U13571 (N_13571,N_11696,N_9431);
nor U13572 (N_13572,N_11697,N_11696);
xnor U13573 (N_13573,N_10886,N_9744);
nor U13574 (N_13574,N_10938,N_10024);
nand U13575 (N_13575,N_10937,N_9112);
nand U13576 (N_13576,N_11342,N_11656);
nand U13577 (N_13577,N_9386,N_11468);
and U13578 (N_13578,N_10878,N_9251);
nor U13579 (N_13579,N_9037,N_10429);
and U13580 (N_13580,N_9497,N_11897);
or U13581 (N_13581,N_11450,N_10400);
or U13582 (N_13582,N_10359,N_11370);
nand U13583 (N_13583,N_9551,N_9065);
nand U13584 (N_13584,N_10602,N_10300);
or U13585 (N_13585,N_11348,N_11576);
or U13586 (N_13586,N_11103,N_11976);
and U13587 (N_13587,N_11581,N_10136);
and U13588 (N_13588,N_11639,N_10031);
xnor U13589 (N_13589,N_11615,N_10044);
nand U13590 (N_13590,N_9936,N_10863);
nor U13591 (N_13591,N_10560,N_9000);
and U13592 (N_13592,N_9040,N_11940);
xnor U13593 (N_13593,N_10282,N_9083);
and U13594 (N_13594,N_9177,N_11223);
nand U13595 (N_13595,N_11034,N_11711);
and U13596 (N_13596,N_11848,N_9012);
and U13597 (N_13597,N_9152,N_10306);
or U13598 (N_13598,N_11891,N_11755);
nand U13599 (N_13599,N_10951,N_10427);
or U13600 (N_13600,N_11198,N_10164);
nand U13601 (N_13601,N_10530,N_11510);
nor U13602 (N_13602,N_11295,N_11907);
and U13603 (N_13603,N_10327,N_11935);
and U13604 (N_13604,N_10553,N_10772);
and U13605 (N_13605,N_11697,N_9663);
and U13606 (N_13606,N_10306,N_11380);
and U13607 (N_13607,N_11224,N_9591);
or U13608 (N_13608,N_9646,N_10169);
and U13609 (N_13609,N_9564,N_9632);
or U13610 (N_13610,N_9393,N_9240);
or U13611 (N_13611,N_11559,N_11034);
nand U13612 (N_13612,N_9345,N_9122);
nor U13613 (N_13613,N_9667,N_11344);
and U13614 (N_13614,N_9516,N_10390);
and U13615 (N_13615,N_9039,N_11306);
or U13616 (N_13616,N_11642,N_10951);
nand U13617 (N_13617,N_9250,N_11605);
nor U13618 (N_13618,N_10731,N_9397);
nand U13619 (N_13619,N_11543,N_10087);
or U13620 (N_13620,N_11456,N_11847);
nor U13621 (N_13621,N_9756,N_9321);
nor U13622 (N_13622,N_9665,N_10431);
nor U13623 (N_13623,N_11260,N_10006);
and U13624 (N_13624,N_9722,N_9010);
nor U13625 (N_13625,N_11164,N_9508);
or U13626 (N_13626,N_10811,N_11268);
xnor U13627 (N_13627,N_11654,N_11419);
and U13628 (N_13628,N_11837,N_11574);
nand U13629 (N_13629,N_9066,N_9838);
nand U13630 (N_13630,N_10261,N_9340);
and U13631 (N_13631,N_11931,N_9808);
and U13632 (N_13632,N_9584,N_9738);
nand U13633 (N_13633,N_9183,N_11794);
nor U13634 (N_13634,N_11576,N_10703);
xnor U13635 (N_13635,N_10244,N_10475);
xnor U13636 (N_13636,N_9539,N_9046);
and U13637 (N_13637,N_11541,N_9509);
nand U13638 (N_13638,N_9642,N_10575);
and U13639 (N_13639,N_11139,N_9814);
and U13640 (N_13640,N_10497,N_9641);
nor U13641 (N_13641,N_11337,N_9906);
nor U13642 (N_13642,N_10982,N_9681);
nand U13643 (N_13643,N_9619,N_10100);
xor U13644 (N_13644,N_11306,N_11490);
and U13645 (N_13645,N_11770,N_10606);
or U13646 (N_13646,N_9646,N_9081);
and U13647 (N_13647,N_11739,N_9009);
nand U13648 (N_13648,N_11670,N_9618);
or U13649 (N_13649,N_9554,N_11649);
xor U13650 (N_13650,N_10067,N_11536);
nand U13651 (N_13651,N_9447,N_9987);
and U13652 (N_13652,N_11294,N_10437);
or U13653 (N_13653,N_9891,N_11040);
or U13654 (N_13654,N_9266,N_11985);
nor U13655 (N_13655,N_9672,N_11781);
nand U13656 (N_13656,N_11163,N_11893);
or U13657 (N_13657,N_10254,N_10339);
nand U13658 (N_13658,N_9462,N_11967);
nor U13659 (N_13659,N_9714,N_11398);
and U13660 (N_13660,N_9902,N_10902);
and U13661 (N_13661,N_11055,N_10511);
and U13662 (N_13662,N_9114,N_11872);
nor U13663 (N_13663,N_11147,N_10751);
and U13664 (N_13664,N_10050,N_10038);
xor U13665 (N_13665,N_11985,N_11225);
nor U13666 (N_13666,N_11544,N_9224);
xnor U13667 (N_13667,N_9450,N_11096);
or U13668 (N_13668,N_10647,N_10661);
nor U13669 (N_13669,N_11873,N_11728);
xor U13670 (N_13670,N_11915,N_10439);
nor U13671 (N_13671,N_10641,N_11562);
and U13672 (N_13672,N_9491,N_10971);
nor U13673 (N_13673,N_9353,N_11938);
nor U13674 (N_13674,N_9003,N_10329);
nor U13675 (N_13675,N_11058,N_10533);
or U13676 (N_13676,N_11115,N_9019);
and U13677 (N_13677,N_11598,N_11694);
and U13678 (N_13678,N_9462,N_11747);
and U13679 (N_13679,N_9762,N_11037);
or U13680 (N_13680,N_10722,N_9589);
or U13681 (N_13681,N_10710,N_11283);
and U13682 (N_13682,N_11537,N_9328);
and U13683 (N_13683,N_11565,N_10839);
nand U13684 (N_13684,N_11975,N_9109);
and U13685 (N_13685,N_10457,N_10320);
nor U13686 (N_13686,N_9060,N_10435);
or U13687 (N_13687,N_11038,N_9100);
nand U13688 (N_13688,N_10431,N_9243);
nor U13689 (N_13689,N_9333,N_11547);
or U13690 (N_13690,N_9894,N_9740);
nor U13691 (N_13691,N_9809,N_10394);
and U13692 (N_13692,N_10168,N_11726);
or U13693 (N_13693,N_9999,N_9067);
or U13694 (N_13694,N_11526,N_9387);
or U13695 (N_13695,N_10474,N_9102);
nor U13696 (N_13696,N_9059,N_11672);
or U13697 (N_13697,N_9627,N_9204);
or U13698 (N_13698,N_9558,N_9853);
nor U13699 (N_13699,N_11533,N_11543);
nand U13700 (N_13700,N_9618,N_11435);
xnor U13701 (N_13701,N_11425,N_9142);
and U13702 (N_13702,N_10347,N_9359);
nor U13703 (N_13703,N_9288,N_10962);
or U13704 (N_13704,N_10112,N_9854);
nor U13705 (N_13705,N_11555,N_11786);
and U13706 (N_13706,N_11791,N_11360);
or U13707 (N_13707,N_11812,N_10741);
and U13708 (N_13708,N_11575,N_11506);
and U13709 (N_13709,N_11122,N_10247);
and U13710 (N_13710,N_11610,N_9878);
nor U13711 (N_13711,N_10183,N_11487);
xor U13712 (N_13712,N_10742,N_9961);
and U13713 (N_13713,N_11280,N_9307);
or U13714 (N_13714,N_9661,N_10488);
xnor U13715 (N_13715,N_10421,N_9487);
and U13716 (N_13716,N_9750,N_10754);
or U13717 (N_13717,N_11402,N_10449);
nand U13718 (N_13718,N_9304,N_11927);
nand U13719 (N_13719,N_10827,N_10990);
xnor U13720 (N_13720,N_9871,N_10156);
and U13721 (N_13721,N_9860,N_10660);
and U13722 (N_13722,N_10072,N_11075);
nand U13723 (N_13723,N_11566,N_10716);
xnor U13724 (N_13724,N_11572,N_11046);
xor U13725 (N_13725,N_10901,N_11106);
nand U13726 (N_13726,N_11452,N_11567);
nor U13727 (N_13727,N_11453,N_9382);
or U13728 (N_13728,N_11987,N_11758);
or U13729 (N_13729,N_11727,N_9852);
nor U13730 (N_13730,N_11532,N_11107);
nand U13731 (N_13731,N_9104,N_10607);
and U13732 (N_13732,N_9894,N_10616);
nor U13733 (N_13733,N_11083,N_10025);
or U13734 (N_13734,N_10329,N_11627);
xnor U13735 (N_13735,N_9083,N_9799);
and U13736 (N_13736,N_9169,N_9925);
and U13737 (N_13737,N_9024,N_11842);
nand U13738 (N_13738,N_10800,N_11693);
nor U13739 (N_13739,N_11845,N_10492);
or U13740 (N_13740,N_9944,N_11391);
or U13741 (N_13741,N_11893,N_9173);
or U13742 (N_13742,N_11053,N_11941);
nor U13743 (N_13743,N_10733,N_10496);
or U13744 (N_13744,N_11746,N_10253);
nand U13745 (N_13745,N_9970,N_9214);
and U13746 (N_13746,N_9252,N_10852);
and U13747 (N_13747,N_9128,N_9965);
xnor U13748 (N_13748,N_9124,N_11676);
or U13749 (N_13749,N_10892,N_9425);
nor U13750 (N_13750,N_9780,N_9789);
or U13751 (N_13751,N_10476,N_11756);
nand U13752 (N_13752,N_11539,N_10951);
and U13753 (N_13753,N_9470,N_11951);
nor U13754 (N_13754,N_9308,N_9633);
nand U13755 (N_13755,N_10631,N_9536);
and U13756 (N_13756,N_9537,N_10340);
nor U13757 (N_13757,N_9465,N_10710);
or U13758 (N_13758,N_10976,N_11280);
nand U13759 (N_13759,N_11748,N_11820);
and U13760 (N_13760,N_9557,N_11704);
xnor U13761 (N_13761,N_9463,N_10770);
and U13762 (N_13762,N_9237,N_9692);
nand U13763 (N_13763,N_9703,N_9281);
nand U13764 (N_13764,N_11083,N_9865);
or U13765 (N_13765,N_9365,N_11372);
nand U13766 (N_13766,N_11521,N_11616);
or U13767 (N_13767,N_11420,N_11279);
nor U13768 (N_13768,N_10711,N_11145);
or U13769 (N_13769,N_10195,N_9527);
or U13770 (N_13770,N_10435,N_9124);
nor U13771 (N_13771,N_10674,N_11513);
nand U13772 (N_13772,N_10066,N_11315);
and U13773 (N_13773,N_9296,N_9800);
or U13774 (N_13774,N_10003,N_10301);
nand U13775 (N_13775,N_10004,N_9570);
nor U13776 (N_13776,N_10030,N_11763);
or U13777 (N_13777,N_11672,N_9615);
and U13778 (N_13778,N_9064,N_10384);
and U13779 (N_13779,N_9219,N_10690);
and U13780 (N_13780,N_11437,N_11669);
nand U13781 (N_13781,N_10206,N_10521);
nand U13782 (N_13782,N_10017,N_10492);
xnor U13783 (N_13783,N_9196,N_10011);
and U13784 (N_13784,N_11158,N_11853);
and U13785 (N_13785,N_10638,N_9723);
and U13786 (N_13786,N_11617,N_10009);
nand U13787 (N_13787,N_9313,N_10859);
and U13788 (N_13788,N_10865,N_9473);
or U13789 (N_13789,N_9806,N_9143);
and U13790 (N_13790,N_11954,N_11994);
xor U13791 (N_13791,N_11321,N_9615);
xnor U13792 (N_13792,N_11890,N_10305);
and U13793 (N_13793,N_11466,N_10192);
nor U13794 (N_13794,N_9357,N_10484);
or U13795 (N_13795,N_11670,N_10012);
and U13796 (N_13796,N_10080,N_10193);
nand U13797 (N_13797,N_10026,N_10371);
nor U13798 (N_13798,N_11141,N_10855);
nor U13799 (N_13799,N_11924,N_9923);
and U13800 (N_13800,N_10013,N_11583);
and U13801 (N_13801,N_10386,N_10065);
xor U13802 (N_13802,N_11949,N_10497);
or U13803 (N_13803,N_10492,N_9622);
or U13804 (N_13804,N_11941,N_10983);
nor U13805 (N_13805,N_10989,N_10021);
or U13806 (N_13806,N_9142,N_10961);
nand U13807 (N_13807,N_11268,N_9142);
and U13808 (N_13808,N_11622,N_11648);
and U13809 (N_13809,N_11371,N_9519);
nand U13810 (N_13810,N_11762,N_10580);
nor U13811 (N_13811,N_10172,N_9425);
xor U13812 (N_13812,N_11668,N_9976);
nor U13813 (N_13813,N_9198,N_9310);
or U13814 (N_13814,N_9490,N_9362);
nand U13815 (N_13815,N_9539,N_10329);
xor U13816 (N_13816,N_9106,N_9584);
nand U13817 (N_13817,N_11434,N_10892);
and U13818 (N_13818,N_10464,N_11640);
nor U13819 (N_13819,N_11501,N_9844);
nor U13820 (N_13820,N_11417,N_9799);
nand U13821 (N_13821,N_9577,N_11184);
or U13822 (N_13822,N_11597,N_9512);
nand U13823 (N_13823,N_11325,N_10244);
xor U13824 (N_13824,N_11438,N_10043);
nor U13825 (N_13825,N_10830,N_11604);
and U13826 (N_13826,N_10786,N_10524);
or U13827 (N_13827,N_10623,N_10491);
nand U13828 (N_13828,N_11211,N_9859);
and U13829 (N_13829,N_11696,N_9171);
and U13830 (N_13830,N_11476,N_10661);
or U13831 (N_13831,N_9949,N_11644);
nor U13832 (N_13832,N_11351,N_11092);
and U13833 (N_13833,N_9067,N_10410);
or U13834 (N_13834,N_11726,N_9207);
or U13835 (N_13835,N_11920,N_11797);
and U13836 (N_13836,N_11016,N_11810);
nand U13837 (N_13837,N_11449,N_9826);
or U13838 (N_13838,N_9086,N_10861);
or U13839 (N_13839,N_10947,N_10391);
or U13840 (N_13840,N_10326,N_10062);
or U13841 (N_13841,N_10703,N_11381);
nor U13842 (N_13842,N_11127,N_9073);
and U13843 (N_13843,N_11860,N_9274);
or U13844 (N_13844,N_9442,N_10146);
or U13845 (N_13845,N_11905,N_9136);
nand U13846 (N_13846,N_9674,N_11092);
and U13847 (N_13847,N_10544,N_10296);
xor U13848 (N_13848,N_11648,N_10328);
nand U13849 (N_13849,N_11161,N_11360);
or U13850 (N_13850,N_11161,N_10275);
nor U13851 (N_13851,N_11246,N_11175);
or U13852 (N_13852,N_9129,N_9403);
or U13853 (N_13853,N_11040,N_10275);
and U13854 (N_13854,N_9873,N_10483);
nor U13855 (N_13855,N_10222,N_9368);
or U13856 (N_13856,N_9892,N_10652);
nand U13857 (N_13857,N_9642,N_11798);
and U13858 (N_13858,N_10707,N_9518);
xor U13859 (N_13859,N_9647,N_10694);
nand U13860 (N_13860,N_9424,N_10990);
nor U13861 (N_13861,N_11732,N_11467);
or U13862 (N_13862,N_9541,N_11956);
or U13863 (N_13863,N_9626,N_10196);
nor U13864 (N_13864,N_9364,N_11210);
nor U13865 (N_13865,N_11571,N_9628);
nand U13866 (N_13866,N_10435,N_10741);
or U13867 (N_13867,N_10485,N_11204);
nor U13868 (N_13868,N_10505,N_11408);
or U13869 (N_13869,N_11525,N_10889);
nand U13870 (N_13870,N_10313,N_10847);
or U13871 (N_13871,N_10572,N_9208);
or U13872 (N_13872,N_11686,N_11614);
nand U13873 (N_13873,N_11253,N_9378);
nor U13874 (N_13874,N_11051,N_9836);
or U13875 (N_13875,N_9657,N_10660);
and U13876 (N_13876,N_9245,N_11798);
xnor U13877 (N_13877,N_10596,N_9113);
and U13878 (N_13878,N_11083,N_11542);
or U13879 (N_13879,N_11037,N_9834);
and U13880 (N_13880,N_9274,N_9048);
nor U13881 (N_13881,N_11040,N_11766);
xnor U13882 (N_13882,N_10750,N_10574);
nand U13883 (N_13883,N_11737,N_11979);
and U13884 (N_13884,N_11872,N_11245);
nand U13885 (N_13885,N_11727,N_9370);
nand U13886 (N_13886,N_9175,N_10605);
or U13887 (N_13887,N_10692,N_10394);
and U13888 (N_13888,N_10333,N_11881);
or U13889 (N_13889,N_11329,N_11488);
or U13890 (N_13890,N_9579,N_9104);
nand U13891 (N_13891,N_10923,N_10409);
nand U13892 (N_13892,N_10636,N_9074);
and U13893 (N_13893,N_10222,N_11208);
nor U13894 (N_13894,N_11401,N_10309);
or U13895 (N_13895,N_10341,N_10361);
xor U13896 (N_13896,N_11682,N_11097);
nand U13897 (N_13897,N_11352,N_9762);
xnor U13898 (N_13898,N_9256,N_9228);
nor U13899 (N_13899,N_11448,N_9102);
and U13900 (N_13900,N_11170,N_9356);
and U13901 (N_13901,N_11844,N_11732);
or U13902 (N_13902,N_11946,N_9917);
and U13903 (N_13903,N_10541,N_11327);
or U13904 (N_13904,N_9388,N_9627);
and U13905 (N_13905,N_11582,N_9478);
nor U13906 (N_13906,N_11427,N_10270);
nand U13907 (N_13907,N_9879,N_10610);
or U13908 (N_13908,N_9024,N_9769);
and U13909 (N_13909,N_10315,N_9934);
and U13910 (N_13910,N_11936,N_10105);
and U13911 (N_13911,N_11731,N_10520);
or U13912 (N_13912,N_9229,N_9061);
nor U13913 (N_13913,N_10140,N_11386);
nor U13914 (N_13914,N_10596,N_9053);
nor U13915 (N_13915,N_10990,N_9847);
nand U13916 (N_13916,N_9635,N_11296);
or U13917 (N_13917,N_11592,N_11288);
or U13918 (N_13918,N_10680,N_10321);
or U13919 (N_13919,N_9120,N_10160);
or U13920 (N_13920,N_10644,N_11633);
or U13921 (N_13921,N_10572,N_9298);
or U13922 (N_13922,N_9631,N_11471);
nor U13923 (N_13923,N_11037,N_10949);
nand U13924 (N_13924,N_11780,N_10701);
nor U13925 (N_13925,N_11300,N_11294);
nand U13926 (N_13926,N_10213,N_11556);
nor U13927 (N_13927,N_10053,N_9641);
and U13928 (N_13928,N_11699,N_10593);
and U13929 (N_13929,N_9868,N_9177);
nor U13930 (N_13930,N_10107,N_11753);
nor U13931 (N_13931,N_9812,N_10055);
nand U13932 (N_13932,N_9646,N_9507);
and U13933 (N_13933,N_11696,N_11885);
nor U13934 (N_13934,N_9338,N_11965);
and U13935 (N_13935,N_11491,N_11364);
nor U13936 (N_13936,N_10416,N_9844);
or U13937 (N_13937,N_10247,N_9090);
nand U13938 (N_13938,N_11745,N_9133);
xnor U13939 (N_13939,N_9146,N_10502);
and U13940 (N_13940,N_11792,N_11651);
and U13941 (N_13941,N_10817,N_9857);
nand U13942 (N_13942,N_9469,N_10798);
or U13943 (N_13943,N_11277,N_11621);
or U13944 (N_13944,N_10584,N_11049);
or U13945 (N_13945,N_10462,N_9644);
or U13946 (N_13946,N_9913,N_10705);
or U13947 (N_13947,N_9908,N_9978);
and U13948 (N_13948,N_10428,N_11784);
nand U13949 (N_13949,N_10155,N_10226);
and U13950 (N_13950,N_9327,N_9481);
or U13951 (N_13951,N_9119,N_10654);
or U13952 (N_13952,N_9768,N_10570);
or U13953 (N_13953,N_9713,N_11642);
nor U13954 (N_13954,N_11574,N_10386);
nand U13955 (N_13955,N_9413,N_10943);
or U13956 (N_13956,N_11422,N_9652);
nor U13957 (N_13957,N_10926,N_11030);
or U13958 (N_13958,N_9144,N_10864);
or U13959 (N_13959,N_10491,N_9883);
or U13960 (N_13960,N_10008,N_9451);
nand U13961 (N_13961,N_10047,N_9481);
and U13962 (N_13962,N_11793,N_11780);
or U13963 (N_13963,N_9950,N_11455);
or U13964 (N_13964,N_11236,N_11202);
and U13965 (N_13965,N_9729,N_9409);
or U13966 (N_13966,N_10573,N_11031);
nand U13967 (N_13967,N_10261,N_11223);
or U13968 (N_13968,N_9830,N_9918);
or U13969 (N_13969,N_10137,N_10672);
nand U13970 (N_13970,N_10307,N_10807);
nand U13971 (N_13971,N_10741,N_9338);
or U13972 (N_13972,N_11549,N_11168);
nor U13973 (N_13973,N_11442,N_9926);
and U13974 (N_13974,N_9474,N_9618);
and U13975 (N_13975,N_11513,N_9804);
and U13976 (N_13976,N_11715,N_10175);
or U13977 (N_13977,N_9160,N_9957);
or U13978 (N_13978,N_10682,N_9472);
nor U13979 (N_13979,N_11190,N_9519);
nand U13980 (N_13980,N_10376,N_11011);
nor U13981 (N_13981,N_10686,N_10666);
or U13982 (N_13982,N_10201,N_9205);
or U13983 (N_13983,N_9656,N_9925);
nor U13984 (N_13984,N_11693,N_10157);
nor U13985 (N_13985,N_11552,N_10225);
and U13986 (N_13986,N_11316,N_11776);
nand U13987 (N_13987,N_10474,N_11027);
or U13988 (N_13988,N_10911,N_10239);
and U13989 (N_13989,N_9406,N_9859);
nand U13990 (N_13990,N_9021,N_11687);
xor U13991 (N_13991,N_11318,N_10399);
or U13992 (N_13992,N_10554,N_11284);
and U13993 (N_13993,N_9608,N_11152);
or U13994 (N_13994,N_9619,N_11224);
nand U13995 (N_13995,N_9583,N_9058);
or U13996 (N_13996,N_9776,N_9542);
nand U13997 (N_13997,N_10660,N_10591);
and U13998 (N_13998,N_9020,N_9657);
nand U13999 (N_13999,N_9135,N_9820);
or U14000 (N_14000,N_10252,N_10355);
nand U14001 (N_14001,N_9533,N_10209);
nor U14002 (N_14002,N_9109,N_10545);
nor U14003 (N_14003,N_10260,N_11398);
nor U14004 (N_14004,N_11458,N_11463);
or U14005 (N_14005,N_11334,N_11727);
or U14006 (N_14006,N_9814,N_11380);
nand U14007 (N_14007,N_11144,N_10632);
or U14008 (N_14008,N_10565,N_11557);
nand U14009 (N_14009,N_10513,N_11941);
and U14010 (N_14010,N_11116,N_11291);
nor U14011 (N_14011,N_11648,N_10029);
and U14012 (N_14012,N_10002,N_11355);
or U14013 (N_14013,N_9658,N_10664);
xnor U14014 (N_14014,N_9257,N_10099);
and U14015 (N_14015,N_10826,N_10716);
nand U14016 (N_14016,N_9584,N_9776);
nor U14017 (N_14017,N_9322,N_10514);
nor U14018 (N_14018,N_11984,N_9743);
or U14019 (N_14019,N_9360,N_10428);
nand U14020 (N_14020,N_10749,N_11479);
nor U14021 (N_14021,N_11822,N_11526);
or U14022 (N_14022,N_11304,N_10028);
or U14023 (N_14023,N_9650,N_9472);
or U14024 (N_14024,N_11498,N_10078);
nand U14025 (N_14025,N_9837,N_10401);
and U14026 (N_14026,N_9269,N_11628);
and U14027 (N_14027,N_10671,N_11597);
xor U14028 (N_14028,N_11026,N_11146);
nor U14029 (N_14029,N_10404,N_9985);
and U14030 (N_14030,N_9135,N_10235);
or U14031 (N_14031,N_11680,N_10258);
nor U14032 (N_14032,N_10086,N_10343);
xor U14033 (N_14033,N_9795,N_10213);
nor U14034 (N_14034,N_10717,N_11570);
nor U14035 (N_14035,N_11678,N_11344);
and U14036 (N_14036,N_9152,N_9161);
and U14037 (N_14037,N_10727,N_11553);
and U14038 (N_14038,N_9616,N_9149);
and U14039 (N_14039,N_10000,N_10218);
xnor U14040 (N_14040,N_9544,N_11135);
nand U14041 (N_14041,N_9033,N_9914);
and U14042 (N_14042,N_9518,N_9203);
nor U14043 (N_14043,N_9950,N_9721);
and U14044 (N_14044,N_11321,N_9495);
nand U14045 (N_14045,N_10542,N_9856);
or U14046 (N_14046,N_9461,N_10749);
xor U14047 (N_14047,N_9949,N_9853);
or U14048 (N_14048,N_9455,N_11731);
xor U14049 (N_14049,N_10604,N_11975);
nand U14050 (N_14050,N_9210,N_11963);
nor U14051 (N_14051,N_10360,N_10777);
nor U14052 (N_14052,N_10491,N_11986);
or U14053 (N_14053,N_11948,N_9794);
xnor U14054 (N_14054,N_9567,N_11334);
and U14055 (N_14055,N_10692,N_11446);
nor U14056 (N_14056,N_11799,N_9716);
nand U14057 (N_14057,N_11443,N_11013);
nand U14058 (N_14058,N_9661,N_9695);
or U14059 (N_14059,N_11620,N_10794);
nor U14060 (N_14060,N_9372,N_10800);
and U14061 (N_14061,N_10062,N_9932);
and U14062 (N_14062,N_9526,N_11439);
or U14063 (N_14063,N_10342,N_11207);
nor U14064 (N_14064,N_9128,N_10084);
and U14065 (N_14065,N_11150,N_9506);
nor U14066 (N_14066,N_11800,N_9590);
nor U14067 (N_14067,N_10500,N_9645);
nand U14068 (N_14068,N_9194,N_10700);
nor U14069 (N_14069,N_11440,N_10190);
and U14070 (N_14070,N_9784,N_10788);
and U14071 (N_14071,N_10549,N_9348);
nand U14072 (N_14072,N_11402,N_10580);
nand U14073 (N_14073,N_9851,N_9409);
nand U14074 (N_14074,N_9723,N_10091);
nand U14075 (N_14075,N_9459,N_11708);
nor U14076 (N_14076,N_9203,N_11798);
or U14077 (N_14077,N_9200,N_11703);
nand U14078 (N_14078,N_9744,N_9915);
and U14079 (N_14079,N_10629,N_11766);
and U14080 (N_14080,N_9090,N_11313);
or U14081 (N_14081,N_11238,N_11586);
nand U14082 (N_14082,N_11398,N_11384);
nand U14083 (N_14083,N_11581,N_9952);
xnor U14084 (N_14084,N_10086,N_10060);
nand U14085 (N_14085,N_11977,N_10447);
or U14086 (N_14086,N_10224,N_9275);
nand U14087 (N_14087,N_10130,N_11774);
nor U14088 (N_14088,N_10473,N_10069);
or U14089 (N_14089,N_10359,N_9408);
and U14090 (N_14090,N_11797,N_11155);
and U14091 (N_14091,N_11175,N_9457);
or U14092 (N_14092,N_9750,N_10716);
and U14093 (N_14093,N_10988,N_10931);
nand U14094 (N_14094,N_10395,N_9954);
nand U14095 (N_14095,N_10983,N_11976);
nand U14096 (N_14096,N_11888,N_10523);
or U14097 (N_14097,N_11882,N_10648);
nand U14098 (N_14098,N_11015,N_11210);
and U14099 (N_14099,N_9104,N_11604);
and U14100 (N_14100,N_10654,N_10703);
or U14101 (N_14101,N_9394,N_9199);
nand U14102 (N_14102,N_9315,N_11130);
and U14103 (N_14103,N_10188,N_9007);
nor U14104 (N_14104,N_11798,N_10471);
and U14105 (N_14105,N_10219,N_10358);
and U14106 (N_14106,N_11836,N_11130);
nand U14107 (N_14107,N_11629,N_9692);
nor U14108 (N_14108,N_11611,N_10529);
and U14109 (N_14109,N_11761,N_9640);
xnor U14110 (N_14110,N_9756,N_11249);
and U14111 (N_14111,N_9833,N_11800);
nand U14112 (N_14112,N_9840,N_10524);
nand U14113 (N_14113,N_11950,N_9152);
and U14114 (N_14114,N_11303,N_10230);
nand U14115 (N_14115,N_10807,N_10490);
xnor U14116 (N_14116,N_9994,N_10602);
and U14117 (N_14117,N_10729,N_11138);
and U14118 (N_14118,N_11224,N_10117);
nand U14119 (N_14119,N_11884,N_9703);
and U14120 (N_14120,N_9135,N_9769);
nand U14121 (N_14121,N_11608,N_10872);
or U14122 (N_14122,N_9390,N_9896);
nor U14123 (N_14123,N_11338,N_11382);
nand U14124 (N_14124,N_11500,N_10333);
nor U14125 (N_14125,N_11813,N_10752);
nand U14126 (N_14126,N_11439,N_11427);
and U14127 (N_14127,N_11481,N_11756);
and U14128 (N_14128,N_10377,N_11287);
nor U14129 (N_14129,N_9788,N_10326);
nand U14130 (N_14130,N_11581,N_11363);
and U14131 (N_14131,N_11848,N_10620);
nand U14132 (N_14132,N_9092,N_9385);
nand U14133 (N_14133,N_11899,N_9682);
and U14134 (N_14134,N_11971,N_10352);
and U14135 (N_14135,N_9551,N_9525);
and U14136 (N_14136,N_9960,N_11283);
nand U14137 (N_14137,N_9305,N_11556);
and U14138 (N_14138,N_9443,N_9747);
nand U14139 (N_14139,N_11907,N_10252);
and U14140 (N_14140,N_10331,N_11739);
nor U14141 (N_14141,N_10180,N_10243);
nor U14142 (N_14142,N_10537,N_10467);
or U14143 (N_14143,N_11326,N_11817);
and U14144 (N_14144,N_9777,N_10242);
and U14145 (N_14145,N_9258,N_11732);
nand U14146 (N_14146,N_9710,N_11712);
or U14147 (N_14147,N_11915,N_11592);
or U14148 (N_14148,N_10002,N_10142);
xnor U14149 (N_14149,N_10534,N_10252);
nor U14150 (N_14150,N_10523,N_9514);
nand U14151 (N_14151,N_11400,N_9858);
or U14152 (N_14152,N_11242,N_10604);
and U14153 (N_14153,N_9319,N_9354);
xnor U14154 (N_14154,N_10776,N_10767);
nor U14155 (N_14155,N_11731,N_10441);
nand U14156 (N_14156,N_10356,N_11367);
nor U14157 (N_14157,N_9997,N_9781);
and U14158 (N_14158,N_9421,N_9908);
nand U14159 (N_14159,N_10739,N_11540);
or U14160 (N_14160,N_9876,N_11732);
or U14161 (N_14161,N_10217,N_10618);
nand U14162 (N_14162,N_10732,N_9545);
xor U14163 (N_14163,N_11356,N_11726);
and U14164 (N_14164,N_11484,N_11040);
or U14165 (N_14165,N_11833,N_9889);
nor U14166 (N_14166,N_9794,N_10712);
or U14167 (N_14167,N_10954,N_10402);
or U14168 (N_14168,N_9392,N_11808);
nand U14169 (N_14169,N_10044,N_10226);
xnor U14170 (N_14170,N_9024,N_10028);
nand U14171 (N_14171,N_9237,N_9127);
nand U14172 (N_14172,N_10189,N_9089);
nor U14173 (N_14173,N_9941,N_9674);
xor U14174 (N_14174,N_10857,N_11636);
nand U14175 (N_14175,N_10092,N_9878);
and U14176 (N_14176,N_11933,N_10780);
or U14177 (N_14177,N_10544,N_9160);
xnor U14178 (N_14178,N_10491,N_11098);
nand U14179 (N_14179,N_11212,N_9685);
and U14180 (N_14180,N_9914,N_11198);
or U14181 (N_14181,N_9070,N_9575);
or U14182 (N_14182,N_11258,N_10167);
or U14183 (N_14183,N_10379,N_11142);
nor U14184 (N_14184,N_9994,N_10917);
xor U14185 (N_14185,N_10037,N_10935);
nand U14186 (N_14186,N_11320,N_10763);
or U14187 (N_14187,N_11852,N_11517);
and U14188 (N_14188,N_9802,N_11497);
or U14189 (N_14189,N_9017,N_9706);
xnor U14190 (N_14190,N_9248,N_9476);
nand U14191 (N_14191,N_10425,N_9477);
or U14192 (N_14192,N_9592,N_10844);
nand U14193 (N_14193,N_9316,N_11984);
nand U14194 (N_14194,N_10680,N_10655);
nor U14195 (N_14195,N_11132,N_11767);
nor U14196 (N_14196,N_11114,N_10045);
and U14197 (N_14197,N_10238,N_9422);
nor U14198 (N_14198,N_11234,N_9917);
and U14199 (N_14199,N_9097,N_9663);
or U14200 (N_14200,N_11769,N_10399);
nor U14201 (N_14201,N_11496,N_9384);
nand U14202 (N_14202,N_9048,N_11318);
or U14203 (N_14203,N_9962,N_10412);
nor U14204 (N_14204,N_10579,N_10443);
and U14205 (N_14205,N_9081,N_9139);
or U14206 (N_14206,N_9046,N_9732);
or U14207 (N_14207,N_11445,N_9807);
nand U14208 (N_14208,N_10680,N_11617);
nand U14209 (N_14209,N_10995,N_11392);
or U14210 (N_14210,N_9442,N_11133);
nand U14211 (N_14211,N_11549,N_9384);
and U14212 (N_14212,N_10638,N_10903);
nand U14213 (N_14213,N_9597,N_9353);
or U14214 (N_14214,N_10877,N_10107);
xnor U14215 (N_14215,N_11334,N_10779);
xnor U14216 (N_14216,N_10971,N_9100);
nand U14217 (N_14217,N_11880,N_11110);
nand U14218 (N_14218,N_9735,N_11116);
nand U14219 (N_14219,N_10249,N_11410);
and U14220 (N_14220,N_9996,N_10039);
and U14221 (N_14221,N_10698,N_11085);
and U14222 (N_14222,N_11014,N_9950);
nor U14223 (N_14223,N_11814,N_9388);
nand U14224 (N_14224,N_10646,N_11051);
nor U14225 (N_14225,N_9526,N_11894);
and U14226 (N_14226,N_10120,N_11153);
nor U14227 (N_14227,N_9234,N_9256);
nor U14228 (N_14228,N_10099,N_10740);
and U14229 (N_14229,N_9477,N_9280);
nor U14230 (N_14230,N_11273,N_11574);
or U14231 (N_14231,N_11764,N_9635);
xor U14232 (N_14232,N_11981,N_10732);
and U14233 (N_14233,N_9200,N_11694);
and U14234 (N_14234,N_11371,N_11207);
nor U14235 (N_14235,N_10779,N_10359);
and U14236 (N_14236,N_11899,N_10781);
and U14237 (N_14237,N_10969,N_11769);
and U14238 (N_14238,N_10260,N_11648);
or U14239 (N_14239,N_9811,N_11196);
and U14240 (N_14240,N_9426,N_10890);
nand U14241 (N_14241,N_10133,N_11914);
xnor U14242 (N_14242,N_9948,N_11279);
or U14243 (N_14243,N_11495,N_11948);
and U14244 (N_14244,N_9550,N_10397);
nand U14245 (N_14245,N_11951,N_11363);
and U14246 (N_14246,N_11506,N_11365);
nor U14247 (N_14247,N_11421,N_11051);
nand U14248 (N_14248,N_9645,N_10761);
nor U14249 (N_14249,N_9581,N_10751);
nand U14250 (N_14250,N_11283,N_10508);
xnor U14251 (N_14251,N_9553,N_9045);
nor U14252 (N_14252,N_11882,N_11646);
or U14253 (N_14253,N_11543,N_11336);
or U14254 (N_14254,N_9010,N_11117);
nor U14255 (N_14255,N_9192,N_9202);
and U14256 (N_14256,N_11023,N_11308);
or U14257 (N_14257,N_9567,N_11536);
xnor U14258 (N_14258,N_11801,N_9543);
nand U14259 (N_14259,N_11424,N_11182);
and U14260 (N_14260,N_11103,N_10547);
or U14261 (N_14261,N_10968,N_11355);
and U14262 (N_14262,N_10030,N_11425);
nand U14263 (N_14263,N_9846,N_11679);
nor U14264 (N_14264,N_11010,N_10350);
nor U14265 (N_14265,N_9566,N_11201);
or U14266 (N_14266,N_11530,N_11644);
nand U14267 (N_14267,N_9637,N_9912);
and U14268 (N_14268,N_11121,N_10282);
nor U14269 (N_14269,N_9211,N_11201);
nor U14270 (N_14270,N_10325,N_11042);
nand U14271 (N_14271,N_9924,N_10359);
or U14272 (N_14272,N_11651,N_9449);
nor U14273 (N_14273,N_11307,N_9912);
nor U14274 (N_14274,N_11189,N_10017);
nand U14275 (N_14275,N_11354,N_11827);
and U14276 (N_14276,N_9329,N_9000);
nand U14277 (N_14277,N_11824,N_10087);
nand U14278 (N_14278,N_11791,N_9599);
nor U14279 (N_14279,N_9931,N_10798);
and U14280 (N_14280,N_11331,N_11897);
nor U14281 (N_14281,N_10914,N_11747);
or U14282 (N_14282,N_10232,N_11938);
nand U14283 (N_14283,N_10236,N_9976);
nand U14284 (N_14284,N_9792,N_9752);
or U14285 (N_14285,N_10443,N_9102);
xor U14286 (N_14286,N_11027,N_10575);
nand U14287 (N_14287,N_10303,N_9311);
and U14288 (N_14288,N_9137,N_10098);
nor U14289 (N_14289,N_10652,N_9645);
or U14290 (N_14290,N_9126,N_10471);
and U14291 (N_14291,N_10086,N_9081);
nor U14292 (N_14292,N_9668,N_10448);
nor U14293 (N_14293,N_10025,N_10245);
nand U14294 (N_14294,N_10895,N_9345);
and U14295 (N_14295,N_9748,N_11340);
nor U14296 (N_14296,N_10361,N_10138);
nand U14297 (N_14297,N_11960,N_11087);
and U14298 (N_14298,N_9323,N_11509);
nand U14299 (N_14299,N_11900,N_10233);
and U14300 (N_14300,N_11335,N_10640);
nor U14301 (N_14301,N_9327,N_11393);
or U14302 (N_14302,N_9518,N_11185);
or U14303 (N_14303,N_9308,N_10217);
and U14304 (N_14304,N_9136,N_11822);
nor U14305 (N_14305,N_9443,N_10386);
nand U14306 (N_14306,N_10559,N_9184);
nand U14307 (N_14307,N_9839,N_10388);
or U14308 (N_14308,N_11475,N_9584);
and U14309 (N_14309,N_11251,N_10227);
xor U14310 (N_14310,N_10888,N_11864);
nand U14311 (N_14311,N_11529,N_11298);
nand U14312 (N_14312,N_9740,N_10849);
or U14313 (N_14313,N_10506,N_9080);
xnor U14314 (N_14314,N_9089,N_11692);
nor U14315 (N_14315,N_9140,N_11397);
and U14316 (N_14316,N_9639,N_9609);
and U14317 (N_14317,N_10369,N_11484);
xor U14318 (N_14318,N_11080,N_11975);
nand U14319 (N_14319,N_11122,N_11951);
and U14320 (N_14320,N_10347,N_10943);
nand U14321 (N_14321,N_10911,N_11951);
nand U14322 (N_14322,N_10213,N_11042);
nand U14323 (N_14323,N_9173,N_10687);
or U14324 (N_14324,N_11210,N_11026);
nor U14325 (N_14325,N_9572,N_9623);
or U14326 (N_14326,N_11866,N_11061);
or U14327 (N_14327,N_11939,N_11271);
xnor U14328 (N_14328,N_10318,N_11474);
and U14329 (N_14329,N_11202,N_10045);
xnor U14330 (N_14330,N_10489,N_11987);
or U14331 (N_14331,N_10274,N_10739);
nand U14332 (N_14332,N_9657,N_10828);
and U14333 (N_14333,N_9651,N_9880);
nor U14334 (N_14334,N_9915,N_9931);
nand U14335 (N_14335,N_10027,N_9312);
or U14336 (N_14336,N_10188,N_11323);
nor U14337 (N_14337,N_11611,N_11783);
nor U14338 (N_14338,N_11137,N_10600);
or U14339 (N_14339,N_10693,N_11727);
xnor U14340 (N_14340,N_11577,N_9234);
nand U14341 (N_14341,N_9739,N_11997);
or U14342 (N_14342,N_9072,N_10005);
nor U14343 (N_14343,N_10702,N_10165);
or U14344 (N_14344,N_11118,N_11472);
nand U14345 (N_14345,N_10514,N_10475);
or U14346 (N_14346,N_11751,N_9426);
and U14347 (N_14347,N_9268,N_11299);
nand U14348 (N_14348,N_11995,N_9540);
or U14349 (N_14349,N_11741,N_9517);
nor U14350 (N_14350,N_9597,N_11566);
xnor U14351 (N_14351,N_11925,N_9945);
xor U14352 (N_14352,N_11600,N_9691);
and U14353 (N_14353,N_11877,N_9898);
and U14354 (N_14354,N_11750,N_10819);
or U14355 (N_14355,N_9457,N_9805);
and U14356 (N_14356,N_10841,N_11685);
or U14357 (N_14357,N_9367,N_11627);
and U14358 (N_14358,N_10646,N_9987);
or U14359 (N_14359,N_10864,N_11204);
or U14360 (N_14360,N_10581,N_10883);
or U14361 (N_14361,N_11431,N_10135);
or U14362 (N_14362,N_10544,N_11143);
or U14363 (N_14363,N_9000,N_11200);
or U14364 (N_14364,N_9322,N_10502);
or U14365 (N_14365,N_11458,N_9333);
or U14366 (N_14366,N_9219,N_10409);
xor U14367 (N_14367,N_9396,N_9626);
or U14368 (N_14368,N_11008,N_9507);
and U14369 (N_14369,N_9049,N_11595);
or U14370 (N_14370,N_10841,N_10353);
nor U14371 (N_14371,N_11509,N_10664);
or U14372 (N_14372,N_11231,N_11781);
nand U14373 (N_14373,N_11314,N_10816);
or U14374 (N_14374,N_9462,N_9060);
xor U14375 (N_14375,N_10200,N_9163);
and U14376 (N_14376,N_9581,N_9782);
or U14377 (N_14377,N_10300,N_10756);
and U14378 (N_14378,N_10606,N_11437);
nor U14379 (N_14379,N_10456,N_9417);
and U14380 (N_14380,N_9037,N_10710);
nand U14381 (N_14381,N_10497,N_9340);
and U14382 (N_14382,N_10547,N_11502);
and U14383 (N_14383,N_9387,N_10062);
nor U14384 (N_14384,N_9099,N_11239);
and U14385 (N_14385,N_9998,N_11049);
xnor U14386 (N_14386,N_9016,N_10486);
or U14387 (N_14387,N_10675,N_9670);
nor U14388 (N_14388,N_10101,N_10629);
or U14389 (N_14389,N_9015,N_11292);
or U14390 (N_14390,N_11362,N_10738);
xor U14391 (N_14391,N_11262,N_10030);
nand U14392 (N_14392,N_10260,N_10852);
and U14393 (N_14393,N_10822,N_9593);
nand U14394 (N_14394,N_10103,N_11142);
and U14395 (N_14395,N_10648,N_10209);
or U14396 (N_14396,N_11244,N_11506);
and U14397 (N_14397,N_9255,N_11170);
and U14398 (N_14398,N_11404,N_10063);
and U14399 (N_14399,N_9453,N_10033);
xnor U14400 (N_14400,N_9094,N_10727);
or U14401 (N_14401,N_9256,N_9998);
or U14402 (N_14402,N_9018,N_11680);
nor U14403 (N_14403,N_11915,N_11724);
or U14404 (N_14404,N_10111,N_11857);
nor U14405 (N_14405,N_9671,N_10427);
or U14406 (N_14406,N_10224,N_9444);
and U14407 (N_14407,N_9637,N_11558);
or U14408 (N_14408,N_9823,N_9858);
and U14409 (N_14409,N_9490,N_10527);
or U14410 (N_14410,N_10890,N_10674);
nand U14411 (N_14411,N_11845,N_11299);
and U14412 (N_14412,N_9658,N_9540);
nor U14413 (N_14413,N_11620,N_11797);
and U14414 (N_14414,N_9450,N_11574);
nor U14415 (N_14415,N_10398,N_9786);
nor U14416 (N_14416,N_9710,N_11676);
xor U14417 (N_14417,N_11355,N_11837);
or U14418 (N_14418,N_10747,N_10685);
or U14419 (N_14419,N_9700,N_11092);
nand U14420 (N_14420,N_9666,N_10961);
xnor U14421 (N_14421,N_11890,N_9211);
and U14422 (N_14422,N_10092,N_9664);
xnor U14423 (N_14423,N_11316,N_10540);
and U14424 (N_14424,N_10600,N_10742);
nand U14425 (N_14425,N_9432,N_11023);
or U14426 (N_14426,N_9438,N_9935);
or U14427 (N_14427,N_10222,N_10590);
xnor U14428 (N_14428,N_10525,N_11666);
nand U14429 (N_14429,N_11484,N_9796);
nand U14430 (N_14430,N_9024,N_10011);
xnor U14431 (N_14431,N_9115,N_11175);
nand U14432 (N_14432,N_9867,N_9940);
nor U14433 (N_14433,N_9900,N_11866);
or U14434 (N_14434,N_10541,N_11807);
and U14435 (N_14435,N_10261,N_9027);
nor U14436 (N_14436,N_9023,N_10028);
nand U14437 (N_14437,N_11167,N_9262);
nand U14438 (N_14438,N_9610,N_10725);
nor U14439 (N_14439,N_9733,N_11452);
nor U14440 (N_14440,N_10716,N_11001);
nand U14441 (N_14441,N_11473,N_9272);
xnor U14442 (N_14442,N_9514,N_11963);
nor U14443 (N_14443,N_11842,N_10829);
nor U14444 (N_14444,N_10915,N_9070);
and U14445 (N_14445,N_11931,N_10686);
nand U14446 (N_14446,N_11424,N_10970);
nand U14447 (N_14447,N_11372,N_9682);
and U14448 (N_14448,N_11954,N_9816);
nand U14449 (N_14449,N_11736,N_10977);
nand U14450 (N_14450,N_9276,N_10331);
and U14451 (N_14451,N_11263,N_10124);
or U14452 (N_14452,N_11503,N_11479);
or U14453 (N_14453,N_11014,N_10782);
nor U14454 (N_14454,N_11273,N_9759);
and U14455 (N_14455,N_9146,N_11446);
or U14456 (N_14456,N_9374,N_11195);
nand U14457 (N_14457,N_9334,N_10433);
nand U14458 (N_14458,N_11310,N_10720);
and U14459 (N_14459,N_10464,N_10421);
nor U14460 (N_14460,N_10400,N_10066);
or U14461 (N_14461,N_10253,N_9307);
and U14462 (N_14462,N_11407,N_11537);
or U14463 (N_14463,N_9011,N_10616);
nand U14464 (N_14464,N_9538,N_11449);
nor U14465 (N_14465,N_10703,N_11986);
and U14466 (N_14466,N_11623,N_11842);
nor U14467 (N_14467,N_11283,N_9851);
or U14468 (N_14468,N_11014,N_10732);
nand U14469 (N_14469,N_9255,N_9829);
nand U14470 (N_14470,N_9652,N_11836);
nor U14471 (N_14471,N_10783,N_11279);
and U14472 (N_14472,N_10378,N_10201);
and U14473 (N_14473,N_11225,N_11432);
nand U14474 (N_14474,N_9900,N_9130);
nor U14475 (N_14475,N_10565,N_9024);
nor U14476 (N_14476,N_11318,N_10521);
and U14477 (N_14477,N_11275,N_9976);
or U14478 (N_14478,N_11320,N_11042);
or U14479 (N_14479,N_9446,N_9208);
nand U14480 (N_14480,N_9268,N_9822);
nand U14481 (N_14481,N_10774,N_11228);
and U14482 (N_14482,N_10160,N_9424);
nand U14483 (N_14483,N_10723,N_10320);
xor U14484 (N_14484,N_9328,N_9983);
nor U14485 (N_14485,N_11631,N_9070);
nor U14486 (N_14486,N_10133,N_11745);
xor U14487 (N_14487,N_9256,N_10854);
or U14488 (N_14488,N_10782,N_9485);
and U14489 (N_14489,N_9132,N_10120);
and U14490 (N_14490,N_9686,N_11398);
nor U14491 (N_14491,N_10486,N_10725);
nor U14492 (N_14492,N_9198,N_10621);
or U14493 (N_14493,N_10386,N_9372);
xor U14494 (N_14494,N_11264,N_10628);
or U14495 (N_14495,N_9455,N_11647);
or U14496 (N_14496,N_9019,N_11912);
and U14497 (N_14497,N_10773,N_10567);
nor U14498 (N_14498,N_10545,N_10640);
or U14499 (N_14499,N_9961,N_11912);
and U14500 (N_14500,N_11964,N_10580);
nor U14501 (N_14501,N_11089,N_10548);
and U14502 (N_14502,N_10856,N_11051);
or U14503 (N_14503,N_10012,N_9800);
nor U14504 (N_14504,N_9683,N_9561);
nor U14505 (N_14505,N_11417,N_11475);
nand U14506 (N_14506,N_11888,N_9308);
nand U14507 (N_14507,N_10664,N_10654);
or U14508 (N_14508,N_9948,N_9914);
and U14509 (N_14509,N_11488,N_10924);
nor U14510 (N_14510,N_9427,N_10231);
nand U14511 (N_14511,N_10154,N_10123);
nand U14512 (N_14512,N_11318,N_9233);
nor U14513 (N_14513,N_11054,N_10741);
nor U14514 (N_14514,N_9290,N_9895);
or U14515 (N_14515,N_9954,N_11036);
or U14516 (N_14516,N_10404,N_11683);
or U14517 (N_14517,N_10887,N_10162);
nor U14518 (N_14518,N_11206,N_9141);
xor U14519 (N_14519,N_9264,N_9773);
or U14520 (N_14520,N_10323,N_11767);
nor U14521 (N_14521,N_11292,N_9167);
nor U14522 (N_14522,N_10765,N_10981);
nor U14523 (N_14523,N_10417,N_11741);
nor U14524 (N_14524,N_11847,N_9534);
nor U14525 (N_14525,N_11582,N_10798);
nor U14526 (N_14526,N_9048,N_10337);
xnor U14527 (N_14527,N_11611,N_9913);
or U14528 (N_14528,N_10525,N_11511);
and U14529 (N_14529,N_10912,N_11329);
nand U14530 (N_14530,N_10121,N_11750);
or U14531 (N_14531,N_10019,N_9832);
and U14532 (N_14532,N_9550,N_9099);
or U14533 (N_14533,N_10050,N_11336);
and U14534 (N_14534,N_11621,N_10170);
and U14535 (N_14535,N_9061,N_10888);
nor U14536 (N_14536,N_11543,N_11660);
or U14537 (N_14537,N_11746,N_9697);
nor U14538 (N_14538,N_11228,N_9778);
or U14539 (N_14539,N_11890,N_11767);
or U14540 (N_14540,N_9367,N_9397);
nor U14541 (N_14541,N_10905,N_10610);
nor U14542 (N_14542,N_9200,N_11282);
nand U14543 (N_14543,N_10246,N_9116);
nand U14544 (N_14544,N_10214,N_9683);
nand U14545 (N_14545,N_11257,N_10946);
or U14546 (N_14546,N_11561,N_11755);
nand U14547 (N_14547,N_10024,N_10376);
and U14548 (N_14548,N_11733,N_9098);
nor U14549 (N_14549,N_9270,N_11231);
and U14550 (N_14550,N_10436,N_11413);
or U14551 (N_14551,N_10092,N_9871);
or U14552 (N_14552,N_9063,N_11169);
or U14553 (N_14553,N_11515,N_11717);
xor U14554 (N_14554,N_11997,N_9397);
and U14555 (N_14555,N_11870,N_10422);
and U14556 (N_14556,N_9075,N_10196);
xor U14557 (N_14557,N_11532,N_11216);
and U14558 (N_14558,N_11717,N_10646);
nor U14559 (N_14559,N_11932,N_10609);
and U14560 (N_14560,N_9804,N_10313);
nor U14561 (N_14561,N_10870,N_9883);
nor U14562 (N_14562,N_10630,N_10294);
xnor U14563 (N_14563,N_9732,N_10408);
nor U14564 (N_14564,N_10648,N_11346);
nor U14565 (N_14565,N_11468,N_11615);
nand U14566 (N_14566,N_10576,N_9538);
nand U14567 (N_14567,N_11260,N_10411);
or U14568 (N_14568,N_9736,N_9697);
nand U14569 (N_14569,N_10955,N_9144);
nand U14570 (N_14570,N_10855,N_10156);
or U14571 (N_14571,N_11601,N_11819);
nand U14572 (N_14572,N_10179,N_11778);
nor U14573 (N_14573,N_10255,N_9880);
and U14574 (N_14574,N_11891,N_11379);
nor U14575 (N_14575,N_10383,N_11997);
nor U14576 (N_14576,N_10891,N_11032);
or U14577 (N_14577,N_10572,N_9283);
and U14578 (N_14578,N_10856,N_9928);
nor U14579 (N_14579,N_11793,N_10091);
nand U14580 (N_14580,N_11762,N_10866);
nand U14581 (N_14581,N_11115,N_10198);
or U14582 (N_14582,N_9038,N_10937);
and U14583 (N_14583,N_9248,N_9570);
nor U14584 (N_14584,N_11472,N_11999);
and U14585 (N_14585,N_11572,N_11253);
or U14586 (N_14586,N_10582,N_11304);
and U14587 (N_14587,N_9611,N_11490);
nand U14588 (N_14588,N_10618,N_11234);
xnor U14589 (N_14589,N_10079,N_9875);
nand U14590 (N_14590,N_10490,N_11546);
nor U14591 (N_14591,N_11732,N_9486);
or U14592 (N_14592,N_11276,N_11097);
or U14593 (N_14593,N_10558,N_9492);
xor U14594 (N_14594,N_11439,N_10018);
nor U14595 (N_14595,N_9535,N_9994);
or U14596 (N_14596,N_9785,N_10089);
xnor U14597 (N_14597,N_11303,N_9144);
xnor U14598 (N_14598,N_10330,N_10743);
nand U14599 (N_14599,N_9509,N_10561);
and U14600 (N_14600,N_10748,N_11498);
or U14601 (N_14601,N_11090,N_9314);
or U14602 (N_14602,N_11536,N_10619);
nand U14603 (N_14603,N_11148,N_10803);
nor U14604 (N_14604,N_11862,N_9319);
and U14605 (N_14605,N_11872,N_10637);
nand U14606 (N_14606,N_11966,N_10845);
nand U14607 (N_14607,N_9245,N_9354);
nand U14608 (N_14608,N_10729,N_9270);
nand U14609 (N_14609,N_10754,N_10636);
or U14610 (N_14610,N_10517,N_9354);
nor U14611 (N_14611,N_11054,N_10636);
or U14612 (N_14612,N_10226,N_9860);
or U14613 (N_14613,N_10067,N_10358);
xor U14614 (N_14614,N_9874,N_9013);
nor U14615 (N_14615,N_9050,N_9042);
and U14616 (N_14616,N_10293,N_9010);
and U14617 (N_14617,N_10699,N_10966);
nand U14618 (N_14618,N_11797,N_11613);
nand U14619 (N_14619,N_11987,N_9411);
and U14620 (N_14620,N_10287,N_9297);
xnor U14621 (N_14621,N_9264,N_11577);
nor U14622 (N_14622,N_11001,N_10462);
nand U14623 (N_14623,N_9931,N_9391);
nand U14624 (N_14624,N_9458,N_11494);
nor U14625 (N_14625,N_9515,N_9672);
nand U14626 (N_14626,N_10194,N_9122);
nand U14627 (N_14627,N_11558,N_11445);
or U14628 (N_14628,N_9425,N_10982);
nor U14629 (N_14629,N_9538,N_10551);
and U14630 (N_14630,N_10699,N_9391);
and U14631 (N_14631,N_10113,N_9064);
and U14632 (N_14632,N_10283,N_11376);
or U14633 (N_14633,N_9436,N_10271);
nor U14634 (N_14634,N_9657,N_9725);
nor U14635 (N_14635,N_11020,N_9184);
and U14636 (N_14636,N_10078,N_10897);
xnor U14637 (N_14637,N_10363,N_11927);
nor U14638 (N_14638,N_11924,N_9999);
nor U14639 (N_14639,N_10960,N_9059);
nor U14640 (N_14640,N_11743,N_10121);
nand U14641 (N_14641,N_11639,N_9290);
nand U14642 (N_14642,N_11870,N_10751);
nor U14643 (N_14643,N_10396,N_11097);
and U14644 (N_14644,N_9196,N_10981);
nor U14645 (N_14645,N_11471,N_9327);
nor U14646 (N_14646,N_11825,N_10541);
nand U14647 (N_14647,N_10812,N_9806);
nand U14648 (N_14648,N_9227,N_10935);
nor U14649 (N_14649,N_11161,N_11670);
xor U14650 (N_14650,N_9522,N_10548);
or U14651 (N_14651,N_9624,N_11068);
or U14652 (N_14652,N_9339,N_9397);
and U14653 (N_14653,N_11888,N_11878);
nand U14654 (N_14654,N_9019,N_11747);
or U14655 (N_14655,N_11744,N_10313);
xor U14656 (N_14656,N_10901,N_9252);
and U14657 (N_14657,N_11641,N_10171);
nand U14658 (N_14658,N_10466,N_9802);
or U14659 (N_14659,N_9531,N_10778);
or U14660 (N_14660,N_9372,N_9834);
nand U14661 (N_14661,N_11687,N_10749);
or U14662 (N_14662,N_9985,N_9387);
and U14663 (N_14663,N_9313,N_10860);
or U14664 (N_14664,N_10139,N_10541);
nand U14665 (N_14665,N_11887,N_10544);
nand U14666 (N_14666,N_11277,N_11094);
nor U14667 (N_14667,N_11328,N_9579);
nor U14668 (N_14668,N_10475,N_11295);
and U14669 (N_14669,N_10033,N_9382);
xnor U14670 (N_14670,N_11051,N_10692);
nor U14671 (N_14671,N_10541,N_11224);
and U14672 (N_14672,N_11983,N_11914);
or U14673 (N_14673,N_9493,N_11588);
nor U14674 (N_14674,N_10224,N_11047);
nand U14675 (N_14675,N_11102,N_9731);
nand U14676 (N_14676,N_9578,N_10069);
xor U14677 (N_14677,N_9317,N_10900);
nor U14678 (N_14678,N_11956,N_9417);
or U14679 (N_14679,N_11746,N_9293);
and U14680 (N_14680,N_11773,N_10328);
or U14681 (N_14681,N_9654,N_10541);
nand U14682 (N_14682,N_10173,N_11805);
and U14683 (N_14683,N_9938,N_11302);
nor U14684 (N_14684,N_11323,N_9769);
nand U14685 (N_14685,N_11286,N_10614);
or U14686 (N_14686,N_11252,N_11630);
nand U14687 (N_14687,N_10890,N_10267);
or U14688 (N_14688,N_11814,N_10012);
xnor U14689 (N_14689,N_10674,N_10669);
nand U14690 (N_14690,N_11953,N_9679);
nor U14691 (N_14691,N_11058,N_11044);
and U14692 (N_14692,N_11687,N_11342);
and U14693 (N_14693,N_11525,N_9032);
or U14694 (N_14694,N_9629,N_11271);
and U14695 (N_14695,N_9284,N_11208);
nand U14696 (N_14696,N_10191,N_11672);
or U14697 (N_14697,N_11292,N_11712);
and U14698 (N_14698,N_10087,N_9950);
nor U14699 (N_14699,N_10726,N_9315);
nand U14700 (N_14700,N_9297,N_11705);
xor U14701 (N_14701,N_10709,N_10583);
or U14702 (N_14702,N_10650,N_9135);
nand U14703 (N_14703,N_10878,N_11187);
nor U14704 (N_14704,N_10549,N_10532);
or U14705 (N_14705,N_10678,N_10123);
or U14706 (N_14706,N_9065,N_11614);
and U14707 (N_14707,N_9330,N_9697);
and U14708 (N_14708,N_10343,N_9851);
and U14709 (N_14709,N_9817,N_11390);
nand U14710 (N_14710,N_10227,N_11348);
nor U14711 (N_14711,N_10003,N_9661);
nor U14712 (N_14712,N_10671,N_9624);
nor U14713 (N_14713,N_10103,N_10952);
and U14714 (N_14714,N_11560,N_11214);
nor U14715 (N_14715,N_9975,N_11798);
nand U14716 (N_14716,N_9017,N_10259);
and U14717 (N_14717,N_9118,N_10937);
and U14718 (N_14718,N_11578,N_10264);
nor U14719 (N_14719,N_11064,N_9815);
nand U14720 (N_14720,N_11996,N_11654);
and U14721 (N_14721,N_10499,N_10914);
nand U14722 (N_14722,N_11163,N_11789);
nand U14723 (N_14723,N_11667,N_10014);
and U14724 (N_14724,N_11643,N_11337);
xnor U14725 (N_14725,N_9719,N_9571);
or U14726 (N_14726,N_11213,N_11211);
or U14727 (N_14727,N_9395,N_10037);
nor U14728 (N_14728,N_11367,N_9799);
nor U14729 (N_14729,N_11815,N_11463);
or U14730 (N_14730,N_11383,N_10710);
nor U14731 (N_14731,N_11847,N_11948);
nor U14732 (N_14732,N_11964,N_10947);
nor U14733 (N_14733,N_11649,N_9015);
and U14734 (N_14734,N_11933,N_10305);
and U14735 (N_14735,N_10804,N_9576);
and U14736 (N_14736,N_11270,N_9122);
nor U14737 (N_14737,N_10224,N_10211);
or U14738 (N_14738,N_10090,N_9874);
nor U14739 (N_14739,N_9225,N_9813);
or U14740 (N_14740,N_9386,N_11489);
nand U14741 (N_14741,N_10619,N_10222);
nor U14742 (N_14742,N_11934,N_11854);
nor U14743 (N_14743,N_9452,N_9376);
nand U14744 (N_14744,N_9484,N_11798);
nor U14745 (N_14745,N_10151,N_11694);
nand U14746 (N_14746,N_9274,N_11764);
and U14747 (N_14747,N_10081,N_10980);
or U14748 (N_14748,N_10319,N_11365);
nand U14749 (N_14749,N_9737,N_11108);
or U14750 (N_14750,N_10136,N_10485);
xnor U14751 (N_14751,N_11444,N_10021);
and U14752 (N_14752,N_10727,N_10788);
xor U14753 (N_14753,N_9755,N_10624);
and U14754 (N_14754,N_10033,N_9982);
nand U14755 (N_14755,N_11956,N_11503);
and U14756 (N_14756,N_9500,N_9777);
or U14757 (N_14757,N_10717,N_10881);
or U14758 (N_14758,N_9058,N_10259);
nor U14759 (N_14759,N_11931,N_9287);
and U14760 (N_14760,N_11243,N_10172);
nand U14761 (N_14761,N_11671,N_10424);
or U14762 (N_14762,N_10731,N_9462);
nand U14763 (N_14763,N_10723,N_11912);
or U14764 (N_14764,N_10412,N_11755);
or U14765 (N_14765,N_9373,N_11695);
or U14766 (N_14766,N_10411,N_11823);
or U14767 (N_14767,N_9823,N_11712);
nor U14768 (N_14768,N_11897,N_11474);
nand U14769 (N_14769,N_9838,N_9904);
or U14770 (N_14770,N_9936,N_10220);
or U14771 (N_14771,N_10132,N_11821);
nand U14772 (N_14772,N_9641,N_9720);
and U14773 (N_14773,N_11841,N_10965);
nand U14774 (N_14774,N_10795,N_11048);
xnor U14775 (N_14775,N_9008,N_10913);
nor U14776 (N_14776,N_10487,N_10282);
and U14777 (N_14777,N_10596,N_9253);
xnor U14778 (N_14778,N_9075,N_11356);
nand U14779 (N_14779,N_9117,N_10473);
xor U14780 (N_14780,N_10856,N_10110);
or U14781 (N_14781,N_10136,N_11035);
or U14782 (N_14782,N_10852,N_9218);
or U14783 (N_14783,N_11128,N_9590);
nand U14784 (N_14784,N_10509,N_11617);
xnor U14785 (N_14785,N_10833,N_9079);
nand U14786 (N_14786,N_11451,N_10104);
nor U14787 (N_14787,N_9769,N_11872);
and U14788 (N_14788,N_9072,N_9103);
or U14789 (N_14789,N_10335,N_10441);
nor U14790 (N_14790,N_10348,N_10240);
and U14791 (N_14791,N_10700,N_10137);
nand U14792 (N_14792,N_10561,N_11732);
and U14793 (N_14793,N_9230,N_11882);
or U14794 (N_14794,N_10969,N_9836);
nor U14795 (N_14795,N_10570,N_9437);
nor U14796 (N_14796,N_11101,N_11671);
nand U14797 (N_14797,N_10813,N_9760);
or U14798 (N_14798,N_11599,N_10598);
nor U14799 (N_14799,N_9643,N_10365);
and U14800 (N_14800,N_9382,N_10933);
xnor U14801 (N_14801,N_9623,N_10418);
or U14802 (N_14802,N_10706,N_11706);
or U14803 (N_14803,N_9292,N_11825);
and U14804 (N_14804,N_10893,N_10897);
xnor U14805 (N_14805,N_10807,N_9003);
nor U14806 (N_14806,N_9724,N_10490);
and U14807 (N_14807,N_11955,N_9878);
nand U14808 (N_14808,N_9449,N_9901);
or U14809 (N_14809,N_10817,N_11485);
and U14810 (N_14810,N_11748,N_10293);
xor U14811 (N_14811,N_9739,N_9979);
nand U14812 (N_14812,N_11729,N_9366);
nand U14813 (N_14813,N_11171,N_9834);
and U14814 (N_14814,N_11823,N_9682);
or U14815 (N_14815,N_11053,N_10482);
nor U14816 (N_14816,N_9093,N_9612);
and U14817 (N_14817,N_11493,N_11792);
and U14818 (N_14818,N_11373,N_9131);
nor U14819 (N_14819,N_9870,N_11448);
nor U14820 (N_14820,N_10685,N_10162);
nor U14821 (N_14821,N_10656,N_9276);
nand U14822 (N_14822,N_9781,N_9139);
nand U14823 (N_14823,N_9836,N_11030);
xnor U14824 (N_14824,N_9386,N_10999);
nand U14825 (N_14825,N_11907,N_9210);
nor U14826 (N_14826,N_10736,N_9107);
xor U14827 (N_14827,N_11620,N_10073);
and U14828 (N_14828,N_10353,N_11124);
xnor U14829 (N_14829,N_11935,N_9851);
nand U14830 (N_14830,N_11996,N_11399);
nor U14831 (N_14831,N_10829,N_9014);
nand U14832 (N_14832,N_11987,N_11019);
and U14833 (N_14833,N_9603,N_10033);
or U14834 (N_14834,N_11138,N_11930);
nor U14835 (N_14835,N_9372,N_11937);
and U14836 (N_14836,N_11854,N_10201);
and U14837 (N_14837,N_9536,N_10282);
nor U14838 (N_14838,N_9628,N_9327);
nand U14839 (N_14839,N_9098,N_11201);
nor U14840 (N_14840,N_9088,N_10976);
and U14841 (N_14841,N_9007,N_10257);
xor U14842 (N_14842,N_9394,N_11479);
nand U14843 (N_14843,N_9777,N_10606);
and U14844 (N_14844,N_10995,N_10790);
nor U14845 (N_14845,N_9807,N_9822);
or U14846 (N_14846,N_10583,N_9260);
nor U14847 (N_14847,N_10613,N_10827);
nor U14848 (N_14848,N_11422,N_11066);
nand U14849 (N_14849,N_11774,N_10755);
and U14850 (N_14850,N_9108,N_9562);
or U14851 (N_14851,N_10899,N_11933);
nand U14852 (N_14852,N_11861,N_11557);
xor U14853 (N_14853,N_11938,N_9842);
nand U14854 (N_14854,N_9824,N_10404);
nand U14855 (N_14855,N_11779,N_10988);
nor U14856 (N_14856,N_10872,N_10153);
nand U14857 (N_14857,N_10068,N_11943);
or U14858 (N_14858,N_9089,N_10141);
nand U14859 (N_14859,N_9491,N_9237);
or U14860 (N_14860,N_11712,N_10809);
or U14861 (N_14861,N_11004,N_9529);
and U14862 (N_14862,N_10045,N_9684);
or U14863 (N_14863,N_9864,N_9154);
nand U14864 (N_14864,N_11388,N_11420);
nand U14865 (N_14865,N_11079,N_11147);
or U14866 (N_14866,N_9953,N_9787);
nand U14867 (N_14867,N_9698,N_9510);
nand U14868 (N_14868,N_10014,N_10500);
xor U14869 (N_14869,N_11218,N_10488);
nor U14870 (N_14870,N_11435,N_11536);
nand U14871 (N_14871,N_11935,N_10068);
and U14872 (N_14872,N_11533,N_9538);
nand U14873 (N_14873,N_9421,N_9220);
nor U14874 (N_14874,N_10671,N_10589);
and U14875 (N_14875,N_10728,N_9733);
or U14876 (N_14876,N_9329,N_11810);
nor U14877 (N_14877,N_10287,N_10126);
and U14878 (N_14878,N_9574,N_9892);
and U14879 (N_14879,N_9802,N_11137);
nor U14880 (N_14880,N_9107,N_11763);
or U14881 (N_14881,N_10603,N_11741);
and U14882 (N_14882,N_10281,N_9562);
and U14883 (N_14883,N_9338,N_9678);
nand U14884 (N_14884,N_11647,N_9539);
or U14885 (N_14885,N_11993,N_11823);
nand U14886 (N_14886,N_10874,N_11870);
nand U14887 (N_14887,N_10687,N_11358);
xnor U14888 (N_14888,N_10547,N_10567);
xor U14889 (N_14889,N_9746,N_10671);
nand U14890 (N_14890,N_9045,N_11129);
or U14891 (N_14891,N_11777,N_11769);
nand U14892 (N_14892,N_9276,N_9132);
or U14893 (N_14893,N_10062,N_9760);
and U14894 (N_14894,N_9023,N_10896);
and U14895 (N_14895,N_9494,N_11414);
nor U14896 (N_14896,N_11330,N_10051);
nor U14897 (N_14897,N_10488,N_10388);
and U14898 (N_14898,N_9825,N_9818);
or U14899 (N_14899,N_11515,N_10770);
and U14900 (N_14900,N_11295,N_9453);
nand U14901 (N_14901,N_11998,N_9648);
nand U14902 (N_14902,N_10515,N_9996);
nand U14903 (N_14903,N_10359,N_11884);
or U14904 (N_14904,N_9092,N_11916);
or U14905 (N_14905,N_11510,N_10845);
nor U14906 (N_14906,N_11888,N_11258);
or U14907 (N_14907,N_11382,N_10212);
xnor U14908 (N_14908,N_11974,N_9888);
or U14909 (N_14909,N_11625,N_10555);
nand U14910 (N_14910,N_10006,N_11595);
nand U14911 (N_14911,N_11919,N_10609);
nand U14912 (N_14912,N_11193,N_11538);
and U14913 (N_14913,N_9907,N_10619);
nand U14914 (N_14914,N_11058,N_10966);
nor U14915 (N_14915,N_11756,N_9167);
nand U14916 (N_14916,N_10315,N_11404);
nand U14917 (N_14917,N_10859,N_10400);
nor U14918 (N_14918,N_11180,N_11223);
or U14919 (N_14919,N_10977,N_10182);
and U14920 (N_14920,N_11236,N_11423);
nand U14921 (N_14921,N_11825,N_9633);
xor U14922 (N_14922,N_10512,N_11221);
nor U14923 (N_14923,N_10761,N_9407);
or U14924 (N_14924,N_10668,N_11539);
nor U14925 (N_14925,N_11639,N_10027);
or U14926 (N_14926,N_11407,N_10067);
or U14927 (N_14927,N_11267,N_10262);
xnor U14928 (N_14928,N_10304,N_11605);
nor U14929 (N_14929,N_9844,N_10477);
nand U14930 (N_14930,N_10033,N_10793);
nor U14931 (N_14931,N_9405,N_10977);
nand U14932 (N_14932,N_11551,N_11543);
and U14933 (N_14933,N_10526,N_9300);
and U14934 (N_14934,N_10890,N_11493);
xor U14935 (N_14935,N_10128,N_11685);
xor U14936 (N_14936,N_10508,N_9200);
nand U14937 (N_14937,N_11112,N_10106);
nor U14938 (N_14938,N_10790,N_10508);
nand U14939 (N_14939,N_10968,N_10401);
or U14940 (N_14940,N_11914,N_11079);
and U14941 (N_14941,N_10738,N_10834);
nand U14942 (N_14942,N_9905,N_10562);
nor U14943 (N_14943,N_9626,N_11506);
nor U14944 (N_14944,N_10183,N_9359);
nand U14945 (N_14945,N_10961,N_10969);
xnor U14946 (N_14946,N_10293,N_10084);
or U14947 (N_14947,N_10659,N_9827);
and U14948 (N_14948,N_9948,N_9049);
nand U14949 (N_14949,N_11431,N_11599);
or U14950 (N_14950,N_10794,N_10217);
nor U14951 (N_14951,N_10188,N_9064);
and U14952 (N_14952,N_11610,N_10220);
nand U14953 (N_14953,N_9866,N_11665);
xor U14954 (N_14954,N_10561,N_10126);
xnor U14955 (N_14955,N_11519,N_11134);
and U14956 (N_14956,N_11785,N_10410);
or U14957 (N_14957,N_9240,N_9941);
or U14958 (N_14958,N_11909,N_10355);
and U14959 (N_14959,N_11929,N_9780);
and U14960 (N_14960,N_9587,N_11999);
and U14961 (N_14961,N_10772,N_10404);
xnor U14962 (N_14962,N_11753,N_10963);
nand U14963 (N_14963,N_9369,N_11517);
or U14964 (N_14964,N_11264,N_10779);
or U14965 (N_14965,N_11914,N_11535);
nor U14966 (N_14966,N_10859,N_9141);
xor U14967 (N_14967,N_11609,N_9744);
nor U14968 (N_14968,N_9678,N_11232);
or U14969 (N_14969,N_9687,N_10673);
nor U14970 (N_14970,N_9565,N_9466);
and U14971 (N_14971,N_10467,N_10864);
nor U14972 (N_14972,N_10923,N_9780);
or U14973 (N_14973,N_11152,N_9935);
nor U14974 (N_14974,N_11248,N_10232);
nand U14975 (N_14975,N_10356,N_9642);
and U14976 (N_14976,N_10998,N_11049);
nor U14977 (N_14977,N_9090,N_11744);
and U14978 (N_14978,N_10699,N_9973);
nand U14979 (N_14979,N_9624,N_9946);
and U14980 (N_14980,N_9030,N_9603);
nor U14981 (N_14981,N_9483,N_10079);
xor U14982 (N_14982,N_11764,N_11744);
nand U14983 (N_14983,N_11929,N_9122);
nor U14984 (N_14984,N_11552,N_11516);
and U14985 (N_14985,N_9879,N_9744);
xor U14986 (N_14986,N_9212,N_9140);
or U14987 (N_14987,N_11450,N_11584);
nor U14988 (N_14988,N_10459,N_10307);
and U14989 (N_14989,N_9116,N_10868);
and U14990 (N_14990,N_11743,N_11825);
and U14991 (N_14991,N_10983,N_11925);
xnor U14992 (N_14992,N_9842,N_10631);
and U14993 (N_14993,N_11893,N_9255);
nor U14994 (N_14994,N_11620,N_9246);
nand U14995 (N_14995,N_9650,N_11345);
nand U14996 (N_14996,N_11938,N_9868);
nand U14997 (N_14997,N_10424,N_10323);
or U14998 (N_14998,N_10673,N_10012);
or U14999 (N_14999,N_9769,N_9549);
and UO_0 (O_0,N_12957,N_13456);
or UO_1 (O_1,N_13934,N_13634);
xnor UO_2 (O_2,N_12015,N_13318);
nor UO_3 (O_3,N_12597,N_14126);
nor UO_4 (O_4,N_14371,N_13404);
and UO_5 (O_5,N_12417,N_13803);
and UO_6 (O_6,N_14636,N_12432);
or UO_7 (O_7,N_14276,N_13664);
nand UO_8 (O_8,N_14350,N_12745);
and UO_9 (O_9,N_13502,N_13773);
nor UO_10 (O_10,N_14867,N_14633);
and UO_11 (O_11,N_12826,N_13589);
or UO_12 (O_12,N_13518,N_14274);
nand UO_13 (O_13,N_14723,N_14556);
nand UO_14 (O_14,N_12727,N_14614);
nor UO_15 (O_15,N_12323,N_12392);
and UO_16 (O_16,N_13470,N_12462);
nand UO_17 (O_17,N_13985,N_13058);
nor UO_18 (O_18,N_13786,N_12492);
and UO_19 (O_19,N_14075,N_14794);
nor UO_20 (O_20,N_13458,N_14256);
nand UO_21 (O_21,N_14626,N_12967);
nand UO_22 (O_22,N_14721,N_14789);
nand UO_23 (O_23,N_12592,N_13876);
or UO_24 (O_24,N_14288,N_14422);
and UO_25 (O_25,N_14325,N_12687);
and UO_26 (O_26,N_12558,N_13667);
or UO_27 (O_27,N_14328,N_13693);
or UO_28 (O_28,N_12916,N_12645);
nor UO_29 (O_29,N_14922,N_14974);
and UO_30 (O_30,N_14404,N_13609);
or UO_31 (O_31,N_13274,N_13959);
nor UO_32 (O_32,N_12758,N_13223);
and UO_33 (O_33,N_12368,N_14216);
nand UO_34 (O_34,N_14188,N_12526);
nand UO_35 (O_35,N_14337,N_13856);
or UO_36 (O_36,N_13270,N_14985);
or UO_37 (O_37,N_14214,N_13428);
nand UO_38 (O_38,N_14012,N_13499);
or UO_39 (O_39,N_12096,N_12282);
and UO_40 (O_40,N_12334,N_14318);
nand UO_41 (O_41,N_12440,N_12494);
or UO_42 (O_42,N_12594,N_12322);
and UO_43 (O_43,N_12667,N_12875);
and UO_44 (O_44,N_12618,N_12636);
and UO_45 (O_45,N_13734,N_14360);
xnor UO_46 (O_46,N_12206,N_13151);
or UO_47 (O_47,N_14650,N_13186);
nor UO_48 (O_48,N_12286,N_12753);
xor UO_49 (O_49,N_13843,N_14973);
nor UO_50 (O_50,N_14174,N_13249);
nor UO_51 (O_51,N_13156,N_14099);
or UO_52 (O_52,N_12883,N_12347);
or UO_53 (O_53,N_12031,N_13036);
nand UO_54 (O_54,N_13874,N_13449);
nand UO_55 (O_55,N_12126,N_13300);
and UO_56 (O_56,N_12847,N_12622);
or UO_57 (O_57,N_12531,N_13132);
xnor UO_58 (O_58,N_13212,N_14811);
xnor UO_59 (O_59,N_12612,N_12128);
xor UO_60 (O_60,N_12375,N_13261);
and UO_61 (O_61,N_14403,N_14374);
nand UO_62 (O_62,N_13415,N_12223);
or UO_63 (O_63,N_13230,N_14107);
nor UO_64 (O_64,N_14200,N_14051);
nand UO_65 (O_65,N_14148,N_13507);
or UO_66 (O_66,N_12398,N_13932);
nor UO_67 (O_67,N_14184,N_13234);
xor UO_68 (O_68,N_14770,N_13878);
xnor UO_69 (O_69,N_12101,N_14815);
xnor UO_70 (O_70,N_13907,N_13911);
and UO_71 (O_71,N_14858,N_14102);
nand UO_72 (O_72,N_14322,N_12291);
nor UO_73 (O_73,N_12729,N_12129);
and UO_74 (O_74,N_12510,N_14895);
and UO_75 (O_75,N_13455,N_12247);
nor UO_76 (O_76,N_13930,N_14097);
nand UO_77 (O_77,N_13015,N_14952);
or UO_78 (O_78,N_12350,N_13776);
xor UO_79 (O_79,N_12751,N_12473);
nor UO_80 (O_80,N_12855,N_12318);
and UO_81 (O_81,N_14740,N_12150);
nand UO_82 (O_82,N_12119,N_14006);
xnor UO_83 (O_83,N_14294,N_14773);
nand UO_84 (O_84,N_13442,N_12045);
or UO_85 (O_85,N_12885,N_14924);
and UO_86 (O_86,N_12098,N_13477);
nor UO_87 (O_87,N_13780,N_13440);
or UO_88 (O_88,N_14571,N_14552);
or UO_89 (O_89,N_13432,N_13100);
or UO_90 (O_90,N_14821,N_13381);
xnor UO_91 (O_91,N_14395,N_12788);
nand UO_92 (O_92,N_13434,N_14824);
nand UO_93 (O_93,N_14275,N_14597);
nand UO_94 (O_94,N_12827,N_13526);
xor UO_95 (O_95,N_13235,N_14730);
nand UO_96 (O_96,N_12979,N_12458);
and UO_97 (O_97,N_14771,N_13850);
and UO_98 (O_98,N_14317,N_12520);
and UO_99 (O_99,N_14508,N_13965);
nor UO_100 (O_100,N_12325,N_12400);
nor UO_101 (O_101,N_14645,N_13338);
nor UO_102 (O_102,N_14084,N_14549);
nand UO_103 (O_103,N_13084,N_13669);
nand UO_104 (O_104,N_12730,N_13691);
and UO_105 (O_105,N_14451,N_14912);
nor UO_106 (O_106,N_12722,N_13747);
nand UO_107 (O_107,N_14864,N_12396);
xnor UO_108 (O_108,N_12770,N_13919);
nand UO_109 (O_109,N_12113,N_13062);
and UO_110 (O_110,N_13884,N_14304);
or UO_111 (O_111,N_14379,N_13943);
nand UO_112 (O_112,N_14843,N_13828);
nor UO_113 (O_113,N_13674,N_13666);
or UO_114 (O_114,N_13183,N_13886);
xnor UO_115 (O_115,N_14505,N_14566);
nor UO_116 (O_116,N_13161,N_12852);
and UO_117 (O_117,N_13574,N_13905);
nor UO_118 (O_118,N_14446,N_14273);
and UO_119 (O_119,N_14072,N_14798);
or UO_120 (O_120,N_13419,N_14070);
or UO_121 (O_121,N_12172,N_14550);
or UO_122 (O_122,N_14632,N_12313);
and UO_123 (O_123,N_12960,N_12507);
nand UO_124 (O_124,N_14932,N_14911);
and UO_125 (O_125,N_14358,N_14164);
or UO_126 (O_126,N_14106,N_13225);
and UO_127 (O_127,N_14837,N_13233);
nor UO_128 (O_128,N_12474,N_12246);
and UO_129 (O_129,N_12600,N_13347);
and UO_130 (O_130,N_14666,N_13559);
nand UO_131 (O_131,N_12429,N_12615);
and UO_132 (O_132,N_14090,N_14417);
nand UO_133 (O_133,N_14477,N_14928);
nor UO_134 (O_134,N_13144,N_13852);
nand UO_135 (O_135,N_12589,N_12424);
xor UO_136 (O_136,N_13054,N_14158);
xnor UO_137 (O_137,N_13475,N_13178);
nand UO_138 (O_138,N_13255,N_12574);
nor UO_139 (O_139,N_13018,N_13775);
nor UO_140 (O_140,N_14617,N_12648);
xor UO_141 (O_141,N_14476,N_14857);
nand UO_142 (O_142,N_14352,N_14363);
or UO_143 (O_143,N_13567,N_12312);
nand UO_144 (O_144,N_12833,N_13414);
and UO_145 (O_145,N_14714,N_14179);
xnor UO_146 (O_146,N_12330,N_12966);
xnor UO_147 (O_147,N_12905,N_14059);
or UO_148 (O_148,N_14865,N_12657);
nand UO_149 (O_149,N_14137,N_13515);
nand UO_150 (O_150,N_13126,N_14676);
nor UO_151 (O_151,N_12794,N_13637);
or UO_152 (O_152,N_12936,N_14988);
nor UO_153 (O_153,N_12864,N_13363);
or UO_154 (O_154,N_12561,N_14035);
nand UO_155 (O_155,N_13158,N_12523);
or UO_156 (O_156,N_13050,N_12351);
and UO_157 (O_157,N_12251,N_13060);
nand UO_158 (O_158,N_12190,N_12217);
and UO_159 (O_159,N_14983,N_12381);
nor UO_160 (O_160,N_12898,N_14224);
xnor UO_161 (O_161,N_13573,N_12656);
or UO_162 (O_162,N_14024,N_14027);
xnor UO_163 (O_163,N_12816,N_12388);
nand UO_164 (O_164,N_12470,N_13057);
or UO_165 (O_165,N_12796,N_14743);
nand UO_166 (O_166,N_13227,N_12066);
and UO_167 (O_167,N_14060,N_14405);
nor UO_168 (O_168,N_14255,N_12352);
and UO_169 (O_169,N_12534,N_13864);
or UO_170 (O_170,N_13582,N_14967);
nand UO_171 (O_171,N_13297,N_14088);
and UO_172 (O_172,N_13308,N_14205);
and UO_173 (O_173,N_14778,N_12203);
nand UO_174 (O_174,N_14194,N_13902);
and UO_175 (O_175,N_13752,N_12506);
nor UO_176 (O_176,N_12359,N_12385);
nor UO_177 (O_177,N_14327,N_13042);
or UO_178 (O_178,N_13447,N_13970);
xor UO_179 (O_179,N_13619,N_12644);
or UO_180 (O_180,N_14578,N_13024);
xnor UO_181 (O_181,N_12902,N_14287);
nor UO_182 (O_182,N_14298,N_14517);
nand UO_183 (O_183,N_13147,N_14885);
nand UO_184 (O_184,N_12938,N_12900);
xor UO_185 (O_185,N_14141,N_13330);
nor UO_186 (O_186,N_14774,N_14217);
nor UO_187 (O_187,N_12586,N_12660);
nor UO_188 (O_188,N_13598,N_14213);
xnor UO_189 (O_189,N_12348,N_12851);
nor UO_190 (O_190,N_14098,N_13554);
and UO_191 (O_191,N_14800,N_12487);
or UO_192 (O_192,N_13772,N_13372);
nand UO_193 (O_193,N_13968,N_12787);
nor UO_194 (O_194,N_12809,N_14277);
nand UO_195 (O_195,N_14863,N_14728);
nand UO_196 (O_196,N_14248,N_12001);
or UO_197 (O_197,N_14025,N_12339);
or UO_198 (O_198,N_12372,N_12465);
or UO_199 (O_199,N_12808,N_12430);
and UO_200 (O_200,N_13903,N_12115);
and UO_201 (O_201,N_13450,N_13185);
nand UO_202 (O_202,N_12909,N_14570);
nor UO_203 (O_203,N_13642,N_14999);
nor UO_204 (O_204,N_14031,N_13676);
nand UO_205 (O_205,N_14877,N_13200);
xnor UO_206 (O_206,N_13189,N_14760);
or UO_207 (O_207,N_14945,N_13472);
nand UO_208 (O_208,N_14943,N_12649);
nand UO_209 (O_209,N_14692,N_13695);
and UO_210 (O_210,N_12894,N_14329);
nand UO_211 (O_211,N_13999,N_13700);
or UO_212 (O_212,N_12479,N_12546);
or UO_213 (O_213,N_13343,N_13239);
and UO_214 (O_214,N_12502,N_13359);
and UO_215 (O_215,N_14268,N_13931);
and UO_216 (O_216,N_12248,N_14125);
xor UO_217 (O_217,N_12994,N_13659);
nor UO_218 (O_218,N_13528,N_14880);
or UO_219 (O_219,N_14267,N_14429);
nand UO_220 (O_220,N_14062,N_12374);
and UO_221 (O_221,N_12838,N_12178);
and UO_222 (O_222,N_12934,N_14584);
or UO_223 (O_223,N_12829,N_13694);
xnor UO_224 (O_224,N_14014,N_14369);
nor UO_225 (O_225,N_13236,N_14028);
nand UO_226 (O_226,N_12965,N_14407);
xor UO_227 (O_227,N_13599,N_13605);
and UO_228 (O_228,N_13867,N_14041);
nand UO_229 (O_229,N_14443,N_13909);
nand UO_230 (O_230,N_13661,N_14131);
and UO_231 (O_231,N_13877,N_13172);
and UO_232 (O_232,N_14900,N_13014);
nor UO_233 (O_233,N_14340,N_13335);
nor UO_234 (O_234,N_13378,N_14687);
xnor UO_235 (O_235,N_14489,N_13379);
nor UO_236 (O_236,N_13882,N_12448);
or UO_237 (O_237,N_13020,N_12873);
xnor UO_238 (O_238,N_14466,N_13096);
nand UO_239 (O_239,N_12877,N_13544);
nand UO_240 (O_240,N_13749,N_12650);
nand UO_241 (O_241,N_14719,N_12005);
and UO_242 (O_242,N_13820,N_13336);
and UO_243 (O_243,N_12870,N_13854);
nor UO_244 (O_244,N_13155,N_13504);
nor UO_245 (O_245,N_14044,N_12114);
nor UO_246 (O_246,N_13006,N_13851);
nand UO_247 (O_247,N_13992,N_12305);
nand UO_248 (O_248,N_13460,N_12270);
nand UO_249 (O_249,N_12509,N_13618);
nor UO_250 (O_250,N_12041,N_14752);
or UO_251 (O_251,N_13461,N_12197);
or UO_252 (O_252,N_13592,N_12680);
or UO_253 (O_253,N_12021,N_14233);
nor UO_254 (O_254,N_14047,N_14828);
nand UO_255 (O_255,N_14221,N_14496);
nand UO_256 (O_256,N_14279,N_12160);
or UO_257 (O_257,N_14039,N_13498);
or UO_258 (O_258,N_14845,N_14670);
and UO_259 (O_259,N_13056,N_14965);
nor UO_260 (O_260,N_14434,N_13658);
nand UO_261 (O_261,N_12969,N_14724);
xor UO_262 (O_262,N_13421,N_12266);
nand UO_263 (O_263,N_13751,N_14534);
and UO_264 (O_264,N_12185,N_14237);
nand UO_265 (O_265,N_13278,N_13352);
nand UO_266 (O_266,N_14426,N_12697);
or UO_267 (O_267,N_12177,N_14452);
nand UO_268 (O_268,N_12602,N_14649);
nand UO_269 (O_269,N_13536,N_13257);
xnor UO_270 (O_270,N_14860,N_14380);
nand UO_271 (O_271,N_13407,N_13037);
xor UO_272 (O_272,N_13304,N_13266);
or UO_273 (O_273,N_14309,N_13310);
nor UO_274 (O_274,N_14034,N_12797);
and UO_275 (O_275,N_14635,N_13153);
and UO_276 (O_276,N_13133,N_13842);
or UO_277 (O_277,N_13229,N_14573);
nor UO_278 (O_278,N_13469,N_14170);
nand UO_279 (O_279,N_12588,N_12775);
xnor UO_280 (O_280,N_14243,N_12846);
nor UO_281 (O_281,N_14618,N_13706);
nand UO_282 (O_282,N_13816,N_12174);
nand UO_283 (O_283,N_14113,N_13248);
or UO_284 (O_284,N_14726,N_13465);
nand UO_285 (O_285,N_14009,N_13433);
nor UO_286 (O_286,N_14907,N_12276);
xnor UO_287 (O_287,N_13958,N_13431);
or UO_288 (O_288,N_14398,N_13991);
and UO_289 (O_289,N_14227,N_12356);
nor UO_290 (O_290,N_13066,N_13832);
nand UO_291 (O_291,N_14167,N_13016);
nor UO_292 (O_292,N_14524,N_13106);
or UO_293 (O_293,N_12414,N_12253);
or UO_294 (O_294,N_14868,N_13323);
and UO_295 (O_295,N_12982,N_12920);
nand UO_296 (O_296,N_13644,N_13840);
xnor UO_297 (O_297,N_14850,N_12881);
nor UO_298 (O_298,N_13400,N_13837);
nor UO_299 (O_299,N_14286,N_12715);
xor UO_300 (O_300,N_13064,N_14450);
nor UO_301 (O_301,N_14874,N_12024);
xor UO_302 (O_302,N_12353,N_12040);
nor UO_303 (O_303,N_12989,N_12263);
and UO_304 (O_304,N_12472,N_13763);
nor UO_305 (O_305,N_14602,N_13730);
or UO_306 (O_306,N_14285,N_13918);
nor UO_307 (O_307,N_14942,N_12858);
and UO_308 (O_308,N_14510,N_13807);
or UO_309 (O_309,N_14947,N_13550);
nand UO_310 (O_310,N_13703,N_12054);
xor UO_311 (O_311,N_13813,N_14261);
nand UO_312 (O_312,N_13929,N_12516);
and UO_313 (O_313,N_12317,N_12383);
nor UO_314 (O_314,N_12605,N_14727);
and UO_315 (O_315,N_13324,N_12252);
xor UO_316 (O_316,N_12078,N_13231);
xor UO_317 (O_317,N_12839,N_12399);
and UO_318 (O_318,N_14690,N_14664);
nand UO_319 (O_319,N_13855,N_14454);
or UO_320 (O_320,N_14753,N_14546);
nor UO_321 (O_321,N_14223,N_13169);
nor UO_322 (O_322,N_14431,N_12964);
nor UO_323 (O_323,N_12933,N_13522);
or UO_324 (O_324,N_13648,N_12111);
nand UO_325 (O_325,N_14219,N_12848);
xnor UO_326 (O_326,N_13862,N_14447);
or UO_327 (O_327,N_14262,N_14756);
nor UO_328 (O_328,N_13289,N_12284);
and UO_329 (O_329,N_14418,N_14409);
and UO_330 (O_330,N_14342,N_12790);
and UO_331 (O_331,N_14581,N_13025);
or UO_332 (O_332,N_13952,N_13756);
nand UO_333 (O_333,N_14608,N_12793);
nand UO_334 (O_334,N_12550,N_13896);
or UO_335 (O_335,N_14893,N_12970);
nand UO_336 (O_336,N_13089,N_12559);
nand UO_337 (O_337,N_12955,N_13416);
or UO_338 (O_338,N_14657,N_13486);
or UO_339 (O_339,N_13569,N_13804);
xor UO_340 (O_340,N_14961,N_14105);
xnor UO_341 (O_341,N_12020,N_14225);
nor UO_342 (O_342,N_12642,N_14118);
or UO_343 (O_343,N_12490,N_12789);
or UO_344 (O_344,N_14343,N_14197);
and UO_345 (O_345,N_13859,N_13602);
and UO_346 (O_346,N_14879,N_12299);
nor UO_347 (O_347,N_12395,N_14604);
nor UO_348 (O_348,N_13360,N_13047);
or UO_349 (O_349,N_12482,N_12382);
nand UO_350 (O_350,N_13979,N_12537);
nor UO_351 (O_351,N_12568,N_13830);
xnor UO_352 (O_352,N_13645,N_14978);
and UO_353 (O_353,N_14071,N_13294);
nor UO_354 (O_354,N_14003,N_13949);
or UO_355 (O_355,N_14781,N_13681);
nor UO_356 (O_356,N_13170,N_13364);
nor UO_357 (O_357,N_13391,N_12918);
nand UO_358 (O_358,N_13821,N_14336);
nor UO_359 (O_359,N_13675,N_12447);
nor UO_360 (O_360,N_14356,N_12195);
or UO_361 (O_361,N_13429,N_13620);
and UO_362 (O_362,N_14751,N_13214);
xnor UO_363 (O_363,N_13596,N_12154);
or UO_364 (O_364,N_12986,N_13192);
nor UO_365 (O_365,N_14842,N_12962);
and UO_366 (O_366,N_12814,N_13105);
nand UO_367 (O_367,N_14143,N_12869);
and UO_368 (O_368,N_13279,N_13779);
nand UO_369 (O_369,N_12607,N_12579);
or UO_370 (O_370,N_14522,N_13941);
and UO_371 (O_371,N_14203,N_14465);
and UO_372 (O_372,N_12521,N_12893);
nor UO_373 (O_373,N_12082,N_12365);
nor UO_374 (O_374,N_12707,N_13789);
nor UO_375 (O_375,N_13412,N_12783);
nor UO_376 (O_376,N_14049,N_13496);
and UO_377 (O_377,N_13370,N_12355);
and UO_378 (O_378,N_14094,N_13549);
or UO_379 (O_379,N_13568,N_12393);
or UO_380 (O_380,N_13485,N_13946);
nor UO_381 (O_381,N_12327,N_14598);
or UO_382 (O_382,N_14580,N_12344);
or UO_383 (O_383,N_13835,N_14852);
nor UO_384 (O_384,N_13535,N_13430);
or UO_385 (O_385,N_13253,N_13474);
nor UO_386 (O_386,N_12407,N_12981);
and UO_387 (O_387,N_13765,N_13626);
or UO_388 (O_388,N_14430,N_14436);
and UO_389 (O_389,N_13514,N_14814);
nand UO_390 (O_390,N_12621,N_12874);
nor UO_391 (O_391,N_14957,N_13295);
nor UO_392 (O_392,N_13892,N_14182);
or UO_393 (O_393,N_13245,N_13858);
nor UO_394 (O_394,N_14272,N_14315);
and UO_395 (O_395,N_14007,N_14717);
nand UO_396 (O_396,N_13221,N_14475);
and UO_397 (O_397,N_14572,N_12678);
and UO_398 (O_398,N_13079,N_12932);
or UO_399 (O_399,N_14930,N_13405);
and UO_400 (O_400,N_12529,N_14045);
and UO_401 (O_401,N_12585,N_12801);
nor UO_402 (O_402,N_12210,N_12686);
nor UO_403 (O_403,N_13530,N_13390);
or UO_404 (O_404,N_12705,N_13376);
nand UO_405 (O_405,N_14545,N_13584);
nor UO_406 (O_406,N_12700,N_14400);
nand UO_407 (O_407,N_14055,N_13898);
nor UO_408 (O_408,N_12362,N_13870);
and UO_409 (O_409,N_13617,N_14242);
and UO_410 (O_410,N_14767,N_13099);
nor UO_411 (O_411,N_14122,N_14758);
or UO_412 (O_412,N_12911,N_14289);
xor UO_413 (O_413,N_14319,N_14801);
nor UO_414 (O_414,N_12153,N_14938);
or UO_415 (O_415,N_14949,N_12019);
nor UO_416 (O_416,N_13829,N_14691);
nand UO_417 (O_417,N_14290,N_13340);
nor UO_418 (O_418,N_12699,N_14816);
nand UO_419 (O_419,N_12739,N_12912);
nand UO_420 (O_420,N_12431,N_13277);
nand UO_421 (O_421,N_12990,N_13662);
and UO_422 (O_422,N_14790,N_12483);
and UO_423 (O_423,N_13216,N_12647);
or UO_424 (O_424,N_13413,N_12202);
and UO_425 (O_425,N_14577,N_12459);
and UO_426 (O_426,N_14392,N_13709);
and UO_427 (O_427,N_13871,N_14755);
nand UO_428 (O_428,N_13122,N_14416);
and UO_429 (O_429,N_12148,N_13962);
or UO_430 (O_430,N_12428,N_14019);
and UO_431 (O_431,N_13385,N_14228);
nand UO_432 (O_432,N_12692,N_12785);
or UO_433 (O_433,N_13800,N_13679);
nand UO_434 (O_434,N_14152,N_13441);
and UO_435 (O_435,N_14338,N_12086);
and UO_436 (O_436,N_12939,N_13040);
nor UO_437 (O_437,N_13796,N_13735);
or UO_438 (O_438,N_12360,N_14296);
nand UO_439 (O_439,N_13994,N_13166);
and UO_440 (O_440,N_12354,N_12209);
nand UO_441 (O_441,N_14487,N_14076);
xor UO_442 (O_442,N_13068,N_13349);
xor UO_443 (O_443,N_12065,N_12922);
nor UO_444 (O_444,N_12199,N_13205);
and UO_445 (O_445,N_12951,N_12403);
and UO_446 (O_446,N_13402,N_12071);
or UO_447 (O_447,N_12501,N_14906);
xor UO_448 (O_448,N_13729,N_13091);
and UO_449 (O_449,N_14054,N_12515);
nor UO_450 (O_450,N_12471,N_12555);
nor UO_451 (O_451,N_12701,N_13345);
and UO_452 (O_452,N_14787,N_12234);
xor UO_453 (O_453,N_12196,N_12243);
nor UO_454 (O_454,N_12110,N_12691);
nor UO_455 (O_455,N_12980,N_14544);
nor UO_456 (O_456,N_12168,N_14469);
and UO_457 (O_457,N_12281,N_14247);
xnor UO_458 (O_458,N_14372,N_12688);
nand UO_459 (O_459,N_14554,N_14722);
nor UO_460 (O_460,N_14791,N_14282);
and UO_461 (O_461,N_13631,N_13409);
xor UO_462 (O_462,N_12378,N_14897);
or UO_463 (O_463,N_12076,N_13947);
or UO_464 (O_464,N_14914,N_13382);
and UO_465 (O_465,N_12774,N_13792);
nand UO_466 (O_466,N_13731,N_14236);
nand UO_467 (O_467,N_12813,N_12135);
nand UO_468 (O_468,N_12614,N_13173);
and UO_469 (O_469,N_14481,N_13680);
nor UO_470 (O_470,N_12630,N_12876);
or UO_471 (O_471,N_14870,N_13553);
nand UO_472 (O_472,N_14810,N_12818);
and UO_473 (O_473,N_14206,N_12624);
nor UO_474 (O_474,N_12169,N_14023);
and UO_475 (O_475,N_14257,N_12498);
or UO_476 (O_476,N_12121,N_12928);
nand UO_477 (O_477,N_13924,N_13090);
or UO_478 (O_478,N_12999,N_12391);
nand UO_479 (O_479,N_14624,N_12485);
or UO_480 (O_480,N_13904,N_12144);
nand UO_481 (O_481,N_13065,N_13027);
nand UO_482 (O_482,N_12320,N_13198);
and UO_483 (O_483,N_12683,N_14799);
nand UO_484 (O_484,N_12401,N_13142);
or UO_485 (O_485,N_12792,N_14330);
or UO_486 (O_486,N_12158,N_12469);
or UO_487 (O_487,N_13080,N_13873);
and UO_488 (O_488,N_13444,N_14745);
and UO_489 (O_489,N_14013,N_12435);
nand UO_490 (O_490,N_12850,N_12930);
nand UO_491 (O_491,N_14630,N_12162);
nor UO_492 (O_492,N_14682,N_12845);
and UO_493 (O_493,N_13206,N_14341);
and UO_494 (O_494,N_13635,N_14887);
xnor UO_495 (O_495,N_12748,N_12496);
nand UO_496 (O_496,N_12231,N_12800);
nand UO_497 (O_497,N_13594,N_12200);
and UO_498 (O_498,N_13031,N_13244);
nand UO_499 (O_499,N_14600,N_12802);
and UO_500 (O_500,N_14929,N_12070);
and UO_501 (O_501,N_14656,N_12118);
and UO_502 (O_502,N_14933,N_12543);
or UO_503 (O_503,N_12508,N_12130);
or UO_504 (O_504,N_13782,N_13463);
and UO_505 (O_505,N_13622,N_13017);
and UO_506 (O_506,N_12861,N_13546);
xnor UO_507 (O_507,N_14565,N_12436);
nor UO_508 (O_508,N_12242,N_14079);
or UO_509 (O_509,N_13831,N_14478);
and UO_510 (O_510,N_12754,N_12068);
nand UO_511 (O_511,N_13000,N_14244);
nor UO_512 (O_512,N_12666,N_12048);
nor UO_513 (O_513,N_14103,N_12361);
nand UO_514 (O_514,N_13791,N_14130);
and UO_515 (O_515,N_13263,N_14994);
nand UO_516 (O_516,N_12386,N_13168);
nor UO_517 (O_517,N_13149,N_13657);
and UO_518 (O_518,N_12191,N_13226);
xor UO_519 (O_519,N_14889,N_14187);
nor UO_520 (O_520,N_12112,N_13583);
nor UO_521 (O_521,N_12868,N_14762);
and UO_522 (O_522,N_14920,N_14514);
nor UO_523 (O_523,N_13201,N_14193);
or UO_524 (O_524,N_14589,N_14504);
nor UO_525 (O_525,N_13910,N_14308);
nand UO_526 (O_526,N_12411,N_13557);
or UO_527 (O_527,N_14181,N_12324);
and UO_528 (O_528,N_13267,N_12817);
nand UO_529 (O_529,N_13111,N_12486);
nand UO_530 (O_530,N_12511,N_13464);
and UO_531 (O_531,N_14218,N_13880);
nand UO_532 (O_532,N_14734,N_13611);
nor UO_533 (O_533,N_13162,N_13808);
and UO_534 (O_534,N_14705,N_14738);
nor UO_535 (O_535,N_12298,N_12079);
nor UO_536 (O_536,N_14264,N_12677);
or UO_537 (O_537,N_12711,N_12890);
nor UO_538 (O_538,N_12819,N_13764);
xnor UO_539 (O_539,N_14110,N_13531);
nand UO_540 (O_540,N_13191,N_14612);
or UO_541 (O_541,N_13944,N_13104);
and UO_542 (O_542,N_14846,N_14512);
or UO_543 (O_543,N_12976,N_14551);
nand UO_544 (O_544,N_13685,N_12953);
nor UO_545 (O_545,N_12342,N_14997);
nand UO_546 (O_546,N_12500,N_14839);
xnor UO_547 (O_547,N_13866,N_14441);
or UO_548 (O_548,N_13606,N_14093);
nand UO_549 (O_549,N_13517,N_12563);
and UO_550 (O_550,N_14861,N_12077);
and UO_551 (O_551,N_13337,N_12632);
nor UO_552 (O_552,N_13788,N_14211);
nor UO_553 (O_553,N_14427,N_12878);
and UO_554 (O_554,N_13019,N_13610);
or UO_555 (O_555,N_13733,N_14526);
and UO_556 (O_556,N_13011,N_12535);
nand UO_557 (O_557,N_12553,N_13059);
and UO_558 (O_558,N_13766,N_14239);
or UO_559 (O_559,N_12651,N_14712);
nand UO_560 (O_560,N_12408,N_12913);
nand UO_561 (O_561,N_14733,N_12944);
nand UO_562 (O_562,N_14083,N_12345);
nor UO_563 (O_563,N_13603,N_13783);
nand UO_564 (O_564,N_12198,N_13002);
nor UO_565 (O_565,N_14827,N_14884);
nand UO_566 (O_566,N_12915,N_14896);
nor UO_567 (O_567,N_14357,N_12226);
or UO_568 (O_568,N_12063,N_13207);
and UO_569 (O_569,N_14796,N_14958);
nor UO_570 (O_570,N_12577,N_12369);
nand UO_571 (O_571,N_13686,N_13238);
nand UO_572 (O_572,N_13714,N_14412);
nand UO_573 (O_573,N_14196,N_13119);
nor UO_574 (O_574,N_12702,N_14804);
or UO_575 (O_575,N_12549,N_13211);
nand UO_576 (O_576,N_12974,N_14586);
and UO_577 (O_577,N_12002,N_14568);
nand UO_578 (O_578,N_12109,N_13978);
nand UO_579 (O_579,N_12917,N_14128);
and UO_580 (O_580,N_12300,N_13129);
nand UO_581 (O_581,N_14923,N_13913);
or UO_582 (O_582,N_13275,N_13491);
nand UO_583 (O_583,N_12409,N_13443);
nor UO_584 (O_584,N_12131,N_14388);
or UO_585 (O_585,N_13542,N_12238);
or UO_586 (O_586,N_13759,N_13801);
and UO_587 (O_587,N_12992,N_12328);
and UO_588 (O_588,N_12825,N_13403);
or UO_589 (O_589,N_13322,N_14312);
nor UO_590 (O_590,N_13092,N_13711);
nand UO_591 (O_591,N_14855,N_13928);
and UO_592 (O_592,N_12562,N_12569);
xor UO_593 (O_593,N_13672,N_14208);
nand UO_594 (O_594,N_12366,N_14872);
nand UO_595 (O_595,N_14866,N_13964);
and UO_596 (O_596,N_13719,N_14095);
nand UO_597 (O_597,N_14809,N_13265);
and UO_598 (O_598,N_14678,N_12204);
nor UO_599 (O_599,N_14960,N_14004);
nor UO_600 (O_600,N_14706,N_13917);
nor UO_601 (O_601,N_13013,N_12638);
or UO_602 (O_602,N_13621,N_14888);
or UO_603 (O_603,N_13476,N_14472);
nor UO_604 (O_604,N_14192,N_14711);
and UO_605 (O_605,N_13136,N_12619);
nand UO_606 (O_606,N_14419,N_14396);
or UO_607 (O_607,N_12937,N_13303);
nand UO_608 (O_608,N_12044,N_12343);
nand UO_609 (O_609,N_13087,N_12467);
or UO_610 (O_610,N_14313,N_13194);
or UO_611 (O_611,N_13509,N_14525);
or UO_612 (O_612,N_14297,N_13586);
xor UO_613 (O_613,N_14591,N_14331);
nor UO_614 (O_614,N_13283,N_14931);
and UO_615 (O_615,N_12724,N_13160);
and UO_616 (O_616,N_13769,N_13001);
xnor UO_617 (O_617,N_14354,N_13237);
nand UO_618 (O_618,N_14067,N_12439);
or UO_619 (O_619,N_14011,N_13446);
and UO_620 (O_620,N_12948,N_12983);
and UO_621 (O_621,N_12461,N_12484);
nor UO_622 (O_622,N_13588,N_13453);
nand UO_623 (O_623,N_12503,N_14953);
xnor UO_624 (O_624,N_14222,N_13298);
or UO_625 (O_625,N_14807,N_13241);
and UO_626 (O_626,N_13607,N_14432);
xor UO_627 (O_627,N_12108,N_12192);
nand UO_628 (O_628,N_14854,N_12228);
and UO_629 (O_629,N_12371,N_14548);
or UO_630 (O_630,N_14471,N_13117);
or UO_631 (O_631,N_13511,N_14520);
and UO_632 (O_632,N_13581,N_12629);
nor UO_633 (O_633,N_14859,N_13737);
xnor UO_634 (O_634,N_13616,N_14016);
and UO_635 (O_635,N_12011,N_13109);
and UO_636 (O_636,N_14826,N_12142);
nor UO_637 (O_637,N_14393,N_13923);
or UO_638 (O_638,N_13145,N_12042);
xnor UO_639 (O_639,N_12259,N_12806);
or UO_640 (O_640,N_14840,N_14500);
or UO_641 (O_641,N_13493,N_13593);
nand UO_642 (O_642,N_14523,N_14259);
nor UO_643 (O_643,N_13448,N_13757);
nand UO_644 (O_644,N_13728,N_14502);
or UO_645 (O_645,N_13551,N_13725);
nor UO_646 (O_646,N_13250,N_14862);
nand UO_647 (O_647,N_12149,N_13795);
and UO_648 (O_648,N_12713,N_12946);
and UO_649 (O_649,N_12294,N_14377);
or UO_650 (O_650,N_14461,N_12106);
nand UO_651 (O_651,N_12942,N_13224);
nand UO_652 (O_652,N_13677,N_14621);
nand UO_653 (O_653,N_14642,N_14043);
nor UO_654 (O_654,N_13328,N_12116);
nor UO_655 (O_655,N_14669,N_14127);
nand UO_656 (O_656,N_14414,N_13762);
or UO_657 (O_657,N_14823,N_14848);
and UO_658 (O_658,N_14903,N_12036);
nor UO_659 (O_659,N_13671,N_13668);
nand UO_660 (O_660,N_12812,N_13955);
or UO_661 (O_661,N_12513,N_13386);
nor UO_662 (O_662,N_14366,N_14937);
nand UO_663 (O_663,N_13125,N_14195);
and UO_664 (O_664,N_13595,N_12961);
or UO_665 (O_665,N_14339,N_13750);
nand UO_666 (O_666,N_13052,N_14702);
nand UO_667 (O_667,N_14479,N_13638);
and UO_668 (O_668,N_12643,N_13371);
and UO_669 (O_669,N_14744,N_12333);
and UO_670 (O_670,N_14449,N_14623);
and UO_671 (O_671,N_13987,N_12567);
or UO_672 (O_672,N_12584,N_14190);
or UO_673 (O_673,N_14644,N_12220);
nand UO_674 (O_674,N_13457,N_12706);
or UO_675 (O_675,N_14806,N_14776);
or UO_676 (O_676,N_14927,N_13745);
and UO_677 (O_677,N_13921,N_13342);
nor UO_678 (O_678,N_14064,N_13118);
nand UO_679 (O_679,N_14010,N_14646);
nand UO_680 (O_680,N_14533,N_13427);
nor UO_681 (O_681,N_14963,N_12147);
nand UO_682 (O_682,N_13778,N_12201);
and UO_683 (O_683,N_13920,N_13687);
or UO_684 (O_684,N_13790,N_12186);
nor UO_685 (O_685,N_12043,N_12427);
nor UO_686 (O_686,N_14444,N_12180);
or UO_687 (O_687,N_12358,N_14081);
or UO_688 (O_688,N_13481,N_12968);
or UO_689 (O_689,N_13861,N_13697);
xnor UO_690 (O_690,N_13196,N_13836);
and UO_691 (O_691,N_12720,N_13576);
and UO_692 (O_692,N_13422,N_13063);
or UO_693 (O_693,N_14119,N_12279);
xor UO_694 (O_694,N_14186,N_14000);
and UO_695 (O_695,N_14672,N_14841);
xor UO_696 (O_696,N_14355,N_14836);
nand UO_697 (O_697,N_14156,N_13417);
and UO_698 (O_698,N_13114,N_13713);
and UO_699 (O_699,N_13654,N_12823);
and UO_700 (O_700,N_12759,N_13067);
or UO_701 (O_701,N_12244,N_12338);
or UO_702 (O_702,N_14497,N_14665);
and UO_703 (O_703,N_12945,N_13314);
nor UO_704 (O_704,N_13998,N_13306);
xor UO_705 (O_705,N_12413,N_13377);
or UO_706 (O_706,N_13954,N_14559);
nor UO_707 (O_707,N_13879,N_12815);
or UO_708 (O_708,N_12766,N_14606);
nor UO_709 (O_709,N_13950,N_12696);
or UO_710 (O_710,N_13411,N_14087);
nand UO_711 (O_711,N_13562,N_13146);
xnor UO_712 (O_712,N_14917,N_12804);
or UO_713 (O_713,N_12213,N_14576);
xnor UO_714 (O_714,N_13960,N_13176);
and UO_715 (O_715,N_14998,N_14833);
nand UO_716 (O_716,N_12446,N_13222);
nand UO_717 (O_717,N_12326,N_12742);
or UO_718 (O_718,N_13088,N_12376);
nand UO_719 (O_719,N_13356,N_14984);
and UO_720 (O_720,N_14324,N_13101);
and UO_721 (O_721,N_13143,N_13438);
nor UO_722 (O_722,N_13956,N_14348);
nor UO_723 (O_723,N_12547,N_12971);
nand UO_724 (O_724,N_12545,N_13321);
nand UO_725 (O_725,N_14486,N_14793);
nor UO_726 (O_726,N_13333,N_14780);
or UO_727 (O_727,N_12927,N_13218);
nand UO_728 (O_728,N_12996,N_12489);
or UO_729 (O_729,N_13344,N_13003);
or UO_730 (O_730,N_12522,N_12122);
or UO_731 (O_731,N_13963,N_12641);
and UO_732 (O_732,N_13007,N_12752);
nor UO_733 (O_733,N_13140,N_12560);
or UO_734 (O_734,N_13811,N_14876);
and UO_735 (O_735,N_13809,N_14519);
nand UO_736 (O_736,N_12184,N_12662);
nand UO_737 (O_737,N_12117,N_13484);
or UO_738 (O_738,N_14513,N_12302);
or UO_739 (O_739,N_14303,N_12684);
and UO_740 (O_740,N_12593,N_14168);
nand UO_741 (O_741,N_13317,N_12099);
and UO_742 (O_742,N_14101,N_14688);
nor UO_743 (O_743,N_14150,N_13311);
nor UO_744 (O_744,N_12987,N_14822);
nor UO_745 (O_745,N_13350,N_12285);
and UO_746 (O_746,N_14401,N_12750);
or UO_747 (O_747,N_12954,N_13927);
nor UO_748 (O_748,N_14299,N_13008);
nand UO_749 (O_749,N_12069,N_14622);
and UO_750 (O_750,N_14271,N_14108);
nor UO_751 (O_751,N_12164,N_14198);
or UO_752 (O_752,N_14601,N_13035);
nand UO_753 (O_753,N_12663,N_12995);
and UO_754 (O_754,N_13260,N_12887);
or UO_755 (O_755,N_13839,N_14516);
nand UO_756 (O_756,N_14663,N_13848);
and UO_757 (O_757,N_13293,N_12437);
nor UO_758 (O_758,N_14467,N_13961);
xor UO_759 (O_759,N_12693,N_12665);
nand UO_760 (O_760,N_14104,N_13702);
and UO_761 (O_761,N_14748,N_12941);
and UO_762 (O_762,N_13665,N_14640);
nor UO_763 (O_763,N_14361,N_14026);
nor UO_764 (O_764,N_14818,N_14610);
or UO_765 (O_765,N_14693,N_12956);
nand UO_766 (O_766,N_14066,N_14492);
or UO_767 (O_767,N_12779,N_13139);
nand UO_768 (O_768,N_13906,N_14629);
or UO_769 (O_769,N_12346,N_12717);
nor UO_770 (O_770,N_14718,N_12309);
or UO_771 (O_771,N_13369,N_13933);
and UO_772 (O_772,N_13467,N_14424);
nor UO_773 (O_773,N_14729,N_14437);
or UO_774 (O_774,N_14232,N_14538);
or UO_775 (O_775,N_13726,N_13157);
or UO_776 (O_776,N_13754,N_12084);
nand UO_777 (O_777,N_14849,N_14121);
nand UO_778 (O_778,N_14485,N_14058);
nand UO_779 (O_779,N_12640,N_13785);
nand UO_780 (O_780,N_13437,N_14935);
and UO_781 (O_781,N_12389,N_12859);
or UO_782 (O_782,N_13826,N_14307);
nor UO_783 (O_783,N_14518,N_13915);
and UO_784 (O_784,N_13215,N_12258);
or UO_785 (O_785,N_14674,N_14503);
nor UO_786 (O_786,N_14695,N_12512);
or UO_787 (O_787,N_12871,N_14391);
or UO_788 (O_788,N_14891,N_13718);
nor UO_789 (O_789,N_13570,N_13655);
xor UO_790 (O_790,N_13563,N_12025);
or UO_791 (O_791,N_13580,N_12073);
or UO_792 (O_792,N_14283,N_13041);
nor UO_793 (O_793,N_14680,N_13121);
nand UO_794 (O_794,N_14310,N_12623);
or UO_795 (O_795,N_12030,N_13516);
nor UO_796 (O_796,N_14291,N_12016);
or UO_797 (O_797,N_13110,N_14112);
or UO_798 (O_798,N_14699,N_13394);
or UO_799 (O_799,N_14241,N_14293);
nor UO_800 (O_800,N_12772,N_14345);
nor UO_801 (O_801,N_13174,N_14406);
nor UO_802 (O_802,N_14749,N_13976);
and UO_803 (O_803,N_12773,N_14709);
nor UO_804 (O_804,N_12580,N_13124);
and UO_805 (O_805,N_13397,N_13810);
and UO_806 (O_806,N_14694,N_14229);
xor UO_807 (O_807,N_14445,N_12714);
or UO_808 (O_808,N_14660,N_14490);
nand UO_809 (O_809,N_13393,N_12003);
xnor UO_810 (O_810,N_13276,N_14038);
or UO_811 (O_811,N_12761,N_12425);
nand UO_812 (O_812,N_14413,N_14609);
or UO_813 (O_813,N_13555,N_13990);
nor UO_814 (O_814,N_12269,N_14782);
or UO_815 (O_815,N_12854,N_12083);
xnor UO_816 (O_816,N_12176,N_14944);
nand UO_817 (O_817,N_12646,N_14529);
nor UO_818 (O_818,N_12769,N_14869);
and UO_819 (O_819,N_12241,N_12734);
and UO_820 (O_820,N_14596,N_13889);
nor UO_821 (O_821,N_12280,N_13232);
nand UO_822 (O_822,N_13534,N_12179);
and UO_823 (O_823,N_12331,N_12821);
nor UO_824 (O_824,N_13942,N_13048);
nor UO_825 (O_825,N_14134,N_14507);
and UO_826 (O_826,N_14382,N_13723);
nand UO_827 (O_827,N_14458,N_12012);
nor UO_828 (O_828,N_12541,N_13937);
or UO_829 (O_829,N_14089,N_13767);
nand UO_830 (O_830,N_14091,N_12527);
nand UO_831 (O_831,N_12006,N_14462);
nor UO_832 (O_832,N_13339,N_12963);
or UO_833 (O_833,N_14527,N_13724);
nand UO_834 (O_834,N_12053,N_12997);
xor UO_835 (O_835,N_12422,N_12193);
or UO_836 (O_836,N_12173,N_12007);
nor UO_837 (O_837,N_13299,N_12914);
or UO_838 (O_838,N_12892,N_12274);
and UO_839 (O_839,N_14667,N_12133);
or UO_840 (O_840,N_12170,N_12364);
nand UO_841 (O_841,N_13738,N_12085);
nor UO_842 (O_842,N_14402,N_12682);
or UO_843 (O_843,N_13647,N_14677);
or UO_844 (O_844,N_14563,N_12155);
and UO_845 (O_845,N_13663,N_12418);
nand UO_846 (O_846,N_14063,N_14036);
and UO_847 (O_847,N_13288,N_14521);
and UO_848 (O_848,N_12767,N_12257);
and UO_849 (O_849,N_14830,N_13558);
and UO_850 (O_850,N_13410,N_14111);
nor UO_851 (O_851,N_14962,N_14739);
or UO_852 (O_852,N_14052,N_12740);
and UO_853 (O_853,N_13868,N_14539);
nand UO_854 (O_854,N_13969,N_12221);
nor UO_855 (O_855,N_13973,N_14590);
or UO_856 (O_856,N_13152,N_14173);
and UO_857 (O_857,N_13758,N_14258);
and UO_858 (O_858,N_12138,N_14741);
nor UO_859 (O_859,N_12950,N_12337);
or UO_860 (O_860,N_12565,N_12314);
xnor UO_861 (O_861,N_14235,N_13210);
and UO_862 (O_862,N_14151,N_13971);
and UO_863 (O_863,N_12124,N_13888);
nor UO_864 (O_864,N_12505,N_13552);
or UO_865 (O_865,N_14701,N_12654);
and UO_866 (O_866,N_13291,N_12857);
and UO_867 (O_867,N_14387,N_14021);
or UO_868 (O_868,N_14311,N_12732);
nor UO_869 (O_869,N_13181,N_13247);
xor UO_870 (O_870,N_14269,N_14553);
or UO_871 (O_871,N_13579,N_13228);
nand UO_872 (O_872,N_13698,N_14939);
and UO_873 (O_873,N_14772,N_12457);
nand UO_874 (O_874,N_12703,N_14161);
xor UO_875 (O_875,N_14558,N_13893);
nand UO_876 (O_876,N_12497,N_12379);
or UO_877 (O_877,N_12637,N_12888);
nor UO_878 (O_878,N_12091,N_13505);
nand UO_879 (O_879,N_14831,N_14231);
nor UO_880 (O_880,N_12095,N_12140);
nor UO_881 (O_881,N_12278,N_14435);
nor UO_882 (O_882,N_13510,N_14708);
and UO_883 (O_883,N_14484,N_12064);
or UO_884 (O_884,N_12704,N_12889);
or UO_885 (O_885,N_14139,N_12661);
xor UO_886 (O_886,N_13900,N_14230);
or UO_887 (O_887,N_14171,N_14746);
or UO_888 (O_888,N_14175,N_14916);
or UO_889 (O_889,N_13327,N_12214);
nor UO_890 (O_890,N_14704,N_13459);
xor UO_891 (O_891,N_13967,N_14316);
nor UO_892 (O_892,N_12867,N_14300);
nand UO_893 (O_893,N_12008,N_14390);
and UO_894 (O_894,N_12161,N_12205);
and UO_895 (O_895,N_12207,N_14189);
or UO_896 (O_896,N_14133,N_12907);
nand UO_897 (O_897,N_14587,N_12763);
and UO_898 (O_898,N_14784,N_13073);
or UO_899 (O_899,N_14883,N_12795);
nor UO_900 (O_900,N_13154,N_14783);
nand UO_901 (O_901,N_13305,N_14234);
nand UO_902 (O_902,N_14731,N_14698);
nor UO_903 (O_903,N_12652,N_14856);
nor UO_904 (O_904,N_14685,N_13175);
or UO_905 (O_905,N_12296,N_12604);
or UO_906 (O_906,N_13190,N_14114);
or UO_907 (O_907,N_13823,N_13717);
xnor UO_908 (O_908,N_12952,N_13578);
or UO_909 (O_909,N_12709,N_12272);
and UO_910 (O_910,N_13332,N_12405);
or UO_911 (O_911,N_12450,N_14292);
and UO_912 (O_912,N_13130,N_13627);
nor UO_913 (O_913,N_13282,N_12896);
nor UO_914 (O_914,N_14941,N_12988);
and UO_915 (O_915,N_14918,N_13891);
nand UO_916 (O_916,N_12052,N_12211);
xnor UO_917 (O_917,N_14162,N_12639);
nand UO_918 (O_918,N_12463,N_12977);
or UO_919 (O_919,N_12227,N_14808);
nand UO_920 (O_920,N_14263,N_12626);
and UO_921 (O_921,N_13953,N_12308);
or UO_922 (O_922,N_14117,N_13727);
or UO_923 (O_923,N_12167,N_12139);
nor UO_924 (O_924,N_12000,N_12387);
or UO_925 (O_925,N_12778,N_12037);
or UO_926 (O_926,N_12477,N_13246);
or UO_927 (O_927,N_13012,N_12499);
nand UO_928 (O_928,N_12551,N_13600);
and UO_929 (O_929,N_12655,N_12055);
nor UO_930 (O_930,N_14613,N_14386);
or UO_931 (O_931,N_13643,N_14116);
and UO_932 (O_932,N_13597,N_13545);
xor UO_933 (O_933,N_14881,N_14619);
nand UO_934 (O_934,N_14593,N_13857);
and UO_935 (O_935,N_14499,N_14819);
nor UO_936 (O_936,N_14056,N_12010);
nand UO_937 (O_937,N_12504,N_13296);
and UO_938 (O_938,N_14191,N_13538);
nor UO_939 (O_939,N_14109,N_12698);
nor UO_940 (O_940,N_14029,N_12570);
nand UO_941 (O_941,N_13532,N_13380);
nor UO_942 (O_942,N_12674,N_13521);
nand UO_943 (O_943,N_13846,N_13494);
nor UO_944 (O_944,N_14488,N_14768);
and UO_945 (O_945,N_13993,N_12218);
nand UO_946 (O_946,N_14802,N_12321);
nor UO_947 (O_947,N_13197,N_13179);
nor UO_948 (O_948,N_14132,N_13102);
or UO_949 (O_949,N_12975,N_13707);
or UO_950 (O_950,N_13495,N_12420);
or UO_951 (O_951,N_13029,N_13972);
nor UO_952 (O_952,N_14375,N_13072);
nor UO_953 (O_953,N_14002,N_14302);
nor UO_954 (O_954,N_13537,N_13784);
nor UO_955 (O_955,N_14306,N_13374);
nand UO_956 (O_956,N_14483,N_14585);
and UO_957 (O_957,N_13252,N_14575);
nor UO_958 (O_958,N_14344,N_12578);
nand UO_959 (O_959,N_12137,N_13529);
nand UO_960 (O_960,N_12764,N_14266);
nand UO_961 (O_961,N_12319,N_13439);
nand UO_962 (O_962,N_14653,N_13033);
and UO_963 (O_963,N_13615,N_12716);
and UO_964 (O_964,N_12837,N_14926);
and UO_965 (O_965,N_12441,N_14018);
xnor UO_966 (O_966,N_14648,N_13290);
nor UO_967 (O_967,N_14470,N_13543);
or UO_968 (O_968,N_13123,N_12476);
nor UO_969 (O_969,N_14428,N_14981);
or UO_970 (O_970,N_13112,N_13399);
nor UO_971 (O_971,N_12056,N_12628);
nor UO_972 (O_972,N_14595,N_14147);
nor UO_973 (O_973,N_13004,N_13392);
or UO_974 (O_974,N_12768,N_12575);
nor UO_975 (O_975,N_13022,N_12183);
nor UO_976 (O_976,N_14875,N_12120);
nor UO_977 (O_977,N_13478,N_14964);
and UO_978 (O_978,N_12668,N_14154);
or UO_979 (O_979,N_14433,N_12616);
and UO_980 (O_980,N_14955,N_14812);
and UO_981 (O_981,N_13670,N_12475);
or UO_982 (O_982,N_14383,N_13220);
xor UO_983 (O_983,N_14641,N_13565);
nor UO_984 (O_984,N_13204,N_13838);
nor UO_985 (O_985,N_12538,N_14989);
nor UO_986 (O_986,N_13912,N_14567);
and UO_987 (O_987,N_13113,N_14792);
or UO_988 (O_988,N_13082,N_13167);
xnor UO_989 (O_989,N_12884,N_14178);
xnor UO_990 (O_990,N_12777,N_12601);
or UO_991 (O_991,N_14163,N_14180);
and UO_992 (O_992,N_14683,N_13794);
nand UO_993 (O_993,N_13078,N_13629);
and UO_994 (O_994,N_13083,N_12250);
nand UO_995 (O_995,N_12542,N_14913);
nor UO_996 (O_996,N_12288,N_13712);
nand UO_997 (O_997,N_12136,N_14910);
nor UO_998 (O_998,N_12728,N_12719);
nand UO_999 (O_999,N_14638,N_14415);
nor UO_1000 (O_1000,N_13512,N_12921);
nand UO_1001 (O_1001,N_12256,N_14564);
or UO_1002 (O_1002,N_13046,N_12514);
or UO_1003 (O_1003,N_12596,N_12212);
or UO_1004 (O_1004,N_12233,N_12303);
or UO_1005 (O_1005,N_13503,N_13740);
and UO_1006 (O_1006,N_13895,N_13590);
nor UO_1007 (O_1007,N_14115,N_12018);
and UO_1008 (O_1008,N_13639,N_13164);
nand UO_1009 (O_1009,N_13280,N_13319);
nand UO_1010 (O_1010,N_13897,N_12239);
and UO_1011 (O_1011,N_13793,N_12060);
or UO_1012 (O_1012,N_14144,N_12958);
nand UO_1013 (O_1013,N_13781,N_13650);
or UO_1014 (O_1014,N_14995,N_12679);
nand UO_1015 (O_1015,N_14976,N_12306);
or UO_1016 (O_1016,N_13075,N_12891);
nand UO_1017 (O_1017,N_14599,N_13701);
xnor UO_1018 (O_1018,N_12406,N_12225);
nand UO_1019 (O_1019,N_14971,N_14046);
and UO_1020 (O_1020,N_14332,N_14871);
nor UO_1021 (O_1021,N_12478,N_13032);
or UO_1022 (O_1022,N_12820,N_13986);
nand UO_1023 (O_1023,N_13256,N_12442);
and UO_1024 (O_1024,N_12710,N_14140);
and UO_1025 (O_1025,N_14611,N_12416);
nor UO_1026 (O_1026,N_14684,N_14160);
xnor UO_1027 (O_1027,N_12488,N_13043);
or UO_1028 (O_1028,N_13743,N_13690);
nand UO_1029 (O_1029,N_13471,N_14226);
and UO_1030 (O_1030,N_13085,N_12620);
and UO_1031 (O_1031,N_13366,N_14238);
nand UO_1032 (O_1032,N_14716,N_13150);
or UO_1033 (O_1033,N_13732,N_13948);
and UO_1034 (O_1034,N_13540,N_13682);
and UO_1035 (O_1035,N_13744,N_14169);
and UO_1036 (O_1036,N_12292,N_14651);
xnor UO_1037 (O_1037,N_14639,N_14561);
and UO_1038 (O_1038,N_14440,N_13454);
or UO_1039 (O_1039,N_12034,N_12237);
or UO_1040 (O_1040,N_12843,N_13329);
or UO_1041 (O_1041,N_13787,N_14157);
nand UO_1042 (O_1042,N_13134,N_12978);
nand UO_1043 (O_1043,N_12171,N_12830);
nor UO_1044 (O_1044,N_13375,N_14700);
and UO_1045 (O_1045,N_13420,N_12879);
and UO_1046 (O_1046,N_14786,N_12175);
xor UO_1047 (O_1047,N_13575,N_13689);
nor UO_1048 (O_1048,N_13482,N_13199);
xnor UO_1049 (O_1049,N_14250,N_13890);
nand UO_1050 (O_1050,N_12984,N_13489);
xnor UO_1051 (O_1051,N_13389,N_12943);
or UO_1052 (O_1052,N_13488,N_14323);
nor UO_1053 (O_1053,N_12023,N_13899);
nand UO_1054 (O_1054,N_12603,N_13049);
xnor UO_1055 (O_1055,N_12092,N_12232);
or UO_1056 (O_1056,N_14439,N_12438);
and UO_1057 (O_1057,N_14210,N_13302);
and UO_1058 (O_1058,N_13539,N_13865);
nor UO_1059 (O_1059,N_12690,N_13883);
nor UO_1060 (O_1060,N_14777,N_12842);
nor UO_1061 (O_1061,N_12582,N_13396);
nor UO_1062 (O_1062,N_13423,N_13069);
nor UO_1063 (O_1063,N_14142,N_12017);
nor UO_1064 (O_1064,N_13699,N_14251);
or UO_1065 (O_1065,N_14803,N_13989);
xor UO_1066 (O_1066,N_13171,N_13827);
nor UO_1067 (O_1067,N_14788,N_14951);
nor UO_1068 (O_1068,N_13849,N_13320);
nand UO_1069 (O_1069,N_14463,N_12576);
nor UO_1070 (O_1070,N_14456,N_12072);
xnor UO_1071 (O_1071,N_14817,N_12685);
or UO_1072 (O_1072,N_14155,N_12631);
or UO_1073 (O_1073,N_12156,N_13331);
nand UO_1074 (O_1074,N_12610,N_13524);
or UO_1075 (O_1075,N_13716,N_14321);
nand UO_1076 (O_1076,N_12824,N_13268);
or UO_1077 (O_1077,N_14365,N_13451);
and UO_1078 (O_1078,N_12495,N_12776);
and UO_1079 (O_1079,N_12673,N_12132);
or UO_1080 (O_1080,N_13982,N_12712);
or UO_1081 (O_1081,N_14085,N_13922);
and UO_1082 (O_1082,N_13653,N_13914);
nand UO_1083 (O_1083,N_12349,N_13894);
and UO_1084 (O_1084,N_13487,N_12081);
and UO_1085 (O_1085,N_12277,N_13354);
and UO_1086 (O_1086,N_12765,N_13026);
nor UO_1087 (O_1087,N_12782,N_13462);
or UO_1088 (O_1088,N_13269,N_12723);
nand UO_1089 (O_1089,N_12762,N_12240);
nor UO_1090 (O_1090,N_12028,N_14785);
or UO_1091 (O_1091,N_12419,N_12182);
and UO_1092 (O_1092,N_12840,N_13135);
xnor UO_1093 (O_1093,N_14346,N_13869);
or UO_1094 (O_1094,N_14399,N_14353);
nand UO_1095 (O_1095,N_12102,N_14425);
nor UO_1096 (O_1096,N_13984,N_14509);
nor UO_1097 (O_1097,N_12080,N_12454);
or UO_1098 (O_1098,N_13541,N_13287);
and UO_1099 (O_1099,N_12444,N_12061);
and UO_1100 (O_1100,N_14954,N_13797);
and UO_1101 (O_1101,N_13103,N_13281);
nor UO_1102 (O_1102,N_12412,N_14389);
and UO_1103 (O_1103,N_12756,N_12341);
nand UO_1104 (O_1104,N_12090,N_12552);
nand UO_1105 (O_1105,N_14847,N_12718);
and UO_1106 (O_1106,N_14579,N_14681);
nand UO_1107 (O_1107,N_14703,N_13513);
nand UO_1108 (O_1108,N_13988,N_12127);
nand UO_1109 (O_1109,N_12088,N_14659);
nor UO_1110 (O_1110,N_13070,N_12163);
or UO_1111 (O_1111,N_13326,N_14574);
nor UO_1112 (O_1112,N_14086,N_12835);
and UO_1113 (O_1113,N_14825,N_14813);
or UO_1114 (O_1114,N_14829,N_13887);
nor UO_1115 (O_1115,N_13209,N_12026);
nand UO_1116 (O_1116,N_14940,N_13120);
nor UO_1117 (O_1117,N_13180,N_14878);
and UO_1118 (O_1118,N_13587,N_13313);
and UO_1119 (O_1119,N_14040,N_12760);
and UO_1120 (O_1120,N_14838,N_12836);
or UO_1121 (O_1121,N_14397,N_14742);
xor UO_1122 (O_1122,N_12853,N_13137);
nand UO_1123 (O_1123,N_14073,N_14757);
and UO_1124 (O_1124,N_13564,N_12828);
and UO_1125 (O_1125,N_12973,N_13916);
and UO_1126 (O_1126,N_13863,N_12681);
xnor UO_1127 (O_1127,N_14607,N_12397);
and UO_1128 (O_1128,N_14212,N_14634);
and UO_1129 (O_1129,N_14246,N_13720);
nand UO_1130 (O_1130,N_14270,N_12544);
nand UO_1131 (O_1131,N_12721,N_12157);
or UO_1132 (O_1132,N_12449,N_13107);
or UO_1133 (O_1133,N_12810,N_12336);
nor UO_1134 (O_1134,N_12107,N_13213);
nor UO_1135 (O_1135,N_12583,N_13408);
and UO_1136 (O_1136,N_12062,N_13480);
nand UO_1137 (O_1137,N_12089,N_14373);
nor UO_1138 (O_1138,N_13116,N_12901);
and UO_1139 (O_1139,N_13501,N_13548);
or UO_1140 (O_1140,N_14754,N_13966);
or UO_1141 (O_1141,N_14265,N_13760);
xor UO_1142 (O_1142,N_12807,N_13074);
nor UO_1143 (O_1143,N_12781,N_13812);
or UO_1144 (O_1144,N_13346,N_12059);
or UO_1145 (O_1145,N_13817,N_14096);
nand UO_1146 (O_1146,N_13081,N_14370);
xor UO_1147 (O_1147,N_14411,N_14069);
and UO_1148 (O_1148,N_13005,N_13138);
nor UO_1149 (O_1149,N_13497,N_13613);
and UO_1150 (O_1150,N_12658,N_12746);
nand UO_1151 (O_1151,N_12249,N_12557);
or UO_1152 (O_1152,N_14378,N_13094);
nor UO_1153 (O_1153,N_12771,N_12991);
xor UO_1154 (O_1154,N_14410,N_13710);
nand UO_1155 (O_1155,N_12947,N_14245);
nand UO_1156 (O_1156,N_14153,N_14351);
nand UO_1157 (O_1157,N_13715,N_14805);
nor UO_1158 (O_1158,N_12735,N_14844);
xnor UO_1159 (O_1159,N_14582,N_14763);
nand UO_1160 (O_1160,N_13872,N_14124);
and UO_1161 (O_1161,N_13805,N_13184);
or UO_1162 (O_1162,N_13753,N_14359);
and UO_1163 (O_1163,N_12786,N_14689);
and UO_1164 (O_1164,N_13802,N_13021);
and UO_1165 (O_1165,N_13799,N_14460);
xnor UO_1166 (O_1166,N_13395,N_12453);
and UO_1167 (O_1167,N_14468,N_12390);
xnor UO_1168 (O_1168,N_12301,N_14491);
nor UO_1169 (O_1169,N_14423,N_13981);
xor UO_1170 (O_1170,N_13814,N_14252);
nor UO_1171 (O_1171,N_13755,N_13577);
nor UO_1172 (O_1172,N_14530,N_12254);
or UO_1173 (O_1173,N_13361,N_13051);
nand UO_1174 (O_1174,N_13030,N_12737);
nand UO_1175 (O_1175,N_12047,N_13061);
and UO_1176 (O_1176,N_13875,N_14696);
xor UO_1177 (O_1177,N_13315,N_14647);
and UO_1178 (O_1178,N_12929,N_14686);
nor UO_1179 (O_1179,N_12590,N_13881);
nor UO_1180 (O_1180,N_14996,N_14240);
and UO_1181 (O_1181,N_13527,N_14655);
and UO_1182 (O_1182,N_12599,N_12566);
or UO_1183 (O_1183,N_14050,N_13351);
xor UO_1184 (O_1184,N_14201,N_14882);
nor UO_1185 (O_1185,N_14149,N_14146);
nor UO_1186 (O_1186,N_13479,N_13038);
or UO_1187 (O_1187,N_14421,N_12152);
and UO_1188 (O_1188,N_12670,N_12726);
and UO_1189 (O_1189,N_12022,N_14515);
nor UO_1190 (O_1190,N_13571,N_12571);
nand UO_1191 (O_1191,N_12694,N_13187);
and UO_1192 (O_1192,N_14120,N_14899);
nor UO_1193 (O_1193,N_12260,N_13547);
and UO_1194 (O_1194,N_12035,N_12803);
nand UO_1195 (O_1195,N_12540,N_12736);
and UO_1196 (O_1196,N_12075,N_13202);
nand UO_1197 (O_1197,N_13365,N_14908);
or UO_1198 (O_1198,N_14384,N_13980);
or UO_1199 (O_1199,N_14901,N_14915);
nor UO_1200 (O_1200,N_14020,N_13977);
nor UO_1201 (O_1201,N_14394,N_14969);
nand UO_1202 (O_1202,N_13483,N_12027);
nor UO_1203 (O_1203,N_12100,N_14005);
or UO_1204 (O_1204,N_14775,N_12865);
and UO_1205 (O_1205,N_14832,N_14725);
or UO_1206 (O_1206,N_14562,N_12159);
nor UO_1207 (O_1207,N_12261,N_13771);
or UO_1208 (O_1208,N_13721,N_13844);
nor UO_1209 (O_1209,N_14747,N_14367);
nand UO_1210 (O_1210,N_13128,N_14668);
and UO_1211 (O_1211,N_12998,N_13741);
nor UO_1212 (O_1212,N_12923,N_13822);
nor UO_1213 (O_1213,N_14183,N_14675);
xor UO_1214 (O_1214,N_13401,N_12695);
nand UO_1215 (O_1215,N_12455,N_13935);
xor UO_1216 (O_1216,N_14199,N_13165);
or UO_1217 (O_1217,N_12731,N_12822);
and UO_1218 (O_1218,N_12402,N_14030);
or UO_1219 (O_1219,N_12524,N_12307);
nand UO_1220 (O_1220,N_14284,N_12798);
nand UO_1221 (O_1221,N_14008,N_12895);
or UO_1222 (O_1222,N_13243,N_13939);
xor UO_1223 (O_1223,N_12311,N_14820);
nand UO_1224 (O_1224,N_13996,N_12434);
nor UO_1225 (O_1225,N_12067,N_14934);
nand UO_1226 (O_1226,N_14215,N_12749);
nor UO_1227 (O_1227,N_13656,N_14123);
or UO_1228 (O_1228,N_13325,N_14536);
nand UO_1229 (O_1229,N_14453,N_12295);
and UO_1230 (O_1230,N_13975,N_12264);
nand UO_1231 (O_1231,N_14501,N_13115);
nor UO_1232 (O_1232,N_13240,N_14991);
xnor UO_1233 (O_1233,N_13926,N_12959);
nand UO_1234 (O_1234,N_12491,N_13722);
or UO_1235 (O_1235,N_12564,N_12165);
nand UO_1236 (O_1236,N_14735,N_14498);
xnor UO_1237 (O_1237,N_13818,N_12151);
and UO_1238 (O_1238,N_13572,N_12290);
nor UO_1239 (O_1239,N_12468,N_13309);
nor UO_1240 (O_1240,N_13708,N_14779);
nor UO_1241 (O_1241,N_14894,N_12332);
nor UO_1242 (O_1242,N_12224,N_14057);
and UO_1243 (O_1243,N_14720,N_14202);
nand UO_1244 (O_1244,N_12262,N_13940);
and UO_1245 (O_1245,N_12784,N_12811);
or UO_1246 (O_1246,N_14616,N_13908);
nand UO_1247 (O_1247,N_14061,N_12834);
and UO_1248 (O_1248,N_14165,N_13633);
nand UO_1249 (O_1249,N_12525,N_14592);
xor UO_1250 (O_1250,N_14959,N_14074);
xor UO_1251 (O_1251,N_12316,N_13614);
or UO_1252 (O_1252,N_13646,N_12268);
nand UO_1253 (O_1253,N_13632,N_14022);
nor UO_1254 (O_1254,N_13819,N_12532);
nor UO_1255 (O_1255,N_13761,N_12103);
or UO_1256 (O_1256,N_13039,N_12480);
xnor UO_1257 (O_1257,N_12097,N_12123);
or UO_1258 (O_1258,N_13251,N_12039);
nand UO_1259 (O_1259,N_14904,N_13436);
nand UO_1260 (O_1260,N_13885,N_14506);
nor UO_1261 (O_1261,N_13825,N_13806);
nor UO_1262 (O_1262,N_12926,N_14979);
and UO_1263 (O_1263,N_12013,N_12367);
or UO_1264 (O_1264,N_13847,N_12906);
and UO_1265 (O_1265,N_13660,N_13525);
nor UO_1266 (O_1266,N_12181,N_12304);
nand UO_1267 (O_1267,N_12554,N_14605);
xnor UO_1268 (O_1268,N_12493,N_12009);
nor UO_1269 (O_1269,N_14925,N_12528);
nor UO_1270 (O_1270,N_14368,N_13770);
and UO_1271 (O_1271,N_12613,N_12675);
and UO_1272 (O_1272,N_13383,N_14457);
nand UO_1273 (O_1273,N_13936,N_12189);
or UO_1274 (O_1274,N_14715,N_14438);
or UO_1275 (O_1275,N_14658,N_13163);
nor UO_1276 (O_1276,N_14092,N_12046);
nor UO_1277 (O_1277,N_12229,N_13983);
nand UO_1278 (O_1278,N_12572,N_13217);
xnor UO_1279 (O_1279,N_14732,N_12519);
xor UO_1280 (O_1280,N_12271,N_12669);
nand UO_1281 (O_1281,N_12897,N_14835);
xor UO_1282 (O_1282,N_12844,N_13853);
nand UO_1283 (O_1283,N_14541,N_13307);
and UO_1284 (O_1284,N_13636,N_13774);
nand UO_1285 (O_1285,N_14032,N_13159);
nor UO_1286 (O_1286,N_14902,N_13098);
nor UO_1287 (O_1287,N_14077,N_14207);
nand UO_1288 (O_1288,N_14921,N_12394);
or UO_1289 (O_1289,N_14543,N_12595);
nor UO_1290 (O_1290,N_14053,N_13426);
nand UO_1291 (O_1291,N_14557,N_14972);
nand UO_1292 (O_1292,N_14892,N_13452);
or UO_1293 (O_1293,N_14713,N_13108);
nand UO_1294 (O_1294,N_12443,N_13506);
nor UO_1295 (O_1295,N_13860,N_12335);
or UO_1296 (O_1296,N_12460,N_13468);
and UO_1297 (O_1297,N_12860,N_13841);
nand UO_1298 (O_1298,N_12862,N_12384);
and UO_1299 (O_1299,N_13045,N_14254);
or UO_1300 (O_1300,N_14946,N_14511);
or UO_1301 (O_1301,N_12141,N_13641);
or UO_1302 (O_1302,N_13673,N_14966);
xnor UO_1303 (O_1303,N_14547,N_14588);
or UO_1304 (O_1304,N_12733,N_12791);
xor UO_1305 (O_1305,N_12275,N_14459);
nand UO_1306 (O_1306,N_12404,N_14992);
nand UO_1307 (O_1307,N_12410,N_12676);
or UO_1308 (O_1308,N_12380,N_13591);
or UO_1309 (O_1309,N_13435,N_13640);
and UO_1310 (O_1310,N_12672,N_14919);
and UO_1311 (O_1311,N_13053,N_14138);
and UO_1312 (O_1312,N_13034,N_12886);
nor UO_1313 (O_1313,N_12245,N_14628);
nand UO_1314 (O_1314,N_12145,N_12757);
and UO_1315 (O_1315,N_14766,N_12051);
or UO_1316 (O_1316,N_14673,N_13316);
or UO_1317 (O_1317,N_13705,N_13071);
xor UO_1318 (O_1318,N_14970,N_12598);
nor UO_1319 (O_1319,N_12880,N_13262);
nand UO_1320 (O_1320,N_13561,N_13519);
nand UO_1321 (O_1321,N_12014,N_12653);
xnor UO_1322 (O_1322,N_14661,N_13254);
nand UO_1323 (O_1323,N_13777,N_13612);
nand UO_1324 (O_1324,N_14736,N_14851);
nand UO_1325 (O_1325,N_14537,N_12146);
xnor UO_1326 (O_1326,N_12634,N_14129);
or UO_1327 (O_1327,N_13341,N_14455);
nand UO_1328 (O_1328,N_14950,N_13097);
xor UO_1329 (O_1329,N_12841,N_13623);
xnor UO_1330 (O_1330,N_13077,N_13264);
xor UO_1331 (O_1331,N_12370,N_13739);
nand UO_1332 (O_1332,N_12993,N_13523);
nor UO_1333 (O_1333,N_14528,N_12134);
or UO_1334 (O_1334,N_12985,N_14333);
or UO_1335 (O_1335,N_14349,N_12940);
nand UO_1336 (O_1336,N_12166,N_13258);
or UO_1337 (O_1337,N_14697,N_13353);
xnor UO_1338 (O_1338,N_12050,N_14662);
nor UO_1339 (O_1339,N_14314,N_12741);
nand UO_1340 (O_1340,N_13997,N_13500);
xor UO_1341 (O_1341,N_12105,N_12518);
or UO_1342 (O_1342,N_14975,N_12882);
xnor UO_1343 (O_1343,N_13177,N_12451);
nand UO_1344 (O_1344,N_13692,N_12533);
or UO_1345 (O_1345,N_12057,N_12315);
nor UO_1346 (O_1346,N_12215,N_12049);
nor UO_1347 (O_1347,N_14542,N_12094);
or UO_1348 (O_1348,N_14671,N_12287);
nand UO_1349 (O_1349,N_12924,N_12235);
nand UO_1350 (O_1350,N_14555,N_13095);
or UO_1351 (O_1351,N_12340,N_14909);
and UO_1352 (O_1352,N_12423,N_12466);
nor UO_1353 (O_1353,N_13076,N_12293);
xor UO_1354 (O_1354,N_14797,N_12187);
nand UO_1355 (O_1355,N_12609,N_13388);
or UO_1356 (O_1356,N_13492,N_13748);
nor UO_1357 (O_1357,N_12872,N_14873);
and UO_1358 (O_1358,N_13357,N_13742);
nor UO_1359 (O_1359,N_12743,N_13974);
xor UO_1360 (O_1360,N_12297,N_14159);
nand UO_1361 (O_1361,N_14764,N_14048);
nand UO_1362 (O_1362,N_14710,N_13649);
and UO_1363 (O_1363,N_13995,N_12671);
nand UO_1364 (O_1364,N_13010,N_14652);
xnor UO_1365 (O_1365,N_12627,N_12029);
nand UO_1366 (O_1366,N_13824,N_14068);
xnor UO_1367 (O_1367,N_14890,N_13208);
nor UO_1368 (O_1368,N_14448,N_13023);
nand UO_1369 (O_1369,N_13368,N_13141);
nor UO_1370 (O_1370,N_13242,N_13560);
and UO_1371 (O_1371,N_12255,N_12517);
nor UO_1372 (O_1372,N_12377,N_14569);
nand UO_1373 (O_1373,N_12863,N_13901);
and UO_1374 (O_1374,N_13678,N_14065);
nand UO_1375 (O_1375,N_14987,N_12708);
or UO_1376 (O_1376,N_13608,N_12747);
xnor UO_1377 (O_1377,N_14185,N_14376);
or UO_1378 (O_1378,N_13624,N_12456);
and UO_1379 (O_1379,N_12548,N_13312);
nor UO_1380 (O_1380,N_14037,N_12033);
nand UO_1381 (O_1381,N_13585,N_14166);
and UO_1382 (O_1382,N_14278,N_14637);
nor UO_1383 (O_1383,N_14474,N_12452);
or UO_1384 (O_1384,N_12363,N_14795);
or UO_1385 (O_1385,N_13131,N_13292);
and UO_1386 (O_1386,N_12004,N_13348);
nor UO_1387 (O_1387,N_13285,N_12536);
or UO_1388 (O_1388,N_13286,N_13398);
and UO_1389 (O_1389,N_13334,N_12799);
and UO_1390 (O_1390,N_14993,N_14625);
and UO_1391 (O_1391,N_12899,N_13601);
or UO_1392 (O_1392,N_14364,N_14295);
nand UO_1393 (O_1393,N_12573,N_14334);
nand UO_1394 (O_1394,N_12949,N_14707);
nor UO_1395 (O_1395,N_12329,N_14532);
nor UO_1396 (O_1396,N_13490,N_13704);
or UO_1397 (O_1397,N_14408,N_12935);
nor UO_1398 (O_1398,N_13406,N_12931);
and UO_1399 (O_1399,N_14100,N_13688);
and UO_1400 (O_1400,N_14627,N_12725);
or UO_1401 (O_1401,N_12093,N_12755);
or UO_1402 (O_1402,N_12230,N_13628);
nand UO_1403 (O_1403,N_13009,N_13384);
and UO_1404 (O_1404,N_13625,N_14898);
and UO_1405 (O_1405,N_14420,N_13044);
xnor UO_1406 (O_1406,N_14362,N_12464);
and UO_1407 (O_1407,N_12581,N_14603);
and UO_1408 (O_1408,N_14654,N_14482);
nor UO_1409 (O_1409,N_14765,N_14015);
and UO_1410 (O_1410,N_13055,N_14750);
nor UO_1411 (O_1411,N_12265,N_14305);
and UO_1412 (O_1412,N_12866,N_14078);
and UO_1413 (O_1413,N_13373,N_13367);
or UO_1414 (O_1414,N_12087,N_12421);
nand UO_1415 (O_1415,N_13193,N_14281);
or UO_1416 (O_1416,N_14209,N_14977);
nand UO_1417 (O_1417,N_14968,N_14326);
and UO_1418 (O_1418,N_14172,N_14594);
nand UO_1419 (O_1419,N_13203,N_14001);
nand UO_1420 (O_1420,N_12635,N_13284);
xnor UO_1421 (O_1421,N_14761,N_13815);
xnor UO_1422 (O_1422,N_12539,N_13798);
nor UO_1423 (O_1423,N_13358,N_13259);
and UO_1424 (O_1424,N_12208,N_14531);
nor UO_1425 (O_1425,N_12283,N_12611);
or UO_1426 (O_1426,N_13148,N_12273);
and UO_1427 (O_1427,N_12910,N_13684);
nand UO_1428 (O_1428,N_13746,N_12606);
or UO_1429 (O_1429,N_13736,N_14769);
and UO_1430 (O_1430,N_12426,N_14301);
nor UO_1431 (O_1431,N_13473,N_12104);
nor UO_1432 (O_1432,N_12689,N_13195);
and UO_1433 (O_1433,N_12267,N_12591);
nor UO_1434 (O_1434,N_12445,N_14560);
or UO_1435 (O_1435,N_12289,N_14956);
nand UO_1436 (O_1436,N_12530,N_12972);
nand UO_1437 (O_1437,N_13556,N_13833);
or UO_1438 (O_1438,N_12222,N_14204);
nor UO_1439 (O_1439,N_12236,N_14493);
and UO_1440 (O_1440,N_14631,N_14615);
nor UO_1441 (O_1441,N_14948,N_13630);
or UO_1442 (O_1442,N_14320,N_14679);
or UO_1443 (O_1443,N_13362,N_14495);
nor UO_1444 (O_1444,N_14473,N_14385);
or UO_1445 (O_1445,N_13951,N_12216);
nand UO_1446 (O_1446,N_12415,N_13387);
nand UO_1447 (O_1447,N_13533,N_13925);
and UO_1448 (O_1448,N_13834,N_12925);
nand UO_1449 (O_1449,N_12664,N_13093);
nor UO_1450 (O_1450,N_14737,N_14136);
nor UO_1451 (O_1451,N_14643,N_14082);
and UO_1452 (O_1452,N_13520,N_14220);
nor UO_1453 (O_1453,N_12856,N_13271);
nor UO_1454 (O_1454,N_12659,N_13957);
nor UO_1455 (O_1455,N_14017,N_12832);
or UO_1456 (O_1456,N_13272,N_13445);
nor UO_1457 (O_1457,N_12625,N_12738);
and UO_1458 (O_1458,N_14620,N_14905);
xnor UO_1459 (O_1459,N_12038,N_14033);
nor UO_1460 (O_1460,N_14480,N_13355);
nor UO_1461 (O_1461,N_12219,N_13127);
nor UO_1462 (O_1462,N_13945,N_13651);
and UO_1463 (O_1463,N_12433,N_13696);
or UO_1464 (O_1464,N_12903,N_14381);
nor UO_1465 (O_1465,N_12831,N_14540);
nand UO_1466 (O_1466,N_14853,N_14583);
xnor UO_1467 (O_1467,N_12608,N_14335);
nor UO_1468 (O_1468,N_14464,N_12849);
nor UO_1469 (O_1469,N_14176,N_12143);
nor UO_1470 (O_1470,N_13273,N_14280);
xor UO_1471 (O_1471,N_13301,N_12556);
and UO_1472 (O_1472,N_14990,N_12904);
or UO_1473 (O_1473,N_12633,N_13652);
nor UO_1474 (O_1474,N_14535,N_12310);
nand UO_1475 (O_1475,N_13424,N_13418);
or UO_1476 (O_1476,N_14135,N_13086);
nor UO_1477 (O_1477,N_14936,N_12188);
nor UO_1478 (O_1478,N_14145,N_14260);
nor UO_1479 (O_1479,N_13466,N_12125);
and UO_1480 (O_1480,N_14494,N_13188);
nand UO_1481 (O_1481,N_13219,N_13028);
nor UO_1482 (O_1482,N_12032,N_13938);
nand UO_1483 (O_1483,N_14982,N_12373);
nand UO_1484 (O_1484,N_12194,N_12908);
and UO_1485 (O_1485,N_13683,N_14886);
nor UO_1486 (O_1486,N_13845,N_12074);
and UO_1487 (O_1487,N_14759,N_12805);
nor UO_1488 (O_1488,N_12058,N_13768);
or UO_1489 (O_1489,N_12744,N_13425);
and UO_1490 (O_1490,N_14347,N_14080);
and UO_1491 (O_1491,N_14042,N_14986);
or UO_1492 (O_1492,N_12587,N_13182);
nor UO_1493 (O_1493,N_12357,N_14253);
and UO_1494 (O_1494,N_12919,N_14177);
nand UO_1495 (O_1495,N_12481,N_12617);
and UO_1496 (O_1496,N_13508,N_14249);
or UO_1497 (O_1497,N_13604,N_14442);
nor UO_1498 (O_1498,N_14834,N_14980);
nand UO_1499 (O_1499,N_13566,N_12780);
nor UO_1500 (O_1500,N_12442,N_12783);
and UO_1501 (O_1501,N_12217,N_12587);
nand UO_1502 (O_1502,N_13050,N_14573);
and UO_1503 (O_1503,N_14068,N_14564);
nand UO_1504 (O_1504,N_12168,N_13276);
nand UO_1505 (O_1505,N_13622,N_13961);
nand UO_1506 (O_1506,N_13142,N_13959);
nand UO_1507 (O_1507,N_14537,N_13310);
nand UO_1508 (O_1508,N_12298,N_13013);
nand UO_1509 (O_1509,N_13853,N_12140);
xnor UO_1510 (O_1510,N_12593,N_13953);
and UO_1511 (O_1511,N_14579,N_13218);
nor UO_1512 (O_1512,N_13555,N_12342);
nand UO_1513 (O_1513,N_13556,N_12336);
and UO_1514 (O_1514,N_14928,N_14577);
nor UO_1515 (O_1515,N_13189,N_12335);
nor UO_1516 (O_1516,N_12113,N_12709);
xnor UO_1517 (O_1517,N_13880,N_14802);
nand UO_1518 (O_1518,N_13949,N_13441);
and UO_1519 (O_1519,N_12824,N_14985);
xor UO_1520 (O_1520,N_13270,N_13960);
xnor UO_1521 (O_1521,N_14705,N_13422);
or UO_1522 (O_1522,N_13583,N_14666);
or UO_1523 (O_1523,N_12001,N_12627);
and UO_1524 (O_1524,N_14046,N_14589);
or UO_1525 (O_1525,N_12447,N_12196);
nor UO_1526 (O_1526,N_13761,N_13847);
nor UO_1527 (O_1527,N_14100,N_14216);
or UO_1528 (O_1528,N_14618,N_12288);
nand UO_1529 (O_1529,N_12866,N_12107);
or UO_1530 (O_1530,N_13178,N_12472);
or UO_1531 (O_1531,N_12759,N_12836);
nor UO_1532 (O_1532,N_12829,N_13249);
and UO_1533 (O_1533,N_12770,N_13858);
and UO_1534 (O_1534,N_14173,N_14560);
nand UO_1535 (O_1535,N_14795,N_14860);
nor UO_1536 (O_1536,N_13736,N_13092);
xnor UO_1537 (O_1537,N_14578,N_12882);
nand UO_1538 (O_1538,N_13271,N_14347);
or UO_1539 (O_1539,N_12117,N_13501);
nand UO_1540 (O_1540,N_13454,N_14209);
or UO_1541 (O_1541,N_13303,N_13154);
nor UO_1542 (O_1542,N_14625,N_12846);
xor UO_1543 (O_1543,N_13448,N_13228);
or UO_1544 (O_1544,N_14550,N_14582);
nor UO_1545 (O_1545,N_13862,N_13426);
and UO_1546 (O_1546,N_13730,N_12343);
and UO_1547 (O_1547,N_13274,N_14158);
nor UO_1548 (O_1548,N_12940,N_14235);
nand UO_1549 (O_1549,N_12291,N_14629);
nor UO_1550 (O_1550,N_14965,N_12499);
xor UO_1551 (O_1551,N_13394,N_12119);
nand UO_1552 (O_1552,N_12106,N_14054);
xor UO_1553 (O_1553,N_12118,N_14955);
nor UO_1554 (O_1554,N_13575,N_13861);
and UO_1555 (O_1555,N_12174,N_12424);
nand UO_1556 (O_1556,N_14932,N_12504);
nand UO_1557 (O_1557,N_13631,N_14141);
or UO_1558 (O_1558,N_14940,N_12591);
nor UO_1559 (O_1559,N_12302,N_14384);
or UO_1560 (O_1560,N_14376,N_14721);
nand UO_1561 (O_1561,N_12675,N_14353);
nor UO_1562 (O_1562,N_14525,N_12171);
nand UO_1563 (O_1563,N_13952,N_13335);
and UO_1564 (O_1564,N_12575,N_13664);
nor UO_1565 (O_1565,N_13416,N_14099);
nand UO_1566 (O_1566,N_14270,N_13034);
nor UO_1567 (O_1567,N_14277,N_13579);
nor UO_1568 (O_1568,N_12885,N_12624);
nand UO_1569 (O_1569,N_14727,N_12641);
and UO_1570 (O_1570,N_14914,N_14646);
nand UO_1571 (O_1571,N_12183,N_13142);
xnor UO_1572 (O_1572,N_14652,N_12643);
or UO_1573 (O_1573,N_13963,N_12504);
nor UO_1574 (O_1574,N_13595,N_13326);
and UO_1575 (O_1575,N_13046,N_12150);
xnor UO_1576 (O_1576,N_14312,N_12208);
or UO_1577 (O_1577,N_13473,N_13142);
nand UO_1578 (O_1578,N_13994,N_12728);
nand UO_1579 (O_1579,N_13812,N_13611);
nand UO_1580 (O_1580,N_14913,N_14954);
or UO_1581 (O_1581,N_14554,N_14933);
and UO_1582 (O_1582,N_14254,N_14537);
nand UO_1583 (O_1583,N_14078,N_12030);
or UO_1584 (O_1584,N_13296,N_12873);
or UO_1585 (O_1585,N_12944,N_12535);
and UO_1586 (O_1586,N_13991,N_12515);
xnor UO_1587 (O_1587,N_13770,N_14817);
or UO_1588 (O_1588,N_12392,N_13034);
nand UO_1589 (O_1589,N_13493,N_13489);
and UO_1590 (O_1590,N_13926,N_12609);
nand UO_1591 (O_1591,N_13091,N_13951);
xor UO_1592 (O_1592,N_14927,N_12483);
nor UO_1593 (O_1593,N_12119,N_14796);
and UO_1594 (O_1594,N_14285,N_12395);
and UO_1595 (O_1595,N_13869,N_12399);
nand UO_1596 (O_1596,N_12004,N_13038);
nor UO_1597 (O_1597,N_12405,N_12017);
nor UO_1598 (O_1598,N_12288,N_13664);
and UO_1599 (O_1599,N_13664,N_12468);
or UO_1600 (O_1600,N_13078,N_13772);
nand UO_1601 (O_1601,N_12102,N_12575);
and UO_1602 (O_1602,N_14401,N_14948);
nor UO_1603 (O_1603,N_13314,N_14058);
nor UO_1604 (O_1604,N_13907,N_12326);
nand UO_1605 (O_1605,N_12831,N_14205);
xor UO_1606 (O_1606,N_13723,N_12315);
nor UO_1607 (O_1607,N_13408,N_12352);
or UO_1608 (O_1608,N_14835,N_12568);
or UO_1609 (O_1609,N_14206,N_14433);
and UO_1610 (O_1610,N_14937,N_14992);
nor UO_1611 (O_1611,N_13681,N_12649);
and UO_1612 (O_1612,N_12490,N_13910);
xnor UO_1613 (O_1613,N_13997,N_13860);
nor UO_1614 (O_1614,N_14465,N_12212);
nor UO_1615 (O_1615,N_14153,N_12092);
and UO_1616 (O_1616,N_14987,N_13557);
or UO_1617 (O_1617,N_14610,N_12185);
and UO_1618 (O_1618,N_14656,N_13967);
xor UO_1619 (O_1619,N_13079,N_14971);
xnor UO_1620 (O_1620,N_13390,N_14302);
and UO_1621 (O_1621,N_12857,N_12454);
nor UO_1622 (O_1622,N_12781,N_14947);
xnor UO_1623 (O_1623,N_14723,N_12677);
or UO_1624 (O_1624,N_13250,N_14341);
nor UO_1625 (O_1625,N_14792,N_14783);
or UO_1626 (O_1626,N_13441,N_12753);
xnor UO_1627 (O_1627,N_12332,N_12650);
nor UO_1628 (O_1628,N_14462,N_14291);
nand UO_1629 (O_1629,N_12972,N_12783);
xor UO_1630 (O_1630,N_14606,N_14586);
and UO_1631 (O_1631,N_14154,N_12315);
xor UO_1632 (O_1632,N_12416,N_13925);
and UO_1633 (O_1633,N_12982,N_12444);
or UO_1634 (O_1634,N_14456,N_14848);
or UO_1635 (O_1635,N_14358,N_12860);
xor UO_1636 (O_1636,N_12515,N_13234);
nand UO_1637 (O_1637,N_14487,N_13029);
nor UO_1638 (O_1638,N_13380,N_12798);
and UO_1639 (O_1639,N_14144,N_12942);
nand UO_1640 (O_1640,N_12668,N_13299);
nand UO_1641 (O_1641,N_12528,N_13050);
nor UO_1642 (O_1642,N_12515,N_13422);
and UO_1643 (O_1643,N_14238,N_12926);
or UO_1644 (O_1644,N_12091,N_14630);
nor UO_1645 (O_1645,N_14080,N_12818);
and UO_1646 (O_1646,N_14431,N_12722);
nor UO_1647 (O_1647,N_13238,N_12774);
and UO_1648 (O_1648,N_13924,N_12048);
nor UO_1649 (O_1649,N_13154,N_12898);
nor UO_1650 (O_1650,N_13732,N_13520);
xor UO_1651 (O_1651,N_13476,N_13279);
nand UO_1652 (O_1652,N_12720,N_12717);
nand UO_1653 (O_1653,N_14037,N_12002);
nor UO_1654 (O_1654,N_12326,N_12933);
nand UO_1655 (O_1655,N_13626,N_14461);
xnor UO_1656 (O_1656,N_12049,N_14616);
nand UO_1657 (O_1657,N_13257,N_12101);
nand UO_1658 (O_1658,N_12001,N_12478);
nand UO_1659 (O_1659,N_13109,N_14363);
and UO_1660 (O_1660,N_12874,N_12194);
or UO_1661 (O_1661,N_13394,N_14895);
and UO_1662 (O_1662,N_13183,N_13360);
and UO_1663 (O_1663,N_14905,N_14130);
nor UO_1664 (O_1664,N_13695,N_14777);
or UO_1665 (O_1665,N_12433,N_13745);
nand UO_1666 (O_1666,N_14916,N_13899);
and UO_1667 (O_1667,N_14047,N_12039);
nor UO_1668 (O_1668,N_13501,N_14573);
nor UO_1669 (O_1669,N_12434,N_13160);
nor UO_1670 (O_1670,N_12369,N_13486);
and UO_1671 (O_1671,N_12116,N_12956);
nor UO_1672 (O_1672,N_14066,N_13987);
and UO_1673 (O_1673,N_13226,N_13779);
or UO_1674 (O_1674,N_13313,N_14012);
nand UO_1675 (O_1675,N_12495,N_14132);
nand UO_1676 (O_1676,N_12979,N_13382);
or UO_1677 (O_1677,N_12528,N_14050);
and UO_1678 (O_1678,N_13991,N_13444);
and UO_1679 (O_1679,N_14653,N_12006);
nand UO_1680 (O_1680,N_12682,N_14586);
nand UO_1681 (O_1681,N_14777,N_13565);
or UO_1682 (O_1682,N_13783,N_14919);
and UO_1683 (O_1683,N_14474,N_13682);
nand UO_1684 (O_1684,N_13659,N_13986);
nor UO_1685 (O_1685,N_12577,N_13688);
nor UO_1686 (O_1686,N_14696,N_12010);
xnor UO_1687 (O_1687,N_14566,N_12232);
nor UO_1688 (O_1688,N_12095,N_13345);
and UO_1689 (O_1689,N_12236,N_12208);
and UO_1690 (O_1690,N_14510,N_13220);
or UO_1691 (O_1691,N_12074,N_12492);
nand UO_1692 (O_1692,N_14933,N_12250);
or UO_1693 (O_1693,N_12790,N_13870);
or UO_1694 (O_1694,N_12794,N_12082);
and UO_1695 (O_1695,N_14794,N_14097);
nor UO_1696 (O_1696,N_13896,N_12229);
or UO_1697 (O_1697,N_14738,N_13809);
xor UO_1698 (O_1698,N_14142,N_12814);
and UO_1699 (O_1699,N_13323,N_14711);
and UO_1700 (O_1700,N_13597,N_14387);
nor UO_1701 (O_1701,N_12315,N_13517);
xor UO_1702 (O_1702,N_12010,N_13057);
nand UO_1703 (O_1703,N_14820,N_14083);
or UO_1704 (O_1704,N_13470,N_13484);
and UO_1705 (O_1705,N_14196,N_14946);
and UO_1706 (O_1706,N_12583,N_13910);
or UO_1707 (O_1707,N_12489,N_14679);
nor UO_1708 (O_1708,N_12454,N_13731);
nand UO_1709 (O_1709,N_14763,N_12998);
or UO_1710 (O_1710,N_14019,N_12159);
or UO_1711 (O_1711,N_13566,N_12199);
nor UO_1712 (O_1712,N_12775,N_14618);
or UO_1713 (O_1713,N_13356,N_12613);
nand UO_1714 (O_1714,N_12932,N_14317);
and UO_1715 (O_1715,N_13865,N_14907);
nor UO_1716 (O_1716,N_13308,N_12443);
or UO_1717 (O_1717,N_13926,N_14845);
and UO_1718 (O_1718,N_14826,N_13433);
and UO_1719 (O_1719,N_12730,N_14836);
nand UO_1720 (O_1720,N_13161,N_13931);
or UO_1721 (O_1721,N_13540,N_13589);
and UO_1722 (O_1722,N_13632,N_12060);
and UO_1723 (O_1723,N_13436,N_13051);
nand UO_1724 (O_1724,N_14175,N_14002);
nor UO_1725 (O_1725,N_12994,N_14560);
nand UO_1726 (O_1726,N_12149,N_14279);
nand UO_1727 (O_1727,N_14104,N_13078);
nand UO_1728 (O_1728,N_13473,N_12428);
nand UO_1729 (O_1729,N_14147,N_14089);
and UO_1730 (O_1730,N_12427,N_13293);
or UO_1731 (O_1731,N_12110,N_14299);
and UO_1732 (O_1732,N_13370,N_13434);
xor UO_1733 (O_1733,N_13333,N_12204);
nor UO_1734 (O_1734,N_13808,N_13983);
xnor UO_1735 (O_1735,N_12803,N_13428);
nand UO_1736 (O_1736,N_12652,N_14458);
nand UO_1737 (O_1737,N_13060,N_14848);
and UO_1738 (O_1738,N_12610,N_13142);
or UO_1739 (O_1739,N_14101,N_13043);
xor UO_1740 (O_1740,N_14920,N_13904);
or UO_1741 (O_1741,N_12292,N_13963);
and UO_1742 (O_1742,N_12129,N_14324);
nor UO_1743 (O_1743,N_12453,N_12412);
or UO_1744 (O_1744,N_12737,N_13458);
xor UO_1745 (O_1745,N_13656,N_13771);
or UO_1746 (O_1746,N_14891,N_14669);
xnor UO_1747 (O_1747,N_13285,N_12481);
and UO_1748 (O_1748,N_12320,N_14083);
nor UO_1749 (O_1749,N_12105,N_14752);
or UO_1750 (O_1750,N_14178,N_12434);
nor UO_1751 (O_1751,N_13323,N_12860);
or UO_1752 (O_1752,N_14599,N_14781);
nand UO_1753 (O_1753,N_12397,N_12521);
xor UO_1754 (O_1754,N_12525,N_12816);
nor UO_1755 (O_1755,N_12932,N_13272);
or UO_1756 (O_1756,N_14913,N_13341);
or UO_1757 (O_1757,N_14797,N_13325);
or UO_1758 (O_1758,N_13819,N_13696);
or UO_1759 (O_1759,N_14859,N_14721);
nor UO_1760 (O_1760,N_14001,N_13217);
nor UO_1761 (O_1761,N_13594,N_14410);
or UO_1762 (O_1762,N_14295,N_13774);
xnor UO_1763 (O_1763,N_13792,N_14562);
nand UO_1764 (O_1764,N_14102,N_12919);
or UO_1765 (O_1765,N_13642,N_14844);
nand UO_1766 (O_1766,N_14146,N_13745);
or UO_1767 (O_1767,N_12827,N_14309);
and UO_1768 (O_1768,N_13039,N_12373);
nand UO_1769 (O_1769,N_12314,N_14317);
xor UO_1770 (O_1770,N_12320,N_14039);
or UO_1771 (O_1771,N_14408,N_14863);
and UO_1772 (O_1772,N_14513,N_13994);
nor UO_1773 (O_1773,N_12065,N_14653);
nand UO_1774 (O_1774,N_14979,N_12683);
nor UO_1775 (O_1775,N_13729,N_12190);
nor UO_1776 (O_1776,N_14550,N_13542);
or UO_1777 (O_1777,N_12632,N_12414);
nand UO_1778 (O_1778,N_12502,N_14395);
and UO_1779 (O_1779,N_14864,N_12999);
xor UO_1780 (O_1780,N_13927,N_14730);
or UO_1781 (O_1781,N_14543,N_14469);
and UO_1782 (O_1782,N_12956,N_14436);
nand UO_1783 (O_1783,N_12215,N_13313);
nor UO_1784 (O_1784,N_13014,N_12299);
or UO_1785 (O_1785,N_14219,N_13308);
or UO_1786 (O_1786,N_13911,N_13423);
and UO_1787 (O_1787,N_12058,N_14011);
xnor UO_1788 (O_1788,N_13339,N_13273);
or UO_1789 (O_1789,N_14348,N_14496);
nand UO_1790 (O_1790,N_12867,N_14062);
nand UO_1791 (O_1791,N_12435,N_14147);
or UO_1792 (O_1792,N_14168,N_13934);
or UO_1793 (O_1793,N_14704,N_12735);
xnor UO_1794 (O_1794,N_14209,N_14505);
and UO_1795 (O_1795,N_14493,N_12723);
and UO_1796 (O_1796,N_14748,N_13830);
nand UO_1797 (O_1797,N_12333,N_14439);
or UO_1798 (O_1798,N_13089,N_13088);
and UO_1799 (O_1799,N_13906,N_14643);
or UO_1800 (O_1800,N_12515,N_13893);
nor UO_1801 (O_1801,N_13314,N_14479);
xor UO_1802 (O_1802,N_13015,N_12109);
nand UO_1803 (O_1803,N_13956,N_13984);
and UO_1804 (O_1804,N_12889,N_13342);
xnor UO_1805 (O_1805,N_13784,N_13740);
xor UO_1806 (O_1806,N_13923,N_14182);
nor UO_1807 (O_1807,N_13234,N_14356);
and UO_1808 (O_1808,N_13143,N_14272);
and UO_1809 (O_1809,N_14677,N_12222);
and UO_1810 (O_1810,N_12100,N_13109);
nor UO_1811 (O_1811,N_13530,N_14042);
nor UO_1812 (O_1812,N_14504,N_14697);
or UO_1813 (O_1813,N_14498,N_13641);
and UO_1814 (O_1814,N_12760,N_13738);
and UO_1815 (O_1815,N_13322,N_12664);
nand UO_1816 (O_1816,N_12699,N_13725);
or UO_1817 (O_1817,N_14741,N_12489);
nand UO_1818 (O_1818,N_14823,N_14969);
nor UO_1819 (O_1819,N_14520,N_13899);
or UO_1820 (O_1820,N_12211,N_14259);
xor UO_1821 (O_1821,N_12710,N_14402);
nand UO_1822 (O_1822,N_14835,N_12107);
nor UO_1823 (O_1823,N_12543,N_14834);
nor UO_1824 (O_1824,N_12122,N_13095);
nand UO_1825 (O_1825,N_14474,N_12392);
nor UO_1826 (O_1826,N_12246,N_12269);
and UO_1827 (O_1827,N_12400,N_14411);
nor UO_1828 (O_1828,N_13067,N_13602);
nand UO_1829 (O_1829,N_13229,N_14718);
and UO_1830 (O_1830,N_14295,N_13892);
nand UO_1831 (O_1831,N_14689,N_13185);
nor UO_1832 (O_1832,N_12781,N_14166);
nor UO_1833 (O_1833,N_12473,N_12086);
nand UO_1834 (O_1834,N_12810,N_13209);
or UO_1835 (O_1835,N_14792,N_14804);
nor UO_1836 (O_1836,N_14800,N_12232);
and UO_1837 (O_1837,N_13659,N_12869);
and UO_1838 (O_1838,N_14858,N_13721);
and UO_1839 (O_1839,N_14792,N_12666);
nand UO_1840 (O_1840,N_12687,N_12263);
and UO_1841 (O_1841,N_12248,N_14141);
nor UO_1842 (O_1842,N_14393,N_14746);
or UO_1843 (O_1843,N_14854,N_13292);
nand UO_1844 (O_1844,N_13045,N_12541);
xor UO_1845 (O_1845,N_14596,N_13235);
or UO_1846 (O_1846,N_14086,N_12243);
nand UO_1847 (O_1847,N_12113,N_14232);
xor UO_1848 (O_1848,N_14653,N_13006);
nand UO_1849 (O_1849,N_14218,N_14398);
nand UO_1850 (O_1850,N_14010,N_12510);
nor UO_1851 (O_1851,N_13103,N_14374);
or UO_1852 (O_1852,N_14533,N_13193);
nor UO_1853 (O_1853,N_14588,N_12155);
or UO_1854 (O_1854,N_13092,N_14397);
nor UO_1855 (O_1855,N_14744,N_13692);
or UO_1856 (O_1856,N_14293,N_14026);
or UO_1857 (O_1857,N_12088,N_13593);
nor UO_1858 (O_1858,N_13475,N_14403);
nand UO_1859 (O_1859,N_14396,N_14010);
nor UO_1860 (O_1860,N_12928,N_13110);
xor UO_1861 (O_1861,N_14428,N_14155);
nand UO_1862 (O_1862,N_14207,N_12935);
nand UO_1863 (O_1863,N_12750,N_14560);
or UO_1864 (O_1864,N_12562,N_13489);
or UO_1865 (O_1865,N_13825,N_14158);
nand UO_1866 (O_1866,N_14930,N_13418);
nor UO_1867 (O_1867,N_12719,N_14247);
nor UO_1868 (O_1868,N_13486,N_12371);
nand UO_1869 (O_1869,N_12047,N_12612);
nor UO_1870 (O_1870,N_12045,N_13344);
and UO_1871 (O_1871,N_14181,N_13625);
nor UO_1872 (O_1872,N_13080,N_12497);
nor UO_1873 (O_1873,N_14722,N_12276);
and UO_1874 (O_1874,N_14790,N_14455);
and UO_1875 (O_1875,N_12446,N_12662);
or UO_1876 (O_1876,N_13533,N_14779);
nand UO_1877 (O_1877,N_13839,N_14698);
nand UO_1878 (O_1878,N_12629,N_12226);
nor UO_1879 (O_1879,N_13973,N_13203);
or UO_1880 (O_1880,N_12157,N_12040);
nor UO_1881 (O_1881,N_13644,N_13449);
or UO_1882 (O_1882,N_13449,N_14456);
nand UO_1883 (O_1883,N_13669,N_13904);
and UO_1884 (O_1884,N_12167,N_12995);
nor UO_1885 (O_1885,N_12585,N_12458);
xnor UO_1886 (O_1886,N_12263,N_13122);
or UO_1887 (O_1887,N_12385,N_14613);
and UO_1888 (O_1888,N_14525,N_13265);
and UO_1889 (O_1889,N_12999,N_12644);
or UO_1890 (O_1890,N_13901,N_13497);
or UO_1891 (O_1891,N_14120,N_13191);
nand UO_1892 (O_1892,N_12795,N_12577);
and UO_1893 (O_1893,N_14255,N_13022);
or UO_1894 (O_1894,N_12972,N_13492);
nor UO_1895 (O_1895,N_13648,N_13169);
nand UO_1896 (O_1896,N_13780,N_12612);
nor UO_1897 (O_1897,N_14299,N_13053);
and UO_1898 (O_1898,N_13675,N_14683);
or UO_1899 (O_1899,N_14935,N_12768);
and UO_1900 (O_1900,N_12377,N_13304);
or UO_1901 (O_1901,N_14339,N_14913);
nor UO_1902 (O_1902,N_12089,N_14195);
nor UO_1903 (O_1903,N_12034,N_12266);
or UO_1904 (O_1904,N_13196,N_13915);
and UO_1905 (O_1905,N_14574,N_13636);
nand UO_1906 (O_1906,N_13875,N_14773);
and UO_1907 (O_1907,N_12852,N_14555);
nand UO_1908 (O_1908,N_13383,N_12838);
nand UO_1909 (O_1909,N_13957,N_12167);
or UO_1910 (O_1910,N_13510,N_13689);
nor UO_1911 (O_1911,N_14438,N_14720);
and UO_1912 (O_1912,N_13318,N_12754);
xnor UO_1913 (O_1913,N_14880,N_12056);
or UO_1914 (O_1914,N_13237,N_13749);
or UO_1915 (O_1915,N_13394,N_12047);
nand UO_1916 (O_1916,N_13448,N_13060);
nor UO_1917 (O_1917,N_14529,N_12563);
nand UO_1918 (O_1918,N_13317,N_12424);
nor UO_1919 (O_1919,N_12384,N_12289);
and UO_1920 (O_1920,N_12956,N_13322);
xor UO_1921 (O_1921,N_14274,N_12828);
or UO_1922 (O_1922,N_14348,N_12119);
nand UO_1923 (O_1923,N_14675,N_12380);
or UO_1924 (O_1924,N_12045,N_12259);
nand UO_1925 (O_1925,N_13679,N_12083);
nand UO_1926 (O_1926,N_13454,N_14950);
nand UO_1927 (O_1927,N_13565,N_12522);
and UO_1928 (O_1928,N_12207,N_14491);
nand UO_1929 (O_1929,N_13244,N_13879);
nand UO_1930 (O_1930,N_12904,N_13003);
and UO_1931 (O_1931,N_14973,N_13102);
nand UO_1932 (O_1932,N_14824,N_14426);
xor UO_1933 (O_1933,N_13919,N_13217);
and UO_1934 (O_1934,N_12132,N_12908);
xnor UO_1935 (O_1935,N_13963,N_12067);
nor UO_1936 (O_1936,N_14383,N_14670);
and UO_1937 (O_1937,N_12974,N_12104);
and UO_1938 (O_1938,N_12385,N_13435);
nand UO_1939 (O_1939,N_14486,N_13775);
nand UO_1940 (O_1940,N_14021,N_14540);
xnor UO_1941 (O_1941,N_14148,N_14913);
nand UO_1942 (O_1942,N_14098,N_12931);
nand UO_1943 (O_1943,N_12523,N_12988);
xor UO_1944 (O_1944,N_12140,N_14612);
or UO_1945 (O_1945,N_12681,N_12927);
nand UO_1946 (O_1946,N_12642,N_13838);
and UO_1947 (O_1947,N_14914,N_13056);
or UO_1948 (O_1948,N_13095,N_13667);
and UO_1949 (O_1949,N_14396,N_14469);
xor UO_1950 (O_1950,N_14740,N_13985);
and UO_1951 (O_1951,N_12731,N_13727);
nor UO_1952 (O_1952,N_12512,N_12338);
or UO_1953 (O_1953,N_12961,N_13061);
nor UO_1954 (O_1954,N_13416,N_12871);
nor UO_1955 (O_1955,N_12162,N_14854);
nand UO_1956 (O_1956,N_13682,N_14348);
nor UO_1957 (O_1957,N_13526,N_13843);
xnor UO_1958 (O_1958,N_13442,N_12330);
or UO_1959 (O_1959,N_12921,N_12014);
or UO_1960 (O_1960,N_14850,N_14534);
nor UO_1961 (O_1961,N_14334,N_13606);
or UO_1962 (O_1962,N_13598,N_12497);
nor UO_1963 (O_1963,N_13131,N_12466);
nand UO_1964 (O_1964,N_12671,N_14681);
and UO_1965 (O_1965,N_14955,N_12632);
nand UO_1966 (O_1966,N_13750,N_12735);
and UO_1967 (O_1967,N_14398,N_12443);
and UO_1968 (O_1968,N_14394,N_12779);
nand UO_1969 (O_1969,N_12095,N_14651);
nand UO_1970 (O_1970,N_13830,N_12339);
nor UO_1971 (O_1971,N_14794,N_13060);
or UO_1972 (O_1972,N_13400,N_12409);
or UO_1973 (O_1973,N_14741,N_12938);
and UO_1974 (O_1974,N_14956,N_12987);
xnor UO_1975 (O_1975,N_12354,N_13515);
nand UO_1976 (O_1976,N_12090,N_14112);
and UO_1977 (O_1977,N_12375,N_12433);
and UO_1978 (O_1978,N_12656,N_14813);
nor UO_1979 (O_1979,N_13430,N_13898);
and UO_1980 (O_1980,N_14158,N_14798);
xnor UO_1981 (O_1981,N_12797,N_13065);
nand UO_1982 (O_1982,N_13751,N_14796);
xor UO_1983 (O_1983,N_13669,N_14212);
or UO_1984 (O_1984,N_14641,N_14006);
or UO_1985 (O_1985,N_13105,N_14525);
nand UO_1986 (O_1986,N_13608,N_13737);
nand UO_1987 (O_1987,N_12807,N_13451);
and UO_1988 (O_1988,N_14016,N_14687);
nand UO_1989 (O_1989,N_14967,N_12467);
and UO_1990 (O_1990,N_13069,N_14149);
or UO_1991 (O_1991,N_14220,N_12107);
or UO_1992 (O_1992,N_13720,N_12663);
nand UO_1993 (O_1993,N_13515,N_13245);
nor UO_1994 (O_1994,N_12767,N_13955);
and UO_1995 (O_1995,N_13741,N_13300);
or UO_1996 (O_1996,N_14383,N_14834);
xor UO_1997 (O_1997,N_12167,N_12328);
or UO_1998 (O_1998,N_14779,N_12954);
nor UO_1999 (O_1999,N_12144,N_13693);
endmodule