module basic_2000_20000_2500_125_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_1120,In_1047);
nand U1 (N_1,In_713,In_710);
nand U2 (N_2,In_783,In_52);
or U3 (N_3,In_458,In_1259);
and U4 (N_4,In_363,In_514);
nor U5 (N_5,In_688,In_1082);
and U6 (N_6,In_167,In_601);
or U7 (N_7,In_271,In_631);
and U8 (N_8,In_324,In_101);
or U9 (N_9,In_1789,In_1270);
and U10 (N_10,In_1786,In_1191);
nor U11 (N_11,In_1842,In_1134);
and U12 (N_12,In_1282,In_655);
nor U13 (N_13,In_574,In_104);
nand U14 (N_14,In_608,In_250);
and U15 (N_15,In_782,In_1336);
and U16 (N_16,In_1998,In_1476);
and U17 (N_17,In_1822,In_1480);
or U18 (N_18,In_1856,In_743);
nor U19 (N_19,In_1668,In_808);
nor U20 (N_20,In_1598,In_1483);
or U21 (N_21,In_235,In_1807);
and U22 (N_22,In_515,In_1803);
nand U23 (N_23,In_448,In_1562);
and U24 (N_24,In_1910,In_1007);
nor U25 (N_25,In_572,In_1566);
and U26 (N_26,In_1564,In_284);
or U27 (N_27,In_1897,In_1982);
nor U28 (N_28,In_1690,In_1416);
nand U29 (N_29,In_1429,In_960);
or U30 (N_30,In_412,In_182);
or U31 (N_31,In_266,In_357);
and U32 (N_32,In_1023,In_168);
nand U33 (N_33,In_599,In_1139);
and U34 (N_34,In_302,In_980);
or U35 (N_35,In_1077,In_1622);
or U36 (N_36,In_468,In_800);
nand U37 (N_37,In_520,In_628);
nor U38 (N_38,In_1300,In_81);
and U39 (N_39,In_280,In_1906);
nand U40 (N_40,In_1316,In_179);
and U41 (N_41,In_508,In_613);
nand U42 (N_42,In_804,In_197);
or U43 (N_43,In_1965,In_680);
nand U44 (N_44,In_140,In_17);
or U45 (N_45,In_13,In_647);
nand U46 (N_46,In_1670,In_1872);
or U47 (N_47,In_1745,In_227);
nor U48 (N_48,In_1680,In_1440);
and U49 (N_49,In_75,In_569);
xor U50 (N_50,In_47,In_927);
or U51 (N_51,In_1891,In_1923);
and U52 (N_52,In_1102,In_625);
nor U53 (N_53,In_546,In_703);
and U54 (N_54,In_822,In_772);
or U55 (N_55,In_1278,In_1359);
or U56 (N_56,In_805,In_1129);
or U57 (N_57,In_1984,In_1116);
xnor U58 (N_58,In_1163,In_1431);
or U59 (N_59,In_764,In_1550);
xnor U60 (N_60,In_941,In_274);
nor U61 (N_61,In_954,In_1708);
nand U62 (N_62,In_1747,In_126);
and U63 (N_63,In_585,In_1530);
and U64 (N_64,In_693,In_490);
nor U65 (N_65,In_1579,In_1949);
nor U66 (N_66,In_1744,In_1655);
nand U67 (N_67,In_650,In_187);
xnor U68 (N_68,In_206,In_1921);
nor U69 (N_69,In_802,In_157);
or U70 (N_70,In_1713,In_603);
and U71 (N_71,In_1337,In_953);
nand U72 (N_72,In_474,In_826);
xnor U73 (N_73,In_1712,In_1348);
and U74 (N_74,In_312,In_1432);
or U75 (N_75,In_1084,In_937);
nand U76 (N_76,In_1449,In_1578);
or U77 (N_77,In_1861,In_753);
xnor U78 (N_78,In_1090,In_1526);
and U79 (N_79,In_1168,In_1013);
nand U80 (N_80,In_624,In_1516);
or U81 (N_81,In_742,In_1182);
nor U82 (N_82,In_1065,In_1800);
nor U83 (N_83,In_355,In_96);
nand U84 (N_84,In_642,In_811);
nand U85 (N_85,In_656,In_1295);
nor U86 (N_86,In_690,In_759);
nor U87 (N_87,In_495,In_1224);
xor U88 (N_88,In_1356,In_63);
nor U89 (N_89,In_1746,In_1044);
nor U90 (N_90,In_887,In_1421);
nor U91 (N_91,In_194,In_921);
and U92 (N_92,In_649,In_1063);
or U93 (N_93,In_697,In_1244);
nand U94 (N_94,In_1836,In_241);
xor U95 (N_95,In_165,In_90);
and U96 (N_96,In_1208,In_427);
xor U97 (N_97,In_4,In_1128);
nor U98 (N_98,In_294,In_113);
or U99 (N_99,In_463,In_1318);
and U100 (N_100,In_1251,In_1413);
nor U101 (N_101,In_1003,In_820);
and U102 (N_102,In_265,In_1952);
or U103 (N_103,In_369,In_1688);
nand U104 (N_104,In_409,In_640);
nand U105 (N_105,In_1238,In_635);
and U106 (N_106,In_1651,In_367);
xor U107 (N_107,In_1617,In_1496);
nand U108 (N_108,In_1927,In_1205);
and U109 (N_109,In_602,In_849);
xor U110 (N_110,In_1437,In_911);
and U111 (N_111,In_23,In_240);
and U112 (N_112,In_1404,In_1078);
nand U113 (N_113,In_659,In_424);
or U114 (N_114,In_721,In_29);
xor U115 (N_115,In_460,In_799);
nand U116 (N_116,In_794,In_14);
and U117 (N_117,In_1430,In_79);
nor U118 (N_118,In_866,In_193);
nor U119 (N_119,In_48,In_1702);
or U120 (N_120,In_1506,In_261);
nand U121 (N_121,In_1871,In_916);
nand U122 (N_122,In_214,In_696);
or U123 (N_123,In_377,In_1743);
and U124 (N_124,In_1727,In_1791);
nand U125 (N_125,In_1170,In_667);
nand U126 (N_126,In_1587,In_1066);
and U127 (N_127,In_1361,In_1847);
or U128 (N_128,In_1592,In_1602);
or U129 (N_129,In_1903,In_1121);
nor U130 (N_130,In_1130,In_1024);
nor U131 (N_131,In_122,In_947);
xnor U132 (N_132,In_1968,In_1286);
and U133 (N_133,In_910,In_762);
and U134 (N_134,In_205,In_19);
or U135 (N_135,In_526,In_1737);
and U136 (N_136,In_718,In_56);
and U137 (N_137,In_971,In_1197);
and U138 (N_138,In_1615,In_778);
nand U139 (N_139,In_408,In_1468);
or U140 (N_140,In_1477,In_1079);
nand U141 (N_141,In_1291,In_1771);
and U142 (N_142,In_1225,In_1433);
xor U143 (N_143,In_547,In_1329);
or U144 (N_144,In_1796,In_597);
nand U145 (N_145,In_1060,In_469);
and U146 (N_146,In_1375,In_269);
and U147 (N_147,In_1654,In_1398);
or U148 (N_148,In_1867,In_488);
nand U149 (N_149,In_1072,In_1344);
and U150 (N_150,In_429,In_1338);
nor U151 (N_151,In_1962,In_1809);
and U152 (N_152,In_632,In_1806);
or U153 (N_153,In_1376,In_1132);
nor U154 (N_154,In_1230,In_1346);
or U155 (N_155,In_1724,In_1040);
and U156 (N_156,In_1798,In_1308);
or U157 (N_157,In_834,In_231);
and U158 (N_158,In_852,In_593);
nand U159 (N_159,In_1080,In_1536);
or U160 (N_160,In_562,In_1817);
or U161 (N_161,In_254,In_108);
nand U162 (N_162,In_1029,In_687);
and U163 (N_163,In_273,In_67);
nor U164 (N_164,In_1025,In_464);
or U165 (N_165,In_1967,In_657);
xnor U166 (N_166,In_1557,In_1884);
nor U167 (N_167,In_1600,In_1932);
nand U168 (N_168,In_1272,In_335);
and U169 (N_169,In_1686,In_532);
nor U170 (N_170,In_1778,In_1151);
nor U171 (N_171,N_7,In_55);
and U172 (N_172,In_1456,In_1123);
or U173 (N_173,In_1647,In_1198);
nand U174 (N_174,In_1497,In_986);
and U175 (N_175,In_391,In_1720);
and U176 (N_176,In_174,In_739);
nor U177 (N_177,N_151,In_117);
and U178 (N_178,N_153,In_612);
or U179 (N_179,In_1083,In_341);
and U180 (N_180,In_1511,In_901);
nand U181 (N_181,In_1262,In_1387);
or U182 (N_182,In_924,In_1898);
nand U183 (N_183,In_1870,In_1169);
nand U184 (N_184,In_933,In_506);
nor U185 (N_185,In_1975,In_15);
and U186 (N_186,In_1500,In_296);
xor U187 (N_187,In_923,N_14);
nand U188 (N_188,In_524,In_1273);
and U189 (N_189,In_342,N_102);
and U190 (N_190,In_1760,In_1000);
nand U191 (N_191,In_112,In_1508);
nor U192 (N_192,In_471,In_816);
nand U193 (N_193,In_1632,In_1604);
xor U194 (N_194,In_955,In_1901);
nand U195 (N_195,In_1877,In_390);
nor U196 (N_196,In_1717,In_1912);
and U197 (N_197,In_1672,In_404);
nor U198 (N_198,In_664,In_548);
or U199 (N_199,N_159,In_1790);
nand U200 (N_200,In_1284,In_479);
nand U201 (N_201,In_1220,In_1926);
nor U202 (N_202,In_172,In_967);
or U203 (N_203,In_677,N_88);
nor U204 (N_204,In_1546,In_51);
or U205 (N_205,In_617,In_1452);
or U206 (N_206,In_1667,In_1695);
nor U207 (N_207,In_1241,In_727);
and U208 (N_208,In_1076,In_436);
nor U209 (N_209,In_1565,In_930);
and U210 (N_210,In_376,In_248);
and U211 (N_211,In_1849,In_1641);
and U212 (N_212,In_1840,In_1075);
and U213 (N_213,In_507,In_1533);
nand U214 (N_214,In_598,In_1769);
nand U215 (N_215,In_24,In_1919);
nand U216 (N_216,In_119,In_496);
nor U217 (N_217,In_1528,N_100);
nor U218 (N_218,In_1772,In_1219);
or U219 (N_219,In_860,N_150);
nand U220 (N_220,N_62,In_929);
and U221 (N_221,In_1648,In_1109);
and U222 (N_222,In_553,In_1733);
and U223 (N_223,In_1249,In_1481);
or U224 (N_224,In_824,N_20);
nor U225 (N_225,In_252,In_1178);
and U226 (N_226,In_843,In_146);
nor U227 (N_227,In_605,In_592);
xnor U228 (N_228,In_210,In_333);
xor U229 (N_229,In_1135,In_1726);
and U230 (N_230,In_1126,In_792);
or U231 (N_231,In_1319,In_567);
nor U232 (N_232,In_1418,In_225);
and U233 (N_233,N_65,In_447);
nor U234 (N_234,In_1218,In_419);
or U235 (N_235,In_1486,In_455);
xnor U236 (N_236,In_1734,N_87);
nand U237 (N_237,In_7,In_827);
nor U238 (N_238,In_1005,In_1749);
and U239 (N_239,In_279,In_503);
nand U240 (N_240,In_1261,In_1174);
xnor U241 (N_241,In_780,In_249);
nand U242 (N_242,In_1770,In_1731);
or U243 (N_243,In_375,In_1704);
and U244 (N_244,In_360,In_576);
and U245 (N_245,In_1401,In_847);
or U246 (N_246,In_1787,In_1860);
or U247 (N_247,In_170,In_606);
and U248 (N_248,In_1845,In_1188);
nand U249 (N_249,In_1523,In_999);
and U250 (N_250,In_1606,In_706);
nor U251 (N_251,N_93,N_26);
nand U252 (N_252,In_666,In_899);
and U253 (N_253,In_556,In_1900);
nor U254 (N_254,In_93,In_1204);
xor U255 (N_255,In_183,In_1988);
nand U256 (N_256,In_141,In_1775);
or U257 (N_257,In_1200,In_856);
or U258 (N_258,N_130,In_1797);
nand U259 (N_259,In_1634,In_1002);
nand U260 (N_260,In_1436,In_178);
nand U261 (N_261,In_350,In_1818);
nand U262 (N_262,In_1888,In_1118);
nand U263 (N_263,In_1794,In_1718);
nor U264 (N_264,In_1246,In_539);
and U265 (N_265,In_337,In_623);
nand U266 (N_266,In_256,In_171);
nor U267 (N_267,In_581,N_10);
and U268 (N_268,In_1274,In_39);
nand U269 (N_269,In_582,In_1265);
nor U270 (N_270,In_867,In_1660);
or U271 (N_271,In_773,In_59);
nand U272 (N_272,N_67,In_566);
and U273 (N_273,In_268,In_906);
nor U274 (N_274,N_3,In_1458);
nor U275 (N_275,In_1347,In_467);
nand U276 (N_276,In_1446,In_1751);
or U277 (N_277,In_485,In_651);
nor U278 (N_278,In_327,In_1100);
and U279 (N_279,In_1367,In_1330);
and U280 (N_280,In_1049,In_968);
nor U281 (N_281,In_217,In_873);
and U282 (N_282,In_1682,N_95);
and U283 (N_283,In_1756,In_1392);
or U284 (N_284,In_30,In_70);
or U285 (N_285,In_1505,In_301);
nor U286 (N_286,In_1362,In_320);
or U287 (N_287,In_482,In_1231);
nor U288 (N_288,In_1678,In_1419);
nor U289 (N_289,In_465,In_133);
and U290 (N_290,N_117,In_1661);
xnor U291 (N_291,In_946,In_1133);
or U292 (N_292,In_875,In_116);
xor U293 (N_293,N_82,In_1824);
nor U294 (N_294,In_1352,In_798);
xor U295 (N_295,In_1091,In_293);
nor U296 (N_296,N_37,In_1184);
or U297 (N_297,In_64,In_821);
nand U298 (N_298,In_671,In_673);
or U299 (N_299,In_1097,N_154);
or U300 (N_300,In_1883,In_1402);
nor U301 (N_301,In_1827,In_646);
nand U302 (N_302,N_68,In_1166);
nand U303 (N_303,In_136,In_43);
nor U304 (N_304,In_151,In_1391);
or U305 (N_305,In_1012,In_1997);
nor U306 (N_306,In_202,In_1753);
nand U307 (N_307,In_578,In_521);
nor U308 (N_308,In_1209,In_1567);
and U309 (N_309,In_300,In_311);
or U310 (N_310,In_452,In_1382);
and U311 (N_311,In_1940,In_1465);
or U312 (N_312,In_344,In_394);
nor U313 (N_313,N_80,In_216);
nand U314 (N_314,In_855,In_444);
nand U315 (N_315,In_1896,In_1774);
nor U316 (N_316,In_470,N_28);
nor U317 (N_317,In_988,In_1955);
nand U318 (N_318,In_1045,In_379);
nand U319 (N_319,In_186,In_1907);
and U320 (N_320,In_1757,In_789);
nand U321 (N_321,In_786,In_1008);
or U322 (N_322,N_244,In_939);
and U323 (N_323,In_694,In_1974);
and U324 (N_324,In_8,In_758);
or U325 (N_325,In_406,N_44);
xnor U326 (N_326,N_301,In_561);
nand U327 (N_327,In_644,In_1524);
nand U328 (N_328,In_1715,In_1155);
xor U329 (N_329,In_619,In_1294);
xor U330 (N_330,N_173,In_152);
xor U331 (N_331,In_1043,In_1485);
nor U332 (N_332,In_627,N_282);
and U333 (N_333,In_1474,In_1313);
and U334 (N_334,In_1138,In_1519);
nand U335 (N_335,N_203,In_332);
and U336 (N_336,In_1351,In_1038);
nor U337 (N_337,In_148,In_83);
nand U338 (N_338,In_1152,In_1607);
nand U339 (N_339,In_258,In_297);
nand U340 (N_340,In_1321,N_241);
and U341 (N_341,In_803,In_20);
and U342 (N_342,N_313,N_156);
and U343 (N_343,In_1180,In_1073);
and U344 (N_344,In_1088,In_373);
xnor U345 (N_345,In_903,In_752);
nor U346 (N_346,In_1944,In_1470);
xor U347 (N_347,In_159,In_1773);
nand U348 (N_348,In_1498,In_1089);
and U349 (N_349,N_164,In_557);
xor U350 (N_350,In_881,In_995);
and U351 (N_351,In_283,In_232);
nor U352 (N_352,In_662,In_641);
or U353 (N_353,In_37,In_9);
nor U354 (N_354,In_1762,In_1288);
nand U355 (N_355,In_563,In_1507);
nand U356 (N_356,In_353,In_568);
nor U357 (N_357,N_219,In_1761);
xor U358 (N_358,In_1192,N_220);
nand U359 (N_359,N_228,In_421);
nand U360 (N_360,In_1640,In_1140);
or U361 (N_361,In_319,In_1014);
xnor U362 (N_362,In_1366,N_92);
nand U363 (N_363,In_1671,In_1142);
nand U364 (N_364,In_872,In_1071);
or U365 (N_365,In_1343,In_487);
and U366 (N_366,In_472,In_1374);
nor U367 (N_367,In_1495,N_312);
nand U368 (N_368,In_904,In_1941);
xnor U369 (N_369,In_990,In_1586);
nand U370 (N_370,In_111,N_299);
and U371 (N_371,In_98,In_1591);
xnor U372 (N_372,N_231,In_1669);
xnor U373 (N_373,In_352,In_768);
nor U374 (N_374,In_1342,In_203);
nor U375 (N_375,N_305,In_1426);
or U376 (N_376,In_1810,N_42);
nor U377 (N_377,In_1582,In_1539);
or U378 (N_378,In_1934,In_538);
nor U379 (N_379,In_1070,In_981);
or U380 (N_380,In_11,N_201);
and U381 (N_381,In_1144,In_103);
nor U382 (N_382,In_1970,N_174);
or U383 (N_383,In_207,N_43);
or U384 (N_384,In_1823,In_1450);
nor U385 (N_385,In_1268,In_1656);
nand U386 (N_386,In_1657,In_1160);
nand U387 (N_387,In_695,N_73);
or U388 (N_388,In_339,In_1302);
nand U389 (N_389,In_813,N_225);
nor U390 (N_390,In_1491,In_1176);
and U391 (N_391,In_10,In_1074);
or U392 (N_392,In_185,In_1222);
nand U393 (N_393,In_1397,In_1518);
and U394 (N_394,In_22,In_1534);
nor U395 (N_395,In_1895,In_1909);
xnor U396 (N_396,In_491,N_303);
and U397 (N_397,N_248,In_728);
nand U398 (N_398,In_16,In_907);
nand U399 (N_399,N_57,N_84);
nor U400 (N_400,N_237,In_173);
or U401 (N_401,N_193,In_1217);
and U402 (N_402,In_1569,In_1150);
nand U403 (N_403,In_305,In_505);
nor U404 (N_404,N_36,In_1257);
nor U405 (N_405,In_1995,In_1517);
nand U406 (N_406,In_876,In_87);
xor U407 (N_407,In_1004,In_443);
nand U408 (N_408,In_1435,In_1514);
nand U409 (N_409,In_964,In_1978);
nand U410 (N_410,In_1529,In_2);
and U411 (N_411,In_1645,In_82);
nor U412 (N_412,N_278,In_1692);
nand U413 (N_413,In_1113,In_1363);
and U414 (N_414,N_176,In_1938);
nor U415 (N_415,In_1414,In_1561);
or U416 (N_416,In_142,In_295);
or U417 (N_417,N_83,N_192);
and U418 (N_418,In_434,In_1190);
xnor U419 (N_419,In_949,N_169);
nand U420 (N_420,In_1427,In_229);
or U421 (N_421,N_317,In_1512);
and U422 (N_422,N_49,In_215);
xnor U423 (N_423,In_155,In_895);
xor U424 (N_424,N_50,In_607);
and U425 (N_425,N_27,N_60);
nor U426 (N_426,In_1396,In_838);
and U427 (N_427,In_21,In_413);
and U428 (N_428,In_1612,In_1301);
or U429 (N_429,In_750,N_120);
or U430 (N_430,In_457,In_264);
nor U431 (N_431,N_267,In_1948);
or U432 (N_432,In_189,In_1032);
and U433 (N_433,In_698,N_75);
or U434 (N_434,In_779,In_1741);
nor U435 (N_435,In_1981,In_801);
xnor U436 (N_436,In_945,In_1153);
and U437 (N_437,N_128,In_1494);
and U438 (N_438,In_1081,In_480);
and U439 (N_439,In_1930,In_430);
and U440 (N_440,In_615,In_1228);
nor U441 (N_441,In_660,N_257);
nand U442 (N_442,In_1985,N_223);
or U443 (N_443,In_164,In_658);
or U444 (N_444,In_983,In_970);
or U445 (N_445,In_670,In_110);
or U446 (N_446,In_1104,N_103);
nand U447 (N_447,In_1444,N_233);
xnor U448 (N_448,N_246,N_284);
or U449 (N_449,In_1463,In_1623);
or U450 (N_450,In_877,In_288);
nand U451 (N_451,In_993,In_1575);
nor U452 (N_452,N_209,In_1580);
or U453 (N_453,In_1122,In_145);
nor U454 (N_454,In_359,In_1694);
and U455 (N_455,In_338,In_1969);
or U456 (N_456,In_131,In_898);
and U457 (N_457,In_1913,In_255);
nand U458 (N_458,In_522,N_6);
nand U459 (N_459,In_323,In_34);
nand U460 (N_460,In_1855,In_1864);
and U461 (N_461,In_1146,In_144);
or U462 (N_462,In_423,In_915);
nand U463 (N_463,In_1851,In_65);
xor U464 (N_464,In_77,In_50);
and U465 (N_465,In_1766,In_497);
or U466 (N_466,N_72,In_291);
nand U467 (N_467,In_912,In_513);
nor U468 (N_468,In_1739,In_40);
and U469 (N_469,In_1475,In_1624);
nand U470 (N_470,In_237,In_1687);
nand U471 (N_471,In_1701,In_1087);
nand U472 (N_472,N_19,In_869);
and U473 (N_473,In_1242,N_175);
and U474 (N_474,In_358,In_411);
or U475 (N_475,N_90,In_1572);
and U476 (N_476,N_242,N_183);
or U477 (N_477,In_416,N_285);
nor U478 (N_478,N_22,N_136);
nand U479 (N_479,In_1571,In_1441);
or U480 (N_480,In_857,In_334);
nor U481 (N_481,In_1054,N_440);
nor U482 (N_482,N_152,In_1924);
nand U483 (N_483,In_1544,In_1537);
nor U484 (N_484,In_889,N_369);
nor U485 (N_485,In_707,In_1714);
or U486 (N_486,N_212,N_371);
or U487 (N_487,In_201,In_1061);
and U488 (N_488,N_185,In_478);
nor U489 (N_489,In_198,In_1738);
nand U490 (N_490,In_719,In_1350);
nand U491 (N_491,In_1173,In_150);
and U492 (N_492,In_236,N_265);
nand U493 (N_493,In_1894,In_1503);
and U494 (N_494,N_406,In_639);
nor U495 (N_495,In_1185,N_295);
and U496 (N_496,N_411,In_1143);
and U497 (N_497,In_163,N_146);
or U498 (N_498,In_1554,N_113);
and U499 (N_499,In_1328,In_853);
and U500 (N_500,In_1015,In_1911);
nand U501 (N_501,In_591,In_1716);
or U502 (N_502,In_962,In_124);
or U503 (N_503,In_386,In_1748);
and U504 (N_504,N_9,In_1357);
and U505 (N_505,In_1247,In_161);
nor U506 (N_506,N_455,In_1335);
nor U507 (N_507,In_61,In_1289);
and U508 (N_508,In_1112,N_172);
and U509 (N_509,In_129,N_394);
xor U510 (N_510,In_1211,In_1740);
and U511 (N_511,In_1378,In_1161);
nor U512 (N_512,N_443,In_95);
and U513 (N_513,In_1684,In_1039);
nor U514 (N_514,In_1725,In_351);
or U515 (N_515,In_689,In_60);
nor U516 (N_516,In_527,In_425);
nor U517 (N_517,In_1889,In_1922);
nor U518 (N_518,In_943,In_1638);
and U519 (N_519,In_1977,N_254);
and U520 (N_520,In_850,In_18);
nand U521 (N_521,In_1385,In_922);
nand U522 (N_522,In_1832,In_1487);
and U523 (N_523,N_413,In_890);
nand U524 (N_524,In_1354,In_675);
xnor U525 (N_525,In_1035,In_1502);
xor U526 (N_526,In_466,In_385);
nand U527 (N_527,N_127,N_262);
nor U528 (N_528,In_1943,In_1058);
and U529 (N_529,In_1882,In_1568);
nand U530 (N_530,In_1548,N_166);
and U531 (N_531,In_326,N_376);
and U532 (N_532,In_787,N_311);
and U533 (N_533,In_1627,In_407);
and U534 (N_534,N_452,In_1904);
nand U535 (N_535,In_1171,In_1545);
and U536 (N_536,N_232,In_1196);
or U537 (N_537,In_836,N_343);
xnor U538 (N_538,In_1086,In_1454);
nor U539 (N_539,In_512,In_1095);
or U540 (N_540,In_1018,N_359);
nor U541 (N_541,In_1467,In_1400);
xnor U542 (N_542,In_629,N_155);
or U543 (N_543,In_846,In_1101);
or U544 (N_544,In_709,N_61);
and U545 (N_545,In_1125,In_931);
and U546 (N_546,N_327,N_363);
or U547 (N_547,In_1799,In_243);
nand U548 (N_548,In_41,In_861);
nor U549 (N_549,In_1233,N_399);
or U550 (N_550,N_450,N_119);
xnor U551 (N_551,In_1255,In_1538);
nor U552 (N_552,In_1619,In_1858);
nor U553 (N_553,In_1866,In_741);
xnor U554 (N_554,In_1666,N_336);
nor U555 (N_555,N_180,In_275);
nand U556 (N_556,In_432,In_1681);
nor U557 (N_557,N_252,In_473);
nand U558 (N_558,In_1263,In_829);
nor U559 (N_559,In_823,In_982);
or U560 (N_560,In_1117,In_1814);
and U561 (N_561,In_1172,N_122);
nor U562 (N_562,N_23,In_1960);
nor U563 (N_563,In_1473,N_439);
nor U564 (N_564,In_298,In_761);
xor U565 (N_565,N_29,In_1553);
and U566 (N_566,In_1267,In_621);
or U567 (N_567,In_1275,In_1448);
and U568 (N_568,In_534,In_1828);
xnor U569 (N_569,In_1324,In_49);
nor U570 (N_570,N_457,In_863);
and U571 (N_571,In_858,N_1);
or U572 (N_572,In_257,In_1068);
nand U573 (N_573,N_38,N_390);
or U574 (N_574,In_184,In_1311);
nand U575 (N_575,In_1552,In_1353);
nand U576 (N_576,In_218,In_1051);
and U577 (N_577,N_379,In_1811);
or U578 (N_578,In_1826,N_213);
nand U579 (N_579,In_1177,In_735);
nand U580 (N_580,In_53,In_208);
or U581 (N_581,In_25,In_976);
nor U582 (N_582,In_809,In_1094);
xnor U583 (N_583,N_341,In_1795);
or U584 (N_584,In_1420,In_57);
and U585 (N_585,In_361,In_908);
and U586 (N_586,In_510,In_1408);
nor U587 (N_587,In_384,In_1812);
and U588 (N_588,N_437,In_1371);
or U589 (N_589,In_746,In_1287);
or U590 (N_590,N_391,In_851);
and U591 (N_591,N_427,N_304);
nand U592 (N_592,In_1373,In_951);
nand U593 (N_593,In_1521,N_393);
nand U594 (N_594,In_842,In_107);
nor U595 (N_595,In_1221,N_125);
or U596 (N_596,In_433,N_45);
nor U597 (N_597,In_1620,N_294);
nor U598 (N_598,In_730,In_620);
nand U599 (N_599,In_1410,In_364);
or U600 (N_600,In_940,In_1466);
or U601 (N_601,In_382,N_419);
or U602 (N_602,N_468,N_47);
nor U603 (N_603,In_1464,In_1986);
or U604 (N_604,N_250,In_1341);
nand U605 (N_605,In_1779,In_1556);
or U606 (N_606,In_1250,In_751);
and U607 (N_607,In_328,N_58);
and U608 (N_608,In_1976,N_91);
xor U609 (N_609,In_1469,In_492);
or U610 (N_610,In_790,In_1603);
nor U611 (N_611,N_196,In_678);
and U612 (N_612,In_905,In_1406);
and U613 (N_613,In_756,In_1611);
or U614 (N_614,N_147,N_142);
and U615 (N_615,N_401,In_1525);
nand U616 (N_616,In_1629,In_897);
nor U617 (N_617,In_1281,In_1560);
nor U618 (N_618,In_1048,In_1588);
nor U619 (N_619,In_935,In_397);
nand U620 (N_620,In_387,In_975);
nand U621 (N_621,In_1990,In_1555);
nand U622 (N_622,In_1710,In_1403);
nand U623 (N_623,In_676,N_326);
nor U624 (N_624,In_127,In_1159);
nor U625 (N_625,N_199,N_308);
nor U626 (N_626,N_187,In_1793);
xor U627 (N_627,N_86,In_1237);
nor U628 (N_628,In_1331,In_486);
nor U629 (N_629,In_1407,In_1258);
and U630 (N_630,In_1482,In_1735);
nand U631 (N_631,In_154,In_1207);
xor U632 (N_632,In_426,In_160);
nand U633 (N_633,N_429,In_732);
and U634 (N_634,In_819,N_438);
xnor U635 (N_635,In_106,In_956);
xor U636 (N_636,In_1893,In_1711);
or U637 (N_637,N_55,N_230);
nor U638 (N_638,In_1277,In_1835);
and U639 (N_639,In_1179,In_1951);
nand U640 (N_640,N_462,In_1917);
and U641 (N_641,N_536,In_1876);
and U642 (N_642,In_1046,In_865);
and U643 (N_643,In_1443,In_1973);
nor U644 (N_644,N_194,N_467);
nor U645 (N_645,In_1355,In_277);
nor U646 (N_646,In_1758,In_299);
nand U647 (N_647,In_389,In_383);
and U648 (N_648,In_734,In_1905);
nand U649 (N_649,In_306,In_893);
or U650 (N_650,In_845,In_149);
and U651 (N_651,N_527,In_1559);
nor U652 (N_652,In_948,N_217);
or U653 (N_653,In_1618,In_936);
or U654 (N_654,In_1665,In_253);
nor U655 (N_655,In_630,In_1232);
or U656 (N_656,In_399,In_481);
nand U657 (N_657,In_551,In_475);
xor U658 (N_658,N_524,N_492);
nand U659 (N_659,In_1377,N_2);
xnor U660 (N_660,In_286,N_280);
nand U661 (N_661,In_220,N_446);
nand U662 (N_662,N_30,N_382);
nor U663 (N_663,N_335,In_1563);
and U664 (N_664,In_1547,N_310);
and U665 (N_665,In_1056,In_1417);
nand U666 (N_666,In_1461,In_1605);
or U667 (N_667,In_1558,In_1243);
nor U668 (N_668,In_86,N_546);
and U669 (N_669,In_177,In_1635);
or U670 (N_670,In_604,N_12);
nand U671 (N_671,In_1050,In_1785);
and U672 (N_672,N_460,In_331);
and U673 (N_673,N_240,N_485);
nand U674 (N_674,N_271,In_226);
and U675 (N_675,In_1158,In_35);
nand U676 (N_676,In_885,N_66);
or U677 (N_677,In_814,N_99);
xor U678 (N_678,In_726,N_386);
xnor U679 (N_679,In_477,In_343);
xnor U680 (N_680,In_1652,In_1399);
nand U681 (N_681,N_81,In_1110);
nor U682 (N_682,In_1381,In_1833);
nor U683 (N_683,N_625,In_1280);
and U684 (N_684,In_711,N_222);
nor U685 (N_685,N_116,In_1928);
nor U686 (N_686,In_1549,In_868);
or U687 (N_687,N_249,N_259);
nand U688 (N_688,In_745,In_1092);
nor U689 (N_689,In_362,In_686);
and U690 (N_690,N_177,In_528);
nor U691 (N_691,N_275,In_105);
or U692 (N_692,N_85,In_1540);
nand U693 (N_693,In_1030,N_566);
nand U694 (N_694,N_604,N_325);
nor U695 (N_695,N_434,N_261);
nand U696 (N_696,N_506,N_355);
nor U697 (N_697,In_1223,N_459);
nand U698 (N_698,In_330,N_56);
nor U699 (N_699,In_242,In_1384);
and U700 (N_700,N_529,N_13);
nand U701 (N_701,N_417,In_449);
nand U702 (N_702,In_115,In_1315);
and U703 (N_703,N_622,In_1878);
and U704 (N_704,In_71,In_702);
nor U705 (N_705,N_300,In_1202);
nand U706 (N_706,In_340,In_221);
xnor U707 (N_707,N_320,In_1676);
nor U708 (N_708,In_176,In_1235);
or U709 (N_709,N_581,N_549);
or U710 (N_710,In_276,N_392);
nand U711 (N_711,In_1689,In_777);
and U712 (N_712,In_1393,In_844);
nor U713 (N_713,In_989,In_440);
nand U714 (N_714,In_1945,In_1886);
nand U715 (N_715,N_89,In_99);
and U716 (N_716,In_618,In_454);
or U717 (N_717,In_1788,N_123);
or U718 (N_718,In_493,In_442);
xor U719 (N_719,In_1358,N_121);
xor U720 (N_720,N_495,In_1115);
nor U721 (N_721,N_34,In_1260);
nor U722 (N_722,In_701,N_441);
nor U723 (N_723,N_512,In_181);
nor U724 (N_724,N_227,N_555);
and U725 (N_725,In_806,In_1195);
and U726 (N_726,N_540,In_1931);
or U727 (N_727,N_559,N_366);
xnor U728 (N_728,In_1131,In_1959);
or U729 (N_729,N_534,In_73);
nor U730 (N_730,In_549,In_1963);
xnor U731 (N_731,N_170,In_1297);
and U732 (N_732,N_428,In_1719);
xor U733 (N_733,In_1194,In_292);
or U734 (N_734,In_1386,In_1994);
nand U735 (N_735,In_633,In_1423);
nor U736 (N_736,In_316,In_977);
and U737 (N_737,N_354,In_1108);
nand U738 (N_738,In_415,N_4);
or U739 (N_739,N_409,In_281);
nand U740 (N_740,In_1723,In_1453);
nand U741 (N_741,N_631,In_871);
nand U742 (N_742,N_41,N_515);
xor U743 (N_743,In_1424,In_648);
nand U744 (N_744,In_586,N_583);
nand U745 (N_745,N_163,In_290);
or U746 (N_746,In_1098,N_109);
nor U747 (N_747,N_533,N_617);
or U748 (N_748,N_211,In_795);
or U749 (N_749,In_346,In_1379);
nor U750 (N_750,N_202,In_729);
nor U751 (N_751,N_567,In_531);
nand U752 (N_752,In_1881,In_247);
or U753 (N_753,In_1415,In_166);
nand U754 (N_754,N_520,N_627);
or U755 (N_755,In_812,In_445);
nand U756 (N_756,N_612,In_519);
nand U757 (N_757,In_1042,N_207);
and U758 (N_758,In_325,In_1036);
and U759 (N_759,N_332,In_1698);
nand U760 (N_760,N_258,In_717);
or U761 (N_761,In_1479,In_1370);
nor U762 (N_762,In_1157,In_1365);
or U763 (N_763,In_830,In_1631);
and U764 (N_764,In_1203,In_1034);
nand U765 (N_765,In_1099,In_942);
or U766 (N_766,N_578,In_501);
and U767 (N_767,N_607,In_1879);
nor U768 (N_768,N_532,N_53);
nand U769 (N_769,In_1784,In_1862);
or U770 (N_770,In_1966,In_12);
nand U771 (N_771,N_245,In_450);
and U772 (N_772,N_613,N_190);
or U773 (N_773,In_1821,In_1920);
and U774 (N_774,In_1053,In_5);
and U775 (N_775,In_1830,In_200);
or U776 (N_776,In_722,In_1697);
and U777 (N_777,N_472,N_281);
or U778 (N_778,In_32,N_426);
nor U779 (N_779,In_1535,In_972);
xnor U780 (N_780,N_454,In_1543);
nand U781 (N_781,N_256,In_725);
xnor U782 (N_782,In_438,In_733);
nand U783 (N_783,In_1947,N_531);
or U784 (N_784,In_1802,N_104);
and U785 (N_785,In_692,N_168);
and U786 (N_786,In_894,In_533);
nand U787 (N_787,In_1857,In_879);
nor U788 (N_788,In_691,N_568);
and U789 (N_789,In_402,N_274);
or U790 (N_790,In_1499,In_1780);
or U791 (N_791,N_357,In_554);
and U792 (N_792,In_1193,In_1216);
nor U793 (N_793,In_740,In_228);
and U794 (N_794,N_96,In_1206);
and U795 (N_795,In_278,In_388);
nand U796 (N_796,In_1340,In_1501);
and U797 (N_797,In_88,In_1915);
and U798 (N_798,N_35,N_255);
and U799 (N_799,In_1442,In_1577);
and U800 (N_800,In_595,In_28);
and U801 (N_801,In_708,N_46);
nand U802 (N_802,In_476,In_1993);
xnor U803 (N_803,N_686,In_920);
xnor U804 (N_804,N_18,In_1462);
and U805 (N_805,In_420,N_449);
xnor U806 (N_806,N_640,In_238);
xor U807 (N_807,N_577,In_1052);
or U808 (N_808,In_1069,In_994);
nand U809 (N_809,In_1162,N_630);
nand U810 (N_810,N_402,N_624);
xor U811 (N_811,In_1691,In_410);
and U812 (N_812,In_1700,N_105);
nor U813 (N_813,N_509,In_188);
nor U814 (N_814,N_269,In_400);
and U815 (N_815,In_1992,In_870);
nand U816 (N_816,In_1768,N_652);
nand U817 (N_817,In_626,In_354);
nor U818 (N_818,N_648,N_651);
or U819 (N_819,In_1609,In_704);
nor U820 (N_820,In_1614,In_1405);
and U821 (N_821,In_349,N_204);
and U822 (N_822,N_528,In_123);
nand U823 (N_823,N_774,In_1542);
nor U824 (N_824,In_1961,In_1409);
nor U825 (N_825,N_425,In_356);
nor U826 (N_826,In_1865,In_886);
or U827 (N_827,In_1504,In_1010);
xor U828 (N_828,N_674,In_1320);
or U829 (N_829,In_765,N_610);
nor U830 (N_830,N_356,N_51);
or U831 (N_831,N_157,In_1599);
nor U832 (N_832,In_1628,In_128);
or U833 (N_833,In_1642,In_1859);
and U834 (N_834,N_76,N_106);
or U835 (N_835,N_650,N_330);
or U836 (N_836,N_307,N_139);
or U837 (N_837,In_775,N_605);
nor U838 (N_838,In_1037,N_699);
xnor U839 (N_839,In_1850,N_340);
or U840 (N_840,N_235,In_195);
and U841 (N_841,N_602,N_611);
nor U842 (N_842,N_293,N_636);
or U843 (N_843,N_380,In_748);
nor U844 (N_844,In_959,In_190);
nand U845 (N_845,N_266,N_451);
and U846 (N_846,N_345,N_702);
xnor U847 (N_847,In_1659,In_1);
nor U848 (N_848,In_6,N_291);
or U849 (N_849,In_1957,In_1658);
or U850 (N_850,N_491,In_1210);
or U851 (N_851,N_759,In_1509);
or U852 (N_852,N_561,N_705);
nor U853 (N_853,N_764,N_306);
or U854 (N_854,In_130,In_1428);
nor U855 (N_855,In_211,In_1899);
and U856 (N_856,N_576,N_562);
nor U857 (N_857,N_138,In_1447);
nand U858 (N_858,N_783,In_175);
or U859 (N_859,In_776,In_1312);
nor U860 (N_860,In_321,N_253);
nor U861 (N_861,In_928,In_1460);
nor U862 (N_862,N_251,In_1583);
or U863 (N_863,N_350,In_1819);
and U864 (N_864,In_1908,N_0);
or U865 (N_865,In_212,In_500);
nor U866 (N_866,In_1136,N_706);
and U867 (N_867,N_556,In_888);
nand U868 (N_868,In_36,N_339);
nor U869 (N_869,N_731,In_1471);
or U870 (N_870,N_161,In_848);
and U871 (N_871,In_1165,N_700);
nor U872 (N_872,In_1673,N_395);
or U873 (N_873,N_445,N_552);
and U874 (N_874,In_137,N_621);
or U875 (N_875,In_754,N_608);
and U876 (N_876,N_688,N_550);
or U877 (N_877,N_132,N_564);
nand U878 (N_878,In_763,In_1493);
or U879 (N_879,N_689,N_135);
nor U880 (N_880,N_596,In_245);
xnor U881 (N_881,In_1594,In_502);
nor U882 (N_882,In_230,In_1939);
or U883 (N_883,N_186,N_720);
nand U884 (N_884,N_690,In_985);
and U885 (N_885,N_171,In_1581);
nand U886 (N_886,N_17,N_479);
nor U887 (N_887,In_405,In_966);
xnor U888 (N_888,N_618,In_831);
and U889 (N_889,N_594,In_609);
xnor U890 (N_890,N_197,In_825);
nand U891 (N_891,In_1699,In_1964);
and U892 (N_892,In_303,In_1532);
and U893 (N_893,In_839,N_544);
nor U894 (N_894,In_1643,In_536);
or U895 (N_895,In_1999,In_1625);
nand U896 (N_896,N_718,N_368);
or U897 (N_897,In_1253,In_1305);
nor U898 (N_898,In_610,N_557);
and U899 (N_899,In_1887,N_158);
nand U900 (N_900,N_210,In_1245);
or U901 (N_901,In_1279,N_496);
xnor U902 (N_902,N_733,In_1264);
nor U903 (N_903,In_1369,N_595);
xor U904 (N_904,In_1360,N_358);
nor U905 (N_905,In_308,N_571);
nor U906 (N_906,N_713,In_1933);
nor U907 (N_907,N_649,N_768);
nor U908 (N_908,In_246,In_1815);
or U909 (N_909,In_462,In_1616);
and U910 (N_910,N_537,N_198);
nor U911 (N_911,N_758,In_1515);
nand U912 (N_912,N_569,In_322);
or U913 (N_913,In_1839,N_701);
or U914 (N_914,N_39,N_133);
or U915 (N_915,N_456,N_279);
nor U916 (N_916,In_558,N_667);
and U917 (N_917,N_779,In_1875);
nand U918 (N_918,N_474,In_138);
xnor U919 (N_919,In_1980,N_765);
or U920 (N_920,N_337,In_1484);
nor U921 (N_921,In_46,In_565);
nor U922 (N_922,In_1953,N_791);
xor U923 (N_923,N_372,N_389);
nand U924 (N_924,In_1323,N_342);
nor U925 (N_925,In_1310,N_458);
nor U926 (N_926,N_760,N_761);
and U927 (N_927,In_336,N_205);
nor U928 (N_928,In_587,N_582);
nor U929 (N_929,In_1527,N_547);
xnor U930 (N_930,In_368,In_791);
and U931 (N_931,N_448,N_16);
xor U932 (N_932,N_638,In_1813);
and U933 (N_933,In_1390,In_1777);
and U934 (N_934,N_493,N_563);
nand U935 (N_935,N_346,In_44);
nor U936 (N_936,N_780,In_1041);
nand U937 (N_937,In_370,N_497);
nor U938 (N_938,In_1199,N_668);
or U939 (N_939,In_705,In_1754);
nor U940 (N_940,N_710,N_698);
xnor U941 (N_941,N_25,In_1646);
nor U942 (N_942,N_684,N_276);
xnor U943 (N_943,In_1016,N_349);
and U944 (N_944,In_1838,In_590);
and U945 (N_945,N_697,In_374);
nor U946 (N_946,In_244,In_1326);
nor U947 (N_947,N_108,In_84);
nor U948 (N_948,In_287,N_666);
nor U949 (N_949,In_781,N_499);
or U950 (N_950,In_1763,N_148);
xor U951 (N_951,In_1732,N_226);
or U952 (N_952,N_687,In_54);
nor U953 (N_953,In_525,N_772);
nor U954 (N_954,N_778,In_282);
xnor U955 (N_955,N_530,In_121);
xnor U956 (N_956,In_653,In_1422);
or U957 (N_957,N_510,N_542);
nand U958 (N_958,N_344,N_482);
nand U959 (N_959,In_950,N_696);
and U960 (N_960,In_1333,In_31);
nor U961 (N_961,N_929,In_997);
nand U962 (N_962,In_1972,In_600);
nand U963 (N_963,In_209,In_1317);
and U964 (N_964,N_738,In_1240);
nor U965 (N_965,N_959,N_918);
nor U966 (N_966,In_1705,In_1996);
nand U967 (N_967,In_1472,N_518);
or U968 (N_968,In_0,N_954);
and U969 (N_969,N_817,N_717);
nand U970 (N_970,N_691,In_926);
nand U971 (N_971,N_815,N_755);
nand U972 (N_972,N_430,N_184);
and U973 (N_973,In_307,In_1395);
nor U974 (N_974,In_1721,In_540);
nand U975 (N_975,N_642,N_586);
or U976 (N_976,N_785,In_665);
or U977 (N_977,In_1156,In_1380);
nand U978 (N_978,N_59,N_263);
xnor U979 (N_979,In_62,In_1765);
or U980 (N_980,N_97,In_1332);
nand U981 (N_981,N_870,In_91);
nand U982 (N_982,In_1026,In_1759);
nor U983 (N_983,N_673,In_418);
or U984 (N_984,In_318,In_222);
nand U985 (N_985,In_1327,N_129);
or U986 (N_986,In_1776,In_674);
nand U987 (N_987,N_516,In_1925);
nor U988 (N_988,N_64,In_784);
or U989 (N_989,In_132,In_196);
nand U990 (N_990,N_722,N_911);
nand U991 (N_991,In_969,N_829);
xnor U992 (N_992,N_752,N_178);
nand U993 (N_993,In_1892,N_887);
and U994 (N_994,N_903,N_734);
or U995 (N_995,In_428,In_1389);
nand U996 (N_996,In_1011,N_353);
nand U997 (N_997,N_937,In_66);
nor U998 (N_998,In_1677,In_978);
and U999 (N_999,In_979,In_213);
nand U1000 (N_1000,N_554,In_191);
or U1001 (N_1001,N_498,N_494);
or U1002 (N_1002,N_756,In_74);
and U1003 (N_1003,In_987,N_385);
nand U1004 (N_1004,In_1736,In_1621);
nand U1005 (N_1005,N_78,N_838);
and U1006 (N_1006,In_998,In_1675);
and U1007 (N_1007,In_1663,In_1781);
and U1008 (N_1008,In_1584,N_331);
or U1009 (N_1009,In_1175,In_1942);
nand U1010 (N_1010,N_115,In_965);
nor U1011 (N_1011,N_247,N_724);
nand U1012 (N_1012,In_1457,In_961);
and U1013 (N_1013,N_857,N_404);
nor U1014 (N_1014,In_841,In_1916);
nor U1015 (N_1015,N_827,In_883);
or U1016 (N_1016,N_896,In_118);
or U1017 (N_1017,In_1293,N_910);
or U1018 (N_1018,N_521,In_712);
nand U1019 (N_1019,In_684,In_380);
or U1020 (N_1020,In_1455,N_763);
xnor U1021 (N_1021,In_518,In_1127);
nor U1022 (N_1022,N_188,In_1520);
xnor U1023 (N_1023,In_304,In_114);
nand U1024 (N_1024,N_899,N_716);
nor U1025 (N_1025,In_1057,N_802);
and U1026 (N_1026,N_801,In_1439);
xnor U1027 (N_1027,In_1685,N_297);
nand U1028 (N_1028,In_571,N_634);
nor U1029 (N_1029,N_934,N_735);
and U1030 (N_1030,N_162,In_1239);
nand U1031 (N_1031,N_408,In_1304);
nor U1032 (N_1032,In_736,N_925);
and U1033 (N_1033,N_858,In_1388);
nor U1034 (N_1034,N_743,N_939);
nor U1035 (N_1035,N_360,In_1085);
nor U1036 (N_1036,In_900,N_900);
and U1037 (N_1037,N_420,N_264);
nand U1038 (N_1038,N_110,In_403);
and U1039 (N_1039,N_898,In_459);
nor U1040 (N_1040,N_200,In_80);
and U1041 (N_1041,In_1742,N_729);
and U1042 (N_1042,In_1946,In_530);
or U1043 (N_1043,N_737,In_345);
nand U1044 (N_1044,In_329,In_1059);
nor U1045 (N_1045,N_676,N_626);
nor U1046 (N_1046,N_381,N_69);
nand U1047 (N_1047,N_664,N_414);
and U1048 (N_1048,In_1653,N_268);
nor U1049 (N_1049,In_1412,N_721);
nor U1050 (N_1050,In_1306,In_832);
nand U1051 (N_1051,N_936,N_868);
and U1052 (N_1052,In_45,N_238);
nor U1053 (N_1053,In_1601,In_902);
nor U1054 (N_1054,N_519,In_1590);
nand U1055 (N_1055,In_575,In_637);
nor U1056 (N_1056,N_526,N_677);
and U1057 (N_1057,In_984,In_952);
nand U1058 (N_1058,N_893,N_736);
or U1059 (N_1059,In_1269,N_850);
nand U1060 (N_1060,N_902,In_1792);
nor U1061 (N_1061,In_1729,In_807);
nand U1062 (N_1062,In_679,N_599);
and U1063 (N_1063,N_767,In_973);
and U1064 (N_1064,In_1434,N_847);
or U1065 (N_1065,N_589,In_683);
and U1066 (N_1066,N_315,N_747);
or U1067 (N_1067,In_543,In_645);
and U1068 (N_1068,N_505,N_63);
or U1069 (N_1069,In_1869,In_489);
and U1070 (N_1070,In_1693,N_852);
nand U1071 (N_1071,In_437,N_292);
nor U1072 (N_1072,In_1478,In_1236);
or U1073 (N_1073,In_884,In_139);
nor U1074 (N_1074,N_591,N_844);
nor U1075 (N_1075,N_432,N_814);
nand U1076 (N_1076,In_537,N_504);
xnor U1077 (N_1077,In_1626,N_616);
nand U1078 (N_1078,In_125,In_636);
and U1079 (N_1079,N_453,In_192);
nor U1080 (N_1080,N_742,N_769);
and U1081 (N_1081,N_74,N_416);
or U1082 (N_1082,In_957,In_1703);
nand U1083 (N_1083,In_1296,N_21);
or U1084 (N_1084,In_263,In_1119);
or U1085 (N_1085,In_1105,In_1808);
and U1086 (N_1086,In_272,In_723);
xor U1087 (N_1087,N_601,In_392);
or U1088 (N_1088,N_661,In_580);
or U1089 (N_1089,N_370,In_26);
nand U1090 (N_1090,N_397,In_1019);
or U1091 (N_1091,N_447,In_1212);
and U1092 (N_1092,In_925,In_314);
nor U1093 (N_1093,In_1064,In_550);
and U1094 (N_1094,N_655,N_575);
nor U1095 (N_1095,N_926,In_499);
nor U1096 (N_1096,N_421,In_914);
nand U1097 (N_1097,In_516,In_262);
nand U1098 (N_1098,N_881,N_165);
xnor U1099 (N_1099,In_366,In_992);
nand U1100 (N_1100,N_855,In_1234);
or U1101 (N_1101,In_1816,N_270);
xor U1102 (N_1102,N_913,In_1709);
nand U1103 (N_1103,N_730,N_879);
nor U1104 (N_1104,N_319,In_1303);
nor U1105 (N_1105,N_384,In_1644);
nand U1106 (N_1106,In_909,In_451);
and U1107 (N_1107,In_835,N_892);
or U1108 (N_1108,In_1880,In_414);
and U1109 (N_1109,In_158,In_1154);
or U1110 (N_1110,N_229,In_1918);
or U1111 (N_1111,In_38,In_854);
and U1112 (N_1112,N_680,In_102);
or U1113 (N_1113,N_866,In_199);
nor U1114 (N_1114,In_1027,In_313);
nor U1115 (N_1115,N_833,N_853);
and U1116 (N_1116,In_1141,In_1339);
nor U1117 (N_1117,In_919,N_906);
nor U1118 (N_1118,N_403,N_283);
nand U1119 (N_1119,N_71,In_594);
or U1120 (N_1120,In_1783,N_580);
nand U1121 (N_1121,In_682,In_757);
nor U1122 (N_1122,N_8,In_1950);
or U1123 (N_1123,In_1093,In_1256);
or U1124 (N_1124,N_860,N_816);
or U1125 (N_1125,N_480,N_1097);
or U1126 (N_1126,In_1488,N_1056);
or U1127 (N_1127,N_901,N_886);
and U1128 (N_1128,In_1055,N_1046);
xnor U1129 (N_1129,N_598,In_1062);
and U1130 (N_1130,N_1016,In_483);
and U1131 (N_1131,In_309,In_643);
nand U1132 (N_1132,N_989,N_11);
nor U1133 (N_1133,In_1214,N_114);
and U1134 (N_1134,N_728,In_1936);
nand U1135 (N_1135,N_912,In_934);
or U1136 (N_1136,In_1349,N_410);
and U1137 (N_1137,N_484,N_465);
and U1138 (N_1138,In_1831,N_992);
or U1139 (N_1139,In_378,N_681);
or U1140 (N_1140,N_749,N_863);
nand U1141 (N_1141,In_134,N_966);
nand U1142 (N_1142,In_1009,In_766);
or U1143 (N_1143,In_1593,N_1109);
and U1144 (N_1144,In_348,In_372);
and U1145 (N_1145,N_654,N_1116);
or U1146 (N_1146,In_1633,In_891);
nor U1147 (N_1147,N_373,N_782);
or U1148 (N_1148,N_221,N_236);
and U1149 (N_1149,In_1595,In_396);
and U1150 (N_1150,In_94,N_1062);
nor U1151 (N_1151,In_1825,N_646);
nand U1152 (N_1152,In_1935,N_723);
and U1153 (N_1153,N_849,N_131);
nand U1154 (N_1154,N_991,N_593);
xor U1155 (N_1155,N_1000,N_775);
nand U1156 (N_1156,N_398,N_1034);
nor U1157 (N_1157,In_1639,N_920);
or U1158 (N_1158,In_1383,N_107);
nor U1159 (N_1159,N_977,N_541);
nand U1160 (N_1160,In_92,N_865);
and U1161 (N_1161,In_1513,N_797);
and U1162 (N_1162,In_771,In_769);
nand U1163 (N_1163,In_892,In_918);
nand U1164 (N_1164,In_453,N_422);
xor U1165 (N_1165,In_731,In_461);
or U1166 (N_1166,N_808,In_1820);
and U1167 (N_1167,N_776,N_1054);
nand U1168 (N_1168,N_660,N_490);
or U1169 (N_1169,N_864,N_314);
or U1170 (N_1170,In_27,In_267);
nand U1171 (N_1171,In_1510,In_85);
or U1172 (N_1172,N_804,N_1017);
and U1173 (N_1173,N_635,In_1706);
nand U1174 (N_1174,In_1285,N_1029);
xor U1175 (N_1175,In_669,In_1853);
nor U1176 (N_1176,In_395,In_78);
nand U1177 (N_1177,In_1345,N_968);
or U1178 (N_1178,N_1110,N_412);
or U1179 (N_1179,In_1445,N_1040);
nand U1180 (N_1180,N_1027,N_514);
and U1181 (N_1181,N_600,In_42);
or U1182 (N_1182,In_577,In_661);
or U1183 (N_1183,In_498,In_974);
nand U1184 (N_1184,N_945,N_218);
and U1185 (N_1185,N_216,N_208);
nor U1186 (N_1186,In_1531,N_732);
nor U1187 (N_1187,N_585,In_579);
nand U1188 (N_1188,In_932,N_1112);
or U1189 (N_1189,N_659,In_1394);
nor U1190 (N_1190,In_1574,In_289);
nand U1191 (N_1191,N_994,N_538);
nor U1192 (N_1192,N_835,N_675);
nand U1193 (N_1193,N_488,N_1071);
and U1194 (N_1194,N_243,N_805);
nor U1195 (N_1195,N_1095,In_859);
or U1196 (N_1196,N_1105,In_68);
or U1197 (N_1197,In_169,In_1890);
and U1198 (N_1198,N_1038,N_708);
and U1199 (N_1199,N_967,N_272);
or U1200 (N_1200,In_219,In_1551);
and U1201 (N_1201,N_770,In_714);
or U1202 (N_1202,N_657,N_1072);
xor U1203 (N_1203,N_574,In_417);
nor U1204 (N_1204,N_1119,N_941);
or U1205 (N_1205,N_77,In_1801);
nor U1206 (N_1206,N_753,N_1004);
nor U1207 (N_1207,N_1007,N_859);
and U1208 (N_1208,In_616,In_401);
or U1209 (N_1209,N_615,N_592);
xnor U1210 (N_1210,N_1094,N_523);
or U1211 (N_1211,In_347,In_1929);
nor U1212 (N_1212,In_1630,N_1013);
nand U1213 (N_1213,N_895,N_980);
and U1214 (N_1214,In_535,In_913);
nor U1215 (N_1215,In_833,N_828);
nand U1216 (N_1216,N_1009,N_1088);
and U1217 (N_1217,In_810,N_707);
nand U1218 (N_1218,In_744,N_665);
nand U1219 (N_1219,N_1079,In_381);
xnor U1220 (N_1220,In_584,N_663);
nand U1221 (N_1221,In_162,In_223);
nand U1222 (N_1222,In_1541,In_668);
nand U1223 (N_1223,N_1068,In_1368);
or U1224 (N_1224,N_773,N_1055);
nand U1225 (N_1225,N_990,N_365);
nand U1226 (N_1226,In_484,N_826);
nor U1227 (N_1227,In_1991,N_682);
or U1228 (N_1228,N_418,N_501);
and U1229 (N_1229,N_1106,N_141);
xor U1230 (N_1230,N_914,In_638);
or U1231 (N_1231,In_1490,N_639);
and U1232 (N_1232,N_400,N_633);
xor U1233 (N_1233,N_522,In_1215);
nor U1234 (N_1234,In_774,N_794);
and U1235 (N_1235,In_880,N_1051);
nand U1236 (N_1236,In_560,N_909);
nor U1237 (N_1237,In_1124,N_587);
or U1238 (N_1238,In_818,N_983);
or U1239 (N_1239,N_375,N_1043);
xnor U1240 (N_1240,In_1276,In_1451);
and U1241 (N_1241,N_629,N_1026);
xnor U1242 (N_1242,N_880,N_70);
nand U1243 (N_1243,N_848,In_559);
and U1244 (N_1244,N_930,In_1804);
or U1245 (N_1245,N_924,N_962);
nand U1246 (N_1246,In_511,In_1764);
and U1247 (N_1247,In_1683,N_54);
nand U1248 (N_1248,N_641,N_1035);
and U1249 (N_1249,N_565,N_124);
nand U1250 (N_1250,N_324,N_140);
nor U1251 (N_1251,N_821,N_995);
nor U1252 (N_1252,N_1083,N_579);
nor U1253 (N_1253,N_1100,N_692);
xor U1254 (N_1254,N_979,N_40);
nor U1255 (N_1255,In_1989,N_52);
and U1256 (N_1256,N_374,N_803);
nor U1257 (N_1257,N_500,N_94);
and U1258 (N_1258,N_101,N_975);
or U1259 (N_1259,In_737,N_572);
and U1260 (N_1260,N_1005,N_810);
nand U1261 (N_1261,In_509,In_1722);
or U1262 (N_1262,In_1111,N_333);
and U1263 (N_1263,N_669,N_933);
nor U1264 (N_1264,N_145,In_1492);
and U1265 (N_1265,In_1248,N_1076);
nand U1266 (N_1266,In_760,In_1608);
nor U1267 (N_1267,N_470,N_796);
and U1268 (N_1268,N_787,N_407);
and U1269 (N_1269,N_644,In_1987);
and U1270 (N_1270,N_118,In_896);
or U1271 (N_1271,In_523,In_1914);
or U1272 (N_1272,N_405,N_693);
and U1273 (N_1273,N_685,In_611);
nand U1274 (N_1274,In_654,In_1021);
or U1275 (N_1275,In_1307,In_672);
nor U1276 (N_1276,N_415,N_1025);
nor U1277 (N_1277,N_750,In_1187);
xor U1278 (N_1278,In_1372,N_988);
nand U1279 (N_1279,N_781,In_1873);
nor U1280 (N_1280,In_589,N_1254);
nand U1281 (N_1281,N_377,N_834);
nor U1282 (N_1282,N_1150,In_544);
nand U1283 (N_1283,N_539,N_466);
nand U1284 (N_1284,N_969,N_1265);
and U1285 (N_1285,N_998,N_1264);
xor U1286 (N_1286,N_1224,N_545);
or U1287 (N_1287,N_1202,N_548);
and U1288 (N_1288,N_957,N_1180);
and U1289 (N_1289,N_1015,N_435);
nor U1290 (N_1290,N_928,N_619);
nor U1291 (N_1291,N_1214,In_1290);
or U1292 (N_1292,In_770,N_1234);
xnor U1293 (N_1293,N_1036,N_1213);
nand U1294 (N_1294,N_921,N_1081);
nor U1295 (N_1295,N_442,N_189);
and U1296 (N_1296,N_792,N_1063);
or U1297 (N_1297,N_1102,N_1065);
and U1298 (N_1298,N_812,N_1259);
or U1299 (N_1299,N_1111,N_1172);
nor U1300 (N_1300,In_963,In_720);
and U1301 (N_1301,N_273,N_1080);
nor U1302 (N_1302,N_823,N_584);
or U1303 (N_1303,In_259,N_609);
nand U1304 (N_1304,N_679,N_1127);
or U1305 (N_1305,In_1958,N_1053);
and U1306 (N_1306,In_944,In_1438);
and U1307 (N_1307,N_961,N_352);
and U1308 (N_1308,N_329,N_206);
and U1309 (N_1309,N_1126,In_1298);
and U1310 (N_1310,N_822,N_671);
nand U1311 (N_1311,In_724,In_840);
nor U1312 (N_1312,N_1185,In_614);
xnor U1313 (N_1313,N_963,N_987);
xor U1314 (N_1314,In_1107,In_1183);
xnor U1315 (N_1315,N_1260,In_681);
nor U1316 (N_1316,N_766,N_1266);
xor U1317 (N_1317,In_1570,In_874);
xnor U1318 (N_1318,N_321,N_553);
and U1319 (N_1319,N_179,N_1033);
xor U1320 (N_1320,In_1254,N_469);
nand U1321 (N_1321,In_545,In_260);
or U1322 (N_1322,N_383,N_1248);
nor U1323 (N_1323,N_486,In_1031);
nand U1324 (N_1324,N_1183,N_943);
nand U1325 (N_1325,In_435,In_1585);
nand U1326 (N_1326,In_1902,N_1153);
nand U1327 (N_1327,In_1937,N_1175);
nand U1328 (N_1328,N_837,N_1022);
nand U1329 (N_1329,N_1028,In_864);
nand U1330 (N_1330,In_1954,N_1147);
or U1331 (N_1331,N_1276,In_797);
nor U1332 (N_1332,N_809,N_862);
or U1333 (N_1333,In_715,N_748);
nor U1334 (N_1334,N_167,N_800);
or U1335 (N_1335,In_1854,In_788);
nor U1336 (N_1336,N_1121,In_1597);
nor U1337 (N_1337,N_1156,In_570);
nand U1338 (N_1338,N_1052,N_543);
nor U1339 (N_1339,N_1124,N_1162);
nor U1340 (N_1340,N_1212,N_1251);
nor U1341 (N_1341,N_1209,N_1232);
and U1342 (N_1342,N_726,In_1020);
nand U1343 (N_1343,N_1160,N_1268);
or U1344 (N_1344,N_1012,N_143);
and U1345 (N_1345,N_972,N_513);
nor U1346 (N_1346,In_747,N_1130);
xor U1347 (N_1347,N_234,N_364);
nor U1348 (N_1348,In_1213,N_952);
and U1349 (N_1349,N_1001,N_1082);
nor U1350 (N_1350,N_1242,N_944);
or U1351 (N_1351,N_1257,N_1178);
nor U1352 (N_1352,N_224,N_1271);
or U1353 (N_1353,N_1075,In_315);
and U1354 (N_1354,N_790,In_1006);
xnor U1355 (N_1355,N_739,N_1023);
nand U1356 (N_1356,N_678,N_875);
or U1357 (N_1357,N_725,N_653);
xor U1358 (N_1358,In_1189,N_1006);
xnor U1359 (N_1359,In_431,In_1843);
nand U1360 (N_1360,N_1216,N_289);
or U1361 (N_1361,N_658,N_935);
and U1362 (N_1362,In_862,N_1142);
nand U1363 (N_1363,N_424,N_894);
and U1364 (N_1364,N_191,N_917);
and U1365 (N_1365,N_134,N_588);
and U1366 (N_1366,N_714,N_877);
or U1367 (N_1367,N_1227,N_1118);
and U1368 (N_1368,N_1148,N_1151);
xnor U1369 (N_1369,N_328,N_694);
and U1370 (N_1370,In_1149,In_310);
and U1371 (N_1371,In_1096,N_851);
xnor U1372 (N_1372,In_1411,In_1730);
or U1373 (N_1373,N_1140,N_215);
or U1374 (N_1374,N_1169,In_1848);
nand U1375 (N_1375,N_628,In_755);
nand U1376 (N_1376,N_1070,In_1229);
nand U1377 (N_1377,In_1852,N_316);
and U1378 (N_1378,N_1218,N_1019);
nand U1379 (N_1379,In_1017,In_958);
nor U1380 (N_1380,In_1147,N_1073);
nor U1381 (N_1381,N_1186,N_1137);
and U1382 (N_1382,N_239,N_978);
nand U1383 (N_1383,N_1261,In_1613);
nand U1384 (N_1384,In_120,N_986);
or U1385 (N_1385,In_147,N_1278);
or U1386 (N_1386,N_1131,In_663);
nor U1387 (N_1387,N_982,N_709);
nand U1388 (N_1388,In_1767,N_841);
and U1389 (N_1389,N_1164,In_1863);
or U1390 (N_1390,N_302,In_100);
and U1391 (N_1391,In_1885,N_856);
nor U1392 (N_1392,N_290,N_882);
nor U1393 (N_1393,In_1637,N_1114);
or U1394 (N_1394,In_439,N_947);
nand U1395 (N_1395,N_905,N_1152);
and U1396 (N_1396,N_15,N_1117);
and U1397 (N_1397,N_1144,N_444);
nand U1398 (N_1398,In_1489,In_996);
nand U1399 (N_1399,In_233,N_1193);
and U1400 (N_1400,N_985,N_1270);
and U1401 (N_1401,N_632,In_1841);
nor U1402 (N_1402,In_504,N_1179);
nand U1403 (N_1403,N_927,N_1238);
and U1404 (N_1404,N_942,In_1576);
or U1405 (N_1405,N_1215,N_873);
nor U1406 (N_1406,N_861,N_33);
nor U1407 (N_1407,N_1163,N_570);
nor U1408 (N_1408,In_1589,N_744);
or U1409 (N_1409,N_288,N_1165);
or U1410 (N_1410,N_1077,N_277);
and U1411 (N_1411,N_1166,N_1129);
xnor U1412 (N_1412,N_1262,In_180);
xor U1413 (N_1413,In_1573,N_1146);
nand U1414 (N_1414,In_72,N_820);
and U1415 (N_1415,N_1044,In_1314);
nor U1416 (N_1416,In_699,N_1217);
nor U1417 (N_1417,N_1057,In_1334);
or U1418 (N_1418,N_1020,N_525);
nand U1419 (N_1419,In_239,N_387);
or U1420 (N_1420,N_112,N_361);
and U1421 (N_1421,N_1252,N_1198);
nor U1422 (N_1422,N_1208,N_740);
nand U1423 (N_1423,In_1834,N_1256);
xnor U1424 (N_1424,In_1137,In_1186);
nand U1425 (N_1425,N_334,In_58);
nand U1426 (N_1426,N_1176,N_1031);
nor U1427 (N_1427,N_884,N_1219);
xor U1428 (N_1428,N_904,N_956);
or U1429 (N_1429,N_309,In_1837);
or U1430 (N_1430,In_1829,In_552);
nor U1431 (N_1431,N_1098,N_1161);
or U1432 (N_1432,N_378,N_597);
or U1433 (N_1433,In_1364,N_949);
and U1434 (N_1434,N_1190,In_685);
nand U1435 (N_1435,N_832,In_33);
nand U1436 (N_1436,N_286,N_1184);
or U1437 (N_1437,N_476,N_784);
nor U1438 (N_1438,N_1253,N_560);
nor U1439 (N_1439,N_473,N_367);
or U1440 (N_1440,N_111,N_1438);
nor U1441 (N_1441,N_1382,N_1018);
and U1442 (N_1442,In_1696,N_31);
or U1443 (N_1443,In_1164,In_1252);
and U1444 (N_1444,N_1032,N_296);
and U1445 (N_1445,N_1384,N_1375);
nand U1446 (N_1446,N_1360,N_1315);
xor U1447 (N_1447,N_1235,N_1413);
nand U1448 (N_1448,N_1296,N_1376);
nor U1449 (N_1449,N_1255,In_1649);
or U1450 (N_1450,N_1336,N_1368);
or U1451 (N_1451,N_573,N_754);
nand U1452 (N_1452,N_1059,In_393);
or U1453 (N_1453,N_1108,In_652);
nand U1454 (N_1454,In_1636,N_874);
or U1455 (N_1455,N_891,In_1971);
nand U1456 (N_1456,N_1401,In_583);
nand U1457 (N_1457,N_643,N_1286);
or U1458 (N_1458,N_1138,N_1047);
nand U1459 (N_1459,N_1377,N_746);
and U1460 (N_1460,N_922,N_478);
nand U1461 (N_1461,N_1239,In_817);
nand U1462 (N_1462,N_1249,N_946);
nand U1463 (N_1463,N_1233,N_1122);
or U1464 (N_1464,N_287,N_1066);
or U1465 (N_1465,In_371,N_845);
and U1466 (N_1466,N_1403,N_1419);
nor U1467 (N_1467,In_837,In_270);
nor U1468 (N_1468,In_1459,N_1010);
nand U1469 (N_1469,N_1399,N_1086);
nand U1470 (N_1470,In_1752,N_487);
or U1471 (N_1471,In_422,N_1101);
nand U1472 (N_1472,N_1199,N_1220);
nor U1473 (N_1473,N_1245,N_1246);
or U1474 (N_1474,In_878,N_1415);
nor U1475 (N_1475,N_1359,N_1096);
and U1476 (N_1476,N_1042,N_1201);
and U1477 (N_1477,N_1349,N_1223);
or U1478 (N_1478,N_1338,N_502);
or U1479 (N_1479,N_1087,N_1300);
or U1480 (N_1480,N_711,N_1274);
xnor U1481 (N_1481,N_950,In_1750);
nand U1482 (N_1482,N_1352,In_456);
and U1483 (N_1483,N_1340,N_1240);
nor U1484 (N_1484,N_871,N_1409);
nand U1485 (N_1485,N_965,In_1227);
nor U1486 (N_1486,In_555,N_1341);
xnor U1487 (N_1487,N_1210,In_446);
nor U1488 (N_1488,N_1103,N_5);
nor U1489 (N_1489,N_788,N_1361);
and U1490 (N_1490,N_1344,N_948);
nand U1491 (N_1491,N_1289,N_953);
nand U1492 (N_1492,N_1132,N_1041);
nor U1493 (N_1493,In_204,N_1312);
nand U1494 (N_1494,N_1133,In_494);
nor U1495 (N_1495,N_916,N_463);
nand U1496 (N_1496,N_1330,N_620);
or U1497 (N_1497,N_1241,N_1374);
nand U1498 (N_1498,In_573,In_1596);
or U1499 (N_1499,In_1425,In_1874);
or U1500 (N_1500,N_1405,In_1844);
nand U1501 (N_1501,N_1356,N_1093);
nand U1502 (N_1502,N_1431,N_1362);
nand U1503 (N_1503,In_1674,N_1250);
nor U1504 (N_1504,N_431,N_1370);
or U1505 (N_1505,N_1074,N_1143);
nand U1506 (N_1506,In_1271,In_700);
nor U1507 (N_1507,N_1427,In_767);
or U1508 (N_1508,N_351,N_1191);
nand U1509 (N_1509,N_1408,In_1650);
xor U1510 (N_1510,N_1115,N_1203);
nor U1511 (N_1511,N_1372,N_973);
nor U1512 (N_1512,In_1782,N_806);
nand U1513 (N_1513,N_1302,N_1367);
and U1514 (N_1514,N_1328,N_931);
and U1515 (N_1515,N_1434,In_815);
xor U1516 (N_1516,N_908,N_1426);
nor U1517 (N_1517,N_1275,In_1167);
nand U1518 (N_1518,N_889,N_1171);
and U1519 (N_1519,N_1343,N_1348);
xor U1520 (N_1520,N_614,N_1371);
nand U1521 (N_1521,N_1335,N_1424);
and U1522 (N_1522,N_1326,N_503);
and U1523 (N_1523,N_1295,N_1406);
or U1524 (N_1524,N_872,N_1339);
nor U1525 (N_1525,N_670,N_48);
nor U1526 (N_1526,N_704,N_1411);
nand U1527 (N_1527,In_156,In_828);
nor U1528 (N_1528,N_1181,N_489);
nor U1529 (N_1529,In_1145,N_1192);
or U1530 (N_1530,N_1273,In_1292);
nor U1531 (N_1531,N_1420,N_1294);
nor U1532 (N_1532,N_888,In_1299);
nand U1533 (N_1533,In_1181,N_1383);
and U1534 (N_1534,N_1436,N_181);
and U1535 (N_1535,N_1272,N_1282);
nand U1536 (N_1536,In_1201,N_1159);
nand U1537 (N_1537,N_757,In_1662);
nor U1538 (N_1538,N_1327,N_137);
xnor U1539 (N_1539,N_471,N_798);
and U1540 (N_1540,N_1170,In_441);
and U1541 (N_1541,N_1316,N_1085);
and U1542 (N_1542,N_1267,In_109);
and U1543 (N_1543,N_1287,N_1090);
nor U1544 (N_1544,N_298,N_1321);
and U1545 (N_1545,N_960,N_195);
and U1546 (N_1546,N_1258,N_1393);
xor U1547 (N_1547,N_1078,N_951);
xor U1548 (N_1548,N_1303,N_1024);
nor U1549 (N_1549,In_1103,N_535);
nand U1550 (N_1550,N_1135,N_1347);
nand U1551 (N_1551,N_338,N_79);
nand U1552 (N_1552,N_915,N_1167);
and U1553 (N_1553,N_1342,In_1979);
and U1554 (N_1554,N_662,N_1177);
nor U1555 (N_1555,In_1106,N_1197);
and U1556 (N_1556,N_1236,N_984);
xnor U1557 (N_1557,N_1064,N_811);
xor U1558 (N_1558,N_1423,N_1400);
or U1559 (N_1559,N_1301,N_1003);
nor U1560 (N_1560,N_1398,In_796);
nor U1561 (N_1561,N_511,N_885);
nand U1562 (N_1562,N_799,In_398);
or U1563 (N_1563,N_1205,N_1412);
and U1564 (N_1564,N_1113,In_1956);
nand U1565 (N_1565,N_551,N_1182);
nor U1566 (N_1566,N_1313,N_1206);
nand U1567 (N_1567,N_786,N_1281);
nor U1568 (N_1568,In_76,N_1230);
xor U1569 (N_1569,N_461,N_842);
nand U1570 (N_1570,N_1002,N_964);
nand U1571 (N_1571,N_831,N_1174);
nand U1572 (N_1572,N_1395,N_1263);
or U1573 (N_1573,N_1354,N_182);
nand U1574 (N_1574,N_745,N_1432);
nand U1575 (N_1575,In_529,N_1418);
nor U1576 (N_1576,N_1011,N_703);
and U1577 (N_1577,N_824,In_69);
and U1578 (N_1578,N_1310,In_1755);
or U1579 (N_1579,N_98,N_590);
or U1580 (N_1580,N_839,N_1332);
and U1581 (N_1581,N_1243,In_1325);
xnor U1582 (N_1582,N_1145,In_224);
nor U1583 (N_1583,N_1429,N_1314);
and U1584 (N_1584,N_840,N_1351);
and U1585 (N_1585,N_1067,N_819);
and U1586 (N_1586,N_1439,In_317);
nor U1587 (N_1587,N_1416,N_1391);
nand U1588 (N_1588,N_1318,N_1410);
nor U1589 (N_1589,In_596,N_1280);
nor U1590 (N_1590,N_1430,N_876);
xnor U1591 (N_1591,N_1437,N_1357);
or U1592 (N_1592,N_777,N_1363);
or U1593 (N_1593,N_1417,N_606);
and U1594 (N_1594,N_830,N_1353);
or U1595 (N_1595,N_1157,In_1033);
or U1596 (N_1596,N_1387,In_3);
nand U1597 (N_1597,N_1204,N_1388);
nand U1598 (N_1598,N_1322,N_656);
and U1599 (N_1599,N_1298,N_1333);
nor U1600 (N_1600,N_1188,N_1560);
or U1601 (N_1601,In_135,N_1524);
and U1602 (N_1602,N_1323,N_1511);
nand U1603 (N_1603,In_1868,N_1337);
nor U1604 (N_1604,In_541,N_1311);
xnor U1605 (N_1605,N_1571,N_1448);
nand U1606 (N_1606,N_323,N_1089);
nor U1607 (N_1607,N_715,N_1562);
nand U1608 (N_1608,N_1469,N_1309);
nand U1609 (N_1609,N_1358,In_1707);
nor U1610 (N_1610,N_1445,N_1570);
and U1611 (N_1611,N_1441,N_1465);
nor U1612 (N_1612,N_24,N_433);
and U1613 (N_1613,N_1373,N_1139);
and U1614 (N_1614,N_1522,N_149);
or U1615 (N_1615,N_1450,N_1123);
nand U1616 (N_1616,N_483,N_1195);
nor U1617 (N_1617,N_976,N_1517);
and U1618 (N_1618,In_517,N_1039);
and U1619 (N_1619,In_938,N_1460);
and U1620 (N_1620,N_1211,N_1482);
and U1621 (N_1621,N_974,N_1381);
xnor U1622 (N_1622,N_1575,N_1125);
nand U1623 (N_1623,N_867,In_285);
and U1624 (N_1624,N_1402,N_1529);
and U1625 (N_1625,N_1506,N_727);
nor U1626 (N_1626,N_1451,N_1200);
nor U1627 (N_1627,N_623,N_1589);
xor U1628 (N_1628,N_1503,In_588);
and U1629 (N_1629,N_1060,N_1422);
and U1630 (N_1630,N_1285,N_1237);
or U1631 (N_1631,N_1504,N_1592);
and U1632 (N_1632,N_1455,N_1586);
nand U1633 (N_1633,N_1324,N_1545);
or U1634 (N_1634,N_1535,N_1491);
nor U1635 (N_1635,N_1435,N_1449);
nor U1636 (N_1636,N_1291,N_1173);
or U1637 (N_1637,N_1513,N_1021);
nor U1638 (N_1638,N_813,In_1067);
nor U1639 (N_1639,N_1565,N_1389);
nor U1640 (N_1640,N_1331,In_1226);
and U1641 (N_1641,N_1497,N_1519);
or U1642 (N_1642,N_1290,N_1574);
or U1643 (N_1643,N_1599,In_1664);
xnor U1644 (N_1644,N_1365,N_1134);
nor U1645 (N_1645,N_1099,In_917);
and U1646 (N_1646,N_1472,N_32);
and U1647 (N_1647,N_1292,N_1550);
nor U1648 (N_1648,N_1591,N_1231);
xnor U1649 (N_1649,N_1578,N_464);
nor U1650 (N_1650,N_1556,N_846);
and U1651 (N_1651,N_1092,N_1364);
xor U1652 (N_1652,N_1598,N_1582);
nor U1653 (N_1653,N_1555,N_1168);
nand U1654 (N_1654,N_1478,N_1573);
nand U1655 (N_1655,N_1493,N_869);
nor U1656 (N_1656,N_322,N_1490);
and U1657 (N_1657,N_1444,In_1322);
nor U1658 (N_1658,N_1521,N_347);
nand U1659 (N_1659,N_1483,N_996);
or U1660 (N_1660,N_1136,In_622);
nand U1661 (N_1661,N_1492,In_1983);
nand U1662 (N_1662,N_1452,N_1084);
or U1663 (N_1663,N_672,N_1588);
nor U1664 (N_1664,N_1158,N_1425);
nand U1665 (N_1665,N_1154,In_1283);
nand U1666 (N_1666,In_89,N_1061);
or U1667 (N_1667,N_1104,N_1050);
or U1668 (N_1668,In_1001,N_1583);
nand U1669 (N_1669,N_1421,N_1462);
and U1670 (N_1670,In_365,N_1350);
nor U1671 (N_1671,In_1679,N_1247);
nand U1672 (N_1672,N_1477,N_1307);
nor U1673 (N_1673,N_683,N_1279);
nand U1674 (N_1674,N_981,N_1433);
nor U1675 (N_1675,N_741,N_1014);
and U1676 (N_1676,N_1499,N_1293);
nand U1677 (N_1677,N_558,N_1505);
and U1678 (N_1678,N_1580,N_1541);
and U1679 (N_1679,N_751,In_1846);
xnor U1680 (N_1680,N_436,N_1488);
nand U1681 (N_1681,N_836,N_1554);
and U1682 (N_1682,N_1369,In_634);
nor U1683 (N_1683,N_1141,N_1222);
xnor U1684 (N_1684,N_1501,N_1563);
and U1685 (N_1685,N_1277,In_1028);
and U1686 (N_1686,N_481,N_1496);
and U1687 (N_1687,N_1456,N_932);
and U1688 (N_1688,N_1549,N_1471);
nand U1689 (N_1689,N_1194,N_1468);
nand U1690 (N_1690,N_1149,N_1464);
nor U1691 (N_1691,N_1346,N_825);
xnor U1692 (N_1692,N_1502,N_214);
or U1693 (N_1693,In_749,N_1304);
xor U1694 (N_1694,N_1548,N_1048);
or U1695 (N_1695,N_818,N_1442);
nand U1696 (N_1696,N_1037,N_1543);
nand U1697 (N_1697,N_1596,N_1484);
or U1698 (N_1698,N_1523,N_883);
or U1699 (N_1699,N_1526,N_1525);
and U1700 (N_1700,In_991,N_807);
and U1701 (N_1701,N_1386,N_1446);
nor U1702 (N_1702,N_1551,N_940);
nand U1703 (N_1703,In_1309,N_1485);
nand U1704 (N_1704,N_1049,N_1567);
or U1705 (N_1705,N_1584,In_1266);
nand U1706 (N_1706,In_1022,N_938);
or U1707 (N_1707,N_795,N_762);
or U1708 (N_1708,N_793,N_1308);
nor U1709 (N_1709,N_1537,N_1597);
nand U1710 (N_1710,N_1414,N_955);
nand U1711 (N_1711,N_1510,N_1334);
xor U1712 (N_1712,N_477,N_1229);
nand U1713 (N_1713,In_153,N_1325);
or U1714 (N_1714,N_1475,N_1508);
or U1715 (N_1715,In_1610,N_719);
nand U1716 (N_1716,N_1221,N_1512);
nor U1717 (N_1717,N_919,N_1536);
nor U1718 (N_1718,N_1520,N_1495);
xnor U1719 (N_1719,N_1538,N_1553);
and U1720 (N_1720,N_993,N_1345);
and U1721 (N_1721,N_1461,N_1564);
nand U1722 (N_1722,N_1542,N_1585);
and U1723 (N_1723,N_388,N_971);
or U1724 (N_1724,N_1516,N_997);
nor U1725 (N_1725,N_1527,N_1283);
nand U1726 (N_1726,N_1045,N_645);
nor U1727 (N_1727,N_1288,N_897);
nand U1728 (N_1728,N_1189,N_1539);
xnor U1729 (N_1729,N_1487,In_1114);
nor U1730 (N_1730,N_1489,N_1128);
nand U1731 (N_1731,N_1207,N_603);
xor U1732 (N_1732,N_260,N_1447);
nand U1733 (N_1733,N_1587,N_1396);
and U1734 (N_1734,N_1544,N_878);
or U1735 (N_1735,N_1319,N_1509);
xor U1736 (N_1736,N_1407,N_647);
and U1737 (N_1737,N_1008,N_160);
nor U1738 (N_1738,N_1284,N_970);
or U1739 (N_1739,In_251,N_843);
or U1740 (N_1740,In_1728,N_1561);
xor U1741 (N_1741,N_1559,N_999);
nor U1742 (N_1742,In_785,N_1458);
xor U1743 (N_1743,N_1479,N_1428);
or U1744 (N_1744,N_1390,N_1514);
or U1745 (N_1745,In_1148,N_1355);
nor U1746 (N_1746,N_1385,N_423);
nor U1747 (N_1747,N_1594,N_1568);
nor U1748 (N_1748,N_1228,N_1528);
and U1749 (N_1749,N_1486,N_1225);
nand U1750 (N_1750,N_789,N_712);
and U1751 (N_1751,N_1397,N_1440);
and U1752 (N_1752,N_1069,N_1558);
or U1753 (N_1753,N_923,In_1805);
nor U1754 (N_1754,N_1196,N_1030);
and U1755 (N_1755,N_517,N_1546);
nor U1756 (N_1756,N_637,N_1155);
nor U1757 (N_1757,N_1473,N_1380);
xnor U1758 (N_1758,N_1454,N_771);
nor U1759 (N_1759,N_1269,In_97);
nor U1760 (N_1760,N_1651,N_1672);
nor U1761 (N_1761,N_1624,N_1518);
nand U1762 (N_1762,N_1701,N_1615);
nand U1763 (N_1763,N_854,N_1679);
and U1764 (N_1764,N_1632,N_1605);
or U1765 (N_1765,N_348,N_1718);
nor U1766 (N_1766,N_1692,N_1653);
nand U1767 (N_1767,N_1700,N_1547);
or U1768 (N_1768,N_1498,N_1712);
xor U1769 (N_1769,N_1663,N_1611);
or U1770 (N_1770,N_144,N_1719);
or U1771 (N_1771,N_1674,N_1757);
nand U1772 (N_1772,N_1639,N_1566);
nand U1773 (N_1773,N_1733,N_1515);
nor U1774 (N_1774,N_1730,N_890);
and U1775 (N_1775,N_1691,N_1443);
nor U1776 (N_1776,N_1695,N_1645);
nor U1777 (N_1777,N_1646,In_1522);
nor U1778 (N_1778,N_1626,N_1657);
nand U1779 (N_1779,N_1647,N_1740);
or U1780 (N_1780,N_1572,N_1638);
xnor U1781 (N_1781,N_1621,N_1552);
and U1782 (N_1782,N_1658,N_1661);
or U1783 (N_1783,N_1713,N_1736);
nand U1784 (N_1784,N_1481,N_1737);
nand U1785 (N_1785,N_1680,N_1577);
nor U1786 (N_1786,N_1453,In_234);
nand U1787 (N_1787,N_1637,N_1748);
nand U1788 (N_1788,N_1751,N_1531);
or U1789 (N_1789,N_1727,N_1494);
and U1790 (N_1790,N_1619,N_1540);
xnor U1791 (N_1791,N_1728,N_1620);
xor U1792 (N_1792,N_1636,N_1606);
nand U1793 (N_1793,N_958,N_1187);
and U1794 (N_1794,N_1530,N_1603);
nand U1795 (N_1795,N_1709,N_1557);
nor U1796 (N_1796,N_1532,In_564);
nand U1797 (N_1797,N_1629,N_1649);
and U1798 (N_1798,N_1699,N_1742);
nor U1799 (N_1799,N_1724,N_1617);
or U1800 (N_1800,N_1297,N_1660);
nor U1801 (N_1801,N_318,N_1533);
nor U1802 (N_1802,N_1648,N_1725);
xnor U1803 (N_1803,N_1689,N_1627);
and U1804 (N_1804,N_1379,N_1507);
nor U1805 (N_1805,N_1470,N_1688);
nor U1806 (N_1806,N_1459,N_1749);
and U1807 (N_1807,N_1669,N_1595);
and U1808 (N_1808,N_1642,N_1392);
or U1809 (N_1809,N_396,N_1635);
or U1810 (N_1810,In_143,N_1690);
and U1811 (N_1811,N_1593,N_1656);
nand U1812 (N_1812,N_1731,N_1404);
xor U1813 (N_1813,N_1576,N_1618);
and U1814 (N_1814,N_1745,N_1683);
xnor U1815 (N_1815,N_508,N_1675);
and U1816 (N_1816,N_1682,N_1650);
xnor U1817 (N_1817,N_1581,N_1750);
nor U1818 (N_1818,N_1467,N_1305);
or U1819 (N_1819,N_362,N_1655);
or U1820 (N_1820,N_1667,N_1608);
and U1821 (N_1821,N_1744,N_1625);
nand U1822 (N_1822,N_1609,N_1630);
nand U1823 (N_1823,N_1466,N_1659);
nand U1824 (N_1824,N_1678,N_1614);
or U1825 (N_1825,N_1569,N_1706);
nor U1826 (N_1826,N_1747,N_1631);
xor U1827 (N_1827,N_1457,N_1604);
nor U1828 (N_1828,N_1721,N_1634);
and U1829 (N_1829,N_907,N_1710);
or U1830 (N_1830,N_1697,N_1476);
or U1831 (N_1831,N_1107,N_1601);
nor U1832 (N_1832,N_1622,N_1590);
nand U1833 (N_1833,N_1668,N_1716);
nand U1834 (N_1834,N_1058,N_1378);
nor U1835 (N_1835,N_1756,N_1752);
and U1836 (N_1836,N_1746,N_1628);
or U1837 (N_1837,In_738,N_1394);
nor U1838 (N_1838,N_1743,N_1681);
nand U1839 (N_1839,N_1705,N_1670);
nor U1840 (N_1840,N_1600,N_1687);
nand U1841 (N_1841,N_695,In_542);
and U1842 (N_1842,N_1120,N_1722);
nand U1843 (N_1843,N_1696,N_1707);
or U1844 (N_1844,N_1317,N_1366);
nand U1845 (N_1845,N_1720,N_1693);
and U1846 (N_1846,N_1732,N_1644);
nand U1847 (N_1847,N_1607,N_1734);
nor U1848 (N_1848,N_1677,N_1703);
xor U1849 (N_1849,N_1463,N_1474);
and U1850 (N_1850,N_1534,N_1612);
or U1851 (N_1851,N_1729,N_126);
and U1852 (N_1852,N_1723,N_1755);
nand U1853 (N_1853,N_1643,N_1299);
or U1854 (N_1854,N_1704,N_1684);
xnor U1855 (N_1855,In_882,N_1686);
or U1856 (N_1856,N_1673,In_793);
nor U1857 (N_1857,N_1702,N_1244);
nand U1858 (N_1858,N_1662,N_1711);
nand U1859 (N_1859,N_1738,N_1685);
xor U1860 (N_1860,N_1633,N_1715);
and U1861 (N_1861,N_1616,N_1739);
nor U1862 (N_1862,N_1671,N_1579);
nor U1863 (N_1863,N_1664,N_1623);
nand U1864 (N_1864,N_1741,N_1694);
nand U1865 (N_1865,N_1759,N_1735);
xnor U1866 (N_1866,N_1602,N_1500);
and U1867 (N_1867,N_475,N_1320);
nor U1868 (N_1868,N_1758,N_1652);
nor U1869 (N_1869,N_507,N_1640);
xnor U1870 (N_1870,In_716,N_1754);
nor U1871 (N_1871,N_1717,N_1226);
and U1872 (N_1872,N_1091,N_1480);
nand U1873 (N_1873,N_1613,N_1714);
or U1874 (N_1874,N_1708,N_1753);
and U1875 (N_1875,N_1676,N_1329);
and U1876 (N_1876,N_1641,N_1666);
or U1877 (N_1877,N_1698,N_1654);
and U1878 (N_1878,N_1665,N_1726);
or U1879 (N_1879,N_1610,N_1306);
and U1880 (N_1880,In_882,N_126);
and U1881 (N_1881,N_1707,N_1748);
nor U1882 (N_1882,N_1605,N_1726);
nor U1883 (N_1883,N_1656,N_1746);
nor U1884 (N_1884,N_1655,N_1507);
nor U1885 (N_1885,N_1605,N_1714);
and U1886 (N_1886,N_1692,N_1729);
or U1887 (N_1887,N_1569,N_1682);
xnor U1888 (N_1888,N_1752,N_1625);
nand U1889 (N_1889,N_1576,N_1306);
or U1890 (N_1890,N_1532,N_1602);
xor U1891 (N_1891,N_1715,N_1651);
nand U1892 (N_1892,N_1107,In_234);
and U1893 (N_1893,N_1683,N_1457);
nor U1894 (N_1894,N_1742,In_716);
xor U1895 (N_1895,N_1320,N_1607);
nand U1896 (N_1896,N_1617,N_1620);
xor U1897 (N_1897,N_508,N_318);
nor U1898 (N_1898,N_1737,N_1706);
or U1899 (N_1899,In_1522,N_1755);
and U1900 (N_1900,N_1616,N_1602);
xor U1901 (N_1901,N_1692,N_1645);
nand U1902 (N_1902,N_1610,N_1633);
nand U1903 (N_1903,N_1682,N_1476);
or U1904 (N_1904,N_1533,N_475);
and U1905 (N_1905,N_1659,N_1681);
or U1906 (N_1906,N_1680,N_1654);
and U1907 (N_1907,N_1673,N_1317);
or U1908 (N_1908,N_854,N_144);
nor U1909 (N_1909,N_1716,N_1673);
and U1910 (N_1910,N_1533,N_1662);
and U1911 (N_1911,N_1715,N_1647);
nand U1912 (N_1912,N_1091,N_1661);
or U1913 (N_1913,N_1630,N_1606);
or U1914 (N_1914,N_1518,N_1470);
and U1915 (N_1915,N_1656,N_1750);
xor U1916 (N_1916,N_1621,N_1727);
and U1917 (N_1917,N_1641,N_1320);
nand U1918 (N_1918,N_1642,N_1320);
nand U1919 (N_1919,N_1605,N_1518);
nand U1920 (N_1920,N_1916,N_1874);
nand U1921 (N_1921,N_1849,N_1845);
and U1922 (N_1922,N_1778,N_1832);
and U1923 (N_1923,N_1908,N_1860);
or U1924 (N_1924,N_1790,N_1876);
nand U1925 (N_1925,N_1906,N_1890);
nor U1926 (N_1926,N_1838,N_1883);
nor U1927 (N_1927,N_1850,N_1896);
or U1928 (N_1928,N_1801,N_1810);
or U1929 (N_1929,N_1885,N_1809);
or U1930 (N_1930,N_1872,N_1770);
nand U1931 (N_1931,N_1786,N_1884);
nor U1932 (N_1932,N_1780,N_1904);
nor U1933 (N_1933,N_1829,N_1805);
nor U1934 (N_1934,N_1917,N_1888);
and U1935 (N_1935,N_1919,N_1867);
and U1936 (N_1936,N_1865,N_1882);
and U1937 (N_1937,N_1763,N_1783);
nand U1938 (N_1938,N_1762,N_1858);
nand U1939 (N_1939,N_1913,N_1843);
or U1940 (N_1940,N_1837,N_1821);
nor U1941 (N_1941,N_1866,N_1902);
nor U1942 (N_1942,N_1879,N_1828);
or U1943 (N_1943,N_1765,N_1803);
xnor U1944 (N_1944,N_1835,N_1825);
nand U1945 (N_1945,N_1871,N_1855);
nor U1946 (N_1946,N_1862,N_1831);
nor U1947 (N_1947,N_1771,N_1901);
nor U1948 (N_1948,N_1889,N_1859);
nor U1949 (N_1949,N_1905,N_1877);
xnor U1950 (N_1950,N_1861,N_1903);
nand U1951 (N_1951,N_1851,N_1784);
nor U1952 (N_1952,N_1873,N_1820);
or U1953 (N_1953,N_1819,N_1769);
nand U1954 (N_1954,N_1775,N_1918);
nand U1955 (N_1955,N_1785,N_1823);
and U1956 (N_1956,N_1791,N_1764);
and U1957 (N_1957,N_1800,N_1878);
nor U1958 (N_1958,N_1774,N_1782);
and U1959 (N_1959,N_1911,N_1847);
nand U1960 (N_1960,N_1909,N_1779);
and U1961 (N_1961,N_1907,N_1836);
nor U1962 (N_1962,N_1893,N_1793);
xnor U1963 (N_1963,N_1814,N_1864);
and U1964 (N_1964,N_1772,N_1834);
or U1965 (N_1965,N_1813,N_1797);
and U1966 (N_1966,N_1806,N_1846);
nand U1967 (N_1967,N_1799,N_1811);
or U1968 (N_1968,N_1760,N_1854);
nor U1969 (N_1969,N_1768,N_1856);
xor U1970 (N_1970,N_1776,N_1766);
nor U1971 (N_1971,N_1857,N_1826);
nand U1972 (N_1972,N_1841,N_1898);
or U1973 (N_1973,N_1899,N_1787);
or U1974 (N_1974,N_1794,N_1875);
or U1975 (N_1975,N_1816,N_1912);
nor U1976 (N_1976,N_1822,N_1777);
nor U1977 (N_1977,N_1914,N_1830);
nand U1978 (N_1978,N_1798,N_1870);
xor U1979 (N_1979,N_1804,N_1812);
and U1980 (N_1980,N_1773,N_1792);
nand U1981 (N_1981,N_1895,N_1795);
or U1982 (N_1982,N_1887,N_1852);
nand U1983 (N_1983,N_1767,N_1880);
and U1984 (N_1984,N_1891,N_1808);
and U1985 (N_1985,N_1827,N_1815);
nor U1986 (N_1986,N_1900,N_1892);
or U1987 (N_1987,N_1842,N_1863);
or U1988 (N_1988,N_1789,N_1796);
xnor U1989 (N_1989,N_1781,N_1761);
nor U1990 (N_1990,N_1807,N_1824);
nor U1991 (N_1991,N_1833,N_1844);
and U1992 (N_1992,N_1881,N_1869);
xor U1993 (N_1993,N_1802,N_1853);
or U1994 (N_1994,N_1848,N_1894);
and U1995 (N_1995,N_1839,N_1897);
xnor U1996 (N_1996,N_1818,N_1886);
or U1997 (N_1997,N_1910,N_1868);
and U1998 (N_1998,N_1840,N_1817);
nor U1999 (N_1999,N_1915,N_1788);
xor U2000 (N_2000,N_1794,N_1899);
nand U2001 (N_2001,N_1822,N_1788);
and U2002 (N_2002,N_1857,N_1849);
or U2003 (N_2003,N_1822,N_1845);
nor U2004 (N_2004,N_1901,N_1887);
and U2005 (N_2005,N_1881,N_1840);
xnor U2006 (N_2006,N_1838,N_1891);
nor U2007 (N_2007,N_1893,N_1816);
and U2008 (N_2008,N_1885,N_1830);
nor U2009 (N_2009,N_1778,N_1919);
or U2010 (N_2010,N_1788,N_1807);
or U2011 (N_2011,N_1892,N_1887);
and U2012 (N_2012,N_1900,N_1852);
nor U2013 (N_2013,N_1868,N_1806);
nor U2014 (N_2014,N_1820,N_1911);
xnor U2015 (N_2015,N_1872,N_1806);
xor U2016 (N_2016,N_1788,N_1767);
xor U2017 (N_2017,N_1839,N_1859);
or U2018 (N_2018,N_1859,N_1760);
or U2019 (N_2019,N_1912,N_1842);
nand U2020 (N_2020,N_1861,N_1790);
nand U2021 (N_2021,N_1791,N_1877);
and U2022 (N_2022,N_1872,N_1843);
or U2023 (N_2023,N_1805,N_1775);
nand U2024 (N_2024,N_1882,N_1897);
xor U2025 (N_2025,N_1788,N_1825);
and U2026 (N_2026,N_1852,N_1834);
nand U2027 (N_2027,N_1816,N_1913);
xnor U2028 (N_2028,N_1800,N_1863);
or U2029 (N_2029,N_1829,N_1818);
and U2030 (N_2030,N_1859,N_1853);
nor U2031 (N_2031,N_1840,N_1880);
or U2032 (N_2032,N_1910,N_1830);
or U2033 (N_2033,N_1873,N_1823);
nand U2034 (N_2034,N_1910,N_1912);
xnor U2035 (N_2035,N_1778,N_1859);
nor U2036 (N_2036,N_1858,N_1912);
nor U2037 (N_2037,N_1869,N_1844);
nand U2038 (N_2038,N_1810,N_1829);
nor U2039 (N_2039,N_1898,N_1844);
and U2040 (N_2040,N_1827,N_1839);
nand U2041 (N_2041,N_1894,N_1821);
nand U2042 (N_2042,N_1878,N_1768);
or U2043 (N_2043,N_1775,N_1780);
nor U2044 (N_2044,N_1841,N_1849);
nor U2045 (N_2045,N_1866,N_1807);
or U2046 (N_2046,N_1797,N_1849);
nand U2047 (N_2047,N_1794,N_1863);
nand U2048 (N_2048,N_1836,N_1840);
nand U2049 (N_2049,N_1780,N_1888);
xor U2050 (N_2050,N_1815,N_1764);
nand U2051 (N_2051,N_1875,N_1867);
and U2052 (N_2052,N_1773,N_1787);
xor U2053 (N_2053,N_1765,N_1805);
nand U2054 (N_2054,N_1866,N_1786);
xor U2055 (N_2055,N_1818,N_1880);
and U2056 (N_2056,N_1867,N_1786);
nor U2057 (N_2057,N_1781,N_1794);
and U2058 (N_2058,N_1839,N_1843);
xnor U2059 (N_2059,N_1873,N_1829);
or U2060 (N_2060,N_1881,N_1795);
and U2061 (N_2061,N_1767,N_1815);
nor U2062 (N_2062,N_1776,N_1800);
and U2063 (N_2063,N_1770,N_1884);
nand U2064 (N_2064,N_1879,N_1823);
nand U2065 (N_2065,N_1765,N_1777);
nor U2066 (N_2066,N_1800,N_1837);
xnor U2067 (N_2067,N_1894,N_1803);
nor U2068 (N_2068,N_1892,N_1819);
nor U2069 (N_2069,N_1784,N_1892);
xnor U2070 (N_2070,N_1805,N_1889);
nor U2071 (N_2071,N_1894,N_1842);
and U2072 (N_2072,N_1816,N_1856);
or U2073 (N_2073,N_1875,N_1863);
or U2074 (N_2074,N_1849,N_1855);
or U2075 (N_2075,N_1901,N_1795);
or U2076 (N_2076,N_1785,N_1766);
or U2077 (N_2077,N_1788,N_1823);
nor U2078 (N_2078,N_1770,N_1781);
or U2079 (N_2079,N_1894,N_1891);
nor U2080 (N_2080,N_2055,N_2019);
or U2081 (N_2081,N_2002,N_2066);
nor U2082 (N_2082,N_1928,N_1984);
and U2083 (N_2083,N_1952,N_2021);
nand U2084 (N_2084,N_2007,N_1982);
nor U2085 (N_2085,N_1948,N_1976);
nand U2086 (N_2086,N_2011,N_1967);
nand U2087 (N_2087,N_1995,N_1961);
nor U2088 (N_2088,N_2067,N_1968);
and U2089 (N_2089,N_1947,N_2005);
or U2090 (N_2090,N_1973,N_2076);
or U2091 (N_2091,N_1991,N_1970);
and U2092 (N_2092,N_2023,N_2030);
nor U2093 (N_2093,N_2042,N_2008);
nand U2094 (N_2094,N_2041,N_1944);
nor U2095 (N_2095,N_2012,N_1939);
xor U2096 (N_2096,N_2026,N_2040);
nand U2097 (N_2097,N_1953,N_1972);
nor U2098 (N_2098,N_1931,N_1974);
nand U2099 (N_2099,N_2025,N_2001);
nor U2100 (N_2100,N_1927,N_1997);
nand U2101 (N_2101,N_1996,N_1942);
nor U2102 (N_2102,N_2075,N_1966);
xor U2103 (N_2103,N_2061,N_1987);
nor U2104 (N_2104,N_1988,N_1920);
or U2105 (N_2105,N_1922,N_2064);
nor U2106 (N_2106,N_1955,N_1975);
and U2107 (N_2107,N_2060,N_1949);
nor U2108 (N_2108,N_2078,N_2053);
or U2109 (N_2109,N_1945,N_1921);
and U2110 (N_2110,N_2070,N_1999);
nand U2111 (N_2111,N_2014,N_2054);
nand U2112 (N_2112,N_2047,N_2029);
and U2113 (N_2113,N_2079,N_2032);
and U2114 (N_2114,N_2015,N_2057);
and U2115 (N_2115,N_1941,N_1924);
and U2116 (N_2116,N_1986,N_1960);
nor U2117 (N_2117,N_2036,N_2000);
xnor U2118 (N_2118,N_2038,N_2044);
or U2119 (N_2119,N_2059,N_2065);
and U2120 (N_2120,N_1940,N_1978);
nor U2121 (N_2121,N_1990,N_2051);
or U2122 (N_2122,N_1933,N_1925);
or U2123 (N_2123,N_2033,N_1958);
or U2124 (N_2124,N_2052,N_1923);
nor U2125 (N_2125,N_2056,N_2073);
xnor U2126 (N_2126,N_2024,N_2072);
nand U2127 (N_2127,N_1956,N_1929);
or U2128 (N_2128,N_2020,N_1964);
nand U2129 (N_2129,N_1957,N_2074);
nand U2130 (N_2130,N_1926,N_1937);
or U2131 (N_2131,N_2037,N_2068);
nor U2132 (N_2132,N_1983,N_2063);
nor U2133 (N_2133,N_1963,N_2035);
xor U2134 (N_2134,N_1989,N_2043);
xor U2135 (N_2135,N_1992,N_2016);
or U2136 (N_2136,N_1950,N_1932);
nand U2137 (N_2137,N_2010,N_2069);
and U2138 (N_2138,N_2028,N_1930);
nand U2139 (N_2139,N_2058,N_2004);
nor U2140 (N_2140,N_2013,N_2009);
nand U2141 (N_2141,N_1935,N_2027);
nand U2142 (N_2142,N_2046,N_1938);
or U2143 (N_2143,N_1943,N_1981);
and U2144 (N_2144,N_2006,N_2045);
nor U2145 (N_2145,N_1934,N_1969);
nor U2146 (N_2146,N_2050,N_2039);
or U2147 (N_2147,N_1994,N_1993);
or U2148 (N_2148,N_1965,N_2017);
xor U2149 (N_2149,N_1977,N_1980);
or U2150 (N_2150,N_1946,N_1962);
or U2151 (N_2151,N_1985,N_1951);
nor U2152 (N_2152,N_2003,N_2031);
nand U2153 (N_2153,N_1959,N_1954);
and U2154 (N_2154,N_1998,N_1971);
nor U2155 (N_2155,N_2048,N_1936);
and U2156 (N_2156,N_1979,N_2077);
nand U2157 (N_2157,N_2049,N_2018);
xnor U2158 (N_2158,N_2022,N_2034);
or U2159 (N_2159,N_2062,N_2071);
or U2160 (N_2160,N_1946,N_2018);
nor U2161 (N_2161,N_1974,N_1952);
nand U2162 (N_2162,N_2061,N_2039);
nor U2163 (N_2163,N_2063,N_2039);
nor U2164 (N_2164,N_1957,N_1999);
and U2165 (N_2165,N_1928,N_1976);
or U2166 (N_2166,N_1920,N_2051);
or U2167 (N_2167,N_2020,N_2061);
nand U2168 (N_2168,N_1992,N_2042);
nor U2169 (N_2169,N_1920,N_2075);
nor U2170 (N_2170,N_1976,N_2058);
or U2171 (N_2171,N_1978,N_1988);
nor U2172 (N_2172,N_2050,N_1982);
nor U2173 (N_2173,N_1976,N_1975);
nand U2174 (N_2174,N_1931,N_1935);
and U2175 (N_2175,N_2072,N_2009);
and U2176 (N_2176,N_2007,N_1937);
nor U2177 (N_2177,N_1923,N_1984);
nor U2178 (N_2178,N_1981,N_2036);
nor U2179 (N_2179,N_2051,N_1994);
and U2180 (N_2180,N_2008,N_1995);
nor U2181 (N_2181,N_2001,N_2047);
xor U2182 (N_2182,N_1924,N_2024);
or U2183 (N_2183,N_2047,N_2042);
or U2184 (N_2184,N_2052,N_1960);
nand U2185 (N_2185,N_2078,N_1942);
or U2186 (N_2186,N_2057,N_1956);
nor U2187 (N_2187,N_1958,N_1971);
or U2188 (N_2188,N_1955,N_2035);
and U2189 (N_2189,N_2013,N_1932);
nand U2190 (N_2190,N_2021,N_2070);
nand U2191 (N_2191,N_2009,N_1977);
and U2192 (N_2192,N_2061,N_2058);
nor U2193 (N_2193,N_1949,N_1930);
and U2194 (N_2194,N_1941,N_1955);
nand U2195 (N_2195,N_1931,N_2054);
nor U2196 (N_2196,N_2049,N_1970);
and U2197 (N_2197,N_1971,N_1947);
nor U2198 (N_2198,N_1934,N_1977);
and U2199 (N_2199,N_1932,N_1928);
nand U2200 (N_2200,N_1939,N_2004);
xor U2201 (N_2201,N_1975,N_2017);
xnor U2202 (N_2202,N_2068,N_1972);
xor U2203 (N_2203,N_1977,N_1989);
nor U2204 (N_2204,N_1982,N_2078);
nand U2205 (N_2205,N_2072,N_2002);
and U2206 (N_2206,N_2062,N_1925);
and U2207 (N_2207,N_1931,N_1948);
nor U2208 (N_2208,N_2075,N_1982);
and U2209 (N_2209,N_1973,N_1999);
and U2210 (N_2210,N_1986,N_2079);
or U2211 (N_2211,N_1929,N_1941);
xnor U2212 (N_2212,N_1994,N_2063);
nor U2213 (N_2213,N_1947,N_2047);
or U2214 (N_2214,N_1946,N_2045);
nand U2215 (N_2215,N_1990,N_1976);
nand U2216 (N_2216,N_1996,N_1997);
nand U2217 (N_2217,N_2008,N_2048);
and U2218 (N_2218,N_2023,N_1996);
nand U2219 (N_2219,N_2071,N_2001);
or U2220 (N_2220,N_2068,N_1970);
nor U2221 (N_2221,N_1923,N_1927);
nand U2222 (N_2222,N_1984,N_2075);
nand U2223 (N_2223,N_1964,N_2048);
and U2224 (N_2224,N_2014,N_1954);
xor U2225 (N_2225,N_2039,N_1995);
and U2226 (N_2226,N_2016,N_2005);
or U2227 (N_2227,N_2040,N_1950);
or U2228 (N_2228,N_2019,N_1996);
nor U2229 (N_2229,N_1977,N_2052);
and U2230 (N_2230,N_2048,N_1992);
nor U2231 (N_2231,N_2024,N_2077);
and U2232 (N_2232,N_2023,N_2025);
and U2233 (N_2233,N_1990,N_1955);
or U2234 (N_2234,N_1952,N_1953);
nor U2235 (N_2235,N_2049,N_1996);
xnor U2236 (N_2236,N_2069,N_2062);
or U2237 (N_2237,N_2032,N_1925);
or U2238 (N_2238,N_2022,N_1984);
nor U2239 (N_2239,N_1929,N_2048);
or U2240 (N_2240,N_2234,N_2220);
nor U2241 (N_2241,N_2210,N_2090);
nor U2242 (N_2242,N_2116,N_2228);
and U2243 (N_2243,N_2157,N_2097);
nand U2244 (N_2244,N_2204,N_2185);
nor U2245 (N_2245,N_2232,N_2093);
or U2246 (N_2246,N_2155,N_2239);
nor U2247 (N_2247,N_2181,N_2126);
xnor U2248 (N_2248,N_2151,N_2190);
or U2249 (N_2249,N_2131,N_2182);
or U2250 (N_2250,N_2225,N_2132);
nor U2251 (N_2251,N_2160,N_2121);
or U2252 (N_2252,N_2146,N_2209);
nand U2253 (N_2253,N_2180,N_2148);
or U2254 (N_2254,N_2211,N_2149);
nand U2255 (N_2255,N_2134,N_2125);
xnor U2256 (N_2256,N_2189,N_2138);
and U2257 (N_2257,N_2178,N_2224);
and U2258 (N_2258,N_2222,N_2122);
and U2259 (N_2259,N_2082,N_2176);
nor U2260 (N_2260,N_2144,N_2111);
and U2261 (N_2261,N_2092,N_2199);
nor U2262 (N_2262,N_2161,N_2215);
and U2263 (N_2263,N_2153,N_2127);
and U2264 (N_2264,N_2172,N_2229);
or U2265 (N_2265,N_2103,N_2231);
nand U2266 (N_2266,N_2113,N_2163);
xor U2267 (N_2267,N_2091,N_2080);
and U2268 (N_2268,N_2100,N_2164);
nand U2269 (N_2269,N_2105,N_2133);
or U2270 (N_2270,N_2217,N_2142);
nor U2271 (N_2271,N_2193,N_2118);
and U2272 (N_2272,N_2086,N_2084);
nor U2273 (N_2273,N_2154,N_2117);
nand U2274 (N_2274,N_2129,N_2089);
nor U2275 (N_2275,N_2227,N_2085);
nand U2276 (N_2276,N_2198,N_2194);
nand U2277 (N_2277,N_2088,N_2177);
nor U2278 (N_2278,N_2166,N_2192);
nand U2279 (N_2279,N_2207,N_2120);
and U2280 (N_2280,N_2159,N_2099);
and U2281 (N_2281,N_2141,N_2137);
and U2282 (N_2282,N_2112,N_2179);
and U2283 (N_2283,N_2104,N_2094);
xnor U2284 (N_2284,N_2226,N_2223);
nor U2285 (N_2285,N_2200,N_2081);
nand U2286 (N_2286,N_2098,N_2119);
nand U2287 (N_2287,N_2124,N_2167);
nor U2288 (N_2288,N_2087,N_2102);
nor U2289 (N_2289,N_2165,N_2216);
and U2290 (N_2290,N_2196,N_2237);
xnor U2291 (N_2291,N_2213,N_2173);
or U2292 (N_2292,N_2096,N_2123);
nand U2293 (N_2293,N_2109,N_2147);
nor U2294 (N_2294,N_2107,N_2230);
nor U2295 (N_2295,N_2171,N_2203);
xnor U2296 (N_2296,N_2083,N_2197);
and U2297 (N_2297,N_2191,N_2170);
nor U2298 (N_2298,N_2136,N_2233);
nand U2299 (N_2299,N_2158,N_2114);
nand U2300 (N_2300,N_2168,N_2152);
nor U2301 (N_2301,N_2184,N_2235);
nand U2302 (N_2302,N_2169,N_2106);
nand U2303 (N_2303,N_2188,N_2101);
nand U2304 (N_2304,N_2202,N_2110);
nor U2305 (N_2305,N_2175,N_2206);
nand U2306 (N_2306,N_2139,N_2221);
or U2307 (N_2307,N_2186,N_2183);
nand U2308 (N_2308,N_2205,N_2219);
nor U2309 (N_2309,N_2135,N_2201);
or U2310 (N_2310,N_2140,N_2208);
nand U2311 (N_2311,N_2174,N_2115);
nand U2312 (N_2312,N_2095,N_2130);
or U2313 (N_2313,N_2145,N_2108);
nand U2314 (N_2314,N_2218,N_2238);
nor U2315 (N_2315,N_2150,N_2195);
xor U2316 (N_2316,N_2187,N_2212);
nand U2317 (N_2317,N_2128,N_2214);
or U2318 (N_2318,N_2236,N_2143);
or U2319 (N_2319,N_2162,N_2156);
nand U2320 (N_2320,N_2165,N_2114);
nand U2321 (N_2321,N_2210,N_2087);
xor U2322 (N_2322,N_2125,N_2160);
or U2323 (N_2323,N_2206,N_2188);
and U2324 (N_2324,N_2085,N_2136);
nor U2325 (N_2325,N_2212,N_2213);
nand U2326 (N_2326,N_2082,N_2134);
nor U2327 (N_2327,N_2230,N_2208);
or U2328 (N_2328,N_2187,N_2100);
and U2329 (N_2329,N_2190,N_2150);
or U2330 (N_2330,N_2174,N_2184);
nor U2331 (N_2331,N_2090,N_2140);
nor U2332 (N_2332,N_2142,N_2160);
nor U2333 (N_2333,N_2139,N_2230);
and U2334 (N_2334,N_2162,N_2088);
nor U2335 (N_2335,N_2191,N_2172);
and U2336 (N_2336,N_2096,N_2187);
nand U2337 (N_2337,N_2186,N_2239);
and U2338 (N_2338,N_2092,N_2138);
nand U2339 (N_2339,N_2200,N_2163);
nand U2340 (N_2340,N_2208,N_2109);
and U2341 (N_2341,N_2148,N_2094);
nand U2342 (N_2342,N_2112,N_2084);
and U2343 (N_2343,N_2128,N_2127);
or U2344 (N_2344,N_2136,N_2082);
nand U2345 (N_2345,N_2087,N_2130);
nand U2346 (N_2346,N_2169,N_2154);
nand U2347 (N_2347,N_2165,N_2179);
and U2348 (N_2348,N_2235,N_2166);
and U2349 (N_2349,N_2089,N_2148);
xor U2350 (N_2350,N_2205,N_2232);
nand U2351 (N_2351,N_2115,N_2229);
or U2352 (N_2352,N_2165,N_2196);
nor U2353 (N_2353,N_2092,N_2150);
and U2354 (N_2354,N_2158,N_2234);
or U2355 (N_2355,N_2119,N_2097);
xor U2356 (N_2356,N_2135,N_2199);
or U2357 (N_2357,N_2197,N_2186);
nor U2358 (N_2358,N_2138,N_2211);
or U2359 (N_2359,N_2222,N_2238);
nor U2360 (N_2360,N_2177,N_2210);
nand U2361 (N_2361,N_2106,N_2164);
nand U2362 (N_2362,N_2196,N_2109);
nand U2363 (N_2363,N_2223,N_2129);
nand U2364 (N_2364,N_2206,N_2120);
nand U2365 (N_2365,N_2147,N_2099);
nand U2366 (N_2366,N_2177,N_2165);
nor U2367 (N_2367,N_2187,N_2177);
and U2368 (N_2368,N_2140,N_2084);
nor U2369 (N_2369,N_2133,N_2153);
xor U2370 (N_2370,N_2163,N_2123);
and U2371 (N_2371,N_2136,N_2178);
nand U2372 (N_2372,N_2115,N_2192);
and U2373 (N_2373,N_2225,N_2168);
nand U2374 (N_2374,N_2163,N_2093);
and U2375 (N_2375,N_2123,N_2169);
and U2376 (N_2376,N_2213,N_2164);
and U2377 (N_2377,N_2237,N_2085);
nand U2378 (N_2378,N_2120,N_2178);
xnor U2379 (N_2379,N_2217,N_2127);
nand U2380 (N_2380,N_2228,N_2160);
nand U2381 (N_2381,N_2100,N_2184);
or U2382 (N_2382,N_2114,N_2235);
nand U2383 (N_2383,N_2086,N_2146);
and U2384 (N_2384,N_2119,N_2103);
nor U2385 (N_2385,N_2091,N_2141);
or U2386 (N_2386,N_2144,N_2231);
and U2387 (N_2387,N_2221,N_2194);
nand U2388 (N_2388,N_2211,N_2207);
or U2389 (N_2389,N_2221,N_2231);
nor U2390 (N_2390,N_2134,N_2133);
nand U2391 (N_2391,N_2189,N_2208);
xnor U2392 (N_2392,N_2177,N_2117);
or U2393 (N_2393,N_2238,N_2086);
or U2394 (N_2394,N_2090,N_2236);
or U2395 (N_2395,N_2168,N_2096);
or U2396 (N_2396,N_2225,N_2100);
or U2397 (N_2397,N_2228,N_2212);
nor U2398 (N_2398,N_2192,N_2214);
or U2399 (N_2399,N_2203,N_2204);
nand U2400 (N_2400,N_2260,N_2378);
and U2401 (N_2401,N_2343,N_2375);
nand U2402 (N_2402,N_2295,N_2391);
nor U2403 (N_2403,N_2326,N_2372);
and U2404 (N_2404,N_2257,N_2386);
xor U2405 (N_2405,N_2342,N_2323);
and U2406 (N_2406,N_2368,N_2317);
or U2407 (N_2407,N_2265,N_2259);
or U2408 (N_2408,N_2356,N_2252);
xor U2409 (N_2409,N_2262,N_2369);
nand U2410 (N_2410,N_2333,N_2397);
nor U2411 (N_2411,N_2286,N_2240);
or U2412 (N_2412,N_2297,N_2388);
or U2413 (N_2413,N_2264,N_2266);
nand U2414 (N_2414,N_2296,N_2334);
nor U2415 (N_2415,N_2390,N_2360);
or U2416 (N_2416,N_2355,N_2327);
nand U2417 (N_2417,N_2352,N_2269);
and U2418 (N_2418,N_2306,N_2324);
nor U2419 (N_2419,N_2381,N_2344);
and U2420 (N_2420,N_2307,N_2330);
or U2421 (N_2421,N_2394,N_2384);
xor U2422 (N_2422,N_2396,N_2312);
or U2423 (N_2423,N_2332,N_2276);
and U2424 (N_2424,N_2316,N_2271);
or U2425 (N_2425,N_2305,N_2294);
or U2426 (N_2426,N_2383,N_2284);
or U2427 (N_2427,N_2353,N_2299);
or U2428 (N_2428,N_2398,N_2242);
nor U2429 (N_2429,N_2329,N_2359);
nor U2430 (N_2430,N_2349,N_2361);
and U2431 (N_2431,N_2335,N_2277);
or U2432 (N_2432,N_2251,N_2354);
nand U2433 (N_2433,N_2365,N_2301);
nand U2434 (N_2434,N_2279,N_2382);
xnor U2435 (N_2435,N_2337,N_2395);
and U2436 (N_2436,N_2300,N_2308);
nor U2437 (N_2437,N_2345,N_2275);
or U2438 (N_2438,N_2392,N_2298);
nor U2439 (N_2439,N_2374,N_2253);
nor U2440 (N_2440,N_2315,N_2274);
or U2441 (N_2441,N_2371,N_2320);
and U2442 (N_2442,N_2281,N_2272);
or U2443 (N_2443,N_2250,N_2325);
nand U2444 (N_2444,N_2263,N_2363);
nand U2445 (N_2445,N_2318,N_2373);
nor U2446 (N_2446,N_2322,N_2319);
or U2447 (N_2447,N_2243,N_2287);
and U2448 (N_2448,N_2358,N_2350);
nand U2449 (N_2449,N_2247,N_2389);
nor U2450 (N_2450,N_2283,N_2310);
or U2451 (N_2451,N_2289,N_2248);
nor U2452 (N_2452,N_2254,N_2270);
nand U2453 (N_2453,N_2246,N_2336);
or U2454 (N_2454,N_2244,N_2303);
nor U2455 (N_2455,N_2314,N_2348);
nor U2456 (N_2456,N_2258,N_2346);
nor U2457 (N_2457,N_2311,N_2367);
or U2458 (N_2458,N_2328,N_2321);
and U2459 (N_2459,N_2347,N_2282);
or U2460 (N_2460,N_2302,N_2357);
or U2461 (N_2461,N_2341,N_2278);
nand U2462 (N_2462,N_2364,N_2267);
or U2463 (N_2463,N_2331,N_2340);
xnor U2464 (N_2464,N_2273,N_2288);
nand U2465 (N_2465,N_2338,N_2256);
or U2466 (N_2466,N_2380,N_2376);
or U2467 (N_2467,N_2387,N_2385);
nor U2468 (N_2468,N_2285,N_2255);
xnor U2469 (N_2469,N_2377,N_2339);
nor U2470 (N_2470,N_2393,N_2291);
or U2471 (N_2471,N_2261,N_2293);
nor U2472 (N_2472,N_2399,N_2249);
nor U2473 (N_2473,N_2366,N_2313);
xor U2474 (N_2474,N_2362,N_2370);
or U2475 (N_2475,N_2379,N_2268);
nor U2476 (N_2476,N_2351,N_2304);
xnor U2477 (N_2477,N_2245,N_2280);
xnor U2478 (N_2478,N_2309,N_2292);
nor U2479 (N_2479,N_2290,N_2241);
xnor U2480 (N_2480,N_2292,N_2370);
nor U2481 (N_2481,N_2249,N_2370);
nor U2482 (N_2482,N_2361,N_2326);
or U2483 (N_2483,N_2255,N_2288);
nand U2484 (N_2484,N_2326,N_2355);
xnor U2485 (N_2485,N_2254,N_2323);
nor U2486 (N_2486,N_2390,N_2284);
or U2487 (N_2487,N_2290,N_2387);
and U2488 (N_2488,N_2334,N_2298);
and U2489 (N_2489,N_2347,N_2340);
or U2490 (N_2490,N_2277,N_2394);
nand U2491 (N_2491,N_2329,N_2252);
nor U2492 (N_2492,N_2322,N_2391);
xnor U2493 (N_2493,N_2287,N_2308);
nor U2494 (N_2494,N_2359,N_2320);
xnor U2495 (N_2495,N_2397,N_2302);
nand U2496 (N_2496,N_2265,N_2367);
nor U2497 (N_2497,N_2242,N_2305);
nor U2498 (N_2498,N_2280,N_2308);
and U2499 (N_2499,N_2360,N_2370);
nor U2500 (N_2500,N_2267,N_2326);
nand U2501 (N_2501,N_2303,N_2292);
nand U2502 (N_2502,N_2349,N_2375);
nor U2503 (N_2503,N_2393,N_2350);
and U2504 (N_2504,N_2248,N_2347);
nand U2505 (N_2505,N_2356,N_2274);
or U2506 (N_2506,N_2350,N_2268);
xnor U2507 (N_2507,N_2316,N_2365);
and U2508 (N_2508,N_2285,N_2258);
xor U2509 (N_2509,N_2370,N_2302);
and U2510 (N_2510,N_2273,N_2283);
nand U2511 (N_2511,N_2396,N_2318);
or U2512 (N_2512,N_2389,N_2381);
and U2513 (N_2513,N_2255,N_2321);
and U2514 (N_2514,N_2241,N_2298);
and U2515 (N_2515,N_2300,N_2394);
nand U2516 (N_2516,N_2348,N_2266);
and U2517 (N_2517,N_2297,N_2399);
nor U2518 (N_2518,N_2378,N_2246);
or U2519 (N_2519,N_2382,N_2280);
xor U2520 (N_2520,N_2257,N_2287);
nor U2521 (N_2521,N_2302,N_2297);
and U2522 (N_2522,N_2267,N_2266);
or U2523 (N_2523,N_2369,N_2304);
or U2524 (N_2524,N_2364,N_2381);
nand U2525 (N_2525,N_2345,N_2297);
and U2526 (N_2526,N_2241,N_2389);
nor U2527 (N_2527,N_2311,N_2382);
nand U2528 (N_2528,N_2390,N_2307);
nor U2529 (N_2529,N_2278,N_2288);
or U2530 (N_2530,N_2303,N_2359);
or U2531 (N_2531,N_2252,N_2271);
and U2532 (N_2532,N_2244,N_2376);
xnor U2533 (N_2533,N_2245,N_2385);
nand U2534 (N_2534,N_2398,N_2270);
nor U2535 (N_2535,N_2379,N_2294);
nand U2536 (N_2536,N_2391,N_2371);
and U2537 (N_2537,N_2282,N_2399);
or U2538 (N_2538,N_2296,N_2295);
or U2539 (N_2539,N_2284,N_2311);
or U2540 (N_2540,N_2255,N_2249);
and U2541 (N_2541,N_2323,N_2305);
nand U2542 (N_2542,N_2398,N_2397);
and U2543 (N_2543,N_2243,N_2291);
and U2544 (N_2544,N_2335,N_2329);
nor U2545 (N_2545,N_2333,N_2365);
nand U2546 (N_2546,N_2365,N_2323);
nand U2547 (N_2547,N_2327,N_2259);
xnor U2548 (N_2548,N_2296,N_2355);
nor U2549 (N_2549,N_2397,N_2362);
or U2550 (N_2550,N_2297,N_2277);
nor U2551 (N_2551,N_2259,N_2370);
nand U2552 (N_2552,N_2279,N_2344);
nor U2553 (N_2553,N_2318,N_2391);
and U2554 (N_2554,N_2257,N_2360);
or U2555 (N_2555,N_2283,N_2395);
nand U2556 (N_2556,N_2263,N_2385);
nor U2557 (N_2557,N_2295,N_2279);
and U2558 (N_2558,N_2319,N_2269);
nor U2559 (N_2559,N_2304,N_2320);
and U2560 (N_2560,N_2439,N_2432);
or U2561 (N_2561,N_2498,N_2525);
nand U2562 (N_2562,N_2552,N_2543);
xor U2563 (N_2563,N_2468,N_2408);
nand U2564 (N_2564,N_2433,N_2524);
or U2565 (N_2565,N_2440,N_2500);
or U2566 (N_2566,N_2503,N_2512);
and U2567 (N_2567,N_2413,N_2518);
and U2568 (N_2568,N_2435,N_2534);
nand U2569 (N_2569,N_2409,N_2508);
nand U2570 (N_2570,N_2422,N_2463);
and U2571 (N_2571,N_2427,N_2404);
nor U2572 (N_2572,N_2482,N_2532);
xor U2573 (N_2573,N_2541,N_2459);
nand U2574 (N_2574,N_2481,N_2506);
and U2575 (N_2575,N_2489,N_2494);
nor U2576 (N_2576,N_2436,N_2464);
or U2577 (N_2577,N_2507,N_2537);
or U2578 (N_2578,N_2502,N_2410);
or U2579 (N_2579,N_2495,N_2429);
nor U2580 (N_2580,N_2553,N_2545);
nand U2581 (N_2581,N_2505,N_2533);
nor U2582 (N_2582,N_2477,N_2471);
nand U2583 (N_2583,N_2431,N_2401);
nand U2584 (N_2584,N_2423,N_2546);
or U2585 (N_2585,N_2441,N_2529);
and U2586 (N_2586,N_2475,N_2514);
nor U2587 (N_2587,N_2540,N_2419);
or U2588 (N_2588,N_2509,N_2492);
or U2589 (N_2589,N_2536,N_2497);
xnor U2590 (N_2590,N_2415,N_2405);
xnor U2591 (N_2591,N_2466,N_2478);
nor U2592 (N_2592,N_2444,N_2480);
nor U2593 (N_2593,N_2400,N_2544);
or U2594 (N_2594,N_2453,N_2558);
nor U2595 (N_2595,N_2467,N_2548);
or U2596 (N_2596,N_2412,N_2430);
nor U2597 (N_2597,N_2511,N_2556);
or U2598 (N_2598,N_2486,N_2531);
nor U2599 (N_2599,N_2445,N_2442);
nand U2600 (N_2600,N_2474,N_2446);
xnor U2601 (N_2601,N_2451,N_2547);
nor U2602 (N_2602,N_2403,N_2523);
nor U2603 (N_2603,N_2434,N_2559);
and U2604 (N_2604,N_2448,N_2510);
and U2605 (N_2605,N_2490,N_2473);
and U2606 (N_2606,N_2417,N_2484);
and U2607 (N_2607,N_2517,N_2501);
xnor U2608 (N_2608,N_2424,N_2554);
or U2609 (N_2609,N_2407,N_2443);
or U2610 (N_2610,N_2414,N_2499);
or U2611 (N_2611,N_2557,N_2496);
or U2612 (N_2612,N_2425,N_2483);
and U2613 (N_2613,N_2458,N_2455);
and U2614 (N_2614,N_2447,N_2476);
nor U2615 (N_2615,N_2450,N_2462);
and U2616 (N_2616,N_2411,N_2472);
nor U2617 (N_2617,N_2485,N_2526);
and U2618 (N_2618,N_2426,N_2470);
or U2619 (N_2619,N_2521,N_2522);
and U2620 (N_2620,N_2519,N_2515);
and U2621 (N_2621,N_2438,N_2549);
or U2622 (N_2622,N_2420,N_2487);
nor U2623 (N_2623,N_2452,N_2418);
nand U2624 (N_2624,N_2550,N_2504);
nand U2625 (N_2625,N_2555,N_2457);
xnor U2626 (N_2626,N_2479,N_2465);
or U2627 (N_2627,N_2513,N_2535);
and U2628 (N_2628,N_2449,N_2456);
and U2629 (N_2629,N_2539,N_2402);
and U2630 (N_2630,N_2493,N_2491);
nand U2631 (N_2631,N_2542,N_2516);
and U2632 (N_2632,N_2551,N_2428);
and U2633 (N_2633,N_2528,N_2469);
nand U2634 (N_2634,N_2530,N_2538);
xnor U2635 (N_2635,N_2406,N_2488);
nand U2636 (N_2636,N_2520,N_2437);
and U2637 (N_2637,N_2461,N_2460);
xnor U2638 (N_2638,N_2416,N_2454);
nor U2639 (N_2639,N_2527,N_2421);
or U2640 (N_2640,N_2533,N_2463);
xor U2641 (N_2641,N_2527,N_2538);
or U2642 (N_2642,N_2509,N_2522);
and U2643 (N_2643,N_2432,N_2503);
nor U2644 (N_2644,N_2499,N_2455);
nor U2645 (N_2645,N_2519,N_2538);
or U2646 (N_2646,N_2403,N_2437);
nand U2647 (N_2647,N_2412,N_2429);
or U2648 (N_2648,N_2479,N_2440);
nor U2649 (N_2649,N_2447,N_2544);
and U2650 (N_2650,N_2500,N_2545);
and U2651 (N_2651,N_2425,N_2522);
and U2652 (N_2652,N_2412,N_2444);
nor U2653 (N_2653,N_2552,N_2532);
nor U2654 (N_2654,N_2477,N_2404);
nor U2655 (N_2655,N_2512,N_2558);
and U2656 (N_2656,N_2417,N_2477);
nor U2657 (N_2657,N_2495,N_2532);
or U2658 (N_2658,N_2408,N_2531);
or U2659 (N_2659,N_2543,N_2533);
or U2660 (N_2660,N_2524,N_2552);
or U2661 (N_2661,N_2428,N_2460);
and U2662 (N_2662,N_2413,N_2437);
nand U2663 (N_2663,N_2465,N_2544);
nand U2664 (N_2664,N_2541,N_2489);
and U2665 (N_2665,N_2449,N_2467);
nor U2666 (N_2666,N_2528,N_2548);
nor U2667 (N_2667,N_2437,N_2484);
nand U2668 (N_2668,N_2464,N_2493);
and U2669 (N_2669,N_2455,N_2553);
xor U2670 (N_2670,N_2528,N_2430);
or U2671 (N_2671,N_2557,N_2500);
or U2672 (N_2672,N_2541,N_2426);
and U2673 (N_2673,N_2402,N_2490);
or U2674 (N_2674,N_2552,N_2555);
xor U2675 (N_2675,N_2515,N_2545);
nor U2676 (N_2676,N_2493,N_2416);
or U2677 (N_2677,N_2499,N_2470);
and U2678 (N_2678,N_2441,N_2434);
xnor U2679 (N_2679,N_2501,N_2486);
and U2680 (N_2680,N_2458,N_2446);
and U2681 (N_2681,N_2446,N_2476);
or U2682 (N_2682,N_2472,N_2473);
nand U2683 (N_2683,N_2450,N_2479);
and U2684 (N_2684,N_2552,N_2426);
nand U2685 (N_2685,N_2406,N_2407);
nand U2686 (N_2686,N_2525,N_2411);
xnor U2687 (N_2687,N_2420,N_2471);
nand U2688 (N_2688,N_2555,N_2557);
or U2689 (N_2689,N_2524,N_2453);
or U2690 (N_2690,N_2508,N_2510);
nor U2691 (N_2691,N_2421,N_2551);
xor U2692 (N_2692,N_2537,N_2496);
nor U2693 (N_2693,N_2549,N_2521);
or U2694 (N_2694,N_2495,N_2456);
nand U2695 (N_2695,N_2440,N_2547);
nand U2696 (N_2696,N_2408,N_2508);
nand U2697 (N_2697,N_2470,N_2466);
and U2698 (N_2698,N_2486,N_2488);
nand U2699 (N_2699,N_2456,N_2490);
or U2700 (N_2700,N_2539,N_2554);
and U2701 (N_2701,N_2400,N_2558);
or U2702 (N_2702,N_2546,N_2542);
xor U2703 (N_2703,N_2512,N_2475);
nor U2704 (N_2704,N_2481,N_2488);
nor U2705 (N_2705,N_2466,N_2526);
or U2706 (N_2706,N_2453,N_2480);
xor U2707 (N_2707,N_2511,N_2489);
or U2708 (N_2708,N_2517,N_2470);
nor U2709 (N_2709,N_2445,N_2410);
and U2710 (N_2710,N_2478,N_2504);
nor U2711 (N_2711,N_2400,N_2453);
nor U2712 (N_2712,N_2462,N_2476);
nand U2713 (N_2713,N_2516,N_2513);
nand U2714 (N_2714,N_2407,N_2520);
nand U2715 (N_2715,N_2497,N_2530);
nor U2716 (N_2716,N_2530,N_2559);
nor U2717 (N_2717,N_2517,N_2427);
or U2718 (N_2718,N_2535,N_2448);
nor U2719 (N_2719,N_2428,N_2469);
nand U2720 (N_2720,N_2693,N_2587);
and U2721 (N_2721,N_2609,N_2630);
or U2722 (N_2722,N_2703,N_2707);
xnor U2723 (N_2723,N_2667,N_2683);
or U2724 (N_2724,N_2576,N_2579);
nand U2725 (N_2725,N_2689,N_2564);
and U2726 (N_2726,N_2663,N_2623);
nand U2727 (N_2727,N_2662,N_2640);
nor U2728 (N_2728,N_2688,N_2704);
or U2729 (N_2729,N_2652,N_2589);
nor U2730 (N_2730,N_2603,N_2566);
or U2731 (N_2731,N_2573,N_2578);
nand U2732 (N_2732,N_2635,N_2636);
nor U2733 (N_2733,N_2642,N_2694);
nand U2734 (N_2734,N_2601,N_2618);
nand U2735 (N_2735,N_2568,N_2592);
or U2736 (N_2736,N_2697,N_2666);
nand U2737 (N_2737,N_2570,N_2655);
nor U2738 (N_2738,N_2698,N_2677);
and U2739 (N_2739,N_2613,N_2585);
and U2740 (N_2740,N_2617,N_2638);
xor U2741 (N_2741,N_2622,N_2645);
and U2742 (N_2742,N_2639,N_2588);
or U2743 (N_2743,N_2606,N_2672);
xnor U2744 (N_2744,N_2715,N_2658);
nand U2745 (N_2745,N_2614,N_2634);
nand U2746 (N_2746,N_2669,N_2691);
or U2747 (N_2747,N_2612,N_2660);
nand U2748 (N_2748,N_2595,N_2597);
and U2749 (N_2749,N_2629,N_2679);
and U2750 (N_2750,N_2604,N_2586);
and U2751 (N_2751,N_2716,N_2561);
or U2752 (N_2752,N_2583,N_2631);
nand U2753 (N_2753,N_2577,N_2580);
nand U2754 (N_2754,N_2581,N_2690);
xnor U2755 (N_2755,N_2643,N_2661);
and U2756 (N_2756,N_2560,N_2674);
and U2757 (N_2757,N_2650,N_2625);
and U2758 (N_2758,N_2599,N_2685);
or U2759 (N_2759,N_2696,N_2572);
nor U2760 (N_2760,N_2719,N_2571);
or U2761 (N_2761,N_2608,N_2590);
nor U2762 (N_2762,N_2648,N_2644);
nor U2763 (N_2763,N_2574,N_2646);
and U2764 (N_2764,N_2712,N_2632);
or U2765 (N_2765,N_2582,N_2705);
xnor U2766 (N_2766,N_2565,N_2651);
or U2767 (N_2767,N_2627,N_2649);
and U2768 (N_2768,N_2600,N_2621);
or U2769 (N_2769,N_2709,N_2708);
and U2770 (N_2770,N_2594,N_2616);
nor U2771 (N_2771,N_2684,N_2717);
or U2772 (N_2772,N_2596,N_2569);
and U2773 (N_2773,N_2605,N_2710);
nand U2774 (N_2774,N_2641,N_2706);
nor U2775 (N_2775,N_2611,N_2633);
and U2776 (N_2776,N_2678,N_2562);
xnor U2777 (N_2777,N_2610,N_2615);
or U2778 (N_2778,N_2619,N_2628);
and U2779 (N_2779,N_2602,N_2702);
nand U2780 (N_2780,N_2676,N_2714);
xnor U2781 (N_2781,N_2665,N_2680);
nor U2782 (N_2782,N_2713,N_2584);
and U2783 (N_2783,N_2686,N_2620);
xor U2784 (N_2784,N_2670,N_2626);
nor U2785 (N_2785,N_2575,N_2675);
or U2786 (N_2786,N_2699,N_2664);
or U2787 (N_2787,N_2711,N_2718);
nor U2788 (N_2788,N_2654,N_2659);
nand U2789 (N_2789,N_2700,N_2695);
or U2790 (N_2790,N_2692,N_2668);
nor U2791 (N_2791,N_2591,N_2701);
nor U2792 (N_2792,N_2624,N_2682);
or U2793 (N_2793,N_2563,N_2593);
or U2794 (N_2794,N_2598,N_2567);
or U2795 (N_2795,N_2687,N_2673);
or U2796 (N_2796,N_2671,N_2647);
and U2797 (N_2797,N_2637,N_2656);
xnor U2798 (N_2798,N_2681,N_2653);
nand U2799 (N_2799,N_2607,N_2657);
nand U2800 (N_2800,N_2688,N_2571);
and U2801 (N_2801,N_2631,N_2570);
xnor U2802 (N_2802,N_2619,N_2719);
nor U2803 (N_2803,N_2660,N_2650);
or U2804 (N_2804,N_2594,N_2599);
or U2805 (N_2805,N_2715,N_2616);
and U2806 (N_2806,N_2705,N_2651);
or U2807 (N_2807,N_2654,N_2571);
and U2808 (N_2808,N_2697,N_2564);
nor U2809 (N_2809,N_2699,N_2661);
or U2810 (N_2810,N_2649,N_2671);
and U2811 (N_2811,N_2639,N_2625);
nand U2812 (N_2812,N_2674,N_2691);
nor U2813 (N_2813,N_2712,N_2697);
and U2814 (N_2814,N_2621,N_2618);
or U2815 (N_2815,N_2590,N_2717);
nand U2816 (N_2816,N_2641,N_2579);
or U2817 (N_2817,N_2573,N_2677);
nand U2818 (N_2818,N_2703,N_2592);
nor U2819 (N_2819,N_2674,N_2598);
nor U2820 (N_2820,N_2653,N_2611);
and U2821 (N_2821,N_2686,N_2627);
or U2822 (N_2822,N_2652,N_2648);
nor U2823 (N_2823,N_2668,N_2635);
xnor U2824 (N_2824,N_2660,N_2673);
and U2825 (N_2825,N_2707,N_2696);
nor U2826 (N_2826,N_2571,N_2586);
xor U2827 (N_2827,N_2657,N_2694);
and U2828 (N_2828,N_2568,N_2681);
nor U2829 (N_2829,N_2623,N_2716);
nand U2830 (N_2830,N_2691,N_2677);
and U2831 (N_2831,N_2650,N_2617);
nand U2832 (N_2832,N_2566,N_2586);
or U2833 (N_2833,N_2599,N_2690);
nor U2834 (N_2834,N_2702,N_2664);
nor U2835 (N_2835,N_2663,N_2616);
and U2836 (N_2836,N_2576,N_2617);
and U2837 (N_2837,N_2667,N_2594);
or U2838 (N_2838,N_2573,N_2651);
xnor U2839 (N_2839,N_2581,N_2578);
nor U2840 (N_2840,N_2710,N_2621);
or U2841 (N_2841,N_2579,N_2649);
nand U2842 (N_2842,N_2707,N_2600);
nand U2843 (N_2843,N_2609,N_2649);
xnor U2844 (N_2844,N_2650,N_2587);
or U2845 (N_2845,N_2587,N_2567);
or U2846 (N_2846,N_2635,N_2634);
or U2847 (N_2847,N_2684,N_2667);
and U2848 (N_2848,N_2647,N_2659);
or U2849 (N_2849,N_2639,N_2633);
nand U2850 (N_2850,N_2569,N_2583);
nand U2851 (N_2851,N_2674,N_2563);
xor U2852 (N_2852,N_2712,N_2658);
nor U2853 (N_2853,N_2592,N_2658);
nor U2854 (N_2854,N_2715,N_2570);
and U2855 (N_2855,N_2563,N_2672);
and U2856 (N_2856,N_2664,N_2657);
or U2857 (N_2857,N_2608,N_2607);
nand U2858 (N_2858,N_2702,N_2715);
and U2859 (N_2859,N_2609,N_2616);
or U2860 (N_2860,N_2605,N_2682);
xor U2861 (N_2861,N_2692,N_2710);
and U2862 (N_2862,N_2624,N_2577);
or U2863 (N_2863,N_2611,N_2662);
or U2864 (N_2864,N_2682,N_2610);
nor U2865 (N_2865,N_2712,N_2588);
and U2866 (N_2866,N_2589,N_2715);
or U2867 (N_2867,N_2636,N_2628);
nand U2868 (N_2868,N_2669,N_2642);
and U2869 (N_2869,N_2610,N_2688);
nand U2870 (N_2870,N_2570,N_2699);
xnor U2871 (N_2871,N_2696,N_2678);
nor U2872 (N_2872,N_2578,N_2572);
or U2873 (N_2873,N_2651,N_2719);
or U2874 (N_2874,N_2572,N_2690);
nand U2875 (N_2875,N_2583,N_2712);
nand U2876 (N_2876,N_2664,N_2578);
and U2877 (N_2877,N_2631,N_2560);
nand U2878 (N_2878,N_2716,N_2706);
xnor U2879 (N_2879,N_2575,N_2679);
nand U2880 (N_2880,N_2800,N_2723);
or U2881 (N_2881,N_2796,N_2733);
or U2882 (N_2882,N_2858,N_2829);
xor U2883 (N_2883,N_2758,N_2768);
nand U2884 (N_2884,N_2754,N_2846);
xor U2885 (N_2885,N_2866,N_2817);
nor U2886 (N_2886,N_2832,N_2775);
nand U2887 (N_2887,N_2851,N_2872);
nor U2888 (N_2888,N_2790,N_2864);
nand U2889 (N_2889,N_2773,N_2797);
nor U2890 (N_2890,N_2738,N_2826);
nand U2891 (N_2891,N_2825,N_2743);
or U2892 (N_2892,N_2782,N_2878);
or U2893 (N_2893,N_2794,N_2847);
nor U2894 (N_2894,N_2792,N_2842);
and U2895 (N_2895,N_2857,N_2761);
or U2896 (N_2896,N_2852,N_2757);
nand U2897 (N_2897,N_2816,N_2860);
and U2898 (N_2898,N_2833,N_2821);
nor U2899 (N_2899,N_2807,N_2823);
nor U2900 (N_2900,N_2759,N_2805);
or U2901 (N_2901,N_2784,N_2755);
nand U2902 (N_2902,N_2859,N_2785);
and U2903 (N_2903,N_2813,N_2849);
and U2904 (N_2904,N_2841,N_2787);
or U2905 (N_2905,N_2777,N_2779);
and U2906 (N_2906,N_2786,N_2769);
nor U2907 (N_2907,N_2865,N_2808);
or U2908 (N_2908,N_2802,N_2778);
and U2909 (N_2909,N_2774,N_2728);
nor U2910 (N_2910,N_2831,N_2727);
nand U2911 (N_2911,N_2861,N_2871);
nand U2912 (N_2912,N_2750,N_2875);
and U2913 (N_2913,N_2811,N_2741);
or U2914 (N_2914,N_2873,N_2824);
nand U2915 (N_2915,N_2848,N_2726);
xor U2916 (N_2916,N_2724,N_2850);
xnor U2917 (N_2917,N_2855,N_2736);
nor U2918 (N_2918,N_2765,N_2843);
nand U2919 (N_2919,N_2869,N_2820);
nor U2920 (N_2920,N_2803,N_2828);
nor U2921 (N_2921,N_2791,N_2740);
and U2922 (N_2922,N_2725,N_2809);
nor U2923 (N_2923,N_2834,N_2804);
or U2924 (N_2924,N_2835,N_2801);
and U2925 (N_2925,N_2868,N_2751);
nor U2926 (N_2926,N_2753,N_2763);
xor U2927 (N_2927,N_2799,N_2844);
nor U2928 (N_2928,N_2760,N_2822);
nor U2929 (N_2929,N_2748,N_2722);
or U2930 (N_2930,N_2730,N_2766);
and U2931 (N_2931,N_2854,N_2806);
or U2932 (N_2932,N_2879,N_2840);
nand U2933 (N_2933,N_2781,N_2795);
or U2934 (N_2934,N_2827,N_2734);
and U2935 (N_2935,N_2874,N_2793);
nand U2936 (N_2936,N_2814,N_2810);
and U2937 (N_2937,N_2836,N_2735);
nand U2938 (N_2938,N_2771,N_2856);
nor U2939 (N_2939,N_2749,N_2772);
nor U2940 (N_2940,N_2720,N_2798);
and U2941 (N_2941,N_2739,N_2815);
xor U2942 (N_2942,N_2752,N_2762);
nor U2943 (N_2943,N_2756,N_2830);
or U2944 (N_2944,N_2876,N_2789);
nor U2945 (N_2945,N_2742,N_2764);
nor U2946 (N_2946,N_2783,N_2877);
nor U2947 (N_2947,N_2818,N_2867);
and U2948 (N_2948,N_2780,N_2870);
nor U2949 (N_2949,N_2729,N_2744);
xnor U2950 (N_2950,N_2853,N_2776);
nand U2951 (N_2951,N_2746,N_2862);
nand U2952 (N_2952,N_2837,N_2767);
or U2953 (N_2953,N_2737,N_2732);
nand U2954 (N_2954,N_2812,N_2819);
xnor U2955 (N_2955,N_2745,N_2731);
nand U2956 (N_2956,N_2845,N_2838);
and U2957 (N_2957,N_2721,N_2863);
or U2958 (N_2958,N_2788,N_2839);
and U2959 (N_2959,N_2770,N_2747);
nor U2960 (N_2960,N_2851,N_2793);
xnor U2961 (N_2961,N_2765,N_2767);
nor U2962 (N_2962,N_2828,N_2725);
and U2963 (N_2963,N_2736,N_2838);
nand U2964 (N_2964,N_2806,N_2847);
and U2965 (N_2965,N_2848,N_2814);
nand U2966 (N_2966,N_2782,N_2748);
nor U2967 (N_2967,N_2746,N_2782);
nand U2968 (N_2968,N_2816,N_2863);
nand U2969 (N_2969,N_2872,N_2773);
nor U2970 (N_2970,N_2740,N_2770);
and U2971 (N_2971,N_2731,N_2801);
or U2972 (N_2972,N_2745,N_2767);
or U2973 (N_2973,N_2868,N_2768);
and U2974 (N_2974,N_2795,N_2765);
nor U2975 (N_2975,N_2722,N_2761);
and U2976 (N_2976,N_2740,N_2742);
xor U2977 (N_2977,N_2733,N_2855);
nor U2978 (N_2978,N_2832,N_2769);
nand U2979 (N_2979,N_2808,N_2770);
or U2980 (N_2980,N_2782,N_2768);
and U2981 (N_2981,N_2856,N_2725);
xnor U2982 (N_2982,N_2870,N_2842);
nor U2983 (N_2983,N_2757,N_2798);
nor U2984 (N_2984,N_2842,N_2751);
and U2985 (N_2985,N_2825,N_2770);
or U2986 (N_2986,N_2739,N_2810);
and U2987 (N_2987,N_2802,N_2774);
xor U2988 (N_2988,N_2724,N_2734);
nor U2989 (N_2989,N_2790,N_2871);
and U2990 (N_2990,N_2721,N_2801);
or U2991 (N_2991,N_2782,N_2815);
xor U2992 (N_2992,N_2774,N_2833);
xor U2993 (N_2993,N_2847,N_2831);
nor U2994 (N_2994,N_2811,N_2760);
and U2995 (N_2995,N_2863,N_2727);
xor U2996 (N_2996,N_2728,N_2812);
or U2997 (N_2997,N_2865,N_2786);
nor U2998 (N_2998,N_2758,N_2853);
nor U2999 (N_2999,N_2721,N_2828);
xor U3000 (N_3000,N_2794,N_2774);
and U3001 (N_3001,N_2789,N_2772);
nand U3002 (N_3002,N_2803,N_2804);
or U3003 (N_3003,N_2729,N_2728);
or U3004 (N_3004,N_2740,N_2811);
or U3005 (N_3005,N_2732,N_2878);
and U3006 (N_3006,N_2844,N_2790);
nor U3007 (N_3007,N_2786,N_2737);
or U3008 (N_3008,N_2789,N_2749);
and U3009 (N_3009,N_2742,N_2732);
and U3010 (N_3010,N_2877,N_2765);
or U3011 (N_3011,N_2761,N_2818);
or U3012 (N_3012,N_2862,N_2733);
nand U3013 (N_3013,N_2733,N_2813);
nor U3014 (N_3014,N_2831,N_2755);
or U3015 (N_3015,N_2860,N_2799);
and U3016 (N_3016,N_2869,N_2862);
and U3017 (N_3017,N_2853,N_2860);
nor U3018 (N_3018,N_2785,N_2858);
nor U3019 (N_3019,N_2759,N_2760);
or U3020 (N_3020,N_2779,N_2819);
or U3021 (N_3021,N_2823,N_2809);
nand U3022 (N_3022,N_2747,N_2803);
xor U3023 (N_3023,N_2795,N_2825);
nor U3024 (N_3024,N_2734,N_2864);
nor U3025 (N_3025,N_2867,N_2795);
or U3026 (N_3026,N_2824,N_2736);
nand U3027 (N_3027,N_2776,N_2724);
nand U3028 (N_3028,N_2818,N_2875);
nor U3029 (N_3029,N_2769,N_2874);
and U3030 (N_3030,N_2878,N_2743);
nor U3031 (N_3031,N_2749,N_2850);
nor U3032 (N_3032,N_2776,N_2730);
nand U3033 (N_3033,N_2829,N_2782);
xnor U3034 (N_3034,N_2831,N_2807);
and U3035 (N_3035,N_2795,N_2767);
or U3036 (N_3036,N_2771,N_2733);
nand U3037 (N_3037,N_2774,N_2750);
nor U3038 (N_3038,N_2877,N_2852);
and U3039 (N_3039,N_2795,N_2876);
nor U3040 (N_3040,N_2964,N_3037);
or U3041 (N_3041,N_2932,N_2913);
xnor U3042 (N_3042,N_3004,N_2970);
nor U3043 (N_3043,N_2892,N_2982);
or U3044 (N_3044,N_2974,N_3036);
xor U3045 (N_3045,N_2899,N_2992);
and U3046 (N_3046,N_2907,N_2965);
and U3047 (N_3047,N_2908,N_2914);
and U3048 (N_3048,N_2918,N_2929);
xor U3049 (N_3049,N_2933,N_3032);
and U3050 (N_3050,N_2959,N_2958);
or U3051 (N_3051,N_2939,N_3002);
and U3052 (N_3052,N_2881,N_2937);
and U3053 (N_3053,N_2996,N_3016);
xor U3054 (N_3054,N_2990,N_2954);
nand U3055 (N_3055,N_3005,N_2923);
and U3056 (N_3056,N_3001,N_2943);
or U3057 (N_3057,N_2976,N_2888);
or U3058 (N_3058,N_2945,N_2981);
nand U3059 (N_3059,N_2904,N_2886);
nor U3060 (N_3060,N_2883,N_3031);
and U3061 (N_3061,N_2984,N_3000);
nor U3062 (N_3062,N_3015,N_2893);
and U3063 (N_3063,N_2900,N_3030);
and U3064 (N_3064,N_2885,N_2920);
and U3065 (N_3065,N_2898,N_2991);
nand U3066 (N_3066,N_2950,N_3003);
nand U3067 (N_3067,N_3008,N_2949);
and U3068 (N_3068,N_2942,N_2897);
or U3069 (N_3069,N_2931,N_2997);
nand U3070 (N_3070,N_2989,N_2979);
xor U3071 (N_3071,N_2922,N_2940);
or U3072 (N_3072,N_2919,N_2944);
xnor U3073 (N_3073,N_2911,N_3019);
nand U3074 (N_3074,N_2960,N_2972);
nor U3075 (N_3075,N_2928,N_3007);
nand U3076 (N_3076,N_2917,N_3024);
nand U3077 (N_3077,N_2963,N_2985);
nand U3078 (N_3078,N_2957,N_3025);
and U3079 (N_3079,N_2961,N_2987);
or U3080 (N_3080,N_2905,N_2967);
xor U3081 (N_3081,N_2946,N_2896);
xor U3082 (N_3082,N_3027,N_2887);
nand U3083 (N_3083,N_2968,N_2884);
nor U3084 (N_3084,N_2956,N_2973);
xor U3085 (N_3085,N_2921,N_2890);
and U3086 (N_3086,N_2906,N_2910);
or U3087 (N_3087,N_2977,N_2916);
nand U3088 (N_3088,N_2891,N_2969);
nand U3089 (N_3089,N_2995,N_2966);
xor U3090 (N_3090,N_2926,N_3006);
nor U3091 (N_3091,N_2924,N_2934);
nand U3092 (N_3092,N_2925,N_2902);
and U3093 (N_3093,N_2903,N_2962);
nor U3094 (N_3094,N_2935,N_3029);
nand U3095 (N_3095,N_2894,N_2986);
nand U3096 (N_3096,N_2978,N_2952);
and U3097 (N_3097,N_3022,N_3012);
nor U3098 (N_3098,N_2930,N_3034);
or U3099 (N_3099,N_2980,N_3028);
nor U3100 (N_3100,N_2999,N_2983);
or U3101 (N_3101,N_3038,N_3018);
and U3102 (N_3102,N_2975,N_2998);
or U3103 (N_3103,N_3023,N_3017);
or U3104 (N_3104,N_3026,N_2936);
or U3105 (N_3105,N_3035,N_2889);
and U3106 (N_3106,N_3010,N_2994);
and U3107 (N_3107,N_3013,N_2993);
nor U3108 (N_3108,N_3014,N_3009);
nand U3109 (N_3109,N_3021,N_2955);
nand U3110 (N_3110,N_2953,N_2909);
and U3111 (N_3111,N_2882,N_2941);
xnor U3112 (N_3112,N_2988,N_2938);
nand U3113 (N_3113,N_3020,N_2912);
and U3114 (N_3114,N_2951,N_2915);
or U3115 (N_3115,N_2927,N_2947);
or U3116 (N_3116,N_2901,N_2971);
and U3117 (N_3117,N_3011,N_2948);
and U3118 (N_3118,N_3039,N_3033);
and U3119 (N_3119,N_2880,N_2895);
nand U3120 (N_3120,N_3019,N_2967);
nor U3121 (N_3121,N_3036,N_2897);
nand U3122 (N_3122,N_3000,N_3018);
or U3123 (N_3123,N_2933,N_2973);
or U3124 (N_3124,N_2883,N_3030);
nor U3125 (N_3125,N_2922,N_2888);
and U3126 (N_3126,N_2927,N_2930);
nand U3127 (N_3127,N_2893,N_2990);
or U3128 (N_3128,N_2917,N_2883);
nand U3129 (N_3129,N_3003,N_3033);
xor U3130 (N_3130,N_3029,N_2885);
and U3131 (N_3131,N_2934,N_2981);
nand U3132 (N_3132,N_2891,N_2977);
or U3133 (N_3133,N_2984,N_3014);
and U3134 (N_3134,N_2969,N_2996);
nor U3135 (N_3135,N_2995,N_2984);
or U3136 (N_3136,N_3036,N_3018);
or U3137 (N_3137,N_3039,N_2965);
nand U3138 (N_3138,N_2999,N_2967);
nand U3139 (N_3139,N_3029,N_3015);
and U3140 (N_3140,N_3010,N_2901);
nand U3141 (N_3141,N_2983,N_3015);
or U3142 (N_3142,N_2935,N_2956);
nand U3143 (N_3143,N_3030,N_2945);
nor U3144 (N_3144,N_2895,N_2986);
or U3145 (N_3145,N_2935,N_2886);
nand U3146 (N_3146,N_2933,N_3001);
and U3147 (N_3147,N_2893,N_3027);
nor U3148 (N_3148,N_2940,N_3029);
and U3149 (N_3149,N_2915,N_2910);
nand U3150 (N_3150,N_2985,N_2954);
nand U3151 (N_3151,N_3021,N_3028);
nor U3152 (N_3152,N_2945,N_2939);
and U3153 (N_3153,N_3034,N_2911);
or U3154 (N_3154,N_2924,N_3015);
or U3155 (N_3155,N_2997,N_3034);
xor U3156 (N_3156,N_2936,N_3013);
or U3157 (N_3157,N_2924,N_2931);
and U3158 (N_3158,N_2944,N_2905);
or U3159 (N_3159,N_2898,N_2912);
nand U3160 (N_3160,N_2909,N_2944);
nor U3161 (N_3161,N_2913,N_3010);
nand U3162 (N_3162,N_3022,N_3014);
or U3163 (N_3163,N_2993,N_2964);
nand U3164 (N_3164,N_2976,N_2926);
nand U3165 (N_3165,N_2978,N_2973);
nand U3166 (N_3166,N_2971,N_2886);
nor U3167 (N_3167,N_3024,N_3013);
nand U3168 (N_3168,N_2968,N_2992);
and U3169 (N_3169,N_3003,N_2942);
nand U3170 (N_3170,N_2883,N_2930);
nor U3171 (N_3171,N_2970,N_2903);
xor U3172 (N_3172,N_2894,N_2989);
and U3173 (N_3173,N_2959,N_2980);
nor U3174 (N_3174,N_3017,N_2911);
nand U3175 (N_3175,N_2893,N_2970);
nand U3176 (N_3176,N_2969,N_2948);
and U3177 (N_3177,N_3031,N_2957);
nand U3178 (N_3178,N_2979,N_3018);
and U3179 (N_3179,N_2968,N_3014);
or U3180 (N_3180,N_2973,N_2943);
and U3181 (N_3181,N_2957,N_2943);
nand U3182 (N_3182,N_2993,N_2888);
or U3183 (N_3183,N_2927,N_2967);
or U3184 (N_3184,N_2994,N_2917);
nand U3185 (N_3185,N_2985,N_2896);
or U3186 (N_3186,N_2915,N_2984);
nand U3187 (N_3187,N_2954,N_2941);
and U3188 (N_3188,N_3004,N_3029);
or U3189 (N_3189,N_2882,N_2999);
nor U3190 (N_3190,N_3030,N_2880);
xnor U3191 (N_3191,N_2929,N_3038);
nand U3192 (N_3192,N_2945,N_3001);
nor U3193 (N_3193,N_2947,N_2898);
and U3194 (N_3194,N_2980,N_2945);
nand U3195 (N_3195,N_2944,N_2938);
xnor U3196 (N_3196,N_2917,N_3003);
or U3197 (N_3197,N_2910,N_3018);
and U3198 (N_3198,N_2936,N_2892);
or U3199 (N_3199,N_2931,N_2892);
and U3200 (N_3200,N_3187,N_3087);
and U3201 (N_3201,N_3044,N_3164);
nor U3202 (N_3202,N_3132,N_3048);
and U3203 (N_3203,N_3151,N_3056);
and U3204 (N_3204,N_3193,N_3145);
and U3205 (N_3205,N_3189,N_3139);
nand U3206 (N_3206,N_3176,N_3091);
xor U3207 (N_3207,N_3076,N_3188);
and U3208 (N_3208,N_3062,N_3052);
or U3209 (N_3209,N_3050,N_3088);
and U3210 (N_3210,N_3079,N_3089);
nand U3211 (N_3211,N_3110,N_3143);
nand U3212 (N_3212,N_3136,N_3147);
and U3213 (N_3213,N_3098,N_3179);
nor U3214 (N_3214,N_3158,N_3172);
nand U3215 (N_3215,N_3135,N_3043);
xnor U3216 (N_3216,N_3112,N_3129);
xnor U3217 (N_3217,N_3075,N_3073);
or U3218 (N_3218,N_3102,N_3178);
or U3219 (N_3219,N_3055,N_3183);
or U3220 (N_3220,N_3184,N_3111);
or U3221 (N_3221,N_3161,N_3053);
or U3222 (N_3222,N_3097,N_3197);
or U3223 (N_3223,N_3065,N_3094);
nand U3224 (N_3224,N_3131,N_3173);
or U3225 (N_3225,N_3182,N_3040);
and U3226 (N_3226,N_3051,N_3133);
nor U3227 (N_3227,N_3095,N_3061);
nand U3228 (N_3228,N_3163,N_3198);
xor U3229 (N_3229,N_3054,N_3185);
or U3230 (N_3230,N_3060,N_3066);
nand U3231 (N_3231,N_3138,N_3057);
or U3232 (N_3232,N_3175,N_3186);
or U3233 (N_3233,N_3195,N_3063);
or U3234 (N_3234,N_3083,N_3128);
nand U3235 (N_3235,N_3107,N_3149);
or U3236 (N_3236,N_3117,N_3162);
nor U3237 (N_3237,N_3191,N_3105);
nand U3238 (N_3238,N_3153,N_3096);
and U3239 (N_3239,N_3067,N_3086);
or U3240 (N_3240,N_3152,N_3130);
nor U3241 (N_3241,N_3082,N_3167);
xnor U3242 (N_3242,N_3146,N_3118);
nand U3243 (N_3243,N_3156,N_3114);
or U3244 (N_3244,N_3170,N_3155);
or U3245 (N_3245,N_3042,N_3140);
nand U3246 (N_3246,N_3159,N_3150);
xnor U3247 (N_3247,N_3174,N_3166);
nand U3248 (N_3248,N_3093,N_3092);
nand U3249 (N_3249,N_3119,N_3165);
nor U3250 (N_3250,N_3125,N_3141);
nor U3251 (N_3251,N_3148,N_3064);
or U3252 (N_3252,N_3071,N_3194);
nand U3253 (N_3253,N_3181,N_3134);
nor U3254 (N_3254,N_3122,N_3157);
and U3255 (N_3255,N_3106,N_3180);
nor U3256 (N_3256,N_3113,N_3070);
xor U3257 (N_3257,N_3104,N_3109);
xnor U3258 (N_3258,N_3090,N_3103);
or U3259 (N_3259,N_3099,N_3068);
or U3260 (N_3260,N_3059,N_3081);
and U3261 (N_3261,N_3069,N_3078);
and U3262 (N_3262,N_3137,N_3126);
xor U3263 (N_3263,N_3171,N_3058);
and U3264 (N_3264,N_3085,N_3080);
and U3265 (N_3265,N_3046,N_3123);
or U3266 (N_3266,N_3077,N_3144);
and U3267 (N_3267,N_3168,N_3041);
nor U3268 (N_3268,N_3154,N_3121);
and U3269 (N_3269,N_3124,N_3100);
and U3270 (N_3270,N_3116,N_3074);
xor U3271 (N_3271,N_3160,N_3115);
nor U3272 (N_3272,N_3072,N_3108);
nor U3273 (N_3273,N_3120,N_3196);
or U3274 (N_3274,N_3049,N_3127);
xor U3275 (N_3275,N_3169,N_3199);
nand U3276 (N_3276,N_3047,N_3192);
and U3277 (N_3277,N_3142,N_3101);
nand U3278 (N_3278,N_3190,N_3177);
nand U3279 (N_3279,N_3045,N_3084);
or U3280 (N_3280,N_3117,N_3198);
xnor U3281 (N_3281,N_3066,N_3052);
nand U3282 (N_3282,N_3064,N_3114);
nor U3283 (N_3283,N_3071,N_3129);
or U3284 (N_3284,N_3078,N_3138);
and U3285 (N_3285,N_3074,N_3054);
nor U3286 (N_3286,N_3066,N_3193);
nand U3287 (N_3287,N_3105,N_3125);
xnor U3288 (N_3288,N_3040,N_3099);
and U3289 (N_3289,N_3114,N_3106);
xor U3290 (N_3290,N_3065,N_3195);
nand U3291 (N_3291,N_3172,N_3121);
or U3292 (N_3292,N_3178,N_3041);
nor U3293 (N_3293,N_3174,N_3040);
nor U3294 (N_3294,N_3113,N_3138);
nor U3295 (N_3295,N_3098,N_3101);
nor U3296 (N_3296,N_3111,N_3088);
nand U3297 (N_3297,N_3051,N_3152);
and U3298 (N_3298,N_3143,N_3157);
or U3299 (N_3299,N_3083,N_3127);
nand U3300 (N_3300,N_3120,N_3058);
nor U3301 (N_3301,N_3184,N_3085);
nor U3302 (N_3302,N_3177,N_3127);
and U3303 (N_3303,N_3155,N_3104);
and U3304 (N_3304,N_3123,N_3073);
nand U3305 (N_3305,N_3049,N_3139);
nor U3306 (N_3306,N_3102,N_3073);
xnor U3307 (N_3307,N_3083,N_3087);
nand U3308 (N_3308,N_3092,N_3142);
nand U3309 (N_3309,N_3135,N_3156);
or U3310 (N_3310,N_3159,N_3165);
or U3311 (N_3311,N_3156,N_3053);
and U3312 (N_3312,N_3177,N_3158);
nor U3313 (N_3313,N_3085,N_3193);
nand U3314 (N_3314,N_3109,N_3153);
or U3315 (N_3315,N_3070,N_3059);
and U3316 (N_3316,N_3154,N_3095);
nor U3317 (N_3317,N_3149,N_3067);
or U3318 (N_3318,N_3196,N_3043);
and U3319 (N_3319,N_3063,N_3100);
and U3320 (N_3320,N_3151,N_3177);
and U3321 (N_3321,N_3063,N_3068);
or U3322 (N_3322,N_3095,N_3167);
and U3323 (N_3323,N_3105,N_3197);
nor U3324 (N_3324,N_3166,N_3195);
nand U3325 (N_3325,N_3143,N_3173);
nor U3326 (N_3326,N_3094,N_3149);
or U3327 (N_3327,N_3102,N_3046);
nand U3328 (N_3328,N_3119,N_3125);
nand U3329 (N_3329,N_3099,N_3083);
nor U3330 (N_3330,N_3053,N_3173);
nand U3331 (N_3331,N_3096,N_3117);
nand U3332 (N_3332,N_3057,N_3187);
nand U3333 (N_3333,N_3151,N_3185);
nor U3334 (N_3334,N_3129,N_3080);
nor U3335 (N_3335,N_3180,N_3056);
or U3336 (N_3336,N_3134,N_3071);
nor U3337 (N_3337,N_3072,N_3137);
and U3338 (N_3338,N_3129,N_3181);
nand U3339 (N_3339,N_3057,N_3113);
nor U3340 (N_3340,N_3058,N_3055);
nor U3341 (N_3341,N_3186,N_3194);
nand U3342 (N_3342,N_3141,N_3103);
nand U3343 (N_3343,N_3169,N_3159);
nor U3344 (N_3344,N_3185,N_3081);
nor U3345 (N_3345,N_3172,N_3076);
xnor U3346 (N_3346,N_3115,N_3132);
or U3347 (N_3347,N_3127,N_3159);
or U3348 (N_3348,N_3197,N_3184);
nor U3349 (N_3349,N_3100,N_3051);
nand U3350 (N_3350,N_3126,N_3054);
nor U3351 (N_3351,N_3175,N_3114);
nand U3352 (N_3352,N_3199,N_3085);
nor U3353 (N_3353,N_3072,N_3070);
nor U3354 (N_3354,N_3069,N_3092);
nor U3355 (N_3355,N_3054,N_3094);
or U3356 (N_3356,N_3057,N_3098);
nor U3357 (N_3357,N_3060,N_3125);
and U3358 (N_3358,N_3178,N_3155);
nand U3359 (N_3359,N_3164,N_3059);
or U3360 (N_3360,N_3211,N_3358);
nor U3361 (N_3361,N_3301,N_3205);
and U3362 (N_3362,N_3359,N_3352);
or U3363 (N_3363,N_3323,N_3214);
nand U3364 (N_3364,N_3217,N_3218);
and U3365 (N_3365,N_3200,N_3212);
nand U3366 (N_3366,N_3261,N_3342);
nor U3367 (N_3367,N_3259,N_3206);
xor U3368 (N_3368,N_3278,N_3327);
nor U3369 (N_3369,N_3265,N_3321);
nor U3370 (N_3370,N_3329,N_3247);
and U3371 (N_3371,N_3227,N_3286);
nor U3372 (N_3372,N_3273,N_3223);
xnor U3373 (N_3373,N_3209,N_3279);
nand U3374 (N_3374,N_3277,N_3350);
or U3375 (N_3375,N_3262,N_3233);
nand U3376 (N_3376,N_3220,N_3307);
and U3377 (N_3377,N_3341,N_3309);
nand U3378 (N_3378,N_3242,N_3238);
nor U3379 (N_3379,N_3331,N_3234);
and U3380 (N_3380,N_3231,N_3246);
nand U3381 (N_3381,N_3204,N_3337);
nand U3382 (N_3382,N_3219,N_3325);
and U3383 (N_3383,N_3201,N_3240);
or U3384 (N_3384,N_3208,N_3320);
and U3385 (N_3385,N_3239,N_3275);
or U3386 (N_3386,N_3312,N_3347);
nand U3387 (N_3387,N_3276,N_3272);
nand U3388 (N_3388,N_3299,N_3224);
nor U3389 (N_3389,N_3293,N_3292);
and U3390 (N_3390,N_3260,N_3317);
xnor U3391 (N_3391,N_3330,N_3351);
or U3392 (N_3392,N_3221,N_3213);
or U3393 (N_3393,N_3308,N_3335);
and U3394 (N_3394,N_3315,N_3300);
or U3395 (N_3395,N_3256,N_3289);
or U3396 (N_3396,N_3225,N_3266);
xnor U3397 (N_3397,N_3316,N_3241);
or U3398 (N_3398,N_3328,N_3270);
nor U3399 (N_3399,N_3314,N_3297);
nand U3400 (N_3400,N_3338,N_3343);
xor U3401 (N_3401,N_3303,N_3318);
or U3402 (N_3402,N_3295,N_3237);
and U3403 (N_3403,N_3348,N_3226);
and U3404 (N_3404,N_3228,N_3236);
nand U3405 (N_3405,N_3287,N_3339);
xnor U3406 (N_3406,N_3245,N_3355);
nand U3407 (N_3407,N_3306,N_3230);
or U3408 (N_3408,N_3357,N_3274);
or U3409 (N_3409,N_3305,N_3210);
and U3410 (N_3410,N_3222,N_3249);
nand U3411 (N_3411,N_3332,N_3284);
and U3412 (N_3412,N_3322,N_3254);
nor U3413 (N_3413,N_3294,N_3215);
or U3414 (N_3414,N_3244,N_3336);
and U3415 (N_3415,N_3258,N_3326);
xor U3416 (N_3416,N_3255,N_3288);
and U3417 (N_3417,N_3281,N_3344);
and U3418 (N_3418,N_3264,N_3304);
nand U3419 (N_3419,N_3285,N_3251);
or U3420 (N_3420,N_3229,N_3296);
or U3421 (N_3421,N_3291,N_3283);
and U3422 (N_3422,N_3203,N_3267);
or U3423 (N_3423,N_3356,N_3324);
xnor U3424 (N_3424,N_3302,N_3313);
and U3425 (N_3425,N_3345,N_3248);
nand U3426 (N_3426,N_3280,N_3268);
nand U3427 (N_3427,N_3250,N_3333);
or U3428 (N_3428,N_3319,N_3271);
nand U3429 (N_3429,N_3311,N_3202);
nand U3430 (N_3430,N_3334,N_3282);
and U3431 (N_3431,N_3353,N_3263);
nor U3432 (N_3432,N_3232,N_3257);
nand U3433 (N_3433,N_3346,N_3252);
nand U3434 (N_3434,N_3207,N_3290);
and U3435 (N_3435,N_3354,N_3243);
and U3436 (N_3436,N_3216,N_3340);
and U3437 (N_3437,N_3269,N_3310);
nor U3438 (N_3438,N_3235,N_3298);
nor U3439 (N_3439,N_3349,N_3253);
nand U3440 (N_3440,N_3247,N_3337);
nand U3441 (N_3441,N_3207,N_3238);
nor U3442 (N_3442,N_3288,N_3314);
nand U3443 (N_3443,N_3272,N_3204);
or U3444 (N_3444,N_3257,N_3285);
xnor U3445 (N_3445,N_3338,N_3232);
or U3446 (N_3446,N_3328,N_3243);
nand U3447 (N_3447,N_3286,N_3356);
nand U3448 (N_3448,N_3258,N_3247);
nand U3449 (N_3449,N_3247,N_3320);
or U3450 (N_3450,N_3251,N_3239);
xor U3451 (N_3451,N_3216,N_3257);
and U3452 (N_3452,N_3332,N_3237);
or U3453 (N_3453,N_3238,N_3261);
nand U3454 (N_3454,N_3258,N_3240);
and U3455 (N_3455,N_3307,N_3292);
nor U3456 (N_3456,N_3309,N_3344);
nor U3457 (N_3457,N_3268,N_3338);
or U3458 (N_3458,N_3231,N_3343);
nand U3459 (N_3459,N_3243,N_3349);
and U3460 (N_3460,N_3203,N_3330);
or U3461 (N_3461,N_3297,N_3323);
nor U3462 (N_3462,N_3294,N_3352);
nand U3463 (N_3463,N_3236,N_3266);
or U3464 (N_3464,N_3214,N_3302);
and U3465 (N_3465,N_3211,N_3204);
nor U3466 (N_3466,N_3237,N_3312);
nor U3467 (N_3467,N_3224,N_3316);
or U3468 (N_3468,N_3243,N_3325);
and U3469 (N_3469,N_3245,N_3289);
and U3470 (N_3470,N_3350,N_3270);
or U3471 (N_3471,N_3339,N_3315);
and U3472 (N_3472,N_3354,N_3355);
or U3473 (N_3473,N_3309,N_3204);
nor U3474 (N_3474,N_3311,N_3211);
or U3475 (N_3475,N_3282,N_3304);
and U3476 (N_3476,N_3260,N_3266);
nand U3477 (N_3477,N_3326,N_3346);
xor U3478 (N_3478,N_3217,N_3201);
or U3479 (N_3479,N_3310,N_3359);
nor U3480 (N_3480,N_3222,N_3304);
nor U3481 (N_3481,N_3348,N_3243);
and U3482 (N_3482,N_3292,N_3282);
nor U3483 (N_3483,N_3327,N_3260);
nor U3484 (N_3484,N_3295,N_3234);
xor U3485 (N_3485,N_3315,N_3243);
nand U3486 (N_3486,N_3348,N_3266);
nand U3487 (N_3487,N_3212,N_3221);
xor U3488 (N_3488,N_3354,N_3275);
or U3489 (N_3489,N_3313,N_3240);
nor U3490 (N_3490,N_3251,N_3313);
and U3491 (N_3491,N_3285,N_3302);
nor U3492 (N_3492,N_3267,N_3205);
nand U3493 (N_3493,N_3241,N_3273);
or U3494 (N_3494,N_3277,N_3240);
or U3495 (N_3495,N_3359,N_3235);
nand U3496 (N_3496,N_3323,N_3270);
nor U3497 (N_3497,N_3273,N_3315);
and U3498 (N_3498,N_3284,N_3232);
or U3499 (N_3499,N_3312,N_3336);
nor U3500 (N_3500,N_3314,N_3253);
or U3501 (N_3501,N_3310,N_3282);
nand U3502 (N_3502,N_3359,N_3295);
or U3503 (N_3503,N_3317,N_3211);
nand U3504 (N_3504,N_3317,N_3343);
xor U3505 (N_3505,N_3220,N_3261);
nor U3506 (N_3506,N_3215,N_3314);
nor U3507 (N_3507,N_3219,N_3347);
nand U3508 (N_3508,N_3282,N_3202);
nand U3509 (N_3509,N_3356,N_3219);
and U3510 (N_3510,N_3288,N_3259);
nand U3511 (N_3511,N_3305,N_3234);
or U3512 (N_3512,N_3307,N_3345);
and U3513 (N_3513,N_3235,N_3246);
and U3514 (N_3514,N_3213,N_3325);
nand U3515 (N_3515,N_3337,N_3319);
or U3516 (N_3516,N_3246,N_3234);
nor U3517 (N_3517,N_3339,N_3298);
or U3518 (N_3518,N_3312,N_3330);
nand U3519 (N_3519,N_3300,N_3231);
or U3520 (N_3520,N_3398,N_3484);
or U3521 (N_3521,N_3392,N_3381);
or U3522 (N_3522,N_3414,N_3486);
and U3523 (N_3523,N_3481,N_3434);
nand U3524 (N_3524,N_3431,N_3372);
nand U3525 (N_3525,N_3474,N_3453);
and U3526 (N_3526,N_3464,N_3378);
or U3527 (N_3527,N_3489,N_3497);
or U3528 (N_3528,N_3420,N_3502);
or U3529 (N_3529,N_3402,N_3461);
nor U3530 (N_3530,N_3468,N_3427);
nor U3531 (N_3531,N_3507,N_3360);
xor U3532 (N_3532,N_3394,N_3508);
and U3533 (N_3533,N_3476,N_3463);
or U3534 (N_3534,N_3475,N_3386);
and U3535 (N_3535,N_3487,N_3488);
or U3536 (N_3536,N_3383,N_3517);
nand U3537 (N_3537,N_3439,N_3501);
or U3538 (N_3538,N_3430,N_3495);
xnor U3539 (N_3539,N_3504,N_3388);
nand U3540 (N_3540,N_3365,N_3397);
or U3541 (N_3541,N_3385,N_3366);
nand U3542 (N_3542,N_3422,N_3456);
nor U3543 (N_3543,N_3515,N_3371);
or U3544 (N_3544,N_3432,N_3401);
and U3545 (N_3545,N_3417,N_3496);
nand U3546 (N_3546,N_3462,N_3438);
nand U3547 (N_3547,N_3425,N_3423);
xnor U3548 (N_3548,N_3480,N_3391);
and U3549 (N_3549,N_3406,N_3451);
or U3550 (N_3550,N_3426,N_3412);
nand U3551 (N_3551,N_3411,N_3516);
or U3552 (N_3552,N_3492,N_3369);
nand U3553 (N_3553,N_3446,N_3447);
or U3554 (N_3554,N_3400,N_3440);
nand U3555 (N_3555,N_3419,N_3377);
or U3556 (N_3556,N_3409,N_3498);
or U3557 (N_3557,N_3513,N_3429);
or U3558 (N_3558,N_3408,N_3441);
and U3559 (N_3559,N_3393,N_3465);
or U3560 (N_3560,N_3380,N_3505);
or U3561 (N_3561,N_3494,N_3506);
or U3562 (N_3562,N_3467,N_3473);
and U3563 (N_3563,N_3384,N_3491);
and U3564 (N_3564,N_3483,N_3510);
and U3565 (N_3565,N_3454,N_3477);
nand U3566 (N_3566,N_3458,N_3437);
xor U3567 (N_3567,N_3466,N_3449);
nor U3568 (N_3568,N_3500,N_3367);
or U3569 (N_3569,N_3389,N_3416);
or U3570 (N_3570,N_3485,N_3452);
nand U3571 (N_3571,N_3424,N_3433);
nor U3572 (N_3572,N_3509,N_3403);
or U3573 (N_3573,N_3364,N_3435);
or U3574 (N_3574,N_3373,N_3444);
xnor U3575 (N_3575,N_3404,N_3457);
or U3576 (N_3576,N_3472,N_3442);
nand U3577 (N_3577,N_3436,N_3512);
nand U3578 (N_3578,N_3363,N_3418);
nor U3579 (N_3579,N_3407,N_3514);
nor U3580 (N_3580,N_3382,N_3459);
nor U3581 (N_3581,N_3379,N_3362);
nor U3582 (N_3582,N_3415,N_3375);
nor U3583 (N_3583,N_3519,N_3511);
nand U3584 (N_3584,N_3368,N_3387);
or U3585 (N_3585,N_3503,N_3479);
and U3586 (N_3586,N_3361,N_3490);
nand U3587 (N_3587,N_3443,N_3460);
or U3588 (N_3588,N_3374,N_3499);
nor U3589 (N_3589,N_3395,N_3445);
nor U3590 (N_3590,N_3421,N_3428);
or U3591 (N_3591,N_3448,N_3390);
or U3592 (N_3592,N_3396,N_3471);
or U3593 (N_3593,N_3370,N_3482);
nand U3594 (N_3594,N_3469,N_3450);
and U3595 (N_3595,N_3413,N_3470);
nand U3596 (N_3596,N_3410,N_3376);
and U3597 (N_3597,N_3518,N_3399);
or U3598 (N_3598,N_3478,N_3405);
nand U3599 (N_3599,N_3455,N_3493);
or U3600 (N_3600,N_3506,N_3366);
and U3601 (N_3601,N_3449,N_3512);
and U3602 (N_3602,N_3369,N_3486);
or U3603 (N_3603,N_3463,N_3401);
xnor U3604 (N_3604,N_3440,N_3404);
nor U3605 (N_3605,N_3428,N_3454);
nor U3606 (N_3606,N_3505,N_3444);
nor U3607 (N_3607,N_3514,N_3379);
and U3608 (N_3608,N_3513,N_3442);
xnor U3609 (N_3609,N_3485,N_3429);
nor U3610 (N_3610,N_3466,N_3380);
nor U3611 (N_3611,N_3496,N_3423);
and U3612 (N_3612,N_3390,N_3437);
nand U3613 (N_3613,N_3402,N_3487);
nor U3614 (N_3614,N_3479,N_3445);
nand U3615 (N_3615,N_3420,N_3470);
or U3616 (N_3616,N_3411,N_3492);
nor U3617 (N_3617,N_3519,N_3437);
or U3618 (N_3618,N_3481,N_3376);
nor U3619 (N_3619,N_3463,N_3448);
and U3620 (N_3620,N_3458,N_3469);
nand U3621 (N_3621,N_3471,N_3512);
nand U3622 (N_3622,N_3409,N_3439);
nor U3623 (N_3623,N_3388,N_3392);
and U3624 (N_3624,N_3391,N_3369);
and U3625 (N_3625,N_3414,N_3367);
nand U3626 (N_3626,N_3506,N_3397);
nor U3627 (N_3627,N_3414,N_3364);
nor U3628 (N_3628,N_3516,N_3509);
and U3629 (N_3629,N_3442,N_3383);
nand U3630 (N_3630,N_3518,N_3431);
nand U3631 (N_3631,N_3449,N_3370);
nand U3632 (N_3632,N_3398,N_3427);
nor U3633 (N_3633,N_3463,N_3411);
nor U3634 (N_3634,N_3408,N_3428);
and U3635 (N_3635,N_3426,N_3370);
nor U3636 (N_3636,N_3486,N_3447);
nor U3637 (N_3637,N_3480,N_3518);
xor U3638 (N_3638,N_3483,N_3465);
or U3639 (N_3639,N_3478,N_3402);
nand U3640 (N_3640,N_3511,N_3410);
nor U3641 (N_3641,N_3514,N_3366);
nand U3642 (N_3642,N_3427,N_3445);
xor U3643 (N_3643,N_3446,N_3485);
nand U3644 (N_3644,N_3483,N_3402);
nor U3645 (N_3645,N_3367,N_3438);
or U3646 (N_3646,N_3381,N_3474);
nand U3647 (N_3647,N_3510,N_3414);
and U3648 (N_3648,N_3381,N_3360);
nand U3649 (N_3649,N_3435,N_3379);
nor U3650 (N_3650,N_3413,N_3477);
nand U3651 (N_3651,N_3376,N_3482);
nand U3652 (N_3652,N_3396,N_3498);
nor U3653 (N_3653,N_3495,N_3463);
nand U3654 (N_3654,N_3468,N_3388);
nor U3655 (N_3655,N_3462,N_3366);
nand U3656 (N_3656,N_3500,N_3451);
and U3657 (N_3657,N_3430,N_3403);
nor U3658 (N_3658,N_3490,N_3395);
nand U3659 (N_3659,N_3456,N_3362);
and U3660 (N_3660,N_3392,N_3477);
nor U3661 (N_3661,N_3468,N_3497);
or U3662 (N_3662,N_3501,N_3516);
or U3663 (N_3663,N_3434,N_3424);
and U3664 (N_3664,N_3507,N_3420);
xnor U3665 (N_3665,N_3471,N_3495);
and U3666 (N_3666,N_3363,N_3517);
or U3667 (N_3667,N_3453,N_3402);
nand U3668 (N_3668,N_3416,N_3435);
or U3669 (N_3669,N_3454,N_3516);
nand U3670 (N_3670,N_3436,N_3505);
or U3671 (N_3671,N_3431,N_3435);
nand U3672 (N_3672,N_3476,N_3499);
xnor U3673 (N_3673,N_3407,N_3509);
or U3674 (N_3674,N_3464,N_3441);
nand U3675 (N_3675,N_3448,N_3467);
xor U3676 (N_3676,N_3412,N_3513);
nor U3677 (N_3677,N_3408,N_3378);
nand U3678 (N_3678,N_3377,N_3364);
nor U3679 (N_3679,N_3498,N_3402);
nand U3680 (N_3680,N_3569,N_3532);
or U3681 (N_3681,N_3677,N_3523);
nand U3682 (N_3682,N_3576,N_3587);
nor U3683 (N_3683,N_3536,N_3660);
nor U3684 (N_3684,N_3675,N_3641);
and U3685 (N_3685,N_3570,N_3559);
nor U3686 (N_3686,N_3657,N_3648);
nor U3687 (N_3687,N_3522,N_3527);
nor U3688 (N_3688,N_3666,N_3543);
or U3689 (N_3689,N_3679,N_3628);
nand U3690 (N_3690,N_3602,N_3598);
nand U3691 (N_3691,N_3638,N_3613);
nand U3692 (N_3692,N_3632,N_3573);
or U3693 (N_3693,N_3642,N_3610);
or U3694 (N_3694,N_3562,N_3603);
and U3695 (N_3695,N_3678,N_3564);
xor U3696 (N_3696,N_3647,N_3551);
nand U3697 (N_3697,N_3579,N_3637);
nand U3698 (N_3698,N_3563,N_3634);
nor U3699 (N_3699,N_3618,N_3595);
nor U3700 (N_3700,N_3676,N_3542);
or U3701 (N_3701,N_3663,N_3534);
or U3702 (N_3702,N_3629,N_3670);
and U3703 (N_3703,N_3636,N_3578);
and U3704 (N_3704,N_3599,N_3558);
and U3705 (N_3705,N_3528,N_3565);
or U3706 (N_3706,N_3631,N_3656);
nand U3707 (N_3707,N_3635,N_3549);
xnor U3708 (N_3708,N_3623,N_3651);
and U3709 (N_3709,N_3530,N_3616);
xnor U3710 (N_3710,N_3545,N_3659);
or U3711 (N_3711,N_3667,N_3548);
nor U3712 (N_3712,N_3661,N_3652);
and U3713 (N_3713,N_3557,N_3664);
nand U3714 (N_3714,N_3662,N_3673);
nor U3715 (N_3715,N_3584,N_3571);
nand U3716 (N_3716,N_3553,N_3619);
or U3717 (N_3717,N_3640,N_3669);
xor U3718 (N_3718,N_3531,N_3653);
xor U3719 (N_3719,N_3566,N_3540);
and U3720 (N_3720,N_3655,N_3606);
and U3721 (N_3721,N_3541,N_3555);
nor U3722 (N_3722,N_3521,N_3649);
and U3723 (N_3723,N_3544,N_3538);
nor U3724 (N_3724,N_3581,N_3525);
or U3725 (N_3725,N_3533,N_3547);
nand U3726 (N_3726,N_3630,N_3537);
nand U3727 (N_3727,N_3620,N_3672);
or U3728 (N_3728,N_3665,N_3607);
nor U3729 (N_3729,N_3609,N_3592);
nand U3730 (N_3730,N_3572,N_3526);
or U3731 (N_3731,N_3582,N_3552);
and U3732 (N_3732,N_3535,N_3593);
nand U3733 (N_3733,N_3554,N_3546);
nor U3734 (N_3734,N_3529,N_3600);
nand U3735 (N_3735,N_3626,N_3577);
xnor U3736 (N_3736,N_3646,N_3560);
and U3737 (N_3737,N_3550,N_3575);
nand U3738 (N_3738,N_3596,N_3624);
and U3739 (N_3739,N_3586,N_3633);
or U3740 (N_3740,N_3605,N_3539);
and U3741 (N_3741,N_3621,N_3625);
nand U3742 (N_3742,N_3644,N_3597);
or U3743 (N_3743,N_3561,N_3520);
and U3744 (N_3744,N_3601,N_3583);
or U3745 (N_3745,N_3568,N_3671);
or U3746 (N_3746,N_3574,N_3604);
xnor U3747 (N_3747,N_3611,N_3650);
or U3748 (N_3748,N_3588,N_3591);
xor U3749 (N_3749,N_3654,N_3580);
nor U3750 (N_3750,N_3585,N_3639);
nand U3751 (N_3751,N_3594,N_3617);
nand U3752 (N_3752,N_3556,N_3612);
and U3753 (N_3753,N_3524,N_3614);
nor U3754 (N_3754,N_3590,N_3567);
nand U3755 (N_3755,N_3615,N_3658);
nor U3756 (N_3756,N_3668,N_3622);
or U3757 (N_3757,N_3608,N_3643);
nand U3758 (N_3758,N_3627,N_3645);
nand U3759 (N_3759,N_3589,N_3674);
xnor U3760 (N_3760,N_3607,N_3580);
xnor U3761 (N_3761,N_3534,N_3675);
and U3762 (N_3762,N_3633,N_3530);
nor U3763 (N_3763,N_3555,N_3533);
xor U3764 (N_3764,N_3624,N_3552);
and U3765 (N_3765,N_3520,N_3544);
or U3766 (N_3766,N_3553,N_3650);
or U3767 (N_3767,N_3523,N_3581);
and U3768 (N_3768,N_3632,N_3675);
and U3769 (N_3769,N_3597,N_3661);
nor U3770 (N_3770,N_3554,N_3614);
or U3771 (N_3771,N_3609,N_3570);
or U3772 (N_3772,N_3671,N_3600);
and U3773 (N_3773,N_3569,N_3552);
or U3774 (N_3774,N_3642,N_3592);
nand U3775 (N_3775,N_3601,N_3618);
nor U3776 (N_3776,N_3559,N_3586);
and U3777 (N_3777,N_3660,N_3674);
and U3778 (N_3778,N_3678,N_3590);
nor U3779 (N_3779,N_3570,N_3533);
nand U3780 (N_3780,N_3623,N_3637);
xnor U3781 (N_3781,N_3635,N_3558);
nand U3782 (N_3782,N_3588,N_3558);
nor U3783 (N_3783,N_3670,N_3628);
nor U3784 (N_3784,N_3553,N_3546);
and U3785 (N_3785,N_3529,N_3537);
or U3786 (N_3786,N_3623,N_3572);
nand U3787 (N_3787,N_3633,N_3532);
and U3788 (N_3788,N_3642,N_3525);
and U3789 (N_3789,N_3661,N_3676);
or U3790 (N_3790,N_3535,N_3621);
and U3791 (N_3791,N_3663,N_3564);
and U3792 (N_3792,N_3663,N_3522);
nand U3793 (N_3793,N_3670,N_3586);
xnor U3794 (N_3794,N_3610,N_3677);
nand U3795 (N_3795,N_3615,N_3657);
nor U3796 (N_3796,N_3558,N_3641);
xnor U3797 (N_3797,N_3553,N_3617);
nor U3798 (N_3798,N_3573,N_3663);
xnor U3799 (N_3799,N_3587,N_3549);
nand U3800 (N_3800,N_3521,N_3588);
and U3801 (N_3801,N_3674,N_3656);
or U3802 (N_3802,N_3678,N_3574);
nand U3803 (N_3803,N_3537,N_3602);
nor U3804 (N_3804,N_3577,N_3617);
or U3805 (N_3805,N_3534,N_3624);
or U3806 (N_3806,N_3540,N_3592);
nand U3807 (N_3807,N_3595,N_3626);
nand U3808 (N_3808,N_3616,N_3542);
nor U3809 (N_3809,N_3652,N_3578);
nand U3810 (N_3810,N_3663,N_3571);
nand U3811 (N_3811,N_3595,N_3607);
or U3812 (N_3812,N_3561,N_3671);
or U3813 (N_3813,N_3587,N_3531);
and U3814 (N_3814,N_3647,N_3576);
or U3815 (N_3815,N_3629,N_3575);
nor U3816 (N_3816,N_3555,N_3557);
nor U3817 (N_3817,N_3548,N_3656);
or U3818 (N_3818,N_3630,N_3625);
and U3819 (N_3819,N_3539,N_3631);
or U3820 (N_3820,N_3578,N_3602);
nand U3821 (N_3821,N_3676,N_3574);
nor U3822 (N_3822,N_3544,N_3619);
and U3823 (N_3823,N_3664,N_3537);
nand U3824 (N_3824,N_3637,N_3606);
and U3825 (N_3825,N_3525,N_3539);
nand U3826 (N_3826,N_3663,N_3641);
or U3827 (N_3827,N_3540,N_3647);
or U3828 (N_3828,N_3530,N_3541);
xor U3829 (N_3829,N_3527,N_3669);
and U3830 (N_3830,N_3657,N_3566);
and U3831 (N_3831,N_3548,N_3645);
or U3832 (N_3832,N_3612,N_3575);
and U3833 (N_3833,N_3596,N_3660);
nor U3834 (N_3834,N_3558,N_3637);
nand U3835 (N_3835,N_3645,N_3555);
and U3836 (N_3836,N_3543,N_3566);
nor U3837 (N_3837,N_3594,N_3655);
and U3838 (N_3838,N_3536,N_3610);
nor U3839 (N_3839,N_3555,N_3674);
nand U3840 (N_3840,N_3737,N_3747);
nor U3841 (N_3841,N_3744,N_3755);
and U3842 (N_3842,N_3716,N_3710);
and U3843 (N_3843,N_3812,N_3714);
and U3844 (N_3844,N_3801,N_3767);
or U3845 (N_3845,N_3695,N_3732);
nand U3846 (N_3846,N_3826,N_3785);
or U3847 (N_3847,N_3762,N_3823);
nor U3848 (N_3848,N_3774,N_3795);
nor U3849 (N_3849,N_3736,N_3715);
or U3850 (N_3850,N_3752,N_3698);
nor U3851 (N_3851,N_3775,N_3753);
nand U3852 (N_3852,N_3726,N_3769);
nand U3853 (N_3853,N_3822,N_3798);
nand U3854 (N_3854,N_3711,N_3790);
nand U3855 (N_3855,N_3702,N_3800);
and U3856 (N_3856,N_3838,N_3764);
nand U3857 (N_3857,N_3771,N_3742);
and U3858 (N_3858,N_3814,N_3789);
nor U3859 (N_3859,N_3787,N_3685);
or U3860 (N_3860,N_3799,N_3712);
xor U3861 (N_3861,N_3796,N_3824);
and U3862 (N_3862,N_3827,N_3751);
nand U3863 (N_3863,N_3761,N_3835);
nor U3864 (N_3864,N_3765,N_3797);
nor U3865 (N_3865,N_3692,N_3815);
and U3866 (N_3866,N_3721,N_3779);
or U3867 (N_3867,N_3805,N_3703);
or U3868 (N_3868,N_3707,N_3748);
nor U3869 (N_3869,N_3810,N_3794);
nand U3870 (N_3870,N_3809,N_3719);
nor U3871 (N_3871,N_3836,N_3746);
and U3872 (N_3872,N_3723,N_3689);
or U3873 (N_3873,N_3696,N_3724);
nor U3874 (N_3874,N_3788,N_3777);
xnor U3875 (N_3875,N_3706,N_3701);
nor U3876 (N_3876,N_3727,N_3807);
nor U3877 (N_3877,N_3757,N_3820);
nor U3878 (N_3878,N_3694,N_3704);
or U3879 (N_3879,N_3735,N_3759);
or U3880 (N_3880,N_3828,N_3718);
xnor U3881 (N_3881,N_3816,N_3782);
nand U3882 (N_3882,N_3784,N_3776);
and U3883 (N_3883,N_3722,N_3690);
nor U3884 (N_3884,N_3763,N_3684);
or U3885 (N_3885,N_3803,N_3740);
nor U3886 (N_3886,N_3745,N_3758);
xor U3887 (N_3887,N_3832,N_3766);
nor U3888 (N_3888,N_3756,N_3699);
or U3889 (N_3889,N_3729,N_3708);
nor U3890 (N_3890,N_3697,N_3780);
nand U3891 (N_3891,N_3817,N_3831);
xnor U3892 (N_3892,N_3837,N_3713);
nand U3893 (N_3893,N_3786,N_3773);
nand U3894 (N_3894,N_3686,N_3730);
nor U3895 (N_3895,N_3680,N_3783);
nand U3896 (N_3896,N_3821,N_3739);
and U3897 (N_3897,N_3829,N_3770);
or U3898 (N_3898,N_3772,N_3819);
or U3899 (N_3899,N_3720,N_3808);
xor U3900 (N_3900,N_3833,N_3682);
nor U3901 (N_3901,N_3793,N_3717);
and U3902 (N_3902,N_3728,N_3768);
and U3903 (N_3903,N_3839,N_3693);
xor U3904 (N_3904,N_3749,N_3683);
and U3905 (N_3905,N_3818,N_3802);
and U3906 (N_3906,N_3733,N_3792);
nor U3907 (N_3907,N_3811,N_3806);
or U3908 (N_3908,N_3738,N_3813);
nor U3909 (N_3909,N_3743,N_3754);
nor U3910 (N_3910,N_3700,N_3687);
and U3911 (N_3911,N_3688,N_3830);
nand U3912 (N_3912,N_3705,N_3681);
and U3913 (N_3913,N_3804,N_3781);
xnor U3914 (N_3914,N_3691,N_3760);
and U3915 (N_3915,N_3734,N_3731);
nor U3916 (N_3916,N_3825,N_3750);
or U3917 (N_3917,N_3725,N_3791);
nor U3918 (N_3918,N_3834,N_3778);
nand U3919 (N_3919,N_3741,N_3709);
or U3920 (N_3920,N_3701,N_3760);
or U3921 (N_3921,N_3837,N_3815);
and U3922 (N_3922,N_3698,N_3728);
or U3923 (N_3923,N_3761,N_3823);
and U3924 (N_3924,N_3787,N_3797);
nor U3925 (N_3925,N_3686,N_3774);
and U3926 (N_3926,N_3837,N_3791);
and U3927 (N_3927,N_3680,N_3816);
nor U3928 (N_3928,N_3694,N_3761);
nor U3929 (N_3929,N_3787,N_3721);
xor U3930 (N_3930,N_3839,N_3681);
xnor U3931 (N_3931,N_3778,N_3786);
nand U3932 (N_3932,N_3755,N_3828);
nand U3933 (N_3933,N_3760,N_3784);
nor U3934 (N_3934,N_3836,N_3795);
xor U3935 (N_3935,N_3704,N_3762);
nand U3936 (N_3936,N_3803,N_3719);
nor U3937 (N_3937,N_3773,N_3712);
or U3938 (N_3938,N_3685,N_3690);
nor U3939 (N_3939,N_3753,N_3792);
nor U3940 (N_3940,N_3681,N_3795);
nand U3941 (N_3941,N_3724,N_3770);
nand U3942 (N_3942,N_3789,N_3802);
nor U3943 (N_3943,N_3832,N_3839);
nand U3944 (N_3944,N_3705,N_3751);
or U3945 (N_3945,N_3732,N_3837);
nand U3946 (N_3946,N_3837,N_3783);
xnor U3947 (N_3947,N_3811,N_3707);
xnor U3948 (N_3948,N_3797,N_3810);
xor U3949 (N_3949,N_3764,N_3834);
nand U3950 (N_3950,N_3686,N_3832);
or U3951 (N_3951,N_3702,N_3684);
nand U3952 (N_3952,N_3818,N_3731);
nand U3953 (N_3953,N_3786,N_3771);
and U3954 (N_3954,N_3798,N_3764);
and U3955 (N_3955,N_3819,N_3724);
nor U3956 (N_3956,N_3754,N_3775);
or U3957 (N_3957,N_3801,N_3784);
and U3958 (N_3958,N_3736,N_3831);
nand U3959 (N_3959,N_3820,N_3832);
and U3960 (N_3960,N_3754,N_3777);
nand U3961 (N_3961,N_3814,N_3784);
nor U3962 (N_3962,N_3778,N_3686);
nor U3963 (N_3963,N_3718,N_3687);
and U3964 (N_3964,N_3740,N_3695);
xnor U3965 (N_3965,N_3746,N_3741);
and U3966 (N_3966,N_3736,N_3802);
nand U3967 (N_3967,N_3772,N_3747);
nand U3968 (N_3968,N_3814,N_3728);
or U3969 (N_3969,N_3685,N_3795);
or U3970 (N_3970,N_3785,N_3750);
or U3971 (N_3971,N_3748,N_3811);
or U3972 (N_3972,N_3778,N_3820);
or U3973 (N_3973,N_3716,N_3727);
nor U3974 (N_3974,N_3717,N_3781);
or U3975 (N_3975,N_3743,N_3697);
nor U3976 (N_3976,N_3825,N_3745);
and U3977 (N_3977,N_3783,N_3687);
nor U3978 (N_3978,N_3750,N_3789);
nor U3979 (N_3979,N_3691,N_3806);
nand U3980 (N_3980,N_3743,N_3768);
or U3981 (N_3981,N_3761,N_3759);
nor U3982 (N_3982,N_3704,N_3707);
nand U3983 (N_3983,N_3697,N_3745);
nor U3984 (N_3984,N_3812,N_3735);
nand U3985 (N_3985,N_3686,N_3834);
nand U3986 (N_3986,N_3755,N_3757);
and U3987 (N_3987,N_3749,N_3715);
and U3988 (N_3988,N_3795,N_3827);
nor U3989 (N_3989,N_3697,N_3681);
or U3990 (N_3990,N_3803,N_3819);
or U3991 (N_3991,N_3808,N_3710);
or U3992 (N_3992,N_3723,N_3756);
nor U3993 (N_3993,N_3799,N_3768);
nand U3994 (N_3994,N_3774,N_3740);
nor U3995 (N_3995,N_3686,N_3702);
nor U3996 (N_3996,N_3762,N_3781);
or U3997 (N_3997,N_3804,N_3717);
nand U3998 (N_3998,N_3750,N_3804);
or U3999 (N_3999,N_3708,N_3761);
and U4000 (N_4000,N_3908,N_3850);
or U4001 (N_4001,N_3918,N_3866);
and U4002 (N_4002,N_3916,N_3891);
nor U4003 (N_4003,N_3925,N_3898);
or U4004 (N_4004,N_3893,N_3942);
and U4005 (N_4005,N_3902,N_3894);
or U4006 (N_4006,N_3992,N_3962);
or U4007 (N_4007,N_3959,N_3924);
and U4008 (N_4008,N_3896,N_3871);
or U4009 (N_4009,N_3886,N_3951);
nand U4010 (N_4010,N_3984,N_3989);
or U4011 (N_4011,N_3848,N_3952);
or U4012 (N_4012,N_3980,N_3867);
and U4013 (N_4013,N_3844,N_3999);
and U4014 (N_4014,N_3865,N_3889);
nor U4015 (N_4015,N_3983,N_3993);
nor U4016 (N_4016,N_3953,N_3978);
nor U4017 (N_4017,N_3849,N_3931);
nand U4018 (N_4018,N_3917,N_3900);
and U4019 (N_4019,N_3970,N_3873);
and U4020 (N_4020,N_3846,N_3915);
nand U4021 (N_4021,N_3858,N_3859);
xnor U4022 (N_4022,N_3957,N_3905);
nand U4023 (N_4023,N_3937,N_3897);
nand U4024 (N_4024,N_3960,N_3947);
and U4025 (N_4025,N_3941,N_3964);
nor U4026 (N_4026,N_3996,N_3880);
and U4027 (N_4027,N_3914,N_3876);
nand U4028 (N_4028,N_3990,N_3911);
or U4029 (N_4029,N_3988,N_3856);
and U4030 (N_4030,N_3926,N_3863);
nand U4031 (N_4031,N_3869,N_3855);
and U4032 (N_4032,N_3935,N_3994);
and U4033 (N_4033,N_3982,N_3934);
nor U4034 (N_4034,N_3868,N_3930);
or U4035 (N_4035,N_3861,N_3965);
nand U4036 (N_4036,N_3938,N_3909);
nand U4037 (N_4037,N_3847,N_3963);
nand U4038 (N_4038,N_3946,N_3879);
and U4039 (N_4039,N_3864,N_3899);
or U4040 (N_4040,N_3854,N_3985);
and U4041 (N_4041,N_3885,N_3874);
and U4042 (N_4042,N_3921,N_3969);
nand U4043 (N_4043,N_3943,N_3906);
nor U4044 (N_4044,N_3881,N_3981);
nor U4045 (N_4045,N_3950,N_3961);
and U4046 (N_4046,N_3903,N_3966);
nand U4047 (N_4047,N_3976,N_3878);
or U4048 (N_4048,N_3888,N_3932);
and U4049 (N_4049,N_3842,N_3877);
and U4050 (N_4050,N_3945,N_3927);
nand U4051 (N_4051,N_3928,N_3933);
or U4052 (N_4052,N_3956,N_3910);
or U4053 (N_4053,N_3912,N_3939);
nand U4054 (N_4054,N_3870,N_3901);
nor U4055 (N_4055,N_3954,N_3967);
and U4056 (N_4056,N_3919,N_3944);
nand U4057 (N_4057,N_3958,N_3973);
or U4058 (N_4058,N_3841,N_3920);
and U4059 (N_4059,N_3936,N_3857);
and U4060 (N_4060,N_3860,N_3875);
nand U4061 (N_4061,N_3995,N_3845);
xnor U4062 (N_4062,N_3974,N_3907);
nor U4063 (N_4063,N_3977,N_3840);
and U4064 (N_4064,N_3986,N_3872);
nand U4065 (N_4065,N_3968,N_3923);
nand U4066 (N_4066,N_3987,N_3975);
nand U4067 (N_4067,N_3862,N_3972);
and U4068 (N_4068,N_3929,N_3884);
nor U4069 (N_4069,N_3851,N_3913);
nand U4070 (N_4070,N_3997,N_3979);
and U4071 (N_4071,N_3971,N_3895);
and U4072 (N_4072,N_3887,N_3998);
or U4073 (N_4073,N_3883,N_3991);
nor U4074 (N_4074,N_3940,N_3852);
nand U4075 (N_4075,N_3904,N_3922);
nand U4076 (N_4076,N_3890,N_3955);
or U4077 (N_4077,N_3949,N_3853);
nand U4078 (N_4078,N_3882,N_3843);
nor U4079 (N_4079,N_3892,N_3948);
xor U4080 (N_4080,N_3846,N_3890);
and U4081 (N_4081,N_3898,N_3863);
and U4082 (N_4082,N_3922,N_3899);
or U4083 (N_4083,N_3960,N_3939);
nor U4084 (N_4084,N_3847,N_3869);
nor U4085 (N_4085,N_3992,N_3881);
nand U4086 (N_4086,N_3963,N_3841);
nor U4087 (N_4087,N_3865,N_3870);
nor U4088 (N_4088,N_3952,N_3936);
nand U4089 (N_4089,N_3962,N_3945);
nor U4090 (N_4090,N_3850,N_3897);
or U4091 (N_4091,N_3993,N_3936);
or U4092 (N_4092,N_3895,N_3893);
or U4093 (N_4093,N_3904,N_3867);
or U4094 (N_4094,N_3868,N_3956);
nand U4095 (N_4095,N_3933,N_3876);
xor U4096 (N_4096,N_3872,N_3862);
nor U4097 (N_4097,N_3907,N_3855);
or U4098 (N_4098,N_3862,N_3961);
nand U4099 (N_4099,N_3843,N_3910);
nand U4100 (N_4100,N_3893,N_3948);
or U4101 (N_4101,N_3843,N_3915);
nor U4102 (N_4102,N_3879,N_3866);
or U4103 (N_4103,N_3945,N_3912);
nor U4104 (N_4104,N_3922,N_3849);
nor U4105 (N_4105,N_3946,N_3899);
or U4106 (N_4106,N_3952,N_3964);
and U4107 (N_4107,N_3914,N_3972);
and U4108 (N_4108,N_3851,N_3929);
or U4109 (N_4109,N_3855,N_3850);
xnor U4110 (N_4110,N_3884,N_3994);
and U4111 (N_4111,N_3915,N_3958);
nor U4112 (N_4112,N_3968,N_3901);
nor U4113 (N_4113,N_3867,N_3918);
xnor U4114 (N_4114,N_3934,N_3941);
xnor U4115 (N_4115,N_3894,N_3856);
or U4116 (N_4116,N_3935,N_3984);
nand U4117 (N_4117,N_3990,N_3840);
nor U4118 (N_4118,N_3877,N_3988);
nor U4119 (N_4119,N_3916,N_3969);
or U4120 (N_4120,N_3922,N_3989);
nor U4121 (N_4121,N_3841,N_3857);
xor U4122 (N_4122,N_3940,N_3925);
nand U4123 (N_4123,N_3912,N_3980);
nor U4124 (N_4124,N_3868,N_3900);
or U4125 (N_4125,N_3894,N_3855);
nand U4126 (N_4126,N_3968,N_3876);
nor U4127 (N_4127,N_3947,N_3845);
nor U4128 (N_4128,N_3901,N_3969);
nand U4129 (N_4129,N_3900,N_3990);
and U4130 (N_4130,N_3964,N_3929);
xnor U4131 (N_4131,N_3922,N_3874);
or U4132 (N_4132,N_3962,N_3986);
nand U4133 (N_4133,N_3876,N_3911);
and U4134 (N_4134,N_3899,N_3846);
and U4135 (N_4135,N_3939,N_3937);
and U4136 (N_4136,N_3960,N_3850);
or U4137 (N_4137,N_3938,N_3923);
nor U4138 (N_4138,N_3925,N_3858);
or U4139 (N_4139,N_3891,N_3863);
nor U4140 (N_4140,N_3925,N_3981);
nor U4141 (N_4141,N_3981,N_3965);
or U4142 (N_4142,N_3852,N_3945);
nand U4143 (N_4143,N_3946,N_3887);
and U4144 (N_4144,N_3960,N_3854);
and U4145 (N_4145,N_3991,N_3925);
nor U4146 (N_4146,N_3973,N_3971);
nor U4147 (N_4147,N_3977,N_3901);
or U4148 (N_4148,N_3905,N_3847);
nor U4149 (N_4149,N_3915,N_3947);
or U4150 (N_4150,N_3968,N_3948);
nor U4151 (N_4151,N_3997,N_3938);
xnor U4152 (N_4152,N_3878,N_3855);
nand U4153 (N_4153,N_3860,N_3858);
nor U4154 (N_4154,N_3910,N_3914);
nand U4155 (N_4155,N_3898,N_3963);
nor U4156 (N_4156,N_3917,N_3977);
nor U4157 (N_4157,N_3880,N_3977);
or U4158 (N_4158,N_3995,N_3994);
nand U4159 (N_4159,N_3935,N_3946);
nor U4160 (N_4160,N_4143,N_4073);
or U4161 (N_4161,N_4026,N_4035);
or U4162 (N_4162,N_4136,N_4011);
or U4163 (N_4163,N_4030,N_4079);
and U4164 (N_4164,N_4146,N_4099);
nand U4165 (N_4165,N_4066,N_4008);
nand U4166 (N_4166,N_4129,N_4157);
nor U4167 (N_4167,N_4102,N_4092);
nor U4168 (N_4168,N_4023,N_4012);
and U4169 (N_4169,N_4059,N_4056);
and U4170 (N_4170,N_4044,N_4050);
and U4171 (N_4171,N_4154,N_4126);
and U4172 (N_4172,N_4104,N_4018);
nor U4173 (N_4173,N_4027,N_4013);
and U4174 (N_4174,N_4045,N_4070);
xnor U4175 (N_4175,N_4139,N_4151);
or U4176 (N_4176,N_4114,N_4020);
nand U4177 (N_4177,N_4071,N_4113);
nor U4178 (N_4178,N_4119,N_4004);
or U4179 (N_4179,N_4159,N_4021);
or U4180 (N_4180,N_4082,N_4087);
xor U4181 (N_4181,N_4091,N_4002);
or U4182 (N_4182,N_4097,N_4095);
nor U4183 (N_4183,N_4141,N_4148);
or U4184 (N_4184,N_4064,N_4155);
nand U4185 (N_4185,N_4074,N_4112);
and U4186 (N_4186,N_4131,N_4124);
and U4187 (N_4187,N_4024,N_4081);
and U4188 (N_4188,N_4069,N_4060);
xnor U4189 (N_4189,N_4086,N_4042);
or U4190 (N_4190,N_4083,N_4055);
or U4191 (N_4191,N_4003,N_4110);
nor U4192 (N_4192,N_4103,N_4034);
nand U4193 (N_4193,N_4105,N_4025);
nand U4194 (N_4194,N_4036,N_4138);
nand U4195 (N_4195,N_4137,N_4147);
or U4196 (N_4196,N_4067,N_4153);
nand U4197 (N_4197,N_4098,N_4111);
nor U4198 (N_4198,N_4039,N_4115);
nor U4199 (N_4199,N_4019,N_4028);
nand U4200 (N_4200,N_4051,N_4005);
or U4201 (N_4201,N_4108,N_4109);
nand U4202 (N_4202,N_4096,N_4048);
nor U4203 (N_4203,N_4006,N_4077);
nand U4204 (N_4204,N_4128,N_4057);
or U4205 (N_4205,N_4117,N_4080);
nand U4206 (N_4206,N_4158,N_4014);
and U4207 (N_4207,N_4123,N_4132);
nand U4208 (N_4208,N_4022,N_4134);
and U4209 (N_4209,N_4100,N_4063);
or U4210 (N_4210,N_4061,N_4041);
or U4211 (N_4211,N_4130,N_4016);
nand U4212 (N_4212,N_4135,N_4118);
or U4213 (N_4213,N_4090,N_4127);
nor U4214 (N_4214,N_4094,N_4033);
or U4215 (N_4215,N_4125,N_4043);
and U4216 (N_4216,N_4149,N_4001);
or U4217 (N_4217,N_4054,N_4072);
nand U4218 (N_4218,N_4031,N_4085);
nand U4219 (N_4219,N_4029,N_4009);
nor U4220 (N_4220,N_4140,N_4062);
or U4221 (N_4221,N_4088,N_4156);
nor U4222 (N_4222,N_4152,N_4052);
nand U4223 (N_4223,N_4015,N_4075);
and U4224 (N_4224,N_4116,N_4076);
nand U4225 (N_4225,N_4107,N_4037);
nor U4226 (N_4226,N_4144,N_4145);
xnor U4227 (N_4227,N_4038,N_4084);
or U4228 (N_4228,N_4078,N_4106);
nand U4229 (N_4229,N_4133,N_4101);
or U4230 (N_4230,N_4150,N_4121);
nor U4231 (N_4231,N_4120,N_4122);
and U4232 (N_4232,N_4093,N_4047);
nor U4233 (N_4233,N_4053,N_4068);
and U4234 (N_4234,N_4010,N_4000);
xor U4235 (N_4235,N_4049,N_4065);
and U4236 (N_4236,N_4058,N_4017);
or U4237 (N_4237,N_4046,N_4032);
nor U4238 (N_4238,N_4007,N_4142);
and U4239 (N_4239,N_4089,N_4040);
or U4240 (N_4240,N_4118,N_4035);
or U4241 (N_4241,N_4097,N_4059);
nor U4242 (N_4242,N_4033,N_4106);
nor U4243 (N_4243,N_4123,N_4072);
nand U4244 (N_4244,N_4150,N_4091);
or U4245 (N_4245,N_4107,N_4067);
nand U4246 (N_4246,N_4129,N_4019);
nand U4247 (N_4247,N_4062,N_4122);
nor U4248 (N_4248,N_4110,N_4009);
and U4249 (N_4249,N_4144,N_4158);
and U4250 (N_4250,N_4146,N_4141);
and U4251 (N_4251,N_4087,N_4002);
and U4252 (N_4252,N_4038,N_4156);
and U4253 (N_4253,N_4082,N_4063);
xor U4254 (N_4254,N_4157,N_4029);
nor U4255 (N_4255,N_4042,N_4090);
nand U4256 (N_4256,N_4137,N_4032);
and U4257 (N_4257,N_4101,N_4004);
nand U4258 (N_4258,N_4093,N_4000);
or U4259 (N_4259,N_4096,N_4147);
xnor U4260 (N_4260,N_4025,N_4143);
nand U4261 (N_4261,N_4085,N_4096);
or U4262 (N_4262,N_4138,N_4064);
nor U4263 (N_4263,N_4004,N_4112);
nor U4264 (N_4264,N_4037,N_4060);
nand U4265 (N_4265,N_4151,N_4064);
or U4266 (N_4266,N_4118,N_4069);
xor U4267 (N_4267,N_4002,N_4066);
nand U4268 (N_4268,N_4110,N_4117);
nor U4269 (N_4269,N_4039,N_4092);
or U4270 (N_4270,N_4087,N_4081);
nand U4271 (N_4271,N_4002,N_4053);
and U4272 (N_4272,N_4048,N_4001);
nand U4273 (N_4273,N_4073,N_4082);
xnor U4274 (N_4274,N_4073,N_4050);
nor U4275 (N_4275,N_4154,N_4130);
xnor U4276 (N_4276,N_4130,N_4043);
nor U4277 (N_4277,N_4158,N_4115);
or U4278 (N_4278,N_4013,N_4099);
and U4279 (N_4279,N_4142,N_4061);
xnor U4280 (N_4280,N_4090,N_4064);
nand U4281 (N_4281,N_4133,N_4034);
or U4282 (N_4282,N_4111,N_4042);
nor U4283 (N_4283,N_4030,N_4036);
or U4284 (N_4284,N_4125,N_4084);
or U4285 (N_4285,N_4098,N_4044);
nor U4286 (N_4286,N_4151,N_4034);
or U4287 (N_4287,N_4011,N_4003);
nor U4288 (N_4288,N_4019,N_4009);
nor U4289 (N_4289,N_4013,N_4101);
nand U4290 (N_4290,N_4134,N_4074);
or U4291 (N_4291,N_4047,N_4101);
nand U4292 (N_4292,N_4008,N_4047);
nand U4293 (N_4293,N_4098,N_4027);
xor U4294 (N_4294,N_4070,N_4120);
or U4295 (N_4295,N_4108,N_4131);
nor U4296 (N_4296,N_4103,N_4071);
and U4297 (N_4297,N_4068,N_4007);
nand U4298 (N_4298,N_4146,N_4089);
and U4299 (N_4299,N_4093,N_4072);
nor U4300 (N_4300,N_4061,N_4158);
or U4301 (N_4301,N_4003,N_4056);
nor U4302 (N_4302,N_4090,N_4079);
nor U4303 (N_4303,N_4078,N_4136);
nor U4304 (N_4304,N_4043,N_4019);
or U4305 (N_4305,N_4065,N_4046);
nor U4306 (N_4306,N_4075,N_4116);
and U4307 (N_4307,N_4061,N_4149);
nor U4308 (N_4308,N_4134,N_4141);
nor U4309 (N_4309,N_4127,N_4158);
and U4310 (N_4310,N_4087,N_4044);
nand U4311 (N_4311,N_4137,N_4039);
nor U4312 (N_4312,N_4135,N_4124);
or U4313 (N_4313,N_4088,N_4023);
or U4314 (N_4314,N_4071,N_4116);
or U4315 (N_4315,N_4087,N_4056);
nor U4316 (N_4316,N_4116,N_4012);
nor U4317 (N_4317,N_4131,N_4078);
nor U4318 (N_4318,N_4157,N_4051);
nand U4319 (N_4319,N_4035,N_4143);
nand U4320 (N_4320,N_4243,N_4219);
nand U4321 (N_4321,N_4276,N_4301);
nor U4322 (N_4322,N_4275,N_4298);
xor U4323 (N_4323,N_4259,N_4200);
nand U4324 (N_4324,N_4263,N_4234);
nand U4325 (N_4325,N_4267,N_4260);
nand U4326 (N_4326,N_4305,N_4296);
and U4327 (N_4327,N_4268,N_4164);
or U4328 (N_4328,N_4175,N_4242);
nor U4329 (N_4329,N_4169,N_4312);
or U4330 (N_4330,N_4179,N_4274);
nor U4331 (N_4331,N_4204,N_4177);
xor U4332 (N_4332,N_4247,N_4223);
and U4333 (N_4333,N_4261,N_4187);
or U4334 (N_4334,N_4192,N_4300);
xnor U4335 (N_4335,N_4222,N_4292);
or U4336 (N_4336,N_4174,N_4172);
xor U4337 (N_4337,N_4283,N_4211);
or U4338 (N_4338,N_4304,N_4281);
nor U4339 (N_4339,N_4184,N_4168);
nor U4340 (N_4340,N_4306,N_4162);
nand U4341 (N_4341,N_4183,N_4271);
and U4342 (N_4342,N_4319,N_4289);
nor U4343 (N_4343,N_4270,N_4167);
and U4344 (N_4344,N_4178,N_4256);
and U4345 (N_4345,N_4212,N_4285);
and U4346 (N_4346,N_4303,N_4191);
and U4347 (N_4347,N_4269,N_4241);
xor U4348 (N_4348,N_4196,N_4280);
or U4349 (N_4349,N_4265,N_4288);
nor U4350 (N_4350,N_4213,N_4221);
nor U4351 (N_4351,N_4246,N_4203);
or U4352 (N_4352,N_4205,N_4199);
and U4353 (N_4353,N_4190,N_4166);
xor U4354 (N_4354,N_4311,N_4209);
nand U4355 (N_4355,N_4185,N_4316);
or U4356 (N_4356,N_4201,N_4215);
nand U4357 (N_4357,N_4307,N_4176);
nand U4358 (N_4358,N_4206,N_4231);
nand U4359 (N_4359,N_4229,N_4249);
and U4360 (N_4360,N_4197,N_4313);
and U4361 (N_4361,N_4317,N_4238);
and U4362 (N_4362,N_4297,N_4258);
nor U4363 (N_4363,N_4170,N_4291);
xnor U4364 (N_4364,N_4314,N_4240);
xor U4365 (N_4365,N_4302,N_4236);
and U4366 (N_4366,N_4198,N_4180);
xor U4367 (N_4367,N_4255,N_4315);
or U4368 (N_4368,N_4161,N_4286);
and U4369 (N_4369,N_4273,N_4310);
nand U4370 (N_4370,N_4217,N_4237);
and U4371 (N_4371,N_4186,N_4295);
or U4372 (N_4372,N_4220,N_4171);
nor U4373 (N_4373,N_4309,N_4244);
nor U4374 (N_4374,N_4232,N_4278);
nor U4375 (N_4375,N_4299,N_4235);
nor U4376 (N_4376,N_4252,N_4208);
or U4377 (N_4377,N_4245,N_4182);
nand U4378 (N_4378,N_4251,N_4202);
or U4379 (N_4379,N_4266,N_4188);
xor U4380 (N_4380,N_4207,N_4294);
xor U4381 (N_4381,N_4254,N_4165);
xor U4382 (N_4382,N_4308,N_4277);
or U4383 (N_4383,N_4214,N_4287);
nor U4384 (N_4384,N_4227,N_4318);
or U4385 (N_4385,N_4224,N_4210);
and U4386 (N_4386,N_4262,N_4173);
or U4387 (N_4387,N_4226,N_4282);
and U4388 (N_4388,N_4233,N_4218);
nand U4389 (N_4389,N_4225,N_4257);
nand U4390 (N_4390,N_4279,N_4284);
nand U4391 (N_4391,N_4264,N_4181);
nand U4392 (N_4392,N_4163,N_4293);
nand U4393 (N_4393,N_4216,N_4194);
nand U4394 (N_4394,N_4193,N_4253);
xnor U4395 (N_4395,N_4160,N_4239);
or U4396 (N_4396,N_4228,N_4250);
and U4397 (N_4397,N_4230,N_4272);
nor U4398 (N_4398,N_4189,N_4248);
and U4399 (N_4399,N_4195,N_4290);
and U4400 (N_4400,N_4204,N_4286);
nand U4401 (N_4401,N_4210,N_4209);
or U4402 (N_4402,N_4256,N_4194);
and U4403 (N_4403,N_4254,N_4265);
and U4404 (N_4404,N_4182,N_4186);
nand U4405 (N_4405,N_4197,N_4290);
or U4406 (N_4406,N_4203,N_4208);
nand U4407 (N_4407,N_4249,N_4186);
xnor U4408 (N_4408,N_4171,N_4257);
or U4409 (N_4409,N_4283,N_4202);
xnor U4410 (N_4410,N_4302,N_4168);
nand U4411 (N_4411,N_4160,N_4199);
or U4412 (N_4412,N_4242,N_4286);
nand U4413 (N_4413,N_4248,N_4309);
nand U4414 (N_4414,N_4253,N_4281);
or U4415 (N_4415,N_4286,N_4230);
nor U4416 (N_4416,N_4190,N_4310);
nand U4417 (N_4417,N_4213,N_4253);
nand U4418 (N_4418,N_4304,N_4279);
and U4419 (N_4419,N_4253,N_4264);
xnor U4420 (N_4420,N_4294,N_4181);
nand U4421 (N_4421,N_4229,N_4199);
and U4422 (N_4422,N_4269,N_4220);
or U4423 (N_4423,N_4172,N_4291);
nand U4424 (N_4424,N_4276,N_4282);
and U4425 (N_4425,N_4237,N_4266);
xnor U4426 (N_4426,N_4236,N_4256);
nor U4427 (N_4427,N_4199,N_4307);
xor U4428 (N_4428,N_4283,N_4229);
and U4429 (N_4429,N_4301,N_4212);
and U4430 (N_4430,N_4304,N_4191);
nand U4431 (N_4431,N_4277,N_4190);
or U4432 (N_4432,N_4195,N_4259);
and U4433 (N_4433,N_4304,N_4231);
or U4434 (N_4434,N_4224,N_4265);
or U4435 (N_4435,N_4299,N_4247);
nand U4436 (N_4436,N_4232,N_4163);
nor U4437 (N_4437,N_4263,N_4169);
xnor U4438 (N_4438,N_4219,N_4212);
or U4439 (N_4439,N_4182,N_4301);
or U4440 (N_4440,N_4162,N_4263);
nand U4441 (N_4441,N_4247,N_4167);
nor U4442 (N_4442,N_4231,N_4313);
and U4443 (N_4443,N_4205,N_4288);
and U4444 (N_4444,N_4319,N_4269);
and U4445 (N_4445,N_4282,N_4248);
and U4446 (N_4446,N_4223,N_4184);
nor U4447 (N_4447,N_4277,N_4257);
and U4448 (N_4448,N_4307,N_4309);
nor U4449 (N_4449,N_4170,N_4240);
and U4450 (N_4450,N_4168,N_4211);
nor U4451 (N_4451,N_4254,N_4224);
and U4452 (N_4452,N_4197,N_4201);
nand U4453 (N_4453,N_4209,N_4220);
or U4454 (N_4454,N_4263,N_4213);
or U4455 (N_4455,N_4266,N_4225);
nor U4456 (N_4456,N_4313,N_4319);
or U4457 (N_4457,N_4230,N_4191);
and U4458 (N_4458,N_4318,N_4277);
and U4459 (N_4459,N_4214,N_4296);
or U4460 (N_4460,N_4258,N_4201);
nand U4461 (N_4461,N_4233,N_4310);
nor U4462 (N_4462,N_4314,N_4223);
nor U4463 (N_4463,N_4279,N_4164);
nor U4464 (N_4464,N_4163,N_4271);
nor U4465 (N_4465,N_4178,N_4315);
and U4466 (N_4466,N_4307,N_4166);
xnor U4467 (N_4467,N_4187,N_4211);
and U4468 (N_4468,N_4171,N_4226);
nor U4469 (N_4469,N_4247,N_4259);
and U4470 (N_4470,N_4243,N_4316);
and U4471 (N_4471,N_4317,N_4253);
nor U4472 (N_4472,N_4290,N_4205);
or U4473 (N_4473,N_4228,N_4160);
nand U4474 (N_4474,N_4171,N_4242);
and U4475 (N_4475,N_4194,N_4224);
nand U4476 (N_4476,N_4179,N_4245);
or U4477 (N_4477,N_4300,N_4290);
nand U4478 (N_4478,N_4204,N_4199);
and U4479 (N_4479,N_4193,N_4291);
nor U4480 (N_4480,N_4463,N_4337);
and U4481 (N_4481,N_4341,N_4447);
nand U4482 (N_4482,N_4436,N_4429);
or U4483 (N_4483,N_4324,N_4471);
nand U4484 (N_4484,N_4423,N_4330);
nor U4485 (N_4485,N_4356,N_4446);
or U4486 (N_4486,N_4393,N_4321);
or U4487 (N_4487,N_4460,N_4415);
or U4488 (N_4488,N_4450,N_4365);
nand U4489 (N_4489,N_4430,N_4354);
xor U4490 (N_4490,N_4404,N_4370);
xnor U4491 (N_4491,N_4380,N_4373);
nor U4492 (N_4492,N_4383,N_4374);
xor U4493 (N_4493,N_4382,N_4390);
nand U4494 (N_4494,N_4407,N_4441);
or U4495 (N_4495,N_4357,N_4338);
or U4496 (N_4496,N_4339,N_4386);
nand U4497 (N_4497,N_4372,N_4425);
xnor U4498 (N_4498,N_4433,N_4442);
nor U4499 (N_4499,N_4381,N_4421);
and U4500 (N_4500,N_4392,N_4322);
nand U4501 (N_4501,N_4417,N_4352);
nand U4502 (N_4502,N_4469,N_4431);
or U4503 (N_4503,N_4459,N_4451);
nand U4504 (N_4504,N_4410,N_4377);
and U4505 (N_4505,N_4409,N_4414);
nand U4506 (N_4506,N_4405,N_4473);
nand U4507 (N_4507,N_4364,N_4408);
xnor U4508 (N_4508,N_4478,N_4331);
nand U4509 (N_4509,N_4388,N_4355);
or U4510 (N_4510,N_4419,N_4472);
nand U4511 (N_4511,N_4434,N_4479);
nand U4512 (N_4512,N_4359,N_4468);
and U4513 (N_4513,N_4385,N_4406);
nand U4514 (N_4514,N_4361,N_4444);
or U4515 (N_4515,N_4437,N_4348);
nand U4516 (N_4516,N_4328,N_4477);
or U4517 (N_4517,N_4369,N_4435);
or U4518 (N_4518,N_4350,N_4332);
nor U4519 (N_4519,N_4367,N_4461);
or U4520 (N_4520,N_4395,N_4474);
nor U4521 (N_4521,N_4453,N_4411);
or U4522 (N_4522,N_4362,N_4418);
nand U4523 (N_4523,N_4422,N_4402);
nor U4524 (N_4524,N_4391,N_4449);
nand U4525 (N_4525,N_4432,N_4335);
and U4526 (N_4526,N_4346,N_4379);
nand U4527 (N_4527,N_4376,N_4448);
xnor U4528 (N_4528,N_4467,N_4326);
or U4529 (N_4529,N_4428,N_4366);
nor U4530 (N_4530,N_4476,N_4347);
nor U4531 (N_4531,N_4384,N_4371);
or U4532 (N_4532,N_4445,N_4466);
nor U4533 (N_4533,N_4345,N_4363);
or U4534 (N_4534,N_4440,N_4455);
nor U4535 (N_4535,N_4426,N_4424);
nand U4536 (N_4536,N_4439,N_4378);
xnor U4537 (N_4537,N_4389,N_4368);
and U4538 (N_4538,N_4464,N_4358);
nor U4539 (N_4539,N_4333,N_4413);
xor U4540 (N_4540,N_4454,N_4353);
nand U4541 (N_4541,N_4438,N_4399);
or U4542 (N_4542,N_4344,N_4400);
nor U4543 (N_4543,N_4457,N_4325);
and U4544 (N_4544,N_4443,N_4416);
nor U4545 (N_4545,N_4401,N_4397);
or U4546 (N_4546,N_4470,N_4320);
nor U4547 (N_4547,N_4349,N_4387);
nor U4548 (N_4548,N_4458,N_4343);
nor U4549 (N_4549,N_4456,N_4427);
and U4550 (N_4550,N_4475,N_4360);
xnor U4551 (N_4551,N_4323,N_4465);
xor U4552 (N_4552,N_4420,N_4327);
nor U4553 (N_4553,N_4403,N_4351);
or U4554 (N_4554,N_4342,N_4336);
and U4555 (N_4555,N_4375,N_4394);
or U4556 (N_4556,N_4396,N_4340);
nand U4557 (N_4557,N_4334,N_4412);
and U4558 (N_4558,N_4329,N_4462);
xor U4559 (N_4559,N_4398,N_4452);
nor U4560 (N_4560,N_4337,N_4347);
or U4561 (N_4561,N_4342,N_4437);
xor U4562 (N_4562,N_4324,N_4332);
or U4563 (N_4563,N_4355,N_4394);
or U4564 (N_4564,N_4462,N_4454);
and U4565 (N_4565,N_4401,N_4406);
and U4566 (N_4566,N_4393,N_4461);
nand U4567 (N_4567,N_4338,N_4411);
nand U4568 (N_4568,N_4451,N_4430);
or U4569 (N_4569,N_4421,N_4429);
nand U4570 (N_4570,N_4439,N_4339);
nand U4571 (N_4571,N_4323,N_4357);
nand U4572 (N_4572,N_4433,N_4363);
or U4573 (N_4573,N_4470,N_4450);
nand U4574 (N_4574,N_4425,N_4335);
nor U4575 (N_4575,N_4360,N_4474);
or U4576 (N_4576,N_4463,N_4454);
or U4577 (N_4577,N_4459,N_4452);
nor U4578 (N_4578,N_4378,N_4406);
or U4579 (N_4579,N_4358,N_4351);
nor U4580 (N_4580,N_4415,N_4357);
and U4581 (N_4581,N_4475,N_4453);
nor U4582 (N_4582,N_4434,N_4422);
xnor U4583 (N_4583,N_4425,N_4348);
nand U4584 (N_4584,N_4426,N_4457);
nand U4585 (N_4585,N_4420,N_4469);
and U4586 (N_4586,N_4456,N_4352);
nand U4587 (N_4587,N_4415,N_4356);
nor U4588 (N_4588,N_4380,N_4401);
nand U4589 (N_4589,N_4328,N_4408);
nor U4590 (N_4590,N_4398,N_4361);
and U4591 (N_4591,N_4447,N_4335);
nor U4592 (N_4592,N_4386,N_4358);
and U4593 (N_4593,N_4420,N_4332);
nor U4594 (N_4594,N_4332,N_4421);
nand U4595 (N_4595,N_4399,N_4411);
or U4596 (N_4596,N_4368,N_4450);
or U4597 (N_4597,N_4393,N_4340);
and U4598 (N_4598,N_4343,N_4436);
and U4599 (N_4599,N_4436,N_4452);
nor U4600 (N_4600,N_4376,N_4437);
nor U4601 (N_4601,N_4363,N_4407);
nor U4602 (N_4602,N_4445,N_4405);
and U4603 (N_4603,N_4409,N_4381);
nor U4604 (N_4604,N_4437,N_4412);
nand U4605 (N_4605,N_4326,N_4347);
nand U4606 (N_4606,N_4374,N_4414);
nand U4607 (N_4607,N_4325,N_4344);
nand U4608 (N_4608,N_4358,N_4470);
nor U4609 (N_4609,N_4464,N_4328);
nor U4610 (N_4610,N_4470,N_4428);
nor U4611 (N_4611,N_4413,N_4390);
xor U4612 (N_4612,N_4458,N_4372);
or U4613 (N_4613,N_4350,N_4473);
nor U4614 (N_4614,N_4371,N_4468);
or U4615 (N_4615,N_4473,N_4425);
nor U4616 (N_4616,N_4337,N_4421);
nand U4617 (N_4617,N_4407,N_4409);
and U4618 (N_4618,N_4393,N_4450);
nand U4619 (N_4619,N_4422,N_4438);
and U4620 (N_4620,N_4393,N_4438);
and U4621 (N_4621,N_4375,N_4417);
nor U4622 (N_4622,N_4400,N_4325);
and U4623 (N_4623,N_4337,N_4330);
nor U4624 (N_4624,N_4351,N_4407);
nor U4625 (N_4625,N_4356,N_4385);
nand U4626 (N_4626,N_4479,N_4369);
and U4627 (N_4627,N_4390,N_4416);
or U4628 (N_4628,N_4398,N_4436);
xnor U4629 (N_4629,N_4330,N_4335);
nor U4630 (N_4630,N_4435,N_4341);
nor U4631 (N_4631,N_4436,N_4341);
and U4632 (N_4632,N_4367,N_4327);
or U4633 (N_4633,N_4370,N_4367);
or U4634 (N_4634,N_4393,N_4408);
nor U4635 (N_4635,N_4397,N_4328);
xnor U4636 (N_4636,N_4333,N_4428);
and U4637 (N_4637,N_4337,N_4344);
nor U4638 (N_4638,N_4353,N_4322);
or U4639 (N_4639,N_4465,N_4419);
and U4640 (N_4640,N_4518,N_4612);
xnor U4641 (N_4641,N_4506,N_4514);
or U4642 (N_4642,N_4583,N_4554);
or U4643 (N_4643,N_4580,N_4526);
nor U4644 (N_4644,N_4592,N_4613);
nand U4645 (N_4645,N_4572,N_4523);
nand U4646 (N_4646,N_4582,N_4605);
and U4647 (N_4647,N_4544,N_4566);
and U4648 (N_4648,N_4513,N_4493);
nand U4649 (N_4649,N_4581,N_4524);
or U4650 (N_4650,N_4488,N_4538);
or U4651 (N_4651,N_4496,N_4574);
nand U4652 (N_4652,N_4608,N_4631);
nor U4653 (N_4653,N_4596,N_4499);
nor U4654 (N_4654,N_4490,N_4510);
nor U4655 (N_4655,N_4485,N_4559);
nand U4656 (N_4656,N_4521,N_4576);
or U4657 (N_4657,N_4560,N_4528);
nor U4658 (N_4658,N_4500,N_4532);
or U4659 (N_4659,N_4603,N_4512);
nor U4660 (N_4660,N_4568,N_4563);
nor U4661 (N_4661,N_4517,N_4616);
and U4662 (N_4662,N_4624,N_4534);
or U4663 (N_4663,N_4639,N_4602);
nand U4664 (N_4664,N_4531,N_4626);
nor U4665 (N_4665,N_4491,N_4611);
and U4666 (N_4666,N_4633,N_4509);
and U4667 (N_4667,N_4617,N_4503);
nor U4668 (N_4668,N_4615,N_4607);
nand U4669 (N_4669,N_4587,N_4542);
and U4670 (N_4670,N_4498,N_4609);
nor U4671 (N_4671,N_4635,N_4597);
nor U4672 (N_4672,N_4627,N_4530);
and U4673 (N_4673,N_4557,N_4620);
nand U4674 (N_4674,N_4584,N_4543);
xnor U4675 (N_4675,N_4614,N_4629);
or U4676 (N_4676,N_4480,N_4546);
nor U4677 (N_4677,N_4618,N_4623);
nand U4678 (N_4678,N_4548,N_4489);
or U4679 (N_4679,N_4486,N_4484);
nor U4680 (N_4680,N_4637,N_4621);
nor U4681 (N_4681,N_4634,N_4598);
or U4682 (N_4682,N_4527,N_4520);
or U4683 (N_4683,N_4501,N_4628);
or U4684 (N_4684,N_4558,N_4553);
nand U4685 (N_4685,N_4505,N_4551);
and U4686 (N_4686,N_4535,N_4638);
nor U4687 (N_4687,N_4562,N_4565);
nor U4688 (N_4688,N_4539,N_4636);
nand U4689 (N_4689,N_4625,N_4508);
nor U4690 (N_4690,N_4511,N_4570);
xnor U4691 (N_4691,N_4540,N_4529);
xor U4692 (N_4692,N_4552,N_4507);
xor U4693 (N_4693,N_4589,N_4561);
nor U4694 (N_4694,N_4545,N_4519);
xnor U4695 (N_4695,N_4632,N_4588);
and U4696 (N_4696,N_4537,N_4577);
or U4697 (N_4697,N_4600,N_4578);
and U4698 (N_4698,N_4515,N_4619);
or U4699 (N_4699,N_4482,N_4533);
nand U4700 (N_4700,N_4630,N_4575);
and U4701 (N_4701,N_4504,N_4601);
nor U4702 (N_4702,N_4492,N_4586);
nor U4703 (N_4703,N_4494,N_4604);
nor U4704 (N_4704,N_4573,N_4595);
nor U4705 (N_4705,N_4622,N_4550);
or U4706 (N_4706,N_4516,N_4495);
or U4707 (N_4707,N_4502,N_4497);
nor U4708 (N_4708,N_4594,N_4590);
and U4709 (N_4709,N_4536,N_4569);
and U4710 (N_4710,N_4481,N_4567);
nor U4711 (N_4711,N_4556,N_4522);
nor U4712 (N_4712,N_4599,N_4483);
or U4713 (N_4713,N_4525,N_4541);
nand U4714 (N_4714,N_4585,N_4610);
nor U4715 (N_4715,N_4593,N_4487);
and U4716 (N_4716,N_4579,N_4564);
nand U4717 (N_4717,N_4549,N_4555);
or U4718 (N_4718,N_4571,N_4547);
or U4719 (N_4719,N_4606,N_4591);
nand U4720 (N_4720,N_4568,N_4522);
or U4721 (N_4721,N_4567,N_4608);
or U4722 (N_4722,N_4481,N_4516);
nor U4723 (N_4723,N_4631,N_4522);
or U4724 (N_4724,N_4481,N_4488);
nor U4725 (N_4725,N_4560,N_4563);
nand U4726 (N_4726,N_4633,N_4535);
or U4727 (N_4727,N_4535,N_4604);
nand U4728 (N_4728,N_4615,N_4507);
nor U4729 (N_4729,N_4485,N_4598);
nor U4730 (N_4730,N_4569,N_4614);
and U4731 (N_4731,N_4505,N_4565);
nor U4732 (N_4732,N_4610,N_4538);
nand U4733 (N_4733,N_4525,N_4635);
and U4734 (N_4734,N_4624,N_4530);
or U4735 (N_4735,N_4607,N_4517);
and U4736 (N_4736,N_4600,N_4485);
or U4737 (N_4737,N_4523,N_4518);
nand U4738 (N_4738,N_4536,N_4518);
and U4739 (N_4739,N_4486,N_4587);
or U4740 (N_4740,N_4569,N_4524);
and U4741 (N_4741,N_4497,N_4610);
xor U4742 (N_4742,N_4599,N_4481);
xor U4743 (N_4743,N_4558,N_4594);
or U4744 (N_4744,N_4587,N_4556);
nor U4745 (N_4745,N_4600,N_4575);
and U4746 (N_4746,N_4492,N_4615);
or U4747 (N_4747,N_4579,N_4606);
nor U4748 (N_4748,N_4535,N_4625);
and U4749 (N_4749,N_4557,N_4536);
or U4750 (N_4750,N_4494,N_4506);
or U4751 (N_4751,N_4539,N_4559);
or U4752 (N_4752,N_4591,N_4546);
and U4753 (N_4753,N_4554,N_4490);
nand U4754 (N_4754,N_4556,N_4503);
or U4755 (N_4755,N_4535,N_4599);
xor U4756 (N_4756,N_4542,N_4510);
nor U4757 (N_4757,N_4548,N_4628);
and U4758 (N_4758,N_4509,N_4620);
nor U4759 (N_4759,N_4538,N_4534);
nor U4760 (N_4760,N_4516,N_4639);
and U4761 (N_4761,N_4564,N_4592);
nand U4762 (N_4762,N_4599,N_4532);
nor U4763 (N_4763,N_4492,N_4587);
nor U4764 (N_4764,N_4575,N_4554);
nor U4765 (N_4765,N_4523,N_4522);
or U4766 (N_4766,N_4562,N_4540);
or U4767 (N_4767,N_4492,N_4522);
nor U4768 (N_4768,N_4560,N_4565);
nand U4769 (N_4769,N_4501,N_4623);
nor U4770 (N_4770,N_4635,N_4557);
and U4771 (N_4771,N_4600,N_4549);
nor U4772 (N_4772,N_4633,N_4605);
and U4773 (N_4773,N_4523,N_4589);
or U4774 (N_4774,N_4537,N_4495);
and U4775 (N_4775,N_4631,N_4564);
nand U4776 (N_4776,N_4587,N_4534);
nor U4777 (N_4777,N_4622,N_4590);
or U4778 (N_4778,N_4546,N_4622);
nor U4779 (N_4779,N_4611,N_4637);
xnor U4780 (N_4780,N_4500,N_4579);
or U4781 (N_4781,N_4503,N_4518);
nor U4782 (N_4782,N_4618,N_4593);
or U4783 (N_4783,N_4547,N_4585);
nor U4784 (N_4784,N_4510,N_4588);
and U4785 (N_4785,N_4531,N_4577);
nor U4786 (N_4786,N_4519,N_4596);
nor U4787 (N_4787,N_4496,N_4591);
nand U4788 (N_4788,N_4505,N_4601);
or U4789 (N_4789,N_4616,N_4503);
and U4790 (N_4790,N_4570,N_4557);
nand U4791 (N_4791,N_4529,N_4610);
nor U4792 (N_4792,N_4492,N_4514);
nand U4793 (N_4793,N_4510,N_4552);
and U4794 (N_4794,N_4489,N_4561);
xor U4795 (N_4795,N_4540,N_4586);
or U4796 (N_4796,N_4582,N_4524);
nor U4797 (N_4797,N_4610,N_4555);
nor U4798 (N_4798,N_4621,N_4511);
nor U4799 (N_4799,N_4509,N_4630);
and U4800 (N_4800,N_4781,N_4708);
xor U4801 (N_4801,N_4778,N_4660);
and U4802 (N_4802,N_4678,N_4726);
and U4803 (N_4803,N_4729,N_4718);
and U4804 (N_4804,N_4711,N_4709);
xor U4805 (N_4805,N_4776,N_4694);
xor U4806 (N_4806,N_4769,N_4677);
or U4807 (N_4807,N_4683,N_4754);
or U4808 (N_4808,N_4742,N_4735);
or U4809 (N_4809,N_4731,N_4704);
xor U4810 (N_4810,N_4698,N_4675);
and U4811 (N_4811,N_4744,N_4792);
or U4812 (N_4812,N_4788,N_4775);
and U4813 (N_4813,N_4697,N_4671);
and U4814 (N_4814,N_4746,N_4649);
nor U4815 (N_4815,N_4772,N_4702);
and U4816 (N_4816,N_4695,N_4662);
and U4817 (N_4817,N_4720,N_4663);
nand U4818 (N_4818,N_4689,N_4655);
or U4819 (N_4819,N_4646,N_4787);
xor U4820 (N_4820,N_4757,N_4784);
or U4821 (N_4821,N_4676,N_4668);
or U4822 (N_4822,N_4667,N_4719);
nor U4823 (N_4823,N_4712,N_4796);
and U4824 (N_4824,N_4687,N_4783);
nor U4825 (N_4825,N_4750,N_4798);
nor U4826 (N_4826,N_4713,N_4692);
or U4827 (N_4827,N_4733,N_4717);
or U4828 (N_4828,N_4652,N_4779);
xnor U4829 (N_4829,N_4696,N_4759);
and U4830 (N_4830,N_4764,N_4734);
nand U4831 (N_4831,N_4672,N_4785);
nor U4832 (N_4832,N_4768,N_4640);
or U4833 (N_4833,N_4690,N_4664);
and U4834 (N_4834,N_4722,N_4766);
or U4835 (N_4835,N_4741,N_4705);
nor U4836 (N_4836,N_4786,N_4728);
and U4837 (N_4837,N_4716,N_4730);
or U4838 (N_4838,N_4765,N_4752);
or U4839 (N_4839,N_4763,N_4758);
and U4840 (N_4840,N_4790,N_4762);
xnor U4841 (N_4841,N_4760,N_4701);
nor U4842 (N_4842,N_4721,N_4727);
xnor U4843 (N_4843,N_4691,N_4791);
nor U4844 (N_4844,N_4693,N_4686);
nor U4845 (N_4845,N_4761,N_4795);
and U4846 (N_4846,N_4688,N_4794);
nor U4847 (N_4847,N_4661,N_4771);
nand U4848 (N_4848,N_4782,N_4682);
nor U4849 (N_4849,N_4669,N_4654);
or U4850 (N_4850,N_4651,N_4703);
nor U4851 (N_4851,N_4659,N_4647);
and U4852 (N_4852,N_4753,N_4642);
nand U4853 (N_4853,N_4748,N_4680);
xor U4854 (N_4854,N_4674,N_4645);
nor U4855 (N_4855,N_4685,N_4740);
xor U4856 (N_4856,N_4749,N_4774);
nor U4857 (N_4857,N_4706,N_4745);
nor U4858 (N_4858,N_4797,N_4665);
nor U4859 (N_4859,N_4777,N_4756);
nor U4860 (N_4860,N_4738,N_4684);
or U4861 (N_4861,N_4643,N_4725);
and U4862 (N_4862,N_4773,N_4641);
nand U4863 (N_4863,N_4714,N_4737);
and U4864 (N_4864,N_4780,N_4699);
nor U4865 (N_4865,N_4755,N_4799);
and U4866 (N_4866,N_4681,N_4700);
nand U4867 (N_4867,N_4679,N_4736);
nor U4868 (N_4868,N_4747,N_4707);
xnor U4869 (N_4869,N_4767,N_4644);
or U4870 (N_4870,N_4648,N_4666);
or U4871 (N_4871,N_4724,N_4751);
nor U4872 (N_4872,N_4793,N_4653);
nand U4873 (N_4873,N_4789,N_4650);
nor U4874 (N_4874,N_4723,N_4739);
nand U4875 (N_4875,N_4710,N_4743);
and U4876 (N_4876,N_4770,N_4670);
nor U4877 (N_4877,N_4658,N_4673);
and U4878 (N_4878,N_4732,N_4657);
xor U4879 (N_4879,N_4715,N_4656);
or U4880 (N_4880,N_4648,N_4655);
nand U4881 (N_4881,N_4783,N_4759);
and U4882 (N_4882,N_4779,N_4642);
xor U4883 (N_4883,N_4698,N_4762);
or U4884 (N_4884,N_4665,N_4649);
or U4885 (N_4885,N_4651,N_4694);
nand U4886 (N_4886,N_4796,N_4689);
xor U4887 (N_4887,N_4781,N_4782);
and U4888 (N_4888,N_4649,N_4740);
or U4889 (N_4889,N_4708,N_4744);
nor U4890 (N_4890,N_4780,N_4665);
or U4891 (N_4891,N_4663,N_4647);
nor U4892 (N_4892,N_4646,N_4665);
or U4893 (N_4893,N_4752,N_4709);
nor U4894 (N_4894,N_4698,N_4687);
or U4895 (N_4895,N_4693,N_4758);
xnor U4896 (N_4896,N_4675,N_4770);
nor U4897 (N_4897,N_4670,N_4643);
nor U4898 (N_4898,N_4646,N_4796);
nor U4899 (N_4899,N_4798,N_4657);
nor U4900 (N_4900,N_4764,N_4726);
or U4901 (N_4901,N_4726,N_4729);
nand U4902 (N_4902,N_4662,N_4777);
nor U4903 (N_4903,N_4738,N_4721);
and U4904 (N_4904,N_4691,N_4688);
nor U4905 (N_4905,N_4676,N_4649);
nor U4906 (N_4906,N_4729,N_4736);
nand U4907 (N_4907,N_4687,N_4720);
and U4908 (N_4908,N_4670,N_4701);
nand U4909 (N_4909,N_4733,N_4687);
xnor U4910 (N_4910,N_4695,N_4711);
xnor U4911 (N_4911,N_4670,N_4655);
nand U4912 (N_4912,N_4754,N_4665);
nor U4913 (N_4913,N_4653,N_4770);
nand U4914 (N_4914,N_4663,N_4662);
and U4915 (N_4915,N_4688,N_4713);
and U4916 (N_4916,N_4771,N_4703);
or U4917 (N_4917,N_4797,N_4749);
and U4918 (N_4918,N_4764,N_4674);
nor U4919 (N_4919,N_4735,N_4767);
nor U4920 (N_4920,N_4699,N_4792);
nor U4921 (N_4921,N_4689,N_4790);
or U4922 (N_4922,N_4688,N_4697);
and U4923 (N_4923,N_4641,N_4653);
or U4924 (N_4924,N_4778,N_4775);
or U4925 (N_4925,N_4707,N_4684);
nor U4926 (N_4926,N_4733,N_4707);
or U4927 (N_4927,N_4787,N_4656);
nand U4928 (N_4928,N_4680,N_4683);
or U4929 (N_4929,N_4708,N_4779);
nor U4930 (N_4930,N_4765,N_4663);
xor U4931 (N_4931,N_4691,N_4751);
nand U4932 (N_4932,N_4737,N_4763);
or U4933 (N_4933,N_4686,N_4670);
nor U4934 (N_4934,N_4680,N_4736);
or U4935 (N_4935,N_4705,N_4797);
or U4936 (N_4936,N_4649,N_4685);
and U4937 (N_4937,N_4793,N_4657);
or U4938 (N_4938,N_4724,N_4746);
nand U4939 (N_4939,N_4789,N_4670);
and U4940 (N_4940,N_4785,N_4642);
nor U4941 (N_4941,N_4690,N_4765);
or U4942 (N_4942,N_4762,N_4727);
nor U4943 (N_4943,N_4728,N_4753);
or U4944 (N_4944,N_4749,N_4675);
or U4945 (N_4945,N_4788,N_4785);
and U4946 (N_4946,N_4702,N_4674);
and U4947 (N_4947,N_4707,N_4700);
nor U4948 (N_4948,N_4702,N_4790);
xnor U4949 (N_4949,N_4764,N_4656);
nand U4950 (N_4950,N_4757,N_4722);
nand U4951 (N_4951,N_4702,N_4693);
and U4952 (N_4952,N_4655,N_4694);
xor U4953 (N_4953,N_4658,N_4763);
nand U4954 (N_4954,N_4777,N_4762);
or U4955 (N_4955,N_4685,N_4727);
nand U4956 (N_4956,N_4665,N_4763);
or U4957 (N_4957,N_4784,N_4755);
or U4958 (N_4958,N_4655,N_4697);
nand U4959 (N_4959,N_4765,N_4743);
nand U4960 (N_4960,N_4881,N_4800);
or U4961 (N_4961,N_4857,N_4808);
or U4962 (N_4962,N_4945,N_4935);
xor U4963 (N_4963,N_4913,N_4831);
nor U4964 (N_4964,N_4835,N_4903);
nand U4965 (N_4965,N_4883,N_4830);
nand U4966 (N_4966,N_4871,N_4851);
nand U4967 (N_4967,N_4899,N_4867);
and U4968 (N_4968,N_4863,N_4894);
nor U4969 (N_4969,N_4880,N_4809);
xor U4970 (N_4970,N_4939,N_4820);
or U4971 (N_4971,N_4912,N_4884);
or U4972 (N_4972,N_4914,N_4839);
nor U4973 (N_4973,N_4848,N_4811);
nand U4974 (N_4974,N_4826,N_4910);
and U4975 (N_4975,N_4953,N_4817);
and U4976 (N_4976,N_4898,N_4864);
and U4977 (N_4977,N_4916,N_4933);
and U4978 (N_4978,N_4957,N_4821);
and U4979 (N_4979,N_4918,N_4896);
xor U4980 (N_4980,N_4838,N_4926);
and U4981 (N_4981,N_4888,N_4949);
or U4982 (N_4982,N_4929,N_4909);
xnor U4983 (N_4983,N_4814,N_4802);
and U4984 (N_4984,N_4812,N_4822);
nor U4985 (N_4985,N_4872,N_4927);
nor U4986 (N_4986,N_4829,N_4917);
or U4987 (N_4987,N_4921,N_4944);
nor U4988 (N_4988,N_4869,N_4803);
nor U4989 (N_4989,N_4825,N_4810);
xnor U4990 (N_4990,N_4832,N_4891);
and U4991 (N_4991,N_4805,N_4931);
nand U4992 (N_4992,N_4827,N_4882);
nand U4993 (N_4993,N_4951,N_4950);
and U4994 (N_4994,N_4942,N_4861);
or U4995 (N_4995,N_4816,N_4856);
nor U4996 (N_4996,N_4886,N_4824);
or U4997 (N_4997,N_4895,N_4870);
nor U4998 (N_4998,N_4941,N_4892);
nand U4999 (N_4999,N_4842,N_4905);
or U5000 (N_5000,N_4932,N_4866);
nor U5001 (N_5001,N_4833,N_4801);
or U5002 (N_5002,N_4853,N_4938);
nand U5003 (N_5003,N_4841,N_4876);
nand U5004 (N_5004,N_4890,N_4925);
nand U5005 (N_5005,N_4859,N_4924);
or U5006 (N_5006,N_4947,N_4858);
or U5007 (N_5007,N_4902,N_4855);
and U5008 (N_5008,N_4823,N_4843);
or U5009 (N_5009,N_4923,N_4804);
nand U5010 (N_5010,N_4845,N_4874);
and U5011 (N_5011,N_4958,N_4834);
or U5012 (N_5012,N_4877,N_4850);
or U5013 (N_5013,N_4911,N_4948);
nor U5014 (N_5014,N_4875,N_4908);
and U5015 (N_5015,N_4956,N_4959);
xnor U5016 (N_5016,N_4930,N_4865);
and U5017 (N_5017,N_4828,N_4852);
nor U5018 (N_5018,N_4844,N_4837);
and U5019 (N_5019,N_4954,N_4847);
nand U5020 (N_5020,N_4904,N_4901);
nor U5021 (N_5021,N_4862,N_4849);
nor U5022 (N_5022,N_4920,N_4952);
nand U5023 (N_5023,N_4943,N_4946);
and U5024 (N_5024,N_4806,N_4878);
xnor U5025 (N_5025,N_4889,N_4887);
and U5026 (N_5026,N_4860,N_4815);
nand U5027 (N_5027,N_4936,N_4854);
and U5028 (N_5028,N_4955,N_4840);
or U5029 (N_5029,N_4940,N_4846);
and U5030 (N_5030,N_4897,N_4937);
and U5031 (N_5031,N_4819,N_4818);
nand U5032 (N_5032,N_4934,N_4922);
nor U5033 (N_5033,N_4885,N_4868);
or U5034 (N_5034,N_4907,N_4900);
or U5035 (N_5035,N_4873,N_4807);
and U5036 (N_5036,N_4879,N_4813);
or U5037 (N_5037,N_4928,N_4906);
nor U5038 (N_5038,N_4836,N_4919);
nor U5039 (N_5039,N_4893,N_4915);
nor U5040 (N_5040,N_4861,N_4932);
nand U5041 (N_5041,N_4908,N_4862);
or U5042 (N_5042,N_4942,N_4903);
nor U5043 (N_5043,N_4884,N_4916);
nor U5044 (N_5044,N_4951,N_4956);
nand U5045 (N_5045,N_4838,N_4941);
and U5046 (N_5046,N_4886,N_4850);
nand U5047 (N_5047,N_4906,N_4839);
nor U5048 (N_5048,N_4860,N_4811);
and U5049 (N_5049,N_4823,N_4884);
or U5050 (N_5050,N_4850,N_4864);
and U5051 (N_5051,N_4882,N_4887);
and U5052 (N_5052,N_4942,N_4851);
or U5053 (N_5053,N_4937,N_4948);
or U5054 (N_5054,N_4871,N_4800);
and U5055 (N_5055,N_4829,N_4943);
nand U5056 (N_5056,N_4842,N_4950);
xnor U5057 (N_5057,N_4855,N_4854);
nand U5058 (N_5058,N_4876,N_4827);
or U5059 (N_5059,N_4890,N_4845);
nand U5060 (N_5060,N_4949,N_4870);
and U5061 (N_5061,N_4919,N_4925);
nand U5062 (N_5062,N_4857,N_4950);
nand U5063 (N_5063,N_4904,N_4882);
and U5064 (N_5064,N_4847,N_4849);
or U5065 (N_5065,N_4801,N_4821);
xor U5066 (N_5066,N_4800,N_4950);
nor U5067 (N_5067,N_4894,N_4881);
and U5068 (N_5068,N_4918,N_4923);
or U5069 (N_5069,N_4945,N_4944);
or U5070 (N_5070,N_4924,N_4818);
xnor U5071 (N_5071,N_4841,N_4930);
or U5072 (N_5072,N_4941,N_4844);
nor U5073 (N_5073,N_4944,N_4825);
nand U5074 (N_5074,N_4940,N_4892);
or U5075 (N_5075,N_4832,N_4834);
or U5076 (N_5076,N_4878,N_4884);
or U5077 (N_5077,N_4898,N_4931);
and U5078 (N_5078,N_4930,N_4887);
nand U5079 (N_5079,N_4833,N_4946);
or U5080 (N_5080,N_4833,N_4908);
nand U5081 (N_5081,N_4890,N_4800);
or U5082 (N_5082,N_4903,N_4811);
and U5083 (N_5083,N_4897,N_4805);
nand U5084 (N_5084,N_4877,N_4806);
nand U5085 (N_5085,N_4834,N_4815);
or U5086 (N_5086,N_4929,N_4802);
xor U5087 (N_5087,N_4926,N_4837);
nor U5088 (N_5088,N_4852,N_4945);
or U5089 (N_5089,N_4907,N_4824);
or U5090 (N_5090,N_4903,N_4945);
nand U5091 (N_5091,N_4933,N_4895);
or U5092 (N_5092,N_4889,N_4870);
and U5093 (N_5093,N_4848,N_4825);
and U5094 (N_5094,N_4804,N_4848);
or U5095 (N_5095,N_4898,N_4863);
and U5096 (N_5096,N_4898,N_4836);
or U5097 (N_5097,N_4927,N_4816);
nand U5098 (N_5098,N_4838,N_4861);
or U5099 (N_5099,N_4914,N_4855);
or U5100 (N_5100,N_4870,N_4810);
nor U5101 (N_5101,N_4812,N_4901);
or U5102 (N_5102,N_4859,N_4912);
or U5103 (N_5103,N_4868,N_4930);
xor U5104 (N_5104,N_4889,N_4877);
and U5105 (N_5105,N_4947,N_4834);
or U5106 (N_5106,N_4803,N_4924);
and U5107 (N_5107,N_4917,N_4948);
and U5108 (N_5108,N_4914,N_4952);
and U5109 (N_5109,N_4823,N_4848);
nor U5110 (N_5110,N_4800,N_4912);
xnor U5111 (N_5111,N_4934,N_4818);
xnor U5112 (N_5112,N_4885,N_4938);
or U5113 (N_5113,N_4849,N_4863);
and U5114 (N_5114,N_4864,N_4849);
nor U5115 (N_5115,N_4943,N_4942);
nand U5116 (N_5116,N_4902,N_4845);
nand U5117 (N_5117,N_4904,N_4958);
nor U5118 (N_5118,N_4861,N_4871);
or U5119 (N_5119,N_4829,N_4878);
and U5120 (N_5120,N_5053,N_5056);
and U5121 (N_5121,N_5118,N_5090);
or U5122 (N_5122,N_5041,N_5048);
and U5123 (N_5123,N_5035,N_5094);
nor U5124 (N_5124,N_5075,N_5034);
xnor U5125 (N_5125,N_4995,N_5049);
nand U5126 (N_5126,N_5046,N_4961);
or U5127 (N_5127,N_5055,N_5114);
xnor U5128 (N_5128,N_5087,N_5023);
or U5129 (N_5129,N_5089,N_5047);
nor U5130 (N_5130,N_5044,N_4969);
or U5131 (N_5131,N_4992,N_5017);
and U5132 (N_5132,N_5115,N_5031);
nand U5133 (N_5133,N_5098,N_5107);
nand U5134 (N_5134,N_5038,N_5100);
nand U5135 (N_5135,N_4966,N_5084);
nand U5136 (N_5136,N_5062,N_4982);
or U5137 (N_5137,N_5085,N_5065);
and U5138 (N_5138,N_5099,N_5051);
xor U5139 (N_5139,N_5081,N_4972);
nand U5140 (N_5140,N_5004,N_4985);
and U5141 (N_5141,N_5074,N_5101);
and U5142 (N_5142,N_5095,N_5116);
nor U5143 (N_5143,N_4964,N_5008);
and U5144 (N_5144,N_5014,N_5036);
and U5145 (N_5145,N_5058,N_5016);
nand U5146 (N_5146,N_5104,N_5045);
nor U5147 (N_5147,N_5060,N_4980);
xnor U5148 (N_5148,N_5119,N_5069);
nor U5149 (N_5149,N_5027,N_5002);
nor U5150 (N_5150,N_5079,N_4990);
and U5151 (N_5151,N_5112,N_5109);
nor U5152 (N_5152,N_5037,N_5078);
nand U5153 (N_5153,N_5086,N_5000);
nand U5154 (N_5154,N_4991,N_5040);
nor U5155 (N_5155,N_5082,N_5077);
or U5156 (N_5156,N_4994,N_4963);
xor U5157 (N_5157,N_5018,N_5028);
nand U5158 (N_5158,N_4998,N_5110);
nand U5159 (N_5159,N_4983,N_4988);
and U5160 (N_5160,N_5032,N_5091);
and U5161 (N_5161,N_4977,N_5010);
or U5162 (N_5162,N_5026,N_5024);
or U5163 (N_5163,N_5052,N_5108);
and U5164 (N_5164,N_5092,N_5093);
xor U5165 (N_5165,N_5061,N_4986);
and U5166 (N_5166,N_5012,N_5022);
nand U5167 (N_5167,N_4996,N_5105);
and U5168 (N_5168,N_4989,N_5059);
nand U5169 (N_5169,N_5071,N_5073);
nor U5170 (N_5170,N_5050,N_5011);
nand U5171 (N_5171,N_5043,N_4993);
or U5172 (N_5172,N_5113,N_4975);
or U5173 (N_5173,N_5117,N_5097);
nand U5174 (N_5174,N_5033,N_5080);
and U5175 (N_5175,N_5106,N_4987);
xor U5176 (N_5176,N_4965,N_4967);
or U5177 (N_5177,N_4973,N_5096);
nand U5178 (N_5178,N_5020,N_5013);
and U5179 (N_5179,N_4978,N_5111);
nand U5180 (N_5180,N_5063,N_4971);
nand U5181 (N_5181,N_4976,N_5003);
or U5182 (N_5182,N_4999,N_5076);
xnor U5183 (N_5183,N_4962,N_5070);
nand U5184 (N_5184,N_5042,N_5005);
and U5185 (N_5185,N_5102,N_5009);
nand U5186 (N_5186,N_5068,N_4979);
and U5187 (N_5187,N_5067,N_5054);
or U5188 (N_5188,N_4974,N_4960);
nand U5189 (N_5189,N_5088,N_5001);
and U5190 (N_5190,N_5021,N_5072);
nand U5191 (N_5191,N_5103,N_5083);
and U5192 (N_5192,N_5029,N_5019);
or U5193 (N_5193,N_4997,N_5057);
nand U5194 (N_5194,N_5039,N_4970);
and U5195 (N_5195,N_5064,N_5066);
nor U5196 (N_5196,N_5006,N_5025);
and U5197 (N_5197,N_5030,N_4984);
nand U5198 (N_5198,N_4981,N_5015);
or U5199 (N_5199,N_4968,N_5007);
xnor U5200 (N_5200,N_5049,N_4986);
and U5201 (N_5201,N_4995,N_5078);
or U5202 (N_5202,N_4973,N_5064);
nand U5203 (N_5203,N_5001,N_4964);
or U5204 (N_5204,N_5089,N_5017);
or U5205 (N_5205,N_5107,N_4999);
or U5206 (N_5206,N_5002,N_5087);
or U5207 (N_5207,N_4992,N_5061);
and U5208 (N_5208,N_5002,N_5108);
and U5209 (N_5209,N_5048,N_5057);
xor U5210 (N_5210,N_5019,N_5053);
nor U5211 (N_5211,N_4983,N_5029);
nand U5212 (N_5212,N_5112,N_5045);
or U5213 (N_5213,N_5103,N_5098);
xnor U5214 (N_5214,N_5025,N_5071);
and U5215 (N_5215,N_5029,N_5071);
and U5216 (N_5216,N_4967,N_5119);
nand U5217 (N_5217,N_5119,N_5080);
or U5218 (N_5218,N_4988,N_5082);
nor U5219 (N_5219,N_5102,N_5011);
and U5220 (N_5220,N_5074,N_5039);
xnor U5221 (N_5221,N_4995,N_5033);
and U5222 (N_5222,N_4991,N_5088);
or U5223 (N_5223,N_4997,N_5050);
nor U5224 (N_5224,N_5055,N_5077);
or U5225 (N_5225,N_4973,N_5015);
nand U5226 (N_5226,N_5016,N_5073);
xor U5227 (N_5227,N_5083,N_5073);
nor U5228 (N_5228,N_5081,N_5038);
nand U5229 (N_5229,N_5081,N_4973);
or U5230 (N_5230,N_5001,N_5092);
nand U5231 (N_5231,N_5102,N_5098);
xnor U5232 (N_5232,N_5028,N_5104);
nand U5233 (N_5233,N_4966,N_5111);
nor U5234 (N_5234,N_5076,N_5072);
or U5235 (N_5235,N_5029,N_5020);
and U5236 (N_5236,N_5038,N_5000);
and U5237 (N_5237,N_5054,N_5018);
nor U5238 (N_5238,N_5047,N_5102);
and U5239 (N_5239,N_4961,N_5050);
nor U5240 (N_5240,N_5081,N_5013);
nand U5241 (N_5241,N_4984,N_4971);
and U5242 (N_5242,N_5037,N_5076);
nor U5243 (N_5243,N_5085,N_5089);
or U5244 (N_5244,N_5075,N_4971);
nand U5245 (N_5245,N_4973,N_5110);
nor U5246 (N_5246,N_5046,N_5068);
xnor U5247 (N_5247,N_4960,N_5039);
or U5248 (N_5248,N_5064,N_5112);
nor U5249 (N_5249,N_5043,N_4974);
nor U5250 (N_5250,N_5040,N_5113);
nand U5251 (N_5251,N_4996,N_5068);
or U5252 (N_5252,N_4985,N_5037);
or U5253 (N_5253,N_5020,N_5044);
nor U5254 (N_5254,N_5022,N_5037);
nand U5255 (N_5255,N_5015,N_5111);
and U5256 (N_5256,N_5036,N_5097);
or U5257 (N_5257,N_5007,N_5087);
nor U5258 (N_5258,N_5097,N_5073);
nor U5259 (N_5259,N_5113,N_5033);
or U5260 (N_5260,N_5032,N_4978);
or U5261 (N_5261,N_5093,N_5005);
and U5262 (N_5262,N_5038,N_5027);
nor U5263 (N_5263,N_5054,N_4966);
and U5264 (N_5264,N_5083,N_4974);
and U5265 (N_5265,N_5099,N_5052);
and U5266 (N_5266,N_5044,N_5083);
and U5267 (N_5267,N_4971,N_5043);
nor U5268 (N_5268,N_5093,N_5035);
or U5269 (N_5269,N_5025,N_4972);
nor U5270 (N_5270,N_4970,N_5075);
or U5271 (N_5271,N_5105,N_4980);
or U5272 (N_5272,N_4990,N_5080);
or U5273 (N_5273,N_4972,N_5115);
nand U5274 (N_5274,N_5100,N_5088);
nor U5275 (N_5275,N_5103,N_5084);
nand U5276 (N_5276,N_5082,N_4969);
and U5277 (N_5277,N_5109,N_4994);
nand U5278 (N_5278,N_5046,N_5107);
and U5279 (N_5279,N_5020,N_4966);
or U5280 (N_5280,N_5257,N_5218);
and U5281 (N_5281,N_5207,N_5202);
or U5282 (N_5282,N_5197,N_5128);
or U5283 (N_5283,N_5227,N_5165);
nand U5284 (N_5284,N_5251,N_5185);
nor U5285 (N_5285,N_5245,N_5153);
nor U5286 (N_5286,N_5252,N_5198);
or U5287 (N_5287,N_5130,N_5215);
or U5288 (N_5288,N_5146,N_5135);
nand U5289 (N_5289,N_5125,N_5145);
and U5290 (N_5290,N_5126,N_5138);
xor U5291 (N_5291,N_5271,N_5244);
or U5292 (N_5292,N_5231,N_5166);
nor U5293 (N_5293,N_5256,N_5200);
nor U5294 (N_5294,N_5206,N_5167);
and U5295 (N_5295,N_5176,N_5188);
nand U5296 (N_5296,N_5238,N_5144);
nor U5297 (N_5297,N_5219,N_5246);
nor U5298 (N_5298,N_5234,N_5139);
nor U5299 (N_5299,N_5249,N_5241);
nand U5300 (N_5300,N_5232,N_5154);
or U5301 (N_5301,N_5201,N_5260);
or U5302 (N_5302,N_5225,N_5140);
and U5303 (N_5303,N_5248,N_5132);
nand U5304 (N_5304,N_5278,N_5191);
or U5305 (N_5305,N_5211,N_5272);
or U5306 (N_5306,N_5228,N_5242);
and U5307 (N_5307,N_5254,N_5155);
xnor U5308 (N_5308,N_5216,N_5212);
or U5309 (N_5309,N_5121,N_5157);
or U5310 (N_5310,N_5179,N_5262);
nand U5311 (N_5311,N_5186,N_5269);
or U5312 (N_5312,N_5273,N_5226);
and U5313 (N_5313,N_5168,N_5190);
nor U5314 (N_5314,N_5123,N_5181);
xor U5315 (N_5315,N_5152,N_5265);
nand U5316 (N_5316,N_5214,N_5208);
and U5317 (N_5317,N_5187,N_5134);
nor U5318 (N_5318,N_5131,N_5220);
xor U5319 (N_5319,N_5129,N_5266);
nor U5320 (N_5320,N_5163,N_5259);
xnor U5321 (N_5321,N_5224,N_5173);
and U5322 (N_5322,N_5223,N_5170);
nor U5323 (N_5323,N_5221,N_5268);
or U5324 (N_5324,N_5124,N_5237);
nor U5325 (N_5325,N_5189,N_5160);
nand U5326 (N_5326,N_5171,N_5196);
xnor U5327 (N_5327,N_5164,N_5258);
nand U5328 (N_5328,N_5210,N_5235);
and U5329 (N_5329,N_5137,N_5279);
and U5330 (N_5330,N_5240,N_5239);
nand U5331 (N_5331,N_5120,N_5205);
and U5332 (N_5332,N_5178,N_5243);
nor U5333 (N_5333,N_5275,N_5158);
or U5334 (N_5334,N_5194,N_5172);
and U5335 (N_5335,N_5276,N_5141);
xor U5336 (N_5336,N_5222,N_5270);
or U5337 (N_5337,N_5195,N_5143);
nor U5338 (N_5338,N_5230,N_5149);
and U5339 (N_5339,N_5263,N_5151);
and U5340 (N_5340,N_5236,N_5255);
or U5341 (N_5341,N_5147,N_5133);
and U5342 (N_5342,N_5253,N_5277);
or U5343 (N_5343,N_5209,N_5148);
nor U5344 (N_5344,N_5142,N_5203);
or U5345 (N_5345,N_5156,N_5261);
xnor U5346 (N_5346,N_5182,N_5175);
nor U5347 (N_5347,N_5184,N_5127);
nor U5348 (N_5348,N_5122,N_5250);
nor U5349 (N_5349,N_5183,N_5161);
nor U5350 (N_5350,N_5174,N_5229);
nand U5351 (N_5351,N_5162,N_5233);
nand U5352 (N_5352,N_5264,N_5247);
nor U5353 (N_5353,N_5217,N_5213);
or U5354 (N_5354,N_5199,N_5180);
xnor U5355 (N_5355,N_5193,N_5177);
nor U5356 (N_5356,N_5274,N_5136);
or U5357 (N_5357,N_5267,N_5169);
and U5358 (N_5358,N_5204,N_5150);
nand U5359 (N_5359,N_5159,N_5192);
nand U5360 (N_5360,N_5178,N_5180);
or U5361 (N_5361,N_5211,N_5121);
nand U5362 (N_5362,N_5196,N_5199);
and U5363 (N_5363,N_5194,N_5121);
nand U5364 (N_5364,N_5144,N_5245);
nand U5365 (N_5365,N_5218,N_5251);
or U5366 (N_5366,N_5223,N_5269);
or U5367 (N_5367,N_5157,N_5150);
xor U5368 (N_5368,N_5253,N_5124);
and U5369 (N_5369,N_5132,N_5236);
and U5370 (N_5370,N_5196,N_5233);
nand U5371 (N_5371,N_5142,N_5187);
or U5372 (N_5372,N_5178,N_5254);
and U5373 (N_5373,N_5269,N_5142);
nor U5374 (N_5374,N_5253,N_5130);
nand U5375 (N_5375,N_5166,N_5213);
nand U5376 (N_5376,N_5123,N_5206);
xnor U5377 (N_5377,N_5240,N_5231);
xor U5378 (N_5378,N_5260,N_5253);
and U5379 (N_5379,N_5229,N_5130);
and U5380 (N_5380,N_5233,N_5174);
nand U5381 (N_5381,N_5130,N_5249);
and U5382 (N_5382,N_5144,N_5137);
nand U5383 (N_5383,N_5141,N_5127);
nor U5384 (N_5384,N_5159,N_5271);
nor U5385 (N_5385,N_5150,N_5120);
and U5386 (N_5386,N_5191,N_5164);
or U5387 (N_5387,N_5131,N_5180);
nor U5388 (N_5388,N_5163,N_5121);
nor U5389 (N_5389,N_5192,N_5209);
nand U5390 (N_5390,N_5270,N_5126);
or U5391 (N_5391,N_5237,N_5254);
and U5392 (N_5392,N_5245,N_5195);
or U5393 (N_5393,N_5245,N_5213);
nand U5394 (N_5394,N_5131,N_5135);
xnor U5395 (N_5395,N_5276,N_5236);
or U5396 (N_5396,N_5172,N_5129);
and U5397 (N_5397,N_5171,N_5240);
nor U5398 (N_5398,N_5210,N_5128);
and U5399 (N_5399,N_5198,N_5124);
nor U5400 (N_5400,N_5122,N_5185);
nor U5401 (N_5401,N_5165,N_5180);
nand U5402 (N_5402,N_5189,N_5255);
and U5403 (N_5403,N_5186,N_5169);
nor U5404 (N_5404,N_5224,N_5241);
nand U5405 (N_5405,N_5206,N_5215);
nor U5406 (N_5406,N_5265,N_5262);
and U5407 (N_5407,N_5256,N_5252);
nor U5408 (N_5408,N_5252,N_5148);
and U5409 (N_5409,N_5156,N_5186);
nand U5410 (N_5410,N_5194,N_5128);
nand U5411 (N_5411,N_5138,N_5133);
or U5412 (N_5412,N_5181,N_5182);
nand U5413 (N_5413,N_5220,N_5228);
and U5414 (N_5414,N_5243,N_5262);
nor U5415 (N_5415,N_5238,N_5181);
nor U5416 (N_5416,N_5200,N_5219);
nand U5417 (N_5417,N_5235,N_5209);
nor U5418 (N_5418,N_5198,N_5135);
and U5419 (N_5419,N_5125,N_5194);
nor U5420 (N_5420,N_5171,N_5205);
nor U5421 (N_5421,N_5234,N_5262);
and U5422 (N_5422,N_5154,N_5133);
nor U5423 (N_5423,N_5190,N_5223);
nand U5424 (N_5424,N_5220,N_5147);
and U5425 (N_5425,N_5179,N_5217);
and U5426 (N_5426,N_5206,N_5223);
and U5427 (N_5427,N_5278,N_5201);
and U5428 (N_5428,N_5123,N_5233);
and U5429 (N_5429,N_5198,N_5213);
nor U5430 (N_5430,N_5132,N_5158);
nand U5431 (N_5431,N_5217,N_5192);
and U5432 (N_5432,N_5196,N_5148);
and U5433 (N_5433,N_5189,N_5271);
or U5434 (N_5434,N_5232,N_5127);
or U5435 (N_5435,N_5272,N_5129);
nand U5436 (N_5436,N_5255,N_5192);
nand U5437 (N_5437,N_5216,N_5204);
nor U5438 (N_5438,N_5145,N_5168);
and U5439 (N_5439,N_5236,N_5196);
nand U5440 (N_5440,N_5375,N_5434);
nor U5441 (N_5441,N_5295,N_5344);
or U5442 (N_5442,N_5326,N_5283);
and U5443 (N_5443,N_5370,N_5289);
nand U5444 (N_5444,N_5401,N_5365);
nor U5445 (N_5445,N_5332,N_5406);
or U5446 (N_5446,N_5421,N_5372);
xor U5447 (N_5447,N_5320,N_5296);
or U5448 (N_5448,N_5417,N_5394);
xnor U5449 (N_5449,N_5281,N_5398);
and U5450 (N_5450,N_5363,N_5408);
nand U5451 (N_5451,N_5354,N_5306);
nor U5452 (N_5452,N_5390,N_5369);
nor U5453 (N_5453,N_5403,N_5302);
nor U5454 (N_5454,N_5395,N_5414);
or U5455 (N_5455,N_5437,N_5366);
nor U5456 (N_5456,N_5399,N_5345);
and U5457 (N_5457,N_5282,N_5310);
nand U5458 (N_5458,N_5315,N_5330);
nand U5459 (N_5459,N_5364,N_5386);
nor U5460 (N_5460,N_5341,N_5313);
and U5461 (N_5461,N_5318,N_5329);
nor U5462 (N_5462,N_5409,N_5382);
or U5463 (N_5463,N_5424,N_5284);
or U5464 (N_5464,N_5351,N_5342);
nor U5465 (N_5465,N_5438,N_5361);
xor U5466 (N_5466,N_5359,N_5339);
nand U5467 (N_5467,N_5294,N_5307);
nand U5468 (N_5468,N_5299,N_5391);
xnor U5469 (N_5469,N_5431,N_5348);
and U5470 (N_5470,N_5422,N_5300);
and U5471 (N_5471,N_5298,N_5439);
and U5472 (N_5472,N_5407,N_5380);
nor U5473 (N_5473,N_5353,N_5356);
nor U5474 (N_5474,N_5423,N_5290);
nand U5475 (N_5475,N_5378,N_5385);
xnor U5476 (N_5476,N_5288,N_5362);
nand U5477 (N_5477,N_5387,N_5308);
and U5478 (N_5478,N_5303,N_5349);
nor U5479 (N_5479,N_5384,N_5331);
nor U5480 (N_5480,N_5286,N_5343);
or U5481 (N_5481,N_5413,N_5373);
and U5482 (N_5482,N_5418,N_5396);
and U5483 (N_5483,N_5368,N_5381);
nand U5484 (N_5484,N_5404,N_5425);
xnor U5485 (N_5485,N_5352,N_5435);
xor U5486 (N_5486,N_5350,N_5333);
and U5487 (N_5487,N_5371,N_5293);
or U5488 (N_5488,N_5301,N_5357);
nand U5489 (N_5489,N_5292,N_5327);
nand U5490 (N_5490,N_5383,N_5392);
xnor U5491 (N_5491,N_5374,N_5334);
nand U5492 (N_5492,N_5402,N_5346);
and U5493 (N_5493,N_5416,N_5388);
nand U5494 (N_5494,N_5347,N_5287);
or U5495 (N_5495,N_5328,N_5317);
and U5496 (N_5496,N_5436,N_5410);
and U5497 (N_5497,N_5314,N_5291);
nor U5498 (N_5498,N_5337,N_5311);
xor U5499 (N_5499,N_5304,N_5412);
or U5500 (N_5500,N_5432,N_5325);
and U5501 (N_5501,N_5321,N_5335);
nand U5502 (N_5502,N_5336,N_5367);
nor U5503 (N_5503,N_5309,N_5280);
xor U5504 (N_5504,N_5397,N_5360);
nand U5505 (N_5505,N_5340,N_5322);
nand U5506 (N_5506,N_5324,N_5379);
nand U5507 (N_5507,N_5377,N_5426);
xor U5508 (N_5508,N_5415,N_5419);
nor U5509 (N_5509,N_5323,N_5427);
nor U5510 (N_5510,N_5312,N_5376);
and U5511 (N_5511,N_5411,N_5285);
and U5512 (N_5512,N_5319,N_5433);
or U5513 (N_5513,N_5405,N_5389);
or U5514 (N_5514,N_5393,N_5316);
or U5515 (N_5515,N_5358,N_5355);
and U5516 (N_5516,N_5297,N_5400);
nand U5517 (N_5517,N_5430,N_5338);
and U5518 (N_5518,N_5420,N_5429);
or U5519 (N_5519,N_5305,N_5428);
or U5520 (N_5520,N_5404,N_5413);
nor U5521 (N_5521,N_5417,N_5423);
xor U5522 (N_5522,N_5380,N_5357);
and U5523 (N_5523,N_5421,N_5437);
nor U5524 (N_5524,N_5435,N_5288);
or U5525 (N_5525,N_5380,N_5304);
or U5526 (N_5526,N_5291,N_5364);
nand U5527 (N_5527,N_5420,N_5319);
nor U5528 (N_5528,N_5410,N_5404);
nand U5529 (N_5529,N_5337,N_5363);
nand U5530 (N_5530,N_5287,N_5394);
and U5531 (N_5531,N_5387,N_5285);
nand U5532 (N_5532,N_5425,N_5421);
and U5533 (N_5533,N_5333,N_5410);
or U5534 (N_5534,N_5309,N_5370);
and U5535 (N_5535,N_5336,N_5410);
or U5536 (N_5536,N_5439,N_5384);
nand U5537 (N_5537,N_5424,N_5403);
or U5538 (N_5538,N_5374,N_5409);
and U5539 (N_5539,N_5430,N_5303);
nand U5540 (N_5540,N_5352,N_5385);
nor U5541 (N_5541,N_5439,N_5320);
nand U5542 (N_5542,N_5382,N_5289);
or U5543 (N_5543,N_5427,N_5435);
nor U5544 (N_5544,N_5335,N_5331);
or U5545 (N_5545,N_5364,N_5375);
and U5546 (N_5546,N_5374,N_5390);
nor U5547 (N_5547,N_5329,N_5438);
nor U5548 (N_5548,N_5398,N_5358);
or U5549 (N_5549,N_5411,N_5310);
or U5550 (N_5550,N_5324,N_5354);
or U5551 (N_5551,N_5406,N_5308);
nand U5552 (N_5552,N_5348,N_5374);
nor U5553 (N_5553,N_5398,N_5387);
nand U5554 (N_5554,N_5312,N_5421);
xor U5555 (N_5555,N_5362,N_5330);
nor U5556 (N_5556,N_5356,N_5381);
nor U5557 (N_5557,N_5313,N_5406);
nor U5558 (N_5558,N_5311,N_5374);
or U5559 (N_5559,N_5414,N_5401);
nor U5560 (N_5560,N_5358,N_5357);
nor U5561 (N_5561,N_5397,N_5329);
nand U5562 (N_5562,N_5289,N_5310);
and U5563 (N_5563,N_5413,N_5286);
nor U5564 (N_5564,N_5408,N_5335);
nand U5565 (N_5565,N_5370,N_5402);
xnor U5566 (N_5566,N_5403,N_5379);
and U5567 (N_5567,N_5328,N_5365);
or U5568 (N_5568,N_5371,N_5288);
nand U5569 (N_5569,N_5366,N_5375);
nor U5570 (N_5570,N_5365,N_5402);
or U5571 (N_5571,N_5353,N_5285);
xnor U5572 (N_5572,N_5384,N_5306);
or U5573 (N_5573,N_5297,N_5300);
nor U5574 (N_5574,N_5310,N_5291);
or U5575 (N_5575,N_5309,N_5354);
and U5576 (N_5576,N_5344,N_5328);
or U5577 (N_5577,N_5385,N_5392);
nand U5578 (N_5578,N_5393,N_5290);
xnor U5579 (N_5579,N_5375,N_5423);
and U5580 (N_5580,N_5339,N_5394);
or U5581 (N_5581,N_5422,N_5289);
nor U5582 (N_5582,N_5364,N_5430);
and U5583 (N_5583,N_5374,N_5297);
nand U5584 (N_5584,N_5333,N_5364);
xor U5585 (N_5585,N_5350,N_5407);
xnor U5586 (N_5586,N_5333,N_5433);
and U5587 (N_5587,N_5352,N_5378);
nor U5588 (N_5588,N_5297,N_5394);
and U5589 (N_5589,N_5363,N_5388);
nand U5590 (N_5590,N_5327,N_5419);
and U5591 (N_5591,N_5293,N_5298);
or U5592 (N_5592,N_5373,N_5299);
xor U5593 (N_5593,N_5343,N_5393);
nor U5594 (N_5594,N_5396,N_5413);
or U5595 (N_5595,N_5367,N_5429);
or U5596 (N_5596,N_5299,N_5306);
or U5597 (N_5597,N_5423,N_5320);
and U5598 (N_5598,N_5380,N_5303);
xor U5599 (N_5599,N_5414,N_5314);
xor U5600 (N_5600,N_5571,N_5562);
or U5601 (N_5601,N_5593,N_5485);
or U5602 (N_5602,N_5526,N_5537);
nand U5603 (N_5603,N_5587,N_5583);
nor U5604 (N_5604,N_5547,N_5484);
xnor U5605 (N_5605,N_5440,N_5543);
or U5606 (N_5606,N_5575,N_5464);
and U5607 (N_5607,N_5539,N_5447);
xnor U5608 (N_5608,N_5466,N_5495);
nor U5609 (N_5609,N_5560,N_5565);
or U5610 (N_5610,N_5568,N_5468);
and U5611 (N_5611,N_5445,N_5460);
nand U5612 (N_5612,N_5519,N_5556);
nand U5613 (N_5613,N_5536,N_5553);
and U5614 (N_5614,N_5480,N_5597);
and U5615 (N_5615,N_5554,N_5463);
or U5616 (N_5616,N_5467,N_5598);
or U5617 (N_5617,N_5588,N_5572);
nor U5618 (N_5618,N_5589,N_5532);
nand U5619 (N_5619,N_5591,N_5465);
nor U5620 (N_5620,N_5496,N_5514);
nor U5621 (N_5621,N_5492,N_5599);
nor U5622 (N_5622,N_5549,N_5552);
or U5623 (N_5623,N_5517,N_5444);
and U5624 (N_5624,N_5584,N_5570);
or U5625 (N_5625,N_5513,N_5511);
nand U5626 (N_5626,N_5475,N_5450);
and U5627 (N_5627,N_5566,N_5472);
nor U5628 (N_5628,N_5520,N_5541);
and U5629 (N_5629,N_5500,N_5493);
nor U5630 (N_5630,N_5442,N_5452);
xor U5631 (N_5631,N_5506,N_5594);
nand U5632 (N_5632,N_5557,N_5573);
and U5633 (N_5633,N_5550,N_5479);
and U5634 (N_5634,N_5503,N_5459);
and U5635 (N_5635,N_5592,N_5497);
nand U5636 (N_5636,N_5527,N_5574);
or U5637 (N_5637,N_5544,N_5505);
or U5638 (N_5638,N_5561,N_5596);
nor U5639 (N_5639,N_5462,N_5451);
or U5640 (N_5640,N_5489,N_5457);
nor U5641 (N_5641,N_5579,N_5508);
nor U5642 (N_5642,N_5487,N_5559);
nor U5643 (N_5643,N_5478,N_5454);
or U5644 (N_5644,N_5471,N_5453);
nor U5645 (N_5645,N_5481,N_5538);
or U5646 (N_5646,N_5469,N_5491);
nor U5647 (N_5647,N_5456,N_5576);
and U5648 (N_5648,N_5586,N_5446);
xor U5649 (N_5649,N_5461,N_5585);
xor U5650 (N_5650,N_5515,N_5507);
nor U5651 (N_5651,N_5490,N_5494);
or U5652 (N_5652,N_5521,N_5581);
and U5653 (N_5653,N_5474,N_5595);
nor U5654 (N_5654,N_5533,N_5501);
and U5655 (N_5655,N_5590,N_5545);
and U5656 (N_5656,N_5555,N_5486);
nor U5657 (N_5657,N_5577,N_5523);
or U5658 (N_5658,N_5529,N_5551);
nor U5659 (N_5659,N_5441,N_5516);
and U5660 (N_5660,N_5542,N_5528);
and U5661 (N_5661,N_5499,N_5510);
nor U5662 (N_5662,N_5531,N_5518);
or U5663 (N_5663,N_5455,N_5564);
nor U5664 (N_5664,N_5548,N_5502);
xnor U5665 (N_5665,N_5578,N_5567);
or U5666 (N_5666,N_5558,N_5509);
nor U5667 (N_5667,N_5477,N_5504);
xnor U5668 (N_5668,N_5534,N_5498);
nand U5669 (N_5669,N_5540,N_5473);
xor U5670 (N_5670,N_5470,N_5530);
or U5671 (N_5671,N_5483,N_5522);
nor U5672 (N_5672,N_5582,N_5535);
nor U5673 (N_5673,N_5476,N_5449);
or U5674 (N_5674,N_5546,N_5524);
nand U5675 (N_5675,N_5482,N_5580);
nand U5676 (N_5676,N_5563,N_5448);
or U5677 (N_5677,N_5512,N_5525);
and U5678 (N_5678,N_5458,N_5488);
and U5679 (N_5679,N_5443,N_5569);
nor U5680 (N_5680,N_5502,N_5580);
nand U5681 (N_5681,N_5522,N_5521);
nor U5682 (N_5682,N_5476,N_5573);
xor U5683 (N_5683,N_5589,N_5551);
or U5684 (N_5684,N_5482,N_5450);
and U5685 (N_5685,N_5561,N_5542);
or U5686 (N_5686,N_5599,N_5580);
nor U5687 (N_5687,N_5463,N_5591);
and U5688 (N_5688,N_5519,N_5463);
and U5689 (N_5689,N_5539,N_5564);
nand U5690 (N_5690,N_5546,N_5568);
nor U5691 (N_5691,N_5510,N_5472);
or U5692 (N_5692,N_5594,N_5565);
or U5693 (N_5693,N_5446,N_5482);
and U5694 (N_5694,N_5440,N_5560);
xnor U5695 (N_5695,N_5516,N_5574);
xor U5696 (N_5696,N_5592,N_5501);
nand U5697 (N_5697,N_5507,N_5577);
nor U5698 (N_5698,N_5458,N_5547);
or U5699 (N_5699,N_5476,N_5547);
and U5700 (N_5700,N_5590,N_5457);
and U5701 (N_5701,N_5521,N_5567);
nor U5702 (N_5702,N_5580,N_5520);
or U5703 (N_5703,N_5528,N_5483);
nand U5704 (N_5704,N_5497,N_5530);
and U5705 (N_5705,N_5452,N_5461);
and U5706 (N_5706,N_5478,N_5501);
nor U5707 (N_5707,N_5540,N_5552);
nand U5708 (N_5708,N_5574,N_5531);
nor U5709 (N_5709,N_5488,N_5562);
nor U5710 (N_5710,N_5463,N_5449);
and U5711 (N_5711,N_5556,N_5520);
xor U5712 (N_5712,N_5502,N_5515);
nor U5713 (N_5713,N_5524,N_5503);
and U5714 (N_5714,N_5473,N_5499);
and U5715 (N_5715,N_5492,N_5484);
nor U5716 (N_5716,N_5523,N_5498);
nor U5717 (N_5717,N_5524,N_5543);
nand U5718 (N_5718,N_5583,N_5558);
nor U5719 (N_5719,N_5497,N_5472);
and U5720 (N_5720,N_5447,N_5545);
nand U5721 (N_5721,N_5501,N_5549);
nor U5722 (N_5722,N_5491,N_5554);
or U5723 (N_5723,N_5518,N_5579);
nor U5724 (N_5724,N_5441,N_5577);
xor U5725 (N_5725,N_5452,N_5593);
xnor U5726 (N_5726,N_5503,N_5578);
nand U5727 (N_5727,N_5581,N_5501);
nor U5728 (N_5728,N_5584,N_5491);
nand U5729 (N_5729,N_5469,N_5591);
and U5730 (N_5730,N_5517,N_5552);
or U5731 (N_5731,N_5563,N_5494);
nor U5732 (N_5732,N_5447,N_5592);
nand U5733 (N_5733,N_5595,N_5479);
nand U5734 (N_5734,N_5484,N_5550);
nand U5735 (N_5735,N_5441,N_5466);
nand U5736 (N_5736,N_5523,N_5461);
nor U5737 (N_5737,N_5590,N_5515);
and U5738 (N_5738,N_5461,N_5573);
nand U5739 (N_5739,N_5549,N_5498);
or U5740 (N_5740,N_5564,N_5481);
or U5741 (N_5741,N_5576,N_5445);
xor U5742 (N_5742,N_5529,N_5544);
xnor U5743 (N_5743,N_5517,N_5442);
and U5744 (N_5744,N_5593,N_5509);
or U5745 (N_5745,N_5573,N_5567);
nand U5746 (N_5746,N_5445,N_5522);
nand U5747 (N_5747,N_5585,N_5497);
or U5748 (N_5748,N_5562,N_5568);
or U5749 (N_5749,N_5536,N_5576);
xor U5750 (N_5750,N_5478,N_5489);
xnor U5751 (N_5751,N_5573,N_5520);
and U5752 (N_5752,N_5512,N_5533);
xor U5753 (N_5753,N_5584,N_5450);
or U5754 (N_5754,N_5478,N_5576);
nand U5755 (N_5755,N_5522,N_5459);
nand U5756 (N_5756,N_5455,N_5588);
xnor U5757 (N_5757,N_5510,N_5482);
xor U5758 (N_5758,N_5565,N_5531);
nor U5759 (N_5759,N_5479,N_5443);
and U5760 (N_5760,N_5681,N_5610);
nand U5761 (N_5761,N_5657,N_5615);
nand U5762 (N_5762,N_5653,N_5611);
nand U5763 (N_5763,N_5753,N_5680);
or U5764 (N_5764,N_5658,N_5656);
and U5765 (N_5765,N_5624,N_5743);
nor U5766 (N_5766,N_5660,N_5701);
or U5767 (N_5767,N_5637,N_5634);
or U5768 (N_5768,N_5718,N_5751);
and U5769 (N_5769,N_5729,N_5754);
nand U5770 (N_5770,N_5725,N_5750);
or U5771 (N_5771,N_5709,N_5626);
nor U5772 (N_5772,N_5670,N_5691);
nor U5773 (N_5773,N_5689,N_5647);
or U5774 (N_5774,N_5694,N_5607);
nor U5775 (N_5775,N_5655,N_5742);
and U5776 (N_5776,N_5652,N_5695);
and U5777 (N_5777,N_5744,N_5621);
xor U5778 (N_5778,N_5711,N_5665);
nand U5779 (N_5779,N_5662,N_5667);
nor U5780 (N_5780,N_5757,N_5629);
or U5781 (N_5781,N_5666,N_5697);
nor U5782 (N_5782,N_5622,N_5687);
and U5783 (N_5783,N_5759,N_5685);
and U5784 (N_5784,N_5734,N_5726);
nand U5785 (N_5785,N_5715,N_5678);
or U5786 (N_5786,N_5640,N_5638);
and U5787 (N_5787,N_5616,N_5748);
nor U5788 (N_5788,N_5693,N_5682);
nor U5789 (N_5789,N_5738,N_5749);
nor U5790 (N_5790,N_5641,N_5716);
nor U5791 (N_5791,N_5747,N_5605);
and U5792 (N_5792,N_5730,N_5713);
and U5793 (N_5793,N_5632,N_5603);
nand U5794 (N_5794,N_5746,N_5731);
and U5795 (N_5795,N_5752,N_5609);
nand U5796 (N_5796,N_5645,N_5646);
or U5797 (N_5797,N_5673,N_5704);
nand U5798 (N_5798,N_5740,N_5712);
nor U5799 (N_5799,N_5733,N_5618);
nand U5800 (N_5800,N_5649,N_5698);
nand U5801 (N_5801,N_5699,N_5724);
nand U5802 (N_5802,N_5684,N_5636);
nor U5803 (N_5803,N_5688,N_5700);
or U5804 (N_5804,N_5679,N_5613);
xnor U5805 (N_5805,N_5625,N_5620);
or U5806 (N_5806,N_5735,N_5676);
nor U5807 (N_5807,N_5635,N_5732);
or U5808 (N_5808,N_5614,N_5669);
xnor U5809 (N_5809,N_5722,N_5604);
or U5810 (N_5810,N_5648,N_5756);
nor U5811 (N_5811,N_5642,N_5719);
nor U5812 (N_5812,N_5602,N_5692);
xor U5813 (N_5813,N_5643,N_5674);
and U5814 (N_5814,N_5651,N_5737);
nand U5815 (N_5815,N_5623,N_5714);
nand U5816 (N_5816,N_5686,N_5721);
and U5817 (N_5817,N_5664,N_5675);
xor U5818 (N_5818,N_5755,N_5668);
and U5819 (N_5819,N_5606,N_5612);
or U5820 (N_5820,N_5703,N_5617);
or U5821 (N_5821,N_5627,N_5601);
or U5822 (N_5822,N_5739,N_5663);
nand U5823 (N_5823,N_5671,N_5672);
and U5824 (N_5824,N_5619,N_5723);
and U5825 (N_5825,N_5661,N_5644);
nor U5826 (N_5826,N_5677,N_5720);
and U5827 (N_5827,N_5628,N_5745);
nand U5828 (N_5828,N_5633,N_5728);
nand U5829 (N_5829,N_5631,N_5630);
and U5830 (N_5830,N_5650,N_5710);
nand U5831 (N_5831,N_5727,N_5741);
nand U5832 (N_5832,N_5708,N_5608);
and U5833 (N_5833,N_5702,N_5706);
nor U5834 (N_5834,N_5639,N_5717);
or U5835 (N_5835,N_5690,N_5696);
or U5836 (N_5836,N_5758,N_5683);
or U5837 (N_5837,N_5705,N_5654);
or U5838 (N_5838,N_5600,N_5736);
nor U5839 (N_5839,N_5659,N_5707);
and U5840 (N_5840,N_5610,N_5645);
nand U5841 (N_5841,N_5683,N_5732);
nand U5842 (N_5842,N_5627,N_5689);
nor U5843 (N_5843,N_5718,N_5637);
and U5844 (N_5844,N_5659,N_5684);
or U5845 (N_5845,N_5697,N_5717);
and U5846 (N_5846,N_5645,N_5683);
or U5847 (N_5847,N_5610,N_5601);
or U5848 (N_5848,N_5682,N_5648);
nand U5849 (N_5849,N_5728,N_5758);
and U5850 (N_5850,N_5671,N_5607);
nor U5851 (N_5851,N_5674,N_5675);
and U5852 (N_5852,N_5644,N_5746);
or U5853 (N_5853,N_5645,N_5687);
nand U5854 (N_5854,N_5650,N_5638);
nand U5855 (N_5855,N_5668,N_5752);
nand U5856 (N_5856,N_5657,N_5704);
or U5857 (N_5857,N_5671,N_5708);
nor U5858 (N_5858,N_5734,N_5728);
or U5859 (N_5859,N_5618,N_5743);
nand U5860 (N_5860,N_5706,N_5682);
or U5861 (N_5861,N_5750,N_5615);
nand U5862 (N_5862,N_5658,N_5617);
nand U5863 (N_5863,N_5701,N_5609);
nor U5864 (N_5864,N_5695,N_5685);
and U5865 (N_5865,N_5722,N_5709);
nor U5866 (N_5866,N_5693,N_5743);
and U5867 (N_5867,N_5630,N_5676);
or U5868 (N_5868,N_5739,N_5700);
nand U5869 (N_5869,N_5626,N_5625);
and U5870 (N_5870,N_5679,N_5629);
nand U5871 (N_5871,N_5648,N_5737);
and U5872 (N_5872,N_5662,N_5746);
and U5873 (N_5873,N_5700,N_5713);
nand U5874 (N_5874,N_5634,N_5713);
nand U5875 (N_5875,N_5663,N_5662);
or U5876 (N_5876,N_5684,N_5648);
and U5877 (N_5877,N_5733,N_5608);
nand U5878 (N_5878,N_5735,N_5693);
and U5879 (N_5879,N_5672,N_5738);
nor U5880 (N_5880,N_5681,N_5638);
or U5881 (N_5881,N_5672,N_5702);
or U5882 (N_5882,N_5684,N_5611);
and U5883 (N_5883,N_5685,N_5662);
and U5884 (N_5884,N_5628,N_5734);
nand U5885 (N_5885,N_5657,N_5647);
or U5886 (N_5886,N_5702,N_5719);
or U5887 (N_5887,N_5652,N_5601);
nand U5888 (N_5888,N_5716,N_5632);
and U5889 (N_5889,N_5676,N_5626);
and U5890 (N_5890,N_5658,N_5606);
nor U5891 (N_5891,N_5709,N_5727);
nor U5892 (N_5892,N_5660,N_5726);
xor U5893 (N_5893,N_5606,N_5617);
and U5894 (N_5894,N_5727,N_5634);
xnor U5895 (N_5895,N_5610,N_5618);
and U5896 (N_5896,N_5613,N_5678);
and U5897 (N_5897,N_5682,N_5624);
or U5898 (N_5898,N_5600,N_5652);
or U5899 (N_5899,N_5719,N_5717);
or U5900 (N_5900,N_5668,N_5674);
nand U5901 (N_5901,N_5758,N_5759);
or U5902 (N_5902,N_5621,N_5720);
xor U5903 (N_5903,N_5748,N_5653);
xor U5904 (N_5904,N_5656,N_5679);
xor U5905 (N_5905,N_5637,N_5620);
nor U5906 (N_5906,N_5715,N_5717);
nand U5907 (N_5907,N_5668,N_5642);
or U5908 (N_5908,N_5737,N_5728);
and U5909 (N_5909,N_5672,N_5752);
and U5910 (N_5910,N_5637,N_5644);
nand U5911 (N_5911,N_5609,N_5664);
xnor U5912 (N_5912,N_5661,N_5610);
and U5913 (N_5913,N_5618,N_5604);
nor U5914 (N_5914,N_5674,N_5635);
nand U5915 (N_5915,N_5636,N_5664);
nor U5916 (N_5916,N_5717,N_5735);
xor U5917 (N_5917,N_5757,N_5632);
and U5918 (N_5918,N_5625,N_5753);
and U5919 (N_5919,N_5683,N_5618);
nor U5920 (N_5920,N_5803,N_5788);
nand U5921 (N_5921,N_5894,N_5774);
and U5922 (N_5922,N_5838,N_5886);
nor U5923 (N_5923,N_5876,N_5820);
nor U5924 (N_5924,N_5830,N_5796);
nor U5925 (N_5925,N_5888,N_5871);
or U5926 (N_5926,N_5873,N_5822);
nor U5927 (N_5927,N_5792,N_5835);
and U5928 (N_5928,N_5847,N_5896);
nand U5929 (N_5929,N_5864,N_5891);
or U5930 (N_5930,N_5789,N_5809);
nor U5931 (N_5931,N_5811,N_5904);
nor U5932 (N_5932,N_5780,N_5826);
xor U5933 (N_5933,N_5793,N_5775);
nor U5934 (N_5934,N_5805,N_5797);
or U5935 (N_5935,N_5913,N_5760);
nor U5936 (N_5936,N_5914,N_5808);
or U5937 (N_5937,N_5892,N_5783);
nor U5938 (N_5938,N_5854,N_5860);
nand U5939 (N_5939,N_5846,N_5907);
or U5940 (N_5940,N_5881,N_5802);
and U5941 (N_5941,N_5912,N_5911);
and U5942 (N_5942,N_5762,N_5856);
nand U5943 (N_5943,N_5824,N_5795);
and U5944 (N_5944,N_5867,N_5831);
xnor U5945 (N_5945,N_5767,N_5915);
nand U5946 (N_5946,N_5768,N_5887);
and U5947 (N_5947,N_5816,N_5810);
nand U5948 (N_5948,N_5868,N_5889);
and U5949 (N_5949,N_5885,N_5836);
nand U5950 (N_5950,N_5861,N_5784);
nor U5951 (N_5951,N_5884,N_5776);
nand U5952 (N_5952,N_5895,N_5855);
nor U5953 (N_5953,N_5781,N_5848);
and U5954 (N_5954,N_5770,N_5828);
nand U5955 (N_5955,N_5880,N_5903);
nand U5956 (N_5956,N_5823,N_5817);
nand U5957 (N_5957,N_5813,N_5897);
or U5958 (N_5958,N_5772,N_5844);
or U5959 (N_5959,N_5878,N_5905);
and U5960 (N_5960,N_5778,N_5918);
or U5961 (N_5961,N_5877,N_5839);
or U5962 (N_5962,N_5910,N_5761);
nand U5963 (N_5963,N_5763,N_5827);
or U5964 (N_5964,N_5919,N_5890);
xnor U5965 (N_5965,N_5765,N_5815);
nand U5966 (N_5966,N_5779,N_5842);
and U5967 (N_5967,N_5801,N_5787);
and U5968 (N_5968,N_5832,N_5852);
xnor U5969 (N_5969,N_5840,N_5879);
nand U5970 (N_5970,N_5806,N_5818);
or U5971 (N_5971,N_5804,N_5785);
nand U5972 (N_5972,N_5819,N_5857);
nand U5973 (N_5973,N_5841,N_5814);
xor U5974 (N_5974,N_5851,N_5833);
or U5975 (N_5975,N_5901,N_5917);
and U5976 (N_5976,N_5870,N_5906);
xnor U5977 (N_5977,N_5908,N_5834);
nand U5978 (N_5978,N_5898,N_5859);
nor U5979 (N_5979,N_5798,N_5865);
nor U5980 (N_5980,N_5771,N_5916);
or U5981 (N_5981,N_5862,N_5872);
nor U5982 (N_5982,N_5874,N_5909);
xor U5983 (N_5983,N_5866,N_5821);
nand U5984 (N_5984,N_5863,N_5773);
nand U5985 (N_5985,N_5853,N_5845);
or U5986 (N_5986,N_5858,N_5766);
nand U5987 (N_5987,N_5782,N_5800);
and U5988 (N_5988,N_5882,N_5794);
nor U5989 (N_5989,N_5825,N_5791);
nand U5990 (N_5990,N_5902,N_5843);
nor U5991 (N_5991,N_5893,N_5850);
and U5992 (N_5992,N_5899,N_5777);
xnor U5993 (N_5993,N_5883,N_5812);
nor U5994 (N_5994,N_5799,N_5849);
nand U5995 (N_5995,N_5875,N_5829);
and U5996 (N_5996,N_5869,N_5764);
nand U5997 (N_5997,N_5769,N_5807);
xnor U5998 (N_5998,N_5786,N_5790);
nor U5999 (N_5999,N_5900,N_5837);
and U6000 (N_6000,N_5864,N_5835);
or U6001 (N_6001,N_5831,N_5837);
nor U6002 (N_6002,N_5829,N_5854);
nand U6003 (N_6003,N_5836,N_5887);
or U6004 (N_6004,N_5763,N_5778);
nand U6005 (N_6005,N_5841,N_5851);
xor U6006 (N_6006,N_5776,N_5810);
nor U6007 (N_6007,N_5888,N_5820);
and U6008 (N_6008,N_5804,N_5820);
xnor U6009 (N_6009,N_5850,N_5843);
and U6010 (N_6010,N_5770,N_5818);
and U6011 (N_6011,N_5863,N_5870);
and U6012 (N_6012,N_5776,N_5843);
nor U6013 (N_6013,N_5867,N_5768);
nor U6014 (N_6014,N_5786,N_5854);
nand U6015 (N_6015,N_5839,N_5774);
or U6016 (N_6016,N_5768,N_5823);
and U6017 (N_6017,N_5903,N_5839);
nor U6018 (N_6018,N_5808,N_5861);
and U6019 (N_6019,N_5897,N_5864);
and U6020 (N_6020,N_5867,N_5873);
xor U6021 (N_6021,N_5766,N_5792);
or U6022 (N_6022,N_5875,N_5834);
nand U6023 (N_6023,N_5827,N_5857);
nand U6024 (N_6024,N_5807,N_5888);
nand U6025 (N_6025,N_5809,N_5837);
or U6026 (N_6026,N_5910,N_5847);
and U6027 (N_6027,N_5875,N_5762);
nand U6028 (N_6028,N_5786,N_5897);
and U6029 (N_6029,N_5867,N_5771);
or U6030 (N_6030,N_5830,N_5898);
and U6031 (N_6031,N_5851,N_5891);
and U6032 (N_6032,N_5880,N_5793);
nand U6033 (N_6033,N_5786,N_5855);
or U6034 (N_6034,N_5816,N_5898);
xor U6035 (N_6035,N_5846,N_5914);
nor U6036 (N_6036,N_5795,N_5765);
or U6037 (N_6037,N_5763,N_5856);
and U6038 (N_6038,N_5880,N_5845);
or U6039 (N_6039,N_5918,N_5791);
nor U6040 (N_6040,N_5802,N_5862);
nor U6041 (N_6041,N_5805,N_5760);
and U6042 (N_6042,N_5857,N_5769);
or U6043 (N_6043,N_5891,N_5792);
xnor U6044 (N_6044,N_5864,N_5845);
or U6045 (N_6045,N_5856,N_5877);
and U6046 (N_6046,N_5865,N_5813);
xnor U6047 (N_6047,N_5856,N_5775);
or U6048 (N_6048,N_5868,N_5891);
nor U6049 (N_6049,N_5840,N_5890);
or U6050 (N_6050,N_5780,N_5850);
nand U6051 (N_6051,N_5886,N_5848);
or U6052 (N_6052,N_5865,N_5895);
nand U6053 (N_6053,N_5856,N_5895);
or U6054 (N_6054,N_5887,N_5859);
nand U6055 (N_6055,N_5779,N_5825);
nand U6056 (N_6056,N_5848,N_5795);
nor U6057 (N_6057,N_5827,N_5814);
nand U6058 (N_6058,N_5807,N_5788);
or U6059 (N_6059,N_5796,N_5838);
or U6060 (N_6060,N_5808,N_5863);
or U6061 (N_6061,N_5919,N_5900);
nor U6062 (N_6062,N_5851,N_5795);
and U6063 (N_6063,N_5779,N_5835);
and U6064 (N_6064,N_5817,N_5814);
nand U6065 (N_6065,N_5871,N_5909);
or U6066 (N_6066,N_5799,N_5896);
xor U6067 (N_6067,N_5913,N_5885);
or U6068 (N_6068,N_5807,N_5895);
and U6069 (N_6069,N_5867,N_5887);
or U6070 (N_6070,N_5819,N_5772);
and U6071 (N_6071,N_5782,N_5844);
nor U6072 (N_6072,N_5784,N_5791);
and U6073 (N_6073,N_5823,N_5874);
and U6074 (N_6074,N_5872,N_5805);
nor U6075 (N_6075,N_5817,N_5843);
xnor U6076 (N_6076,N_5887,N_5778);
nor U6077 (N_6077,N_5766,N_5869);
nand U6078 (N_6078,N_5857,N_5878);
and U6079 (N_6079,N_5797,N_5767);
nor U6080 (N_6080,N_5931,N_5942);
nor U6081 (N_6081,N_5996,N_6078);
nand U6082 (N_6082,N_5955,N_6045);
nand U6083 (N_6083,N_6021,N_5971);
nand U6084 (N_6084,N_6015,N_6072);
nand U6085 (N_6085,N_5988,N_5991);
nand U6086 (N_6086,N_5986,N_6044);
or U6087 (N_6087,N_5957,N_6076);
and U6088 (N_6088,N_6057,N_5947);
xnor U6089 (N_6089,N_6056,N_6071);
or U6090 (N_6090,N_5984,N_6037);
nand U6091 (N_6091,N_6011,N_6036);
and U6092 (N_6092,N_5990,N_5946);
or U6093 (N_6093,N_6052,N_6023);
nor U6094 (N_6094,N_6073,N_5983);
or U6095 (N_6095,N_5941,N_5973);
and U6096 (N_6096,N_5970,N_5923);
nor U6097 (N_6097,N_6058,N_5995);
or U6098 (N_6098,N_6001,N_5921);
or U6099 (N_6099,N_6040,N_5920);
or U6100 (N_6100,N_6009,N_5944);
xnor U6101 (N_6101,N_5987,N_6018);
nor U6102 (N_6102,N_6005,N_6019);
xor U6103 (N_6103,N_6033,N_6039);
and U6104 (N_6104,N_5956,N_5963);
nor U6105 (N_6105,N_6065,N_5999);
nor U6106 (N_6106,N_6064,N_6042);
or U6107 (N_6107,N_6074,N_5932);
nor U6108 (N_6108,N_5952,N_5993);
and U6109 (N_6109,N_6066,N_5975);
nand U6110 (N_6110,N_6070,N_6077);
or U6111 (N_6111,N_6026,N_5954);
and U6112 (N_6112,N_6029,N_5969);
xnor U6113 (N_6113,N_5960,N_5974);
xor U6114 (N_6114,N_5994,N_6028);
and U6115 (N_6115,N_6054,N_5981);
nand U6116 (N_6116,N_5989,N_6017);
or U6117 (N_6117,N_6012,N_6038);
nor U6118 (N_6118,N_5937,N_5966);
and U6119 (N_6119,N_6007,N_6079);
xnor U6120 (N_6120,N_6014,N_6030);
and U6121 (N_6121,N_5997,N_6060);
nand U6122 (N_6122,N_6051,N_5951);
xor U6123 (N_6123,N_6003,N_6049);
and U6124 (N_6124,N_5928,N_6069);
nand U6125 (N_6125,N_6025,N_6032);
or U6126 (N_6126,N_6062,N_5934);
nor U6127 (N_6127,N_6020,N_5927);
nor U6128 (N_6128,N_6013,N_5976);
nor U6129 (N_6129,N_5998,N_5948);
nand U6130 (N_6130,N_6024,N_6035);
or U6131 (N_6131,N_6022,N_5992);
and U6132 (N_6132,N_5949,N_6041);
and U6133 (N_6133,N_6048,N_5962);
nand U6134 (N_6134,N_6050,N_5965);
xor U6135 (N_6135,N_6059,N_6006);
nand U6136 (N_6136,N_5939,N_5950);
nand U6137 (N_6137,N_5967,N_6010);
and U6138 (N_6138,N_5925,N_5922);
nand U6139 (N_6139,N_5943,N_5926);
nand U6140 (N_6140,N_6034,N_5929);
nor U6141 (N_6141,N_5935,N_6004);
nand U6142 (N_6142,N_5968,N_5945);
nor U6143 (N_6143,N_5980,N_5978);
or U6144 (N_6144,N_5953,N_6067);
and U6145 (N_6145,N_5930,N_5959);
and U6146 (N_6146,N_5938,N_5936);
nor U6147 (N_6147,N_5977,N_6061);
nand U6148 (N_6148,N_5933,N_6031);
and U6149 (N_6149,N_6075,N_6053);
and U6150 (N_6150,N_5958,N_6046);
xnor U6151 (N_6151,N_6043,N_6002);
nand U6152 (N_6152,N_5972,N_6027);
and U6153 (N_6153,N_5979,N_6068);
xnor U6154 (N_6154,N_6063,N_6008);
and U6155 (N_6155,N_5985,N_5961);
and U6156 (N_6156,N_5982,N_6047);
nand U6157 (N_6157,N_6000,N_5940);
nand U6158 (N_6158,N_5924,N_6055);
and U6159 (N_6159,N_5964,N_6016);
and U6160 (N_6160,N_6045,N_6042);
nor U6161 (N_6161,N_6018,N_5985);
nand U6162 (N_6162,N_6073,N_5991);
and U6163 (N_6163,N_6063,N_6011);
nor U6164 (N_6164,N_5946,N_6015);
or U6165 (N_6165,N_5988,N_6055);
and U6166 (N_6166,N_5944,N_5967);
nand U6167 (N_6167,N_5990,N_5937);
xnor U6168 (N_6168,N_5987,N_5953);
or U6169 (N_6169,N_6053,N_5954);
nor U6170 (N_6170,N_5974,N_5970);
and U6171 (N_6171,N_6079,N_5999);
or U6172 (N_6172,N_6030,N_6063);
nand U6173 (N_6173,N_6043,N_6008);
and U6174 (N_6174,N_6015,N_5937);
nand U6175 (N_6175,N_5921,N_5922);
nand U6176 (N_6176,N_5948,N_6037);
and U6177 (N_6177,N_6054,N_5999);
nor U6178 (N_6178,N_5972,N_5943);
nand U6179 (N_6179,N_5947,N_5989);
and U6180 (N_6180,N_5959,N_6048);
or U6181 (N_6181,N_5995,N_5992);
or U6182 (N_6182,N_6019,N_5957);
or U6183 (N_6183,N_5938,N_6069);
nand U6184 (N_6184,N_5944,N_5956);
and U6185 (N_6185,N_6069,N_6004);
and U6186 (N_6186,N_6040,N_5956);
and U6187 (N_6187,N_5929,N_6038);
nor U6188 (N_6188,N_5966,N_6041);
nor U6189 (N_6189,N_6038,N_6054);
nand U6190 (N_6190,N_5967,N_5926);
and U6191 (N_6191,N_6006,N_6068);
and U6192 (N_6192,N_6004,N_6009);
and U6193 (N_6193,N_6028,N_6006);
and U6194 (N_6194,N_6009,N_5946);
nor U6195 (N_6195,N_6041,N_5993);
or U6196 (N_6196,N_5963,N_5999);
or U6197 (N_6197,N_5980,N_6050);
or U6198 (N_6198,N_5970,N_6078);
or U6199 (N_6199,N_6037,N_5977);
or U6200 (N_6200,N_6015,N_6028);
or U6201 (N_6201,N_5960,N_5949);
xnor U6202 (N_6202,N_6030,N_5956);
nor U6203 (N_6203,N_5940,N_6068);
or U6204 (N_6204,N_6041,N_5959);
and U6205 (N_6205,N_6061,N_5981);
and U6206 (N_6206,N_6058,N_6007);
and U6207 (N_6207,N_6024,N_5936);
or U6208 (N_6208,N_6046,N_6010);
and U6209 (N_6209,N_6009,N_5979);
and U6210 (N_6210,N_5947,N_6036);
nand U6211 (N_6211,N_5982,N_6049);
and U6212 (N_6212,N_5978,N_6001);
and U6213 (N_6213,N_6077,N_5997);
and U6214 (N_6214,N_5976,N_6073);
nand U6215 (N_6215,N_5966,N_6001);
nor U6216 (N_6216,N_6038,N_5969);
nand U6217 (N_6217,N_6036,N_6002);
nand U6218 (N_6218,N_6031,N_5934);
or U6219 (N_6219,N_5925,N_5969);
nor U6220 (N_6220,N_5970,N_6015);
or U6221 (N_6221,N_6049,N_5946);
nor U6222 (N_6222,N_5936,N_6045);
and U6223 (N_6223,N_5947,N_6014);
or U6224 (N_6224,N_6033,N_6046);
nor U6225 (N_6225,N_6070,N_5926);
or U6226 (N_6226,N_5955,N_5987);
or U6227 (N_6227,N_5931,N_5946);
nor U6228 (N_6228,N_6038,N_5952);
and U6229 (N_6229,N_6010,N_5988);
xor U6230 (N_6230,N_6028,N_5937);
nand U6231 (N_6231,N_5936,N_6041);
nand U6232 (N_6232,N_5941,N_6019);
nor U6233 (N_6233,N_5993,N_6000);
nor U6234 (N_6234,N_5992,N_5963);
nor U6235 (N_6235,N_6064,N_5943);
nor U6236 (N_6236,N_6069,N_6007);
nand U6237 (N_6237,N_5990,N_6021);
and U6238 (N_6238,N_6079,N_5975);
and U6239 (N_6239,N_6037,N_5936);
and U6240 (N_6240,N_6161,N_6095);
and U6241 (N_6241,N_6129,N_6156);
nor U6242 (N_6242,N_6206,N_6085);
nor U6243 (N_6243,N_6178,N_6201);
xnor U6244 (N_6244,N_6082,N_6234);
nand U6245 (N_6245,N_6099,N_6080);
or U6246 (N_6246,N_6148,N_6189);
nor U6247 (N_6247,N_6118,N_6170);
nor U6248 (N_6248,N_6153,N_6174);
xor U6249 (N_6249,N_6093,N_6228);
and U6250 (N_6250,N_6226,N_6157);
nand U6251 (N_6251,N_6175,N_6092);
nor U6252 (N_6252,N_6232,N_6114);
nand U6253 (N_6253,N_6151,N_6199);
nand U6254 (N_6254,N_6176,N_6150);
or U6255 (N_6255,N_6113,N_6185);
nand U6256 (N_6256,N_6165,N_6120);
nor U6257 (N_6257,N_6190,N_6211);
nand U6258 (N_6258,N_6193,N_6121);
xor U6259 (N_6259,N_6191,N_6217);
nor U6260 (N_6260,N_6126,N_6103);
and U6261 (N_6261,N_6203,N_6179);
or U6262 (N_6262,N_6171,N_6109);
or U6263 (N_6263,N_6134,N_6160);
or U6264 (N_6264,N_6221,N_6194);
or U6265 (N_6265,N_6119,N_6087);
nor U6266 (N_6266,N_6102,N_6101);
or U6267 (N_6267,N_6158,N_6224);
or U6268 (N_6268,N_6181,N_6186);
or U6269 (N_6269,N_6110,N_6133);
and U6270 (N_6270,N_6184,N_6143);
nor U6271 (N_6271,N_6112,N_6116);
or U6272 (N_6272,N_6083,N_6097);
nor U6273 (N_6273,N_6132,N_6212);
nor U6274 (N_6274,N_6086,N_6198);
nor U6275 (N_6275,N_6104,N_6122);
or U6276 (N_6276,N_6235,N_6200);
or U6277 (N_6277,N_6236,N_6166);
and U6278 (N_6278,N_6209,N_6213);
and U6279 (N_6279,N_6215,N_6229);
nand U6280 (N_6280,N_6131,N_6196);
and U6281 (N_6281,N_6128,N_6239);
or U6282 (N_6282,N_6096,N_6167);
or U6283 (N_6283,N_6202,N_6147);
xnor U6284 (N_6284,N_6145,N_6208);
nand U6285 (N_6285,N_6225,N_6177);
nor U6286 (N_6286,N_6125,N_6168);
nor U6287 (N_6287,N_6088,N_6220);
nor U6288 (N_6288,N_6140,N_6106);
and U6289 (N_6289,N_6136,N_6089);
nor U6290 (N_6290,N_6138,N_6091);
and U6291 (N_6291,N_6216,N_6169);
and U6292 (N_6292,N_6117,N_6182);
nor U6293 (N_6293,N_6149,N_6108);
and U6294 (N_6294,N_6172,N_6192);
and U6295 (N_6295,N_6135,N_6100);
or U6296 (N_6296,N_6231,N_6238);
and U6297 (N_6297,N_6115,N_6214);
nor U6298 (N_6298,N_6207,N_6219);
and U6299 (N_6299,N_6137,N_6084);
nand U6300 (N_6300,N_6195,N_6141);
nand U6301 (N_6301,N_6164,N_6223);
nand U6302 (N_6302,N_6188,N_6210);
nor U6303 (N_6303,N_6098,N_6163);
nor U6304 (N_6304,N_6197,N_6227);
nand U6305 (N_6305,N_6090,N_6218);
and U6306 (N_6306,N_6130,N_6230);
or U6307 (N_6307,N_6154,N_6142);
nor U6308 (N_6308,N_6205,N_6094);
or U6309 (N_6309,N_6105,N_6124);
nand U6310 (N_6310,N_6152,N_6233);
or U6311 (N_6311,N_6081,N_6107);
nand U6312 (N_6312,N_6127,N_6123);
nand U6313 (N_6313,N_6173,N_6155);
or U6314 (N_6314,N_6237,N_6180);
nor U6315 (N_6315,N_6111,N_6159);
or U6316 (N_6316,N_6139,N_6144);
or U6317 (N_6317,N_6204,N_6183);
nand U6318 (N_6318,N_6146,N_6162);
and U6319 (N_6319,N_6222,N_6187);
xor U6320 (N_6320,N_6167,N_6109);
xor U6321 (N_6321,N_6174,N_6206);
xnor U6322 (N_6322,N_6144,N_6166);
nand U6323 (N_6323,N_6081,N_6214);
nor U6324 (N_6324,N_6149,N_6228);
xor U6325 (N_6325,N_6104,N_6124);
xnor U6326 (N_6326,N_6222,N_6159);
nand U6327 (N_6327,N_6169,N_6202);
and U6328 (N_6328,N_6199,N_6095);
xor U6329 (N_6329,N_6171,N_6188);
nor U6330 (N_6330,N_6159,N_6211);
nand U6331 (N_6331,N_6104,N_6090);
xnor U6332 (N_6332,N_6235,N_6165);
nand U6333 (N_6333,N_6087,N_6239);
or U6334 (N_6334,N_6199,N_6089);
and U6335 (N_6335,N_6159,N_6189);
nand U6336 (N_6336,N_6214,N_6162);
or U6337 (N_6337,N_6093,N_6112);
or U6338 (N_6338,N_6107,N_6098);
and U6339 (N_6339,N_6130,N_6095);
nand U6340 (N_6340,N_6119,N_6110);
nor U6341 (N_6341,N_6207,N_6136);
xor U6342 (N_6342,N_6198,N_6182);
nor U6343 (N_6343,N_6157,N_6113);
nand U6344 (N_6344,N_6185,N_6131);
and U6345 (N_6345,N_6131,N_6187);
nor U6346 (N_6346,N_6163,N_6188);
and U6347 (N_6347,N_6232,N_6227);
nand U6348 (N_6348,N_6230,N_6181);
nand U6349 (N_6349,N_6207,N_6171);
nor U6350 (N_6350,N_6202,N_6121);
and U6351 (N_6351,N_6112,N_6232);
and U6352 (N_6352,N_6090,N_6143);
or U6353 (N_6353,N_6085,N_6163);
nand U6354 (N_6354,N_6082,N_6101);
nand U6355 (N_6355,N_6152,N_6185);
nor U6356 (N_6356,N_6162,N_6228);
or U6357 (N_6357,N_6110,N_6176);
nand U6358 (N_6358,N_6123,N_6212);
and U6359 (N_6359,N_6112,N_6157);
nor U6360 (N_6360,N_6151,N_6201);
or U6361 (N_6361,N_6177,N_6190);
and U6362 (N_6362,N_6108,N_6203);
xor U6363 (N_6363,N_6212,N_6230);
or U6364 (N_6364,N_6106,N_6157);
or U6365 (N_6365,N_6085,N_6148);
or U6366 (N_6366,N_6190,N_6201);
or U6367 (N_6367,N_6131,N_6200);
or U6368 (N_6368,N_6123,N_6185);
nor U6369 (N_6369,N_6203,N_6225);
or U6370 (N_6370,N_6141,N_6180);
nor U6371 (N_6371,N_6153,N_6088);
nor U6372 (N_6372,N_6113,N_6206);
nand U6373 (N_6373,N_6212,N_6112);
nand U6374 (N_6374,N_6210,N_6161);
or U6375 (N_6375,N_6224,N_6150);
nand U6376 (N_6376,N_6142,N_6159);
or U6377 (N_6377,N_6183,N_6100);
nand U6378 (N_6378,N_6187,N_6185);
xnor U6379 (N_6379,N_6116,N_6161);
or U6380 (N_6380,N_6136,N_6148);
or U6381 (N_6381,N_6177,N_6098);
nor U6382 (N_6382,N_6230,N_6087);
nor U6383 (N_6383,N_6227,N_6135);
or U6384 (N_6384,N_6228,N_6087);
or U6385 (N_6385,N_6156,N_6238);
and U6386 (N_6386,N_6108,N_6169);
nor U6387 (N_6387,N_6196,N_6134);
nor U6388 (N_6388,N_6117,N_6083);
nor U6389 (N_6389,N_6132,N_6098);
xnor U6390 (N_6390,N_6204,N_6170);
nand U6391 (N_6391,N_6134,N_6093);
nor U6392 (N_6392,N_6152,N_6145);
or U6393 (N_6393,N_6149,N_6196);
or U6394 (N_6394,N_6095,N_6239);
or U6395 (N_6395,N_6162,N_6156);
or U6396 (N_6396,N_6141,N_6167);
xor U6397 (N_6397,N_6180,N_6172);
nor U6398 (N_6398,N_6128,N_6197);
nand U6399 (N_6399,N_6161,N_6195);
or U6400 (N_6400,N_6307,N_6279);
or U6401 (N_6401,N_6385,N_6380);
nand U6402 (N_6402,N_6389,N_6269);
nand U6403 (N_6403,N_6369,N_6393);
nand U6404 (N_6404,N_6293,N_6252);
nand U6405 (N_6405,N_6364,N_6357);
and U6406 (N_6406,N_6317,N_6242);
nand U6407 (N_6407,N_6368,N_6273);
nand U6408 (N_6408,N_6339,N_6251);
xnor U6409 (N_6409,N_6311,N_6322);
nand U6410 (N_6410,N_6271,N_6315);
nand U6411 (N_6411,N_6354,N_6365);
nand U6412 (N_6412,N_6321,N_6394);
nor U6413 (N_6413,N_6360,N_6399);
nand U6414 (N_6414,N_6390,N_6275);
nand U6415 (N_6415,N_6340,N_6287);
and U6416 (N_6416,N_6254,N_6263);
and U6417 (N_6417,N_6362,N_6303);
or U6418 (N_6418,N_6375,N_6374);
and U6419 (N_6419,N_6383,N_6306);
and U6420 (N_6420,N_6260,N_6262);
nand U6421 (N_6421,N_6371,N_6336);
nand U6422 (N_6422,N_6316,N_6396);
nor U6423 (N_6423,N_6257,N_6358);
nor U6424 (N_6424,N_6276,N_6379);
and U6425 (N_6425,N_6265,N_6370);
or U6426 (N_6426,N_6304,N_6284);
xnor U6427 (N_6427,N_6272,N_6298);
and U6428 (N_6428,N_6319,N_6243);
nand U6429 (N_6429,N_6372,N_6289);
nand U6430 (N_6430,N_6245,N_6309);
nor U6431 (N_6431,N_6240,N_6349);
nor U6432 (N_6432,N_6255,N_6384);
nand U6433 (N_6433,N_6333,N_6346);
and U6434 (N_6434,N_6398,N_6288);
nand U6435 (N_6435,N_6348,N_6332);
or U6436 (N_6436,N_6391,N_6294);
and U6437 (N_6437,N_6320,N_6328);
or U6438 (N_6438,N_6325,N_6249);
nand U6439 (N_6439,N_6397,N_6338);
and U6440 (N_6440,N_6378,N_6292);
and U6441 (N_6441,N_6356,N_6241);
nand U6442 (N_6442,N_6367,N_6283);
nor U6443 (N_6443,N_6301,N_6376);
nor U6444 (N_6444,N_6297,N_6310);
or U6445 (N_6445,N_6314,N_6291);
or U6446 (N_6446,N_6313,N_6353);
nand U6447 (N_6447,N_6327,N_6247);
xnor U6448 (N_6448,N_6377,N_6344);
or U6449 (N_6449,N_6258,N_6246);
and U6450 (N_6450,N_6350,N_6388);
and U6451 (N_6451,N_6366,N_6382);
or U6452 (N_6452,N_6278,N_6352);
or U6453 (N_6453,N_6326,N_6266);
and U6454 (N_6454,N_6345,N_6244);
or U6455 (N_6455,N_6363,N_6373);
xnor U6456 (N_6456,N_6361,N_6342);
nand U6457 (N_6457,N_6253,N_6250);
xnor U6458 (N_6458,N_6386,N_6355);
nor U6459 (N_6459,N_6281,N_6343);
nor U6460 (N_6460,N_6286,N_6381);
or U6461 (N_6461,N_6299,N_6324);
and U6462 (N_6462,N_6308,N_6331);
nor U6463 (N_6463,N_6259,N_6274);
nor U6464 (N_6464,N_6341,N_6312);
nand U6465 (N_6465,N_6323,N_6335);
or U6466 (N_6466,N_6268,N_6295);
xnor U6467 (N_6467,N_6280,N_6334);
nand U6468 (N_6468,N_6347,N_6318);
or U6469 (N_6469,N_6392,N_6277);
nor U6470 (N_6470,N_6267,N_6305);
nor U6471 (N_6471,N_6330,N_6248);
and U6472 (N_6472,N_6256,N_6261);
or U6473 (N_6473,N_6296,N_6282);
or U6474 (N_6474,N_6302,N_6387);
xnor U6475 (N_6475,N_6270,N_6264);
or U6476 (N_6476,N_6300,N_6285);
or U6477 (N_6477,N_6395,N_6351);
nor U6478 (N_6478,N_6359,N_6290);
or U6479 (N_6479,N_6337,N_6329);
nand U6480 (N_6480,N_6374,N_6280);
nand U6481 (N_6481,N_6301,N_6246);
or U6482 (N_6482,N_6314,N_6346);
and U6483 (N_6483,N_6268,N_6276);
nor U6484 (N_6484,N_6378,N_6300);
xnor U6485 (N_6485,N_6378,N_6319);
or U6486 (N_6486,N_6358,N_6258);
or U6487 (N_6487,N_6317,N_6365);
nor U6488 (N_6488,N_6297,N_6270);
and U6489 (N_6489,N_6266,N_6323);
nor U6490 (N_6490,N_6324,N_6314);
and U6491 (N_6491,N_6328,N_6381);
or U6492 (N_6492,N_6328,N_6262);
xor U6493 (N_6493,N_6266,N_6331);
nand U6494 (N_6494,N_6317,N_6296);
and U6495 (N_6495,N_6264,N_6301);
and U6496 (N_6496,N_6269,N_6289);
or U6497 (N_6497,N_6249,N_6297);
or U6498 (N_6498,N_6391,N_6283);
nand U6499 (N_6499,N_6334,N_6308);
and U6500 (N_6500,N_6388,N_6301);
nor U6501 (N_6501,N_6256,N_6315);
xor U6502 (N_6502,N_6308,N_6345);
and U6503 (N_6503,N_6247,N_6245);
and U6504 (N_6504,N_6355,N_6332);
and U6505 (N_6505,N_6317,N_6383);
nand U6506 (N_6506,N_6335,N_6256);
and U6507 (N_6507,N_6383,N_6297);
and U6508 (N_6508,N_6372,N_6374);
and U6509 (N_6509,N_6360,N_6249);
and U6510 (N_6510,N_6369,N_6290);
or U6511 (N_6511,N_6392,N_6272);
nor U6512 (N_6512,N_6312,N_6331);
nor U6513 (N_6513,N_6255,N_6328);
and U6514 (N_6514,N_6388,N_6251);
nor U6515 (N_6515,N_6357,N_6243);
nor U6516 (N_6516,N_6309,N_6261);
and U6517 (N_6517,N_6269,N_6381);
nor U6518 (N_6518,N_6354,N_6242);
nor U6519 (N_6519,N_6269,N_6327);
nand U6520 (N_6520,N_6325,N_6257);
nand U6521 (N_6521,N_6384,N_6367);
nor U6522 (N_6522,N_6265,N_6293);
nand U6523 (N_6523,N_6362,N_6325);
nor U6524 (N_6524,N_6345,N_6291);
nor U6525 (N_6525,N_6298,N_6257);
nand U6526 (N_6526,N_6241,N_6335);
nor U6527 (N_6527,N_6320,N_6347);
nand U6528 (N_6528,N_6345,N_6377);
or U6529 (N_6529,N_6291,N_6398);
and U6530 (N_6530,N_6315,N_6308);
or U6531 (N_6531,N_6341,N_6285);
or U6532 (N_6532,N_6266,N_6243);
and U6533 (N_6533,N_6255,N_6342);
nand U6534 (N_6534,N_6390,N_6399);
nand U6535 (N_6535,N_6393,N_6323);
and U6536 (N_6536,N_6365,N_6279);
xor U6537 (N_6537,N_6384,N_6361);
xnor U6538 (N_6538,N_6368,N_6285);
nand U6539 (N_6539,N_6330,N_6308);
xor U6540 (N_6540,N_6273,N_6383);
nor U6541 (N_6541,N_6353,N_6329);
nor U6542 (N_6542,N_6370,N_6278);
nand U6543 (N_6543,N_6272,N_6398);
nand U6544 (N_6544,N_6279,N_6352);
nor U6545 (N_6545,N_6254,N_6353);
nand U6546 (N_6546,N_6277,N_6311);
nor U6547 (N_6547,N_6293,N_6344);
nand U6548 (N_6548,N_6313,N_6309);
nor U6549 (N_6549,N_6315,N_6373);
or U6550 (N_6550,N_6349,N_6254);
nand U6551 (N_6551,N_6333,N_6259);
nand U6552 (N_6552,N_6324,N_6266);
nor U6553 (N_6553,N_6324,N_6379);
nand U6554 (N_6554,N_6342,N_6370);
xor U6555 (N_6555,N_6268,N_6386);
nor U6556 (N_6556,N_6243,N_6363);
nand U6557 (N_6557,N_6326,N_6329);
nand U6558 (N_6558,N_6393,N_6334);
or U6559 (N_6559,N_6333,N_6242);
nand U6560 (N_6560,N_6488,N_6434);
and U6561 (N_6561,N_6523,N_6410);
or U6562 (N_6562,N_6490,N_6412);
and U6563 (N_6563,N_6502,N_6532);
or U6564 (N_6564,N_6526,N_6485);
nand U6565 (N_6565,N_6552,N_6493);
nand U6566 (N_6566,N_6546,N_6466);
nand U6567 (N_6567,N_6508,N_6478);
and U6568 (N_6568,N_6455,N_6510);
nor U6569 (N_6569,N_6432,N_6465);
and U6570 (N_6570,N_6496,N_6469);
nand U6571 (N_6571,N_6421,N_6501);
nor U6572 (N_6572,N_6472,N_6530);
and U6573 (N_6573,N_6457,N_6431);
and U6574 (N_6574,N_6505,N_6429);
nor U6575 (N_6575,N_6442,N_6427);
and U6576 (N_6576,N_6483,N_6436);
or U6577 (N_6577,N_6428,N_6408);
nor U6578 (N_6578,N_6452,N_6444);
and U6579 (N_6579,N_6521,N_6471);
and U6580 (N_6580,N_6467,N_6406);
nand U6581 (N_6581,N_6486,N_6517);
and U6582 (N_6582,N_6401,N_6522);
and U6583 (N_6583,N_6500,N_6464);
and U6584 (N_6584,N_6456,N_6495);
or U6585 (N_6585,N_6476,N_6514);
and U6586 (N_6586,N_6459,N_6559);
and U6587 (N_6587,N_6463,N_6468);
nor U6588 (N_6588,N_6554,N_6503);
and U6589 (N_6589,N_6544,N_6447);
and U6590 (N_6590,N_6541,N_6549);
and U6591 (N_6591,N_6533,N_6402);
nand U6592 (N_6592,N_6460,N_6422);
nand U6593 (N_6593,N_6536,N_6543);
xnor U6594 (N_6594,N_6542,N_6453);
and U6595 (N_6595,N_6420,N_6424);
nand U6596 (N_6596,N_6451,N_6515);
and U6597 (N_6597,N_6531,N_6507);
or U6598 (N_6598,N_6443,N_6509);
or U6599 (N_6599,N_6528,N_6538);
nor U6600 (N_6600,N_6445,N_6419);
xor U6601 (N_6601,N_6491,N_6545);
and U6602 (N_6602,N_6492,N_6518);
nor U6603 (N_6603,N_6477,N_6439);
or U6604 (N_6604,N_6470,N_6407);
and U6605 (N_6605,N_6506,N_6458);
xor U6606 (N_6606,N_6414,N_6512);
nand U6607 (N_6607,N_6409,N_6529);
nor U6608 (N_6608,N_6494,N_6413);
nor U6609 (N_6609,N_6440,N_6558);
or U6610 (N_6610,N_6519,N_6425);
and U6611 (N_6611,N_6513,N_6430);
nand U6612 (N_6612,N_6438,N_6446);
or U6613 (N_6613,N_6524,N_6527);
nor U6614 (N_6614,N_6418,N_6415);
and U6615 (N_6615,N_6534,N_6475);
nand U6616 (N_6616,N_6481,N_6433);
xor U6617 (N_6617,N_6520,N_6416);
nor U6618 (N_6618,N_6482,N_6474);
or U6619 (N_6619,N_6497,N_6487);
xor U6620 (N_6620,N_6499,N_6480);
xor U6621 (N_6621,N_6449,N_6535);
and U6622 (N_6622,N_6540,N_6556);
nor U6623 (N_6623,N_6479,N_6550);
and U6624 (N_6624,N_6539,N_6403);
nor U6625 (N_6625,N_6448,N_6400);
nand U6626 (N_6626,N_6551,N_6547);
nor U6627 (N_6627,N_6553,N_6504);
or U6628 (N_6628,N_6473,N_6484);
and U6629 (N_6629,N_6516,N_6461);
and U6630 (N_6630,N_6511,N_6435);
nand U6631 (N_6631,N_6537,N_6417);
or U6632 (N_6632,N_6557,N_6454);
and U6633 (N_6633,N_6548,N_6405);
nand U6634 (N_6634,N_6489,N_6423);
nand U6635 (N_6635,N_6462,N_6437);
or U6636 (N_6636,N_6411,N_6450);
and U6637 (N_6637,N_6426,N_6525);
or U6638 (N_6638,N_6404,N_6555);
and U6639 (N_6639,N_6441,N_6498);
nand U6640 (N_6640,N_6517,N_6507);
nor U6641 (N_6641,N_6504,N_6519);
nor U6642 (N_6642,N_6514,N_6518);
and U6643 (N_6643,N_6403,N_6485);
nor U6644 (N_6644,N_6496,N_6519);
nor U6645 (N_6645,N_6452,N_6531);
and U6646 (N_6646,N_6453,N_6495);
and U6647 (N_6647,N_6556,N_6515);
or U6648 (N_6648,N_6413,N_6441);
nand U6649 (N_6649,N_6531,N_6537);
nand U6650 (N_6650,N_6410,N_6485);
and U6651 (N_6651,N_6436,N_6555);
nor U6652 (N_6652,N_6447,N_6401);
or U6653 (N_6653,N_6415,N_6437);
and U6654 (N_6654,N_6434,N_6421);
and U6655 (N_6655,N_6508,N_6437);
nor U6656 (N_6656,N_6430,N_6471);
or U6657 (N_6657,N_6451,N_6530);
or U6658 (N_6658,N_6420,N_6461);
or U6659 (N_6659,N_6532,N_6443);
nand U6660 (N_6660,N_6489,N_6499);
xnor U6661 (N_6661,N_6424,N_6522);
and U6662 (N_6662,N_6411,N_6427);
or U6663 (N_6663,N_6459,N_6557);
nor U6664 (N_6664,N_6459,N_6462);
xor U6665 (N_6665,N_6482,N_6513);
or U6666 (N_6666,N_6559,N_6479);
or U6667 (N_6667,N_6435,N_6451);
xor U6668 (N_6668,N_6539,N_6507);
nor U6669 (N_6669,N_6443,N_6414);
nand U6670 (N_6670,N_6453,N_6489);
nand U6671 (N_6671,N_6444,N_6545);
and U6672 (N_6672,N_6483,N_6469);
or U6673 (N_6673,N_6434,N_6443);
and U6674 (N_6674,N_6442,N_6403);
or U6675 (N_6675,N_6504,N_6453);
and U6676 (N_6676,N_6482,N_6555);
or U6677 (N_6677,N_6518,N_6455);
nor U6678 (N_6678,N_6404,N_6546);
and U6679 (N_6679,N_6408,N_6462);
nand U6680 (N_6680,N_6437,N_6484);
nand U6681 (N_6681,N_6524,N_6491);
nand U6682 (N_6682,N_6530,N_6510);
or U6683 (N_6683,N_6464,N_6424);
or U6684 (N_6684,N_6543,N_6413);
nand U6685 (N_6685,N_6472,N_6546);
nor U6686 (N_6686,N_6461,N_6491);
and U6687 (N_6687,N_6491,N_6531);
or U6688 (N_6688,N_6489,N_6430);
nand U6689 (N_6689,N_6435,N_6457);
and U6690 (N_6690,N_6413,N_6435);
nand U6691 (N_6691,N_6556,N_6497);
nor U6692 (N_6692,N_6518,N_6522);
nor U6693 (N_6693,N_6498,N_6437);
or U6694 (N_6694,N_6536,N_6528);
nor U6695 (N_6695,N_6542,N_6504);
and U6696 (N_6696,N_6496,N_6554);
nand U6697 (N_6697,N_6466,N_6469);
nor U6698 (N_6698,N_6531,N_6412);
or U6699 (N_6699,N_6462,N_6478);
or U6700 (N_6700,N_6460,N_6409);
or U6701 (N_6701,N_6487,N_6486);
nand U6702 (N_6702,N_6556,N_6464);
nand U6703 (N_6703,N_6440,N_6537);
xnor U6704 (N_6704,N_6496,N_6438);
and U6705 (N_6705,N_6459,N_6423);
xor U6706 (N_6706,N_6510,N_6539);
or U6707 (N_6707,N_6408,N_6519);
nor U6708 (N_6708,N_6481,N_6478);
nand U6709 (N_6709,N_6493,N_6476);
nand U6710 (N_6710,N_6505,N_6476);
and U6711 (N_6711,N_6473,N_6432);
and U6712 (N_6712,N_6424,N_6502);
and U6713 (N_6713,N_6543,N_6445);
xnor U6714 (N_6714,N_6516,N_6449);
and U6715 (N_6715,N_6452,N_6424);
and U6716 (N_6716,N_6559,N_6406);
nor U6717 (N_6717,N_6433,N_6454);
nor U6718 (N_6718,N_6514,N_6510);
and U6719 (N_6719,N_6545,N_6436);
nand U6720 (N_6720,N_6681,N_6659);
nand U6721 (N_6721,N_6718,N_6593);
or U6722 (N_6722,N_6648,N_6636);
nand U6723 (N_6723,N_6598,N_6680);
and U6724 (N_6724,N_6575,N_6613);
nand U6725 (N_6725,N_6712,N_6705);
nor U6726 (N_6726,N_6661,N_6666);
nand U6727 (N_6727,N_6610,N_6562);
and U6728 (N_6728,N_6563,N_6629);
or U6729 (N_6729,N_6679,N_6677);
nand U6730 (N_6730,N_6709,N_6632);
or U6731 (N_6731,N_6620,N_6588);
xor U6732 (N_6732,N_6650,N_6630);
nor U6733 (N_6733,N_6689,N_6612);
xor U6734 (N_6734,N_6597,N_6635);
and U6735 (N_6735,N_6695,N_6615);
nor U6736 (N_6736,N_6654,N_6702);
xor U6737 (N_6737,N_6655,N_6639);
or U6738 (N_6738,N_6667,N_6578);
nand U6739 (N_6739,N_6652,N_6590);
or U6740 (N_6740,N_6619,N_6645);
nor U6741 (N_6741,N_6599,N_6676);
and U6742 (N_6742,N_6691,N_6678);
and U6743 (N_6743,N_6638,N_6570);
xnor U6744 (N_6744,N_6595,N_6577);
nor U6745 (N_6745,N_6653,N_6605);
nand U6746 (N_6746,N_6617,N_6640);
nand U6747 (N_6747,N_6690,N_6686);
or U6748 (N_6748,N_6576,N_6704);
nor U6749 (N_6749,N_6683,N_6673);
nor U6750 (N_6750,N_6626,N_6637);
nand U6751 (N_6751,N_6649,N_6671);
and U6752 (N_6752,N_6571,N_6658);
or U6753 (N_6753,N_6647,N_6646);
nor U6754 (N_6754,N_6574,N_6567);
xor U6755 (N_6755,N_6684,N_6708);
or U6756 (N_6756,N_6602,N_6565);
nor U6757 (N_6757,N_6642,N_6616);
and U6758 (N_6758,N_6687,N_6641);
nand U6759 (N_6759,N_6611,N_6699);
or U6760 (N_6760,N_6719,N_6663);
or U6761 (N_6761,N_6564,N_6608);
nand U6762 (N_6762,N_6627,N_6614);
and U6763 (N_6763,N_6716,N_6621);
nand U6764 (N_6764,N_6591,N_6566);
nor U6765 (N_6765,N_6698,N_6606);
or U6766 (N_6766,N_6672,N_6584);
nor U6767 (N_6767,N_6625,N_6688);
or U6768 (N_6768,N_6706,N_6657);
or U6769 (N_6769,N_6622,N_6607);
xor U6770 (N_6770,N_6662,N_6582);
nor U6771 (N_6771,N_6568,N_6651);
nor U6772 (N_6772,N_6669,N_6569);
or U6773 (N_6773,N_6618,N_6660);
and U6774 (N_6774,N_6665,N_6596);
and U6775 (N_6775,N_6715,N_6583);
nand U6776 (N_6776,N_6707,N_6628);
or U6777 (N_6777,N_6634,N_6697);
xor U6778 (N_6778,N_6609,N_6717);
and U6779 (N_6779,N_6644,N_6585);
or U6780 (N_6780,N_6694,N_6631);
nor U6781 (N_6781,N_6580,N_6604);
nor U6782 (N_6782,N_6589,N_6703);
nor U6783 (N_6783,N_6560,N_6624);
xnor U6784 (N_6784,N_6601,N_6682);
and U6785 (N_6785,N_6572,N_6594);
nand U6786 (N_6786,N_6623,N_6581);
and U6787 (N_6787,N_6693,N_6579);
nor U6788 (N_6788,N_6696,N_6633);
nand U6789 (N_6789,N_6713,N_6675);
or U6790 (N_6790,N_6674,N_6714);
nor U6791 (N_6791,N_6586,N_6573);
nand U6792 (N_6792,N_6656,N_6710);
and U6793 (N_6793,N_6700,N_6685);
and U6794 (N_6794,N_6701,N_6643);
nand U6795 (N_6795,N_6664,N_6692);
and U6796 (N_6796,N_6561,N_6603);
or U6797 (N_6797,N_6600,N_6711);
xnor U6798 (N_6798,N_6592,N_6587);
xnor U6799 (N_6799,N_6670,N_6668);
nor U6800 (N_6800,N_6705,N_6701);
xor U6801 (N_6801,N_6575,N_6712);
nand U6802 (N_6802,N_6612,N_6598);
and U6803 (N_6803,N_6645,N_6697);
xnor U6804 (N_6804,N_6617,N_6658);
nand U6805 (N_6805,N_6680,N_6663);
and U6806 (N_6806,N_6562,N_6694);
nand U6807 (N_6807,N_6606,N_6646);
or U6808 (N_6808,N_6581,N_6589);
nand U6809 (N_6809,N_6617,N_6668);
and U6810 (N_6810,N_6648,N_6693);
or U6811 (N_6811,N_6601,N_6584);
and U6812 (N_6812,N_6603,N_6666);
nand U6813 (N_6813,N_6592,N_6639);
nand U6814 (N_6814,N_6689,N_6634);
or U6815 (N_6815,N_6630,N_6706);
or U6816 (N_6816,N_6707,N_6596);
and U6817 (N_6817,N_6574,N_6610);
or U6818 (N_6818,N_6711,N_6605);
nand U6819 (N_6819,N_6616,N_6574);
and U6820 (N_6820,N_6570,N_6618);
or U6821 (N_6821,N_6666,N_6679);
nor U6822 (N_6822,N_6583,N_6567);
nand U6823 (N_6823,N_6658,N_6561);
and U6824 (N_6824,N_6571,N_6703);
or U6825 (N_6825,N_6587,N_6605);
xor U6826 (N_6826,N_6607,N_6568);
and U6827 (N_6827,N_6691,N_6665);
and U6828 (N_6828,N_6656,N_6599);
or U6829 (N_6829,N_6611,N_6616);
or U6830 (N_6830,N_6631,N_6675);
and U6831 (N_6831,N_6636,N_6680);
and U6832 (N_6832,N_6650,N_6648);
and U6833 (N_6833,N_6685,N_6647);
nand U6834 (N_6834,N_6613,N_6582);
or U6835 (N_6835,N_6566,N_6683);
nor U6836 (N_6836,N_6696,N_6606);
nor U6837 (N_6837,N_6712,N_6674);
xnor U6838 (N_6838,N_6620,N_6695);
nand U6839 (N_6839,N_6595,N_6631);
nand U6840 (N_6840,N_6601,N_6688);
nand U6841 (N_6841,N_6577,N_6571);
xnor U6842 (N_6842,N_6623,N_6656);
or U6843 (N_6843,N_6569,N_6714);
nand U6844 (N_6844,N_6668,N_6561);
nor U6845 (N_6845,N_6680,N_6571);
and U6846 (N_6846,N_6638,N_6691);
or U6847 (N_6847,N_6668,N_6567);
or U6848 (N_6848,N_6583,N_6582);
nor U6849 (N_6849,N_6592,N_6694);
nor U6850 (N_6850,N_6618,N_6674);
xnor U6851 (N_6851,N_6616,N_6613);
and U6852 (N_6852,N_6631,N_6573);
nand U6853 (N_6853,N_6602,N_6605);
nand U6854 (N_6854,N_6649,N_6588);
or U6855 (N_6855,N_6671,N_6565);
xor U6856 (N_6856,N_6622,N_6658);
or U6857 (N_6857,N_6578,N_6717);
or U6858 (N_6858,N_6676,N_6574);
or U6859 (N_6859,N_6632,N_6573);
nor U6860 (N_6860,N_6650,N_6618);
and U6861 (N_6861,N_6695,N_6674);
nand U6862 (N_6862,N_6634,N_6645);
xor U6863 (N_6863,N_6704,N_6604);
xnor U6864 (N_6864,N_6661,N_6614);
nor U6865 (N_6865,N_6645,N_6696);
or U6866 (N_6866,N_6565,N_6679);
nor U6867 (N_6867,N_6718,N_6717);
nor U6868 (N_6868,N_6704,N_6618);
nand U6869 (N_6869,N_6666,N_6574);
or U6870 (N_6870,N_6562,N_6631);
nand U6871 (N_6871,N_6649,N_6712);
and U6872 (N_6872,N_6688,N_6562);
or U6873 (N_6873,N_6591,N_6702);
nand U6874 (N_6874,N_6702,N_6575);
nand U6875 (N_6875,N_6681,N_6596);
and U6876 (N_6876,N_6570,N_6660);
nand U6877 (N_6877,N_6571,N_6620);
nor U6878 (N_6878,N_6606,N_6595);
nor U6879 (N_6879,N_6636,N_6647);
nand U6880 (N_6880,N_6752,N_6878);
xor U6881 (N_6881,N_6828,N_6823);
nor U6882 (N_6882,N_6818,N_6786);
nand U6883 (N_6883,N_6835,N_6820);
or U6884 (N_6884,N_6766,N_6792);
nor U6885 (N_6885,N_6790,N_6727);
or U6886 (N_6886,N_6769,N_6875);
or U6887 (N_6887,N_6807,N_6805);
nor U6888 (N_6888,N_6771,N_6733);
and U6889 (N_6889,N_6852,N_6840);
or U6890 (N_6890,N_6830,N_6864);
and U6891 (N_6891,N_6778,N_6811);
and U6892 (N_6892,N_6734,N_6851);
nand U6893 (N_6893,N_6874,N_6738);
or U6894 (N_6894,N_6785,N_6845);
xor U6895 (N_6895,N_6755,N_6866);
or U6896 (N_6896,N_6739,N_6741);
nand U6897 (N_6897,N_6789,N_6726);
and U6898 (N_6898,N_6833,N_6831);
xnor U6899 (N_6899,N_6819,N_6736);
nand U6900 (N_6900,N_6856,N_6810);
nor U6901 (N_6901,N_6841,N_6781);
nand U6902 (N_6902,N_6834,N_6776);
nor U6903 (N_6903,N_6723,N_6857);
nor U6904 (N_6904,N_6751,N_6832);
nand U6905 (N_6905,N_6774,N_6744);
nand U6906 (N_6906,N_6872,N_6843);
nand U6907 (N_6907,N_6737,N_6855);
and U6908 (N_6908,N_6853,N_6796);
nand U6909 (N_6909,N_6750,N_6743);
or U6910 (N_6910,N_6762,N_6803);
xnor U6911 (N_6911,N_6787,N_6829);
nand U6912 (N_6912,N_6749,N_6768);
nor U6913 (N_6913,N_6746,N_6816);
nand U6914 (N_6914,N_6784,N_6858);
nand U6915 (N_6915,N_6850,N_6782);
nor U6916 (N_6916,N_6799,N_6868);
and U6917 (N_6917,N_6876,N_6838);
xor U6918 (N_6918,N_6865,N_6842);
nand U6919 (N_6919,N_6724,N_6821);
or U6920 (N_6920,N_6812,N_6775);
nand U6921 (N_6921,N_6773,N_6814);
nand U6922 (N_6922,N_6808,N_6800);
and U6923 (N_6923,N_6753,N_6780);
nor U6924 (N_6924,N_6765,N_6757);
or U6925 (N_6925,N_6815,N_6767);
and U6926 (N_6926,N_6806,N_6793);
xor U6927 (N_6927,N_6754,N_6794);
nor U6928 (N_6928,N_6859,N_6791);
and U6929 (N_6929,N_6863,N_6760);
or U6930 (N_6930,N_6809,N_6735);
nor U6931 (N_6931,N_6827,N_6759);
and U6932 (N_6932,N_6721,N_6836);
nand U6933 (N_6933,N_6720,N_6817);
xor U6934 (N_6934,N_6822,N_6795);
nand U6935 (N_6935,N_6860,N_6861);
and U6936 (N_6936,N_6747,N_6871);
or U6937 (N_6937,N_6730,N_6846);
and U6938 (N_6938,N_6729,N_6725);
nor U6939 (N_6939,N_6844,N_6763);
and U6940 (N_6940,N_6877,N_6745);
and U6941 (N_6941,N_6772,N_6813);
or U6942 (N_6942,N_6764,N_6728);
and U6943 (N_6943,N_6783,N_6837);
nand U6944 (N_6944,N_6797,N_6826);
or U6945 (N_6945,N_6839,N_6869);
nor U6946 (N_6946,N_6758,N_6854);
and U6947 (N_6947,N_6798,N_6722);
nand U6948 (N_6948,N_6740,N_6731);
nand U6949 (N_6949,N_6770,N_6756);
and U6950 (N_6950,N_6848,N_6742);
or U6951 (N_6951,N_6870,N_6825);
nand U6952 (N_6952,N_6801,N_6849);
nand U6953 (N_6953,N_6761,N_6862);
or U6954 (N_6954,N_6779,N_6732);
xnor U6955 (N_6955,N_6788,N_6802);
xnor U6956 (N_6956,N_6873,N_6748);
nor U6957 (N_6957,N_6824,N_6867);
nor U6958 (N_6958,N_6847,N_6879);
nor U6959 (N_6959,N_6804,N_6777);
and U6960 (N_6960,N_6837,N_6798);
and U6961 (N_6961,N_6786,N_6801);
xnor U6962 (N_6962,N_6869,N_6757);
or U6963 (N_6963,N_6773,N_6821);
nand U6964 (N_6964,N_6748,N_6802);
xor U6965 (N_6965,N_6727,N_6729);
or U6966 (N_6966,N_6847,N_6743);
nor U6967 (N_6967,N_6873,N_6855);
xnor U6968 (N_6968,N_6813,N_6799);
or U6969 (N_6969,N_6819,N_6757);
and U6970 (N_6970,N_6771,N_6762);
nor U6971 (N_6971,N_6807,N_6808);
or U6972 (N_6972,N_6832,N_6765);
and U6973 (N_6973,N_6807,N_6801);
nand U6974 (N_6974,N_6849,N_6752);
and U6975 (N_6975,N_6776,N_6859);
and U6976 (N_6976,N_6805,N_6873);
and U6977 (N_6977,N_6826,N_6862);
and U6978 (N_6978,N_6790,N_6777);
nor U6979 (N_6979,N_6797,N_6805);
nor U6980 (N_6980,N_6780,N_6842);
and U6981 (N_6981,N_6750,N_6765);
and U6982 (N_6982,N_6872,N_6756);
nor U6983 (N_6983,N_6752,N_6852);
and U6984 (N_6984,N_6746,N_6817);
nand U6985 (N_6985,N_6879,N_6860);
nand U6986 (N_6986,N_6801,N_6816);
nand U6987 (N_6987,N_6732,N_6877);
or U6988 (N_6988,N_6769,N_6867);
xnor U6989 (N_6989,N_6871,N_6842);
or U6990 (N_6990,N_6773,N_6823);
or U6991 (N_6991,N_6744,N_6762);
or U6992 (N_6992,N_6878,N_6836);
nor U6993 (N_6993,N_6859,N_6799);
and U6994 (N_6994,N_6772,N_6865);
and U6995 (N_6995,N_6734,N_6741);
nor U6996 (N_6996,N_6802,N_6781);
and U6997 (N_6997,N_6794,N_6817);
nand U6998 (N_6998,N_6787,N_6756);
or U6999 (N_6999,N_6874,N_6803);
or U7000 (N_7000,N_6727,N_6730);
nand U7001 (N_7001,N_6857,N_6872);
or U7002 (N_7002,N_6732,N_6820);
nor U7003 (N_7003,N_6778,N_6762);
or U7004 (N_7004,N_6860,N_6859);
nand U7005 (N_7005,N_6792,N_6878);
nor U7006 (N_7006,N_6841,N_6757);
xor U7007 (N_7007,N_6733,N_6829);
nor U7008 (N_7008,N_6790,N_6785);
xor U7009 (N_7009,N_6768,N_6728);
xnor U7010 (N_7010,N_6842,N_6820);
xor U7011 (N_7011,N_6844,N_6849);
and U7012 (N_7012,N_6833,N_6744);
nand U7013 (N_7013,N_6831,N_6870);
nand U7014 (N_7014,N_6744,N_6830);
xnor U7015 (N_7015,N_6736,N_6858);
and U7016 (N_7016,N_6841,N_6756);
and U7017 (N_7017,N_6732,N_6847);
xnor U7018 (N_7018,N_6799,N_6754);
nand U7019 (N_7019,N_6783,N_6829);
nand U7020 (N_7020,N_6845,N_6871);
nand U7021 (N_7021,N_6809,N_6762);
nand U7022 (N_7022,N_6830,N_6811);
or U7023 (N_7023,N_6826,N_6842);
or U7024 (N_7024,N_6739,N_6757);
nand U7025 (N_7025,N_6820,N_6749);
nor U7026 (N_7026,N_6878,N_6858);
or U7027 (N_7027,N_6842,N_6856);
nor U7028 (N_7028,N_6822,N_6776);
or U7029 (N_7029,N_6818,N_6870);
or U7030 (N_7030,N_6807,N_6854);
nand U7031 (N_7031,N_6809,N_6851);
or U7032 (N_7032,N_6749,N_6791);
nor U7033 (N_7033,N_6831,N_6721);
xor U7034 (N_7034,N_6723,N_6732);
nand U7035 (N_7035,N_6873,N_6794);
and U7036 (N_7036,N_6757,N_6838);
nor U7037 (N_7037,N_6722,N_6793);
nor U7038 (N_7038,N_6770,N_6824);
or U7039 (N_7039,N_6789,N_6803);
xnor U7040 (N_7040,N_6935,N_6986);
and U7041 (N_7041,N_7038,N_6950);
and U7042 (N_7042,N_6978,N_7036);
nand U7043 (N_7043,N_6891,N_6906);
or U7044 (N_7044,N_6994,N_7016);
nor U7045 (N_7045,N_6932,N_6968);
nand U7046 (N_7046,N_7002,N_6989);
or U7047 (N_7047,N_7031,N_6916);
nor U7048 (N_7048,N_6911,N_6969);
and U7049 (N_7049,N_7034,N_7015);
and U7050 (N_7050,N_7005,N_6909);
nor U7051 (N_7051,N_6883,N_6940);
or U7052 (N_7052,N_6889,N_6885);
nor U7053 (N_7053,N_7032,N_6997);
nand U7054 (N_7054,N_6992,N_6975);
nand U7055 (N_7055,N_6957,N_6990);
nand U7056 (N_7056,N_6952,N_6896);
or U7057 (N_7057,N_6973,N_6972);
and U7058 (N_7058,N_6980,N_6902);
and U7059 (N_7059,N_6925,N_7010);
xnor U7060 (N_7060,N_6928,N_6919);
xor U7061 (N_7061,N_6893,N_6901);
xnor U7062 (N_7062,N_7025,N_7029);
nand U7063 (N_7063,N_6944,N_6884);
and U7064 (N_7064,N_6941,N_6961);
nand U7065 (N_7065,N_6931,N_7007);
nor U7066 (N_7066,N_7012,N_6965);
xnor U7067 (N_7067,N_7008,N_6886);
and U7068 (N_7068,N_6963,N_6953);
or U7069 (N_7069,N_6881,N_6967);
nor U7070 (N_7070,N_6946,N_6996);
nor U7071 (N_7071,N_6933,N_6993);
and U7072 (N_7072,N_6959,N_6976);
or U7073 (N_7073,N_6949,N_6921);
and U7074 (N_7074,N_6903,N_6951);
and U7075 (N_7075,N_6970,N_6898);
nand U7076 (N_7076,N_6929,N_7024);
or U7077 (N_7077,N_6914,N_6981);
and U7078 (N_7078,N_6904,N_6908);
and U7079 (N_7079,N_7022,N_7023);
nor U7080 (N_7080,N_7033,N_6888);
nor U7081 (N_7081,N_6995,N_6882);
and U7082 (N_7082,N_7026,N_7009);
and U7083 (N_7083,N_6987,N_6890);
or U7084 (N_7084,N_7021,N_6918);
nor U7085 (N_7085,N_6988,N_7030);
nand U7086 (N_7086,N_6985,N_6956);
and U7087 (N_7087,N_6936,N_6982);
or U7088 (N_7088,N_6892,N_7028);
nor U7089 (N_7089,N_6894,N_6905);
and U7090 (N_7090,N_7003,N_6924);
nand U7091 (N_7091,N_6934,N_6979);
and U7092 (N_7092,N_6912,N_6942);
and U7093 (N_7093,N_7014,N_7001);
or U7094 (N_7094,N_7006,N_6964);
nand U7095 (N_7095,N_7039,N_6998);
nor U7096 (N_7096,N_6983,N_6880);
xor U7097 (N_7097,N_6922,N_7037);
or U7098 (N_7098,N_6945,N_6947);
xor U7099 (N_7099,N_6920,N_6960);
nor U7100 (N_7100,N_6939,N_6999);
and U7101 (N_7101,N_6971,N_6917);
or U7102 (N_7102,N_6962,N_7019);
xnor U7103 (N_7103,N_6907,N_7020);
and U7104 (N_7104,N_7000,N_6955);
nand U7105 (N_7105,N_6966,N_7011);
nor U7106 (N_7106,N_6930,N_6943);
nor U7107 (N_7107,N_6913,N_6954);
nand U7108 (N_7108,N_7004,N_7013);
and U7109 (N_7109,N_6958,N_6899);
nand U7110 (N_7110,N_6977,N_7035);
or U7111 (N_7111,N_6938,N_6887);
nand U7112 (N_7112,N_6900,N_6927);
and U7113 (N_7113,N_7017,N_6915);
nand U7114 (N_7114,N_6948,N_7027);
nor U7115 (N_7115,N_6910,N_6895);
nor U7116 (N_7116,N_6923,N_6897);
and U7117 (N_7117,N_6991,N_6937);
xor U7118 (N_7118,N_6926,N_7018);
nor U7119 (N_7119,N_6974,N_6984);
nand U7120 (N_7120,N_7013,N_6901);
or U7121 (N_7121,N_6936,N_6976);
nand U7122 (N_7122,N_6966,N_6905);
and U7123 (N_7123,N_7037,N_7029);
nor U7124 (N_7124,N_6954,N_7030);
and U7125 (N_7125,N_6963,N_6914);
or U7126 (N_7126,N_6974,N_6993);
nand U7127 (N_7127,N_6901,N_6959);
nor U7128 (N_7128,N_6895,N_6969);
nor U7129 (N_7129,N_6979,N_7019);
nand U7130 (N_7130,N_6982,N_6959);
and U7131 (N_7131,N_6899,N_6938);
or U7132 (N_7132,N_6972,N_7024);
and U7133 (N_7133,N_6930,N_6888);
and U7134 (N_7134,N_6986,N_6938);
and U7135 (N_7135,N_6933,N_6919);
and U7136 (N_7136,N_6888,N_6944);
or U7137 (N_7137,N_6980,N_6969);
nand U7138 (N_7138,N_6909,N_6955);
xor U7139 (N_7139,N_6926,N_6978);
xnor U7140 (N_7140,N_7037,N_6960);
or U7141 (N_7141,N_6896,N_7003);
nand U7142 (N_7142,N_7032,N_6930);
and U7143 (N_7143,N_6951,N_6914);
nand U7144 (N_7144,N_7023,N_7026);
and U7145 (N_7145,N_6885,N_6959);
and U7146 (N_7146,N_6891,N_7030);
and U7147 (N_7147,N_6973,N_7025);
and U7148 (N_7148,N_6940,N_6953);
nand U7149 (N_7149,N_6911,N_6995);
or U7150 (N_7150,N_6997,N_6907);
and U7151 (N_7151,N_6999,N_6931);
and U7152 (N_7152,N_7007,N_6928);
nor U7153 (N_7153,N_6892,N_6908);
or U7154 (N_7154,N_7003,N_6951);
xor U7155 (N_7155,N_7005,N_7019);
xnor U7156 (N_7156,N_6955,N_6991);
nor U7157 (N_7157,N_6984,N_6955);
nor U7158 (N_7158,N_7020,N_6895);
or U7159 (N_7159,N_6987,N_6910);
nand U7160 (N_7160,N_7009,N_7014);
xor U7161 (N_7161,N_7012,N_7017);
and U7162 (N_7162,N_6894,N_6940);
and U7163 (N_7163,N_6897,N_6911);
nor U7164 (N_7164,N_7002,N_6972);
and U7165 (N_7165,N_6957,N_7008);
and U7166 (N_7166,N_7000,N_7013);
nand U7167 (N_7167,N_6880,N_7018);
and U7168 (N_7168,N_6957,N_6934);
nor U7169 (N_7169,N_6982,N_7037);
xnor U7170 (N_7170,N_6883,N_6909);
nand U7171 (N_7171,N_6957,N_6896);
nand U7172 (N_7172,N_6990,N_6994);
nor U7173 (N_7173,N_7016,N_6999);
xor U7174 (N_7174,N_6884,N_6984);
xor U7175 (N_7175,N_6995,N_6983);
nor U7176 (N_7176,N_6931,N_6884);
nand U7177 (N_7177,N_7001,N_6916);
and U7178 (N_7178,N_6943,N_7026);
or U7179 (N_7179,N_6929,N_6881);
and U7180 (N_7180,N_6973,N_7015);
nand U7181 (N_7181,N_7018,N_6922);
xnor U7182 (N_7182,N_7008,N_6979);
xor U7183 (N_7183,N_6946,N_6966);
nand U7184 (N_7184,N_6888,N_6987);
nand U7185 (N_7185,N_6956,N_6998);
nor U7186 (N_7186,N_6902,N_6946);
nand U7187 (N_7187,N_6986,N_7037);
nor U7188 (N_7188,N_6916,N_6991);
or U7189 (N_7189,N_6920,N_6988);
and U7190 (N_7190,N_7006,N_7027);
and U7191 (N_7191,N_7008,N_6917);
xor U7192 (N_7192,N_6898,N_7027);
or U7193 (N_7193,N_6923,N_6984);
nor U7194 (N_7194,N_7009,N_6972);
nor U7195 (N_7195,N_6888,N_6968);
or U7196 (N_7196,N_6880,N_7039);
nand U7197 (N_7197,N_7000,N_6897);
xor U7198 (N_7198,N_7020,N_6977);
or U7199 (N_7199,N_7025,N_6912);
or U7200 (N_7200,N_7194,N_7042);
nand U7201 (N_7201,N_7153,N_7142);
nor U7202 (N_7202,N_7047,N_7159);
nand U7203 (N_7203,N_7045,N_7197);
nand U7204 (N_7204,N_7078,N_7163);
nor U7205 (N_7205,N_7129,N_7144);
xor U7206 (N_7206,N_7141,N_7137);
or U7207 (N_7207,N_7139,N_7057);
nand U7208 (N_7208,N_7120,N_7059);
nand U7209 (N_7209,N_7130,N_7048);
nor U7210 (N_7210,N_7068,N_7083);
nor U7211 (N_7211,N_7052,N_7101);
nand U7212 (N_7212,N_7192,N_7094);
or U7213 (N_7213,N_7066,N_7169);
nor U7214 (N_7214,N_7134,N_7140);
and U7215 (N_7215,N_7041,N_7065);
or U7216 (N_7216,N_7196,N_7151);
nor U7217 (N_7217,N_7149,N_7096);
nand U7218 (N_7218,N_7189,N_7084);
xnor U7219 (N_7219,N_7122,N_7186);
nor U7220 (N_7220,N_7127,N_7062);
nand U7221 (N_7221,N_7103,N_7118);
nor U7222 (N_7222,N_7053,N_7050);
nor U7223 (N_7223,N_7131,N_7184);
nor U7224 (N_7224,N_7092,N_7155);
nand U7225 (N_7225,N_7116,N_7162);
or U7226 (N_7226,N_7133,N_7074);
or U7227 (N_7227,N_7176,N_7109);
or U7228 (N_7228,N_7198,N_7181);
nor U7229 (N_7229,N_7051,N_7076);
nand U7230 (N_7230,N_7106,N_7075);
xnor U7231 (N_7231,N_7123,N_7079);
and U7232 (N_7232,N_7040,N_7173);
nand U7233 (N_7233,N_7195,N_7182);
xor U7234 (N_7234,N_7072,N_7070);
nand U7235 (N_7235,N_7188,N_7090);
nor U7236 (N_7236,N_7143,N_7115);
and U7237 (N_7237,N_7113,N_7199);
and U7238 (N_7238,N_7124,N_7126);
and U7239 (N_7239,N_7148,N_7179);
nand U7240 (N_7240,N_7105,N_7069);
nor U7241 (N_7241,N_7104,N_7077);
or U7242 (N_7242,N_7147,N_7168);
nand U7243 (N_7243,N_7170,N_7061);
xor U7244 (N_7244,N_7190,N_7046);
and U7245 (N_7245,N_7099,N_7136);
or U7246 (N_7246,N_7100,N_7154);
and U7247 (N_7247,N_7098,N_7132);
nor U7248 (N_7248,N_7088,N_7044);
and U7249 (N_7249,N_7058,N_7093);
and U7250 (N_7250,N_7102,N_7097);
or U7251 (N_7251,N_7114,N_7187);
nand U7252 (N_7252,N_7089,N_7135);
and U7253 (N_7253,N_7117,N_7121);
xnor U7254 (N_7254,N_7178,N_7081);
and U7255 (N_7255,N_7056,N_7160);
nand U7256 (N_7256,N_7167,N_7180);
nor U7257 (N_7257,N_7174,N_7165);
nand U7258 (N_7258,N_7064,N_7158);
and U7259 (N_7259,N_7156,N_7049);
or U7260 (N_7260,N_7128,N_7157);
or U7261 (N_7261,N_7110,N_7111);
nand U7262 (N_7262,N_7060,N_7043);
and U7263 (N_7263,N_7175,N_7193);
or U7264 (N_7264,N_7108,N_7185);
and U7265 (N_7265,N_7171,N_7067);
nor U7266 (N_7266,N_7095,N_7055);
nor U7267 (N_7267,N_7054,N_7150);
or U7268 (N_7268,N_7172,N_7166);
xor U7269 (N_7269,N_7125,N_7145);
xor U7270 (N_7270,N_7086,N_7063);
and U7271 (N_7271,N_7112,N_7146);
nand U7272 (N_7272,N_7191,N_7177);
nand U7273 (N_7273,N_7152,N_7087);
and U7274 (N_7274,N_7164,N_7073);
nand U7275 (N_7275,N_7085,N_7082);
nor U7276 (N_7276,N_7119,N_7107);
nor U7277 (N_7277,N_7091,N_7080);
nand U7278 (N_7278,N_7161,N_7138);
and U7279 (N_7279,N_7071,N_7183);
and U7280 (N_7280,N_7153,N_7075);
nand U7281 (N_7281,N_7075,N_7110);
and U7282 (N_7282,N_7199,N_7076);
nand U7283 (N_7283,N_7163,N_7162);
nor U7284 (N_7284,N_7191,N_7069);
and U7285 (N_7285,N_7183,N_7093);
or U7286 (N_7286,N_7078,N_7041);
xnor U7287 (N_7287,N_7137,N_7064);
nor U7288 (N_7288,N_7052,N_7113);
nand U7289 (N_7289,N_7077,N_7144);
nand U7290 (N_7290,N_7143,N_7086);
nand U7291 (N_7291,N_7079,N_7101);
and U7292 (N_7292,N_7129,N_7065);
or U7293 (N_7293,N_7065,N_7043);
nand U7294 (N_7294,N_7091,N_7119);
nand U7295 (N_7295,N_7144,N_7186);
or U7296 (N_7296,N_7162,N_7073);
nand U7297 (N_7297,N_7155,N_7127);
xnor U7298 (N_7298,N_7126,N_7059);
nor U7299 (N_7299,N_7049,N_7122);
nand U7300 (N_7300,N_7096,N_7180);
or U7301 (N_7301,N_7134,N_7089);
nand U7302 (N_7302,N_7077,N_7166);
xnor U7303 (N_7303,N_7161,N_7076);
nand U7304 (N_7304,N_7112,N_7192);
and U7305 (N_7305,N_7045,N_7151);
or U7306 (N_7306,N_7093,N_7051);
xor U7307 (N_7307,N_7178,N_7118);
nor U7308 (N_7308,N_7186,N_7194);
or U7309 (N_7309,N_7177,N_7069);
nand U7310 (N_7310,N_7091,N_7071);
nor U7311 (N_7311,N_7197,N_7041);
nand U7312 (N_7312,N_7146,N_7090);
nor U7313 (N_7313,N_7147,N_7125);
nand U7314 (N_7314,N_7145,N_7077);
or U7315 (N_7315,N_7174,N_7160);
nand U7316 (N_7316,N_7049,N_7085);
nand U7317 (N_7317,N_7046,N_7072);
and U7318 (N_7318,N_7184,N_7146);
and U7319 (N_7319,N_7136,N_7165);
and U7320 (N_7320,N_7126,N_7190);
or U7321 (N_7321,N_7164,N_7040);
nor U7322 (N_7322,N_7134,N_7184);
nand U7323 (N_7323,N_7090,N_7087);
and U7324 (N_7324,N_7055,N_7155);
xnor U7325 (N_7325,N_7120,N_7043);
or U7326 (N_7326,N_7089,N_7081);
or U7327 (N_7327,N_7052,N_7103);
and U7328 (N_7328,N_7047,N_7117);
nor U7329 (N_7329,N_7186,N_7141);
nand U7330 (N_7330,N_7188,N_7133);
nand U7331 (N_7331,N_7137,N_7106);
nor U7332 (N_7332,N_7194,N_7151);
nand U7333 (N_7333,N_7135,N_7163);
and U7334 (N_7334,N_7099,N_7057);
and U7335 (N_7335,N_7183,N_7077);
or U7336 (N_7336,N_7093,N_7135);
or U7337 (N_7337,N_7157,N_7109);
or U7338 (N_7338,N_7152,N_7136);
or U7339 (N_7339,N_7170,N_7185);
and U7340 (N_7340,N_7143,N_7052);
nor U7341 (N_7341,N_7191,N_7050);
nor U7342 (N_7342,N_7041,N_7129);
and U7343 (N_7343,N_7157,N_7139);
nand U7344 (N_7344,N_7175,N_7174);
nor U7345 (N_7345,N_7070,N_7159);
and U7346 (N_7346,N_7162,N_7047);
and U7347 (N_7347,N_7048,N_7171);
or U7348 (N_7348,N_7167,N_7160);
and U7349 (N_7349,N_7134,N_7192);
nor U7350 (N_7350,N_7175,N_7114);
and U7351 (N_7351,N_7196,N_7181);
nor U7352 (N_7352,N_7080,N_7150);
or U7353 (N_7353,N_7112,N_7182);
or U7354 (N_7354,N_7140,N_7164);
or U7355 (N_7355,N_7161,N_7164);
nor U7356 (N_7356,N_7195,N_7084);
or U7357 (N_7357,N_7185,N_7117);
nand U7358 (N_7358,N_7064,N_7112);
xor U7359 (N_7359,N_7116,N_7066);
and U7360 (N_7360,N_7358,N_7257);
or U7361 (N_7361,N_7223,N_7217);
or U7362 (N_7362,N_7357,N_7299);
nand U7363 (N_7363,N_7273,N_7230);
nand U7364 (N_7364,N_7337,N_7272);
or U7365 (N_7365,N_7295,N_7234);
and U7366 (N_7366,N_7349,N_7275);
xnor U7367 (N_7367,N_7352,N_7255);
nand U7368 (N_7368,N_7214,N_7228);
nand U7369 (N_7369,N_7329,N_7262);
nand U7370 (N_7370,N_7277,N_7249);
nand U7371 (N_7371,N_7316,N_7248);
xnor U7372 (N_7372,N_7258,N_7333);
and U7373 (N_7373,N_7315,N_7319);
or U7374 (N_7374,N_7274,N_7318);
nor U7375 (N_7375,N_7332,N_7323);
nand U7376 (N_7376,N_7285,N_7331);
xnor U7377 (N_7377,N_7287,N_7336);
or U7378 (N_7378,N_7338,N_7310);
nand U7379 (N_7379,N_7216,N_7350);
or U7380 (N_7380,N_7283,N_7312);
nor U7381 (N_7381,N_7268,N_7313);
and U7382 (N_7382,N_7294,N_7322);
nor U7383 (N_7383,N_7266,N_7259);
or U7384 (N_7384,N_7340,N_7296);
nor U7385 (N_7385,N_7282,N_7244);
nand U7386 (N_7386,N_7229,N_7256);
nand U7387 (N_7387,N_7225,N_7314);
and U7388 (N_7388,N_7231,N_7292);
nor U7389 (N_7389,N_7200,N_7269);
or U7390 (N_7390,N_7250,N_7240);
or U7391 (N_7391,N_7254,N_7267);
nand U7392 (N_7392,N_7220,N_7201);
or U7393 (N_7393,N_7281,N_7236);
or U7394 (N_7394,N_7279,N_7284);
nand U7395 (N_7395,N_7242,N_7245);
and U7396 (N_7396,N_7286,N_7355);
and U7397 (N_7397,N_7289,N_7304);
nor U7398 (N_7398,N_7328,N_7335);
nor U7399 (N_7399,N_7264,N_7306);
nand U7400 (N_7400,N_7345,N_7260);
nand U7401 (N_7401,N_7202,N_7271);
nand U7402 (N_7402,N_7341,N_7243);
and U7403 (N_7403,N_7219,N_7227);
nor U7404 (N_7404,N_7263,N_7239);
or U7405 (N_7405,N_7302,N_7356);
and U7406 (N_7406,N_7359,N_7326);
or U7407 (N_7407,N_7317,N_7209);
nor U7408 (N_7408,N_7207,N_7330);
and U7409 (N_7409,N_7205,N_7252);
nor U7410 (N_7410,N_7253,N_7293);
xor U7411 (N_7411,N_7278,N_7308);
and U7412 (N_7412,N_7307,N_7291);
or U7413 (N_7413,N_7247,N_7343);
nand U7414 (N_7414,N_7224,N_7241);
nand U7415 (N_7415,N_7208,N_7290);
or U7416 (N_7416,N_7211,N_7354);
or U7417 (N_7417,N_7300,N_7246);
nand U7418 (N_7418,N_7238,N_7203);
nand U7419 (N_7419,N_7303,N_7280);
nor U7420 (N_7420,N_7309,N_7213);
nor U7421 (N_7421,N_7347,N_7215);
or U7422 (N_7422,N_7212,N_7251);
and U7423 (N_7423,N_7344,N_7311);
nor U7424 (N_7424,N_7204,N_7233);
and U7425 (N_7425,N_7353,N_7351);
nor U7426 (N_7426,N_7342,N_7232);
or U7427 (N_7427,N_7327,N_7298);
nand U7428 (N_7428,N_7346,N_7235);
nand U7429 (N_7429,N_7348,N_7222);
or U7430 (N_7430,N_7265,N_7276);
or U7431 (N_7431,N_7210,N_7226);
nor U7432 (N_7432,N_7321,N_7339);
nor U7433 (N_7433,N_7237,N_7325);
xor U7434 (N_7434,N_7288,N_7324);
or U7435 (N_7435,N_7320,N_7334);
and U7436 (N_7436,N_7261,N_7221);
and U7437 (N_7437,N_7218,N_7305);
nand U7438 (N_7438,N_7301,N_7206);
nand U7439 (N_7439,N_7270,N_7297);
nand U7440 (N_7440,N_7204,N_7226);
and U7441 (N_7441,N_7273,N_7269);
or U7442 (N_7442,N_7219,N_7357);
nor U7443 (N_7443,N_7353,N_7238);
nand U7444 (N_7444,N_7240,N_7308);
or U7445 (N_7445,N_7222,N_7276);
nand U7446 (N_7446,N_7302,N_7305);
and U7447 (N_7447,N_7245,N_7299);
or U7448 (N_7448,N_7219,N_7235);
or U7449 (N_7449,N_7313,N_7290);
or U7450 (N_7450,N_7325,N_7331);
nor U7451 (N_7451,N_7251,N_7211);
nand U7452 (N_7452,N_7251,N_7208);
nand U7453 (N_7453,N_7257,N_7300);
nand U7454 (N_7454,N_7343,N_7206);
nand U7455 (N_7455,N_7203,N_7339);
nor U7456 (N_7456,N_7213,N_7335);
nand U7457 (N_7457,N_7279,N_7324);
nand U7458 (N_7458,N_7327,N_7241);
and U7459 (N_7459,N_7221,N_7201);
nand U7460 (N_7460,N_7307,N_7241);
nor U7461 (N_7461,N_7356,N_7220);
and U7462 (N_7462,N_7325,N_7265);
or U7463 (N_7463,N_7332,N_7317);
nor U7464 (N_7464,N_7250,N_7302);
or U7465 (N_7465,N_7245,N_7295);
and U7466 (N_7466,N_7334,N_7273);
nand U7467 (N_7467,N_7223,N_7233);
and U7468 (N_7468,N_7302,N_7240);
or U7469 (N_7469,N_7204,N_7264);
and U7470 (N_7470,N_7285,N_7280);
nand U7471 (N_7471,N_7306,N_7205);
or U7472 (N_7472,N_7275,N_7297);
nand U7473 (N_7473,N_7284,N_7230);
nor U7474 (N_7474,N_7238,N_7333);
and U7475 (N_7475,N_7213,N_7260);
nand U7476 (N_7476,N_7325,N_7275);
and U7477 (N_7477,N_7250,N_7262);
or U7478 (N_7478,N_7334,N_7298);
nor U7479 (N_7479,N_7301,N_7303);
nor U7480 (N_7480,N_7240,N_7353);
nand U7481 (N_7481,N_7337,N_7353);
nand U7482 (N_7482,N_7216,N_7221);
nand U7483 (N_7483,N_7299,N_7283);
nor U7484 (N_7484,N_7223,N_7296);
or U7485 (N_7485,N_7240,N_7200);
nor U7486 (N_7486,N_7261,N_7241);
and U7487 (N_7487,N_7318,N_7200);
xor U7488 (N_7488,N_7299,N_7323);
nor U7489 (N_7489,N_7351,N_7291);
or U7490 (N_7490,N_7218,N_7249);
and U7491 (N_7491,N_7204,N_7306);
xnor U7492 (N_7492,N_7326,N_7303);
nor U7493 (N_7493,N_7203,N_7219);
nor U7494 (N_7494,N_7262,N_7291);
xnor U7495 (N_7495,N_7302,N_7296);
nor U7496 (N_7496,N_7351,N_7232);
or U7497 (N_7497,N_7325,N_7312);
nand U7498 (N_7498,N_7218,N_7319);
nand U7499 (N_7499,N_7217,N_7324);
and U7500 (N_7500,N_7323,N_7208);
and U7501 (N_7501,N_7277,N_7233);
nand U7502 (N_7502,N_7226,N_7299);
nand U7503 (N_7503,N_7287,N_7222);
and U7504 (N_7504,N_7220,N_7340);
nand U7505 (N_7505,N_7335,N_7336);
nor U7506 (N_7506,N_7323,N_7306);
nand U7507 (N_7507,N_7274,N_7235);
xor U7508 (N_7508,N_7321,N_7247);
nand U7509 (N_7509,N_7267,N_7272);
nand U7510 (N_7510,N_7233,N_7280);
and U7511 (N_7511,N_7334,N_7314);
and U7512 (N_7512,N_7302,N_7337);
nand U7513 (N_7513,N_7317,N_7346);
nor U7514 (N_7514,N_7272,N_7234);
or U7515 (N_7515,N_7330,N_7307);
nor U7516 (N_7516,N_7249,N_7217);
nor U7517 (N_7517,N_7346,N_7212);
or U7518 (N_7518,N_7243,N_7314);
or U7519 (N_7519,N_7242,N_7359);
nor U7520 (N_7520,N_7416,N_7401);
or U7521 (N_7521,N_7362,N_7410);
and U7522 (N_7522,N_7515,N_7497);
xor U7523 (N_7523,N_7418,N_7361);
nand U7524 (N_7524,N_7481,N_7424);
xnor U7525 (N_7525,N_7514,N_7402);
or U7526 (N_7526,N_7494,N_7399);
and U7527 (N_7527,N_7476,N_7395);
and U7528 (N_7528,N_7383,N_7413);
nor U7529 (N_7529,N_7468,N_7412);
nand U7530 (N_7530,N_7466,N_7512);
nand U7531 (N_7531,N_7495,N_7434);
and U7532 (N_7532,N_7447,N_7427);
xor U7533 (N_7533,N_7386,N_7435);
and U7534 (N_7534,N_7408,N_7465);
nand U7535 (N_7535,N_7450,N_7437);
xnor U7536 (N_7536,N_7398,N_7444);
and U7537 (N_7537,N_7407,N_7365);
nand U7538 (N_7538,N_7460,N_7499);
xor U7539 (N_7539,N_7436,N_7371);
xnor U7540 (N_7540,N_7480,N_7459);
nand U7541 (N_7541,N_7429,N_7380);
and U7542 (N_7542,N_7491,N_7409);
nand U7543 (N_7543,N_7463,N_7461);
xnor U7544 (N_7544,N_7496,N_7502);
or U7545 (N_7545,N_7516,N_7455);
nand U7546 (N_7546,N_7477,N_7379);
nand U7547 (N_7547,N_7475,N_7454);
nand U7548 (N_7548,N_7377,N_7451);
nand U7549 (N_7549,N_7483,N_7414);
nor U7550 (N_7550,N_7430,N_7471);
xnor U7551 (N_7551,N_7397,N_7441);
nand U7552 (N_7552,N_7373,N_7394);
xnor U7553 (N_7553,N_7406,N_7443);
nor U7554 (N_7554,N_7484,N_7506);
nor U7555 (N_7555,N_7464,N_7501);
nand U7556 (N_7556,N_7452,N_7390);
or U7557 (N_7557,N_7510,N_7445);
and U7558 (N_7558,N_7389,N_7367);
or U7559 (N_7559,N_7503,N_7363);
nand U7560 (N_7560,N_7387,N_7498);
and U7561 (N_7561,N_7511,N_7469);
and U7562 (N_7562,N_7405,N_7487);
and U7563 (N_7563,N_7378,N_7369);
nand U7564 (N_7564,N_7372,N_7519);
or U7565 (N_7565,N_7448,N_7384);
nor U7566 (N_7566,N_7360,N_7513);
or U7567 (N_7567,N_7391,N_7400);
and U7568 (N_7568,N_7375,N_7376);
xnor U7569 (N_7569,N_7381,N_7489);
xnor U7570 (N_7570,N_7507,N_7432);
nand U7571 (N_7571,N_7392,N_7508);
and U7572 (N_7572,N_7411,N_7509);
and U7573 (N_7573,N_7396,N_7433);
nand U7574 (N_7574,N_7393,N_7505);
and U7575 (N_7575,N_7456,N_7462);
or U7576 (N_7576,N_7404,N_7492);
nand U7577 (N_7577,N_7486,N_7382);
xnor U7578 (N_7578,N_7431,N_7388);
xnor U7579 (N_7579,N_7490,N_7374);
nand U7580 (N_7580,N_7370,N_7426);
xnor U7581 (N_7581,N_7474,N_7403);
and U7582 (N_7582,N_7439,N_7366);
and U7583 (N_7583,N_7500,N_7421);
or U7584 (N_7584,N_7417,N_7482);
xor U7585 (N_7585,N_7446,N_7504);
xnor U7586 (N_7586,N_7423,N_7518);
nand U7587 (N_7587,N_7470,N_7457);
nor U7588 (N_7588,N_7479,N_7458);
and U7589 (N_7589,N_7442,N_7440);
xor U7590 (N_7590,N_7467,N_7425);
or U7591 (N_7591,N_7438,N_7473);
or U7592 (N_7592,N_7517,N_7488);
nor U7593 (N_7593,N_7449,N_7419);
or U7594 (N_7594,N_7385,N_7472);
nor U7595 (N_7595,N_7478,N_7485);
and U7596 (N_7596,N_7493,N_7428);
xor U7597 (N_7597,N_7415,N_7453);
nor U7598 (N_7598,N_7364,N_7420);
or U7599 (N_7599,N_7368,N_7422);
and U7600 (N_7600,N_7401,N_7474);
or U7601 (N_7601,N_7416,N_7480);
xor U7602 (N_7602,N_7497,N_7437);
and U7603 (N_7603,N_7396,N_7466);
nor U7604 (N_7604,N_7435,N_7511);
nand U7605 (N_7605,N_7376,N_7505);
xnor U7606 (N_7606,N_7508,N_7379);
and U7607 (N_7607,N_7462,N_7402);
nand U7608 (N_7608,N_7452,N_7488);
nand U7609 (N_7609,N_7453,N_7508);
nand U7610 (N_7610,N_7397,N_7469);
nand U7611 (N_7611,N_7385,N_7486);
nor U7612 (N_7612,N_7437,N_7514);
nand U7613 (N_7613,N_7461,N_7410);
nand U7614 (N_7614,N_7381,N_7485);
and U7615 (N_7615,N_7406,N_7476);
or U7616 (N_7616,N_7384,N_7446);
and U7617 (N_7617,N_7498,N_7405);
nor U7618 (N_7618,N_7381,N_7434);
nor U7619 (N_7619,N_7443,N_7516);
nor U7620 (N_7620,N_7364,N_7400);
and U7621 (N_7621,N_7368,N_7398);
xnor U7622 (N_7622,N_7503,N_7467);
or U7623 (N_7623,N_7442,N_7374);
nor U7624 (N_7624,N_7509,N_7366);
xor U7625 (N_7625,N_7480,N_7519);
and U7626 (N_7626,N_7415,N_7428);
or U7627 (N_7627,N_7428,N_7452);
and U7628 (N_7628,N_7371,N_7512);
nand U7629 (N_7629,N_7508,N_7384);
nor U7630 (N_7630,N_7414,N_7502);
nor U7631 (N_7631,N_7380,N_7430);
nand U7632 (N_7632,N_7485,N_7392);
or U7633 (N_7633,N_7484,N_7370);
nor U7634 (N_7634,N_7495,N_7385);
xnor U7635 (N_7635,N_7422,N_7516);
and U7636 (N_7636,N_7487,N_7518);
nor U7637 (N_7637,N_7490,N_7482);
or U7638 (N_7638,N_7450,N_7465);
xnor U7639 (N_7639,N_7478,N_7488);
nand U7640 (N_7640,N_7430,N_7456);
nor U7641 (N_7641,N_7481,N_7477);
nor U7642 (N_7642,N_7384,N_7485);
xor U7643 (N_7643,N_7404,N_7449);
nand U7644 (N_7644,N_7439,N_7477);
xnor U7645 (N_7645,N_7374,N_7431);
and U7646 (N_7646,N_7509,N_7388);
nand U7647 (N_7647,N_7438,N_7489);
and U7648 (N_7648,N_7505,N_7477);
and U7649 (N_7649,N_7514,N_7516);
nor U7650 (N_7650,N_7417,N_7514);
or U7651 (N_7651,N_7494,N_7374);
nand U7652 (N_7652,N_7405,N_7434);
nand U7653 (N_7653,N_7461,N_7448);
nor U7654 (N_7654,N_7457,N_7448);
or U7655 (N_7655,N_7392,N_7380);
or U7656 (N_7656,N_7408,N_7447);
or U7657 (N_7657,N_7422,N_7366);
or U7658 (N_7658,N_7415,N_7456);
and U7659 (N_7659,N_7414,N_7503);
or U7660 (N_7660,N_7377,N_7509);
xor U7661 (N_7661,N_7394,N_7447);
and U7662 (N_7662,N_7457,N_7517);
and U7663 (N_7663,N_7365,N_7516);
nor U7664 (N_7664,N_7414,N_7468);
nor U7665 (N_7665,N_7368,N_7441);
xor U7666 (N_7666,N_7387,N_7391);
nand U7667 (N_7667,N_7498,N_7396);
or U7668 (N_7668,N_7404,N_7505);
and U7669 (N_7669,N_7432,N_7405);
or U7670 (N_7670,N_7370,N_7451);
or U7671 (N_7671,N_7482,N_7371);
nand U7672 (N_7672,N_7376,N_7399);
or U7673 (N_7673,N_7401,N_7434);
nand U7674 (N_7674,N_7519,N_7438);
or U7675 (N_7675,N_7501,N_7462);
or U7676 (N_7676,N_7516,N_7474);
nand U7677 (N_7677,N_7444,N_7388);
and U7678 (N_7678,N_7378,N_7501);
and U7679 (N_7679,N_7476,N_7439);
xor U7680 (N_7680,N_7553,N_7646);
or U7681 (N_7681,N_7659,N_7520);
nor U7682 (N_7682,N_7633,N_7653);
or U7683 (N_7683,N_7639,N_7607);
and U7684 (N_7684,N_7581,N_7565);
xor U7685 (N_7685,N_7675,N_7635);
or U7686 (N_7686,N_7643,N_7587);
or U7687 (N_7687,N_7540,N_7589);
and U7688 (N_7688,N_7615,N_7625);
xnor U7689 (N_7689,N_7661,N_7528);
or U7690 (N_7690,N_7629,N_7627);
or U7691 (N_7691,N_7624,N_7531);
and U7692 (N_7692,N_7673,N_7620);
xor U7693 (N_7693,N_7674,N_7588);
and U7694 (N_7694,N_7601,N_7525);
nor U7695 (N_7695,N_7527,N_7618);
or U7696 (N_7696,N_7546,N_7617);
nor U7697 (N_7697,N_7664,N_7597);
nand U7698 (N_7698,N_7642,N_7539);
or U7699 (N_7699,N_7522,N_7605);
nand U7700 (N_7700,N_7551,N_7543);
xor U7701 (N_7701,N_7591,N_7628);
nand U7702 (N_7702,N_7610,N_7623);
nor U7703 (N_7703,N_7600,N_7614);
or U7704 (N_7704,N_7542,N_7663);
nor U7705 (N_7705,N_7599,N_7652);
and U7706 (N_7706,N_7598,N_7666);
nand U7707 (N_7707,N_7556,N_7622);
or U7708 (N_7708,N_7577,N_7631);
nand U7709 (N_7709,N_7557,N_7541);
nand U7710 (N_7710,N_7651,N_7580);
nor U7711 (N_7711,N_7634,N_7665);
or U7712 (N_7712,N_7604,N_7578);
nand U7713 (N_7713,N_7590,N_7537);
nor U7714 (N_7714,N_7649,N_7611);
nor U7715 (N_7715,N_7535,N_7526);
nor U7716 (N_7716,N_7523,N_7650);
nand U7717 (N_7717,N_7647,N_7552);
or U7718 (N_7718,N_7559,N_7569);
or U7719 (N_7719,N_7658,N_7563);
nand U7720 (N_7720,N_7585,N_7676);
nor U7721 (N_7721,N_7533,N_7637);
nand U7722 (N_7722,N_7626,N_7632);
nand U7723 (N_7723,N_7566,N_7572);
and U7724 (N_7724,N_7677,N_7638);
nor U7725 (N_7725,N_7655,N_7612);
and U7726 (N_7726,N_7583,N_7606);
nand U7727 (N_7727,N_7592,N_7571);
nor U7728 (N_7728,N_7574,N_7561);
or U7729 (N_7729,N_7562,N_7656);
xor U7730 (N_7730,N_7584,N_7550);
nand U7731 (N_7731,N_7660,N_7595);
nor U7732 (N_7732,N_7636,N_7670);
nor U7733 (N_7733,N_7668,N_7544);
nor U7734 (N_7734,N_7640,N_7558);
or U7735 (N_7735,N_7579,N_7679);
and U7736 (N_7736,N_7529,N_7554);
and U7737 (N_7737,N_7573,N_7645);
xor U7738 (N_7738,N_7568,N_7667);
and U7739 (N_7739,N_7586,N_7613);
nor U7740 (N_7740,N_7555,N_7524);
or U7741 (N_7741,N_7570,N_7576);
nor U7742 (N_7742,N_7678,N_7657);
and U7743 (N_7743,N_7582,N_7545);
and U7744 (N_7744,N_7536,N_7654);
nor U7745 (N_7745,N_7648,N_7532);
and U7746 (N_7746,N_7567,N_7547);
xnor U7747 (N_7747,N_7534,N_7575);
or U7748 (N_7748,N_7602,N_7538);
and U7749 (N_7749,N_7630,N_7608);
nand U7750 (N_7750,N_7671,N_7548);
and U7751 (N_7751,N_7560,N_7672);
nor U7752 (N_7752,N_7596,N_7662);
and U7753 (N_7753,N_7549,N_7603);
nor U7754 (N_7754,N_7521,N_7644);
nand U7755 (N_7755,N_7641,N_7593);
or U7756 (N_7756,N_7564,N_7616);
nor U7757 (N_7757,N_7530,N_7621);
xnor U7758 (N_7758,N_7669,N_7609);
nand U7759 (N_7759,N_7619,N_7594);
nor U7760 (N_7760,N_7655,N_7658);
xnor U7761 (N_7761,N_7546,N_7626);
nor U7762 (N_7762,N_7635,N_7638);
nor U7763 (N_7763,N_7604,N_7657);
nor U7764 (N_7764,N_7625,N_7561);
or U7765 (N_7765,N_7536,N_7640);
nor U7766 (N_7766,N_7535,N_7576);
or U7767 (N_7767,N_7624,N_7580);
and U7768 (N_7768,N_7637,N_7530);
nand U7769 (N_7769,N_7562,N_7529);
or U7770 (N_7770,N_7532,N_7651);
or U7771 (N_7771,N_7613,N_7618);
nor U7772 (N_7772,N_7595,N_7613);
nor U7773 (N_7773,N_7612,N_7622);
nor U7774 (N_7774,N_7556,N_7638);
or U7775 (N_7775,N_7656,N_7551);
or U7776 (N_7776,N_7573,N_7580);
nor U7777 (N_7777,N_7679,N_7670);
nor U7778 (N_7778,N_7671,N_7631);
or U7779 (N_7779,N_7601,N_7679);
nand U7780 (N_7780,N_7661,N_7597);
nand U7781 (N_7781,N_7663,N_7528);
nand U7782 (N_7782,N_7663,N_7577);
and U7783 (N_7783,N_7553,N_7591);
xor U7784 (N_7784,N_7572,N_7581);
and U7785 (N_7785,N_7536,N_7565);
nor U7786 (N_7786,N_7566,N_7554);
nand U7787 (N_7787,N_7574,N_7570);
nand U7788 (N_7788,N_7597,N_7592);
and U7789 (N_7789,N_7556,N_7593);
and U7790 (N_7790,N_7602,N_7524);
nor U7791 (N_7791,N_7624,N_7613);
xor U7792 (N_7792,N_7663,N_7529);
nor U7793 (N_7793,N_7626,N_7556);
xor U7794 (N_7794,N_7521,N_7576);
nand U7795 (N_7795,N_7669,N_7557);
or U7796 (N_7796,N_7600,N_7610);
or U7797 (N_7797,N_7658,N_7661);
nand U7798 (N_7798,N_7679,N_7657);
xor U7799 (N_7799,N_7522,N_7576);
nor U7800 (N_7800,N_7642,N_7646);
xnor U7801 (N_7801,N_7617,N_7643);
nor U7802 (N_7802,N_7654,N_7610);
and U7803 (N_7803,N_7592,N_7558);
and U7804 (N_7804,N_7568,N_7663);
nand U7805 (N_7805,N_7652,N_7658);
nor U7806 (N_7806,N_7672,N_7575);
and U7807 (N_7807,N_7662,N_7639);
xnor U7808 (N_7808,N_7637,N_7647);
and U7809 (N_7809,N_7613,N_7577);
nor U7810 (N_7810,N_7527,N_7593);
and U7811 (N_7811,N_7569,N_7589);
nand U7812 (N_7812,N_7536,N_7544);
or U7813 (N_7813,N_7611,N_7653);
nor U7814 (N_7814,N_7629,N_7664);
or U7815 (N_7815,N_7649,N_7603);
and U7816 (N_7816,N_7650,N_7627);
nand U7817 (N_7817,N_7631,N_7648);
or U7818 (N_7818,N_7584,N_7582);
nor U7819 (N_7819,N_7639,N_7610);
nand U7820 (N_7820,N_7587,N_7534);
nor U7821 (N_7821,N_7592,N_7622);
nand U7822 (N_7822,N_7618,N_7565);
nor U7823 (N_7823,N_7566,N_7520);
nor U7824 (N_7824,N_7629,N_7613);
or U7825 (N_7825,N_7611,N_7595);
nand U7826 (N_7826,N_7583,N_7528);
nor U7827 (N_7827,N_7575,N_7625);
nand U7828 (N_7828,N_7567,N_7562);
nor U7829 (N_7829,N_7613,N_7610);
nor U7830 (N_7830,N_7615,N_7598);
nand U7831 (N_7831,N_7640,N_7652);
and U7832 (N_7832,N_7643,N_7613);
xor U7833 (N_7833,N_7669,N_7671);
nor U7834 (N_7834,N_7585,N_7564);
nand U7835 (N_7835,N_7648,N_7545);
nand U7836 (N_7836,N_7621,N_7561);
xnor U7837 (N_7837,N_7597,N_7642);
or U7838 (N_7838,N_7672,N_7679);
nor U7839 (N_7839,N_7534,N_7637);
or U7840 (N_7840,N_7821,N_7833);
nor U7841 (N_7841,N_7766,N_7750);
and U7842 (N_7842,N_7781,N_7744);
nand U7843 (N_7843,N_7724,N_7756);
nand U7844 (N_7844,N_7746,N_7700);
or U7845 (N_7845,N_7776,N_7827);
nor U7846 (N_7846,N_7795,N_7720);
nor U7847 (N_7847,N_7764,N_7823);
and U7848 (N_7848,N_7836,N_7802);
nand U7849 (N_7849,N_7784,N_7765);
or U7850 (N_7850,N_7683,N_7837);
nand U7851 (N_7851,N_7773,N_7811);
nand U7852 (N_7852,N_7785,N_7684);
or U7853 (N_7853,N_7695,N_7754);
and U7854 (N_7854,N_7741,N_7828);
nor U7855 (N_7855,N_7745,N_7796);
nor U7856 (N_7856,N_7838,N_7693);
or U7857 (N_7857,N_7751,N_7787);
or U7858 (N_7858,N_7714,N_7778);
xnor U7859 (N_7859,N_7747,N_7697);
and U7860 (N_7860,N_7688,N_7711);
and U7861 (N_7861,N_7757,N_7723);
nand U7862 (N_7862,N_7780,N_7769);
or U7863 (N_7863,N_7767,N_7791);
or U7864 (N_7864,N_7709,N_7815);
nand U7865 (N_7865,N_7749,N_7702);
nand U7866 (N_7866,N_7812,N_7813);
and U7867 (N_7867,N_7715,N_7771);
and U7868 (N_7868,N_7730,N_7738);
nor U7869 (N_7869,N_7682,N_7835);
nand U7870 (N_7870,N_7699,N_7829);
nand U7871 (N_7871,N_7708,N_7712);
and U7872 (N_7872,N_7731,N_7788);
and U7873 (N_7873,N_7740,N_7736);
and U7874 (N_7874,N_7803,N_7696);
and U7875 (N_7875,N_7820,N_7814);
nand U7876 (N_7876,N_7698,N_7800);
xnor U7877 (N_7877,N_7689,N_7687);
and U7878 (N_7878,N_7799,N_7779);
or U7879 (N_7879,N_7789,N_7830);
and U7880 (N_7880,N_7713,N_7703);
nand U7881 (N_7881,N_7792,N_7735);
nand U7882 (N_7882,N_7806,N_7733);
nor U7883 (N_7883,N_7832,N_7834);
nand U7884 (N_7884,N_7777,N_7692);
nand U7885 (N_7885,N_7755,N_7763);
nand U7886 (N_7886,N_7824,N_7726);
nand U7887 (N_7887,N_7760,N_7772);
xor U7888 (N_7888,N_7797,N_7717);
nand U7889 (N_7889,N_7742,N_7753);
nor U7890 (N_7890,N_7768,N_7818);
xor U7891 (N_7891,N_7707,N_7801);
and U7892 (N_7892,N_7710,N_7743);
and U7893 (N_7893,N_7762,N_7774);
nand U7894 (N_7894,N_7701,N_7732);
nor U7895 (N_7895,N_7825,N_7816);
nand U7896 (N_7896,N_7759,N_7794);
nor U7897 (N_7897,N_7839,N_7783);
and U7898 (N_7898,N_7805,N_7734);
or U7899 (N_7899,N_7685,N_7786);
nand U7900 (N_7900,N_7817,N_7822);
nand U7901 (N_7901,N_7819,N_7719);
or U7902 (N_7902,N_7681,N_7725);
nor U7903 (N_7903,N_7758,N_7770);
and U7904 (N_7904,N_7739,N_7748);
nor U7905 (N_7905,N_7826,N_7807);
nand U7906 (N_7906,N_7686,N_7790);
or U7907 (N_7907,N_7716,N_7808);
and U7908 (N_7908,N_7705,N_7727);
nand U7909 (N_7909,N_7704,N_7804);
nor U7910 (N_7910,N_7809,N_7775);
nor U7911 (N_7911,N_7721,N_7782);
or U7912 (N_7912,N_7694,N_7761);
or U7913 (N_7913,N_7737,N_7718);
and U7914 (N_7914,N_7793,N_7831);
xor U7915 (N_7915,N_7722,N_7691);
or U7916 (N_7916,N_7810,N_7690);
and U7917 (N_7917,N_7752,N_7680);
or U7918 (N_7918,N_7729,N_7798);
and U7919 (N_7919,N_7728,N_7706);
xnor U7920 (N_7920,N_7805,N_7710);
nand U7921 (N_7921,N_7683,N_7743);
and U7922 (N_7922,N_7818,N_7738);
or U7923 (N_7923,N_7692,N_7705);
nor U7924 (N_7924,N_7797,N_7783);
nor U7925 (N_7925,N_7788,N_7711);
xor U7926 (N_7926,N_7690,N_7681);
or U7927 (N_7927,N_7783,N_7786);
nand U7928 (N_7928,N_7740,N_7796);
or U7929 (N_7929,N_7815,N_7767);
nand U7930 (N_7930,N_7762,N_7777);
or U7931 (N_7931,N_7839,N_7772);
nand U7932 (N_7932,N_7814,N_7726);
xor U7933 (N_7933,N_7787,N_7828);
or U7934 (N_7934,N_7787,N_7826);
and U7935 (N_7935,N_7822,N_7688);
or U7936 (N_7936,N_7700,N_7729);
and U7937 (N_7937,N_7734,N_7766);
nor U7938 (N_7938,N_7753,N_7771);
nor U7939 (N_7939,N_7794,N_7771);
or U7940 (N_7940,N_7757,N_7779);
xnor U7941 (N_7941,N_7807,N_7827);
and U7942 (N_7942,N_7765,N_7722);
and U7943 (N_7943,N_7762,N_7824);
nor U7944 (N_7944,N_7805,N_7806);
nor U7945 (N_7945,N_7771,N_7699);
and U7946 (N_7946,N_7765,N_7754);
nand U7947 (N_7947,N_7682,N_7712);
or U7948 (N_7948,N_7778,N_7816);
nor U7949 (N_7949,N_7701,N_7696);
or U7950 (N_7950,N_7797,N_7735);
and U7951 (N_7951,N_7813,N_7729);
nand U7952 (N_7952,N_7697,N_7767);
or U7953 (N_7953,N_7727,N_7747);
nor U7954 (N_7954,N_7770,N_7833);
or U7955 (N_7955,N_7767,N_7740);
or U7956 (N_7956,N_7795,N_7806);
nand U7957 (N_7957,N_7802,N_7821);
nor U7958 (N_7958,N_7711,N_7785);
nand U7959 (N_7959,N_7754,N_7685);
nand U7960 (N_7960,N_7683,N_7818);
or U7961 (N_7961,N_7713,N_7777);
nand U7962 (N_7962,N_7819,N_7837);
nand U7963 (N_7963,N_7725,N_7715);
or U7964 (N_7964,N_7778,N_7815);
xor U7965 (N_7965,N_7775,N_7768);
nand U7966 (N_7966,N_7766,N_7767);
nand U7967 (N_7967,N_7732,N_7715);
or U7968 (N_7968,N_7801,N_7705);
or U7969 (N_7969,N_7789,N_7733);
and U7970 (N_7970,N_7700,N_7763);
or U7971 (N_7971,N_7726,N_7813);
and U7972 (N_7972,N_7803,N_7695);
or U7973 (N_7973,N_7681,N_7717);
nand U7974 (N_7974,N_7749,N_7831);
xnor U7975 (N_7975,N_7762,N_7720);
or U7976 (N_7976,N_7683,N_7714);
nor U7977 (N_7977,N_7816,N_7758);
nor U7978 (N_7978,N_7743,N_7746);
or U7979 (N_7979,N_7831,N_7755);
nand U7980 (N_7980,N_7785,N_7811);
and U7981 (N_7981,N_7820,N_7818);
nand U7982 (N_7982,N_7781,N_7815);
nor U7983 (N_7983,N_7736,N_7715);
nand U7984 (N_7984,N_7752,N_7794);
xor U7985 (N_7985,N_7696,N_7831);
and U7986 (N_7986,N_7752,N_7836);
xor U7987 (N_7987,N_7815,N_7747);
nand U7988 (N_7988,N_7717,N_7706);
xnor U7989 (N_7989,N_7778,N_7804);
xor U7990 (N_7990,N_7760,N_7745);
nand U7991 (N_7991,N_7784,N_7779);
nor U7992 (N_7992,N_7688,N_7698);
nor U7993 (N_7993,N_7817,N_7742);
xor U7994 (N_7994,N_7695,N_7832);
or U7995 (N_7995,N_7789,N_7728);
or U7996 (N_7996,N_7829,N_7683);
or U7997 (N_7997,N_7754,N_7775);
or U7998 (N_7998,N_7813,N_7823);
or U7999 (N_7999,N_7800,N_7793);
nand U8000 (N_8000,N_7856,N_7872);
nor U8001 (N_8001,N_7949,N_7895);
nor U8002 (N_8002,N_7988,N_7889);
nand U8003 (N_8003,N_7984,N_7944);
nor U8004 (N_8004,N_7901,N_7957);
or U8005 (N_8005,N_7867,N_7879);
and U8006 (N_8006,N_7921,N_7919);
nand U8007 (N_8007,N_7977,N_7946);
nor U8008 (N_8008,N_7947,N_7914);
or U8009 (N_8009,N_7854,N_7862);
nand U8010 (N_8010,N_7996,N_7954);
and U8011 (N_8011,N_7878,N_7913);
xor U8012 (N_8012,N_7936,N_7939);
and U8013 (N_8013,N_7871,N_7846);
nand U8014 (N_8014,N_7848,N_7940);
nand U8015 (N_8015,N_7865,N_7916);
and U8016 (N_8016,N_7979,N_7906);
and U8017 (N_8017,N_7986,N_7966);
and U8018 (N_8018,N_7881,N_7942);
nor U8019 (N_8019,N_7853,N_7961);
nand U8020 (N_8020,N_7880,N_7959);
and U8021 (N_8021,N_7841,N_7902);
and U8022 (N_8022,N_7953,N_7859);
nor U8023 (N_8023,N_7993,N_7960);
nor U8024 (N_8024,N_7897,N_7973);
or U8025 (N_8025,N_7999,N_7910);
xnor U8026 (N_8026,N_7900,N_7938);
nor U8027 (N_8027,N_7975,N_7863);
xor U8028 (N_8028,N_7968,N_7912);
xnor U8029 (N_8029,N_7971,N_7886);
nand U8030 (N_8030,N_7903,N_7987);
nor U8031 (N_8031,N_7958,N_7989);
nand U8032 (N_8032,N_7922,N_7969);
nor U8033 (N_8033,N_7941,N_7849);
and U8034 (N_8034,N_7976,N_7924);
and U8035 (N_8035,N_7929,N_7893);
nor U8036 (N_8036,N_7840,N_7930);
or U8037 (N_8037,N_7982,N_7937);
or U8038 (N_8038,N_7847,N_7927);
or U8039 (N_8039,N_7962,N_7928);
nor U8040 (N_8040,N_7844,N_7908);
or U8041 (N_8041,N_7997,N_7875);
xor U8042 (N_8042,N_7967,N_7874);
nand U8043 (N_8043,N_7860,N_7972);
nor U8044 (N_8044,N_7950,N_7985);
and U8045 (N_8045,N_7948,N_7885);
and U8046 (N_8046,N_7995,N_7888);
nand U8047 (N_8047,N_7980,N_7981);
or U8048 (N_8048,N_7945,N_7934);
xnor U8049 (N_8049,N_7898,N_7876);
or U8050 (N_8050,N_7943,N_7843);
nand U8051 (N_8051,N_7915,N_7883);
nand U8052 (N_8052,N_7850,N_7935);
or U8053 (N_8053,N_7917,N_7983);
nor U8054 (N_8054,N_7877,N_7992);
nor U8055 (N_8055,N_7866,N_7890);
nor U8056 (N_8056,N_7964,N_7923);
and U8057 (N_8057,N_7894,N_7884);
nand U8058 (N_8058,N_7994,N_7965);
and U8059 (N_8059,N_7882,N_7991);
xnor U8060 (N_8060,N_7963,N_7868);
or U8061 (N_8061,N_7869,N_7933);
or U8062 (N_8062,N_7931,N_7904);
nor U8063 (N_8063,N_7905,N_7970);
nor U8064 (N_8064,N_7842,N_7887);
or U8065 (N_8065,N_7864,N_7899);
or U8066 (N_8066,N_7951,N_7861);
and U8067 (N_8067,N_7952,N_7956);
or U8068 (N_8068,N_7990,N_7892);
and U8069 (N_8069,N_7974,N_7955);
and U8070 (N_8070,N_7891,N_7932);
nand U8071 (N_8071,N_7855,N_7998);
nand U8072 (N_8072,N_7851,N_7907);
nand U8073 (N_8073,N_7896,N_7873);
or U8074 (N_8074,N_7925,N_7909);
nor U8075 (N_8075,N_7858,N_7918);
nor U8076 (N_8076,N_7926,N_7911);
nand U8077 (N_8077,N_7845,N_7852);
and U8078 (N_8078,N_7857,N_7978);
xor U8079 (N_8079,N_7870,N_7920);
and U8080 (N_8080,N_7968,N_7881);
or U8081 (N_8081,N_7993,N_7946);
and U8082 (N_8082,N_7991,N_7933);
nand U8083 (N_8083,N_7939,N_7900);
xnor U8084 (N_8084,N_7865,N_7975);
or U8085 (N_8085,N_7978,N_7975);
and U8086 (N_8086,N_7872,N_7878);
or U8087 (N_8087,N_7939,N_7927);
nand U8088 (N_8088,N_7893,N_7903);
xnor U8089 (N_8089,N_7961,N_7897);
nand U8090 (N_8090,N_7948,N_7861);
or U8091 (N_8091,N_7923,N_7950);
or U8092 (N_8092,N_7930,N_7913);
xor U8093 (N_8093,N_7951,N_7858);
xnor U8094 (N_8094,N_7958,N_7917);
and U8095 (N_8095,N_7943,N_7869);
or U8096 (N_8096,N_7870,N_7965);
or U8097 (N_8097,N_7913,N_7948);
or U8098 (N_8098,N_7971,N_7964);
xor U8099 (N_8099,N_7917,N_7869);
and U8100 (N_8100,N_7922,N_7958);
xor U8101 (N_8101,N_7953,N_7938);
or U8102 (N_8102,N_7967,N_7887);
xnor U8103 (N_8103,N_7935,N_7910);
and U8104 (N_8104,N_7908,N_7909);
or U8105 (N_8105,N_7903,N_7937);
and U8106 (N_8106,N_7877,N_7967);
nor U8107 (N_8107,N_7942,N_7932);
nor U8108 (N_8108,N_7977,N_7912);
nand U8109 (N_8109,N_7993,N_7864);
nor U8110 (N_8110,N_7858,N_7856);
and U8111 (N_8111,N_7942,N_7951);
nand U8112 (N_8112,N_7992,N_7892);
and U8113 (N_8113,N_7870,N_7996);
nor U8114 (N_8114,N_7942,N_7869);
nor U8115 (N_8115,N_7866,N_7970);
nor U8116 (N_8116,N_7893,N_7879);
or U8117 (N_8117,N_7931,N_7923);
or U8118 (N_8118,N_7857,N_7849);
nand U8119 (N_8119,N_7861,N_7892);
or U8120 (N_8120,N_7872,N_7972);
and U8121 (N_8121,N_7853,N_7906);
and U8122 (N_8122,N_7995,N_7982);
nand U8123 (N_8123,N_7940,N_7959);
or U8124 (N_8124,N_7890,N_7954);
or U8125 (N_8125,N_7974,N_7980);
xor U8126 (N_8126,N_7918,N_7953);
and U8127 (N_8127,N_7904,N_7944);
or U8128 (N_8128,N_7997,N_7854);
and U8129 (N_8129,N_7946,N_7933);
nor U8130 (N_8130,N_7892,N_7847);
and U8131 (N_8131,N_7921,N_7848);
and U8132 (N_8132,N_7857,N_7922);
and U8133 (N_8133,N_7862,N_7873);
and U8134 (N_8134,N_7916,N_7860);
nand U8135 (N_8135,N_7874,N_7973);
nor U8136 (N_8136,N_7884,N_7926);
or U8137 (N_8137,N_7856,N_7950);
xnor U8138 (N_8138,N_7913,N_7923);
nor U8139 (N_8139,N_7851,N_7858);
and U8140 (N_8140,N_7942,N_7852);
nand U8141 (N_8141,N_7979,N_7910);
nand U8142 (N_8142,N_7852,N_7885);
and U8143 (N_8143,N_7931,N_7996);
nor U8144 (N_8144,N_7890,N_7928);
nor U8145 (N_8145,N_7877,N_7936);
or U8146 (N_8146,N_7956,N_7935);
or U8147 (N_8147,N_7842,N_7935);
nor U8148 (N_8148,N_7942,N_7998);
xor U8149 (N_8149,N_7873,N_7886);
and U8150 (N_8150,N_7929,N_7980);
xor U8151 (N_8151,N_7995,N_7962);
and U8152 (N_8152,N_7860,N_7874);
nand U8153 (N_8153,N_7964,N_7844);
and U8154 (N_8154,N_7986,N_7928);
or U8155 (N_8155,N_7997,N_7963);
and U8156 (N_8156,N_7922,N_7909);
and U8157 (N_8157,N_7907,N_7854);
and U8158 (N_8158,N_7855,N_7859);
nand U8159 (N_8159,N_7957,N_7882);
and U8160 (N_8160,N_8009,N_8077);
nor U8161 (N_8161,N_8097,N_8007);
nand U8162 (N_8162,N_8096,N_8157);
or U8163 (N_8163,N_8037,N_8150);
nand U8164 (N_8164,N_8129,N_8004);
nor U8165 (N_8165,N_8021,N_8019);
xnor U8166 (N_8166,N_8047,N_8158);
and U8167 (N_8167,N_8038,N_8045);
nor U8168 (N_8168,N_8029,N_8035);
or U8169 (N_8169,N_8111,N_8136);
nor U8170 (N_8170,N_8008,N_8141);
nor U8171 (N_8171,N_8052,N_8114);
nor U8172 (N_8172,N_8092,N_8018);
or U8173 (N_8173,N_8034,N_8084);
nor U8174 (N_8174,N_8140,N_8022);
nor U8175 (N_8175,N_8054,N_8010);
nand U8176 (N_8176,N_8102,N_8066);
or U8177 (N_8177,N_8119,N_8147);
nor U8178 (N_8178,N_8016,N_8027);
or U8179 (N_8179,N_8134,N_8124);
nand U8180 (N_8180,N_8087,N_8023);
nor U8181 (N_8181,N_8154,N_8030);
nand U8182 (N_8182,N_8053,N_8011);
nand U8183 (N_8183,N_8090,N_8067);
and U8184 (N_8184,N_8131,N_8148);
nor U8185 (N_8185,N_8100,N_8076);
nor U8186 (N_8186,N_8137,N_8159);
nor U8187 (N_8187,N_8062,N_8048);
nand U8188 (N_8188,N_8091,N_8068);
and U8189 (N_8189,N_8138,N_8000);
and U8190 (N_8190,N_8130,N_8003);
and U8191 (N_8191,N_8074,N_8012);
or U8192 (N_8192,N_8046,N_8122);
nand U8193 (N_8193,N_8050,N_8146);
and U8194 (N_8194,N_8020,N_8039);
or U8195 (N_8195,N_8017,N_8115);
nor U8196 (N_8196,N_8069,N_8075);
nand U8197 (N_8197,N_8112,N_8121);
nand U8198 (N_8198,N_8072,N_8151);
or U8199 (N_8199,N_8109,N_8086);
or U8200 (N_8200,N_8058,N_8040);
nand U8201 (N_8201,N_8070,N_8133);
and U8202 (N_8202,N_8107,N_8063);
nand U8203 (N_8203,N_8028,N_8117);
or U8204 (N_8204,N_8155,N_8156);
and U8205 (N_8205,N_8042,N_8057);
nor U8206 (N_8206,N_8025,N_8123);
or U8207 (N_8207,N_8093,N_8031);
and U8208 (N_8208,N_8094,N_8015);
or U8209 (N_8209,N_8079,N_8118);
nor U8210 (N_8210,N_8024,N_8041);
and U8211 (N_8211,N_8005,N_8044);
nand U8212 (N_8212,N_8149,N_8078);
nor U8213 (N_8213,N_8081,N_8055);
and U8214 (N_8214,N_8139,N_8105);
nand U8215 (N_8215,N_8033,N_8145);
xor U8216 (N_8216,N_8059,N_8064);
nor U8217 (N_8217,N_8116,N_8108);
or U8218 (N_8218,N_8002,N_8071);
nand U8219 (N_8219,N_8103,N_8089);
nor U8220 (N_8220,N_8153,N_8099);
nor U8221 (N_8221,N_8061,N_8013);
xor U8222 (N_8222,N_8043,N_8085);
nor U8223 (N_8223,N_8051,N_8080);
nand U8224 (N_8224,N_8128,N_8032);
nand U8225 (N_8225,N_8135,N_8120);
or U8226 (N_8226,N_8095,N_8060);
nor U8227 (N_8227,N_8101,N_8036);
or U8228 (N_8228,N_8127,N_8065);
xnor U8229 (N_8229,N_8088,N_8049);
nor U8230 (N_8230,N_8142,N_8083);
or U8231 (N_8231,N_8026,N_8106);
or U8232 (N_8232,N_8014,N_8104);
and U8233 (N_8233,N_8126,N_8098);
nand U8234 (N_8234,N_8144,N_8056);
or U8235 (N_8235,N_8006,N_8152);
xnor U8236 (N_8236,N_8001,N_8110);
or U8237 (N_8237,N_8113,N_8132);
or U8238 (N_8238,N_8082,N_8073);
nand U8239 (N_8239,N_8125,N_8143);
nor U8240 (N_8240,N_8113,N_8156);
nor U8241 (N_8241,N_8138,N_8149);
nor U8242 (N_8242,N_8079,N_8011);
nor U8243 (N_8243,N_8035,N_8066);
nand U8244 (N_8244,N_8086,N_8135);
xnor U8245 (N_8245,N_8075,N_8012);
nor U8246 (N_8246,N_8040,N_8080);
and U8247 (N_8247,N_8106,N_8049);
nand U8248 (N_8248,N_8113,N_8084);
nor U8249 (N_8249,N_8159,N_8048);
nand U8250 (N_8250,N_8065,N_8147);
or U8251 (N_8251,N_8113,N_8136);
and U8252 (N_8252,N_8132,N_8019);
nor U8253 (N_8253,N_8028,N_8000);
or U8254 (N_8254,N_8036,N_8085);
or U8255 (N_8255,N_8109,N_8114);
or U8256 (N_8256,N_8109,N_8104);
nand U8257 (N_8257,N_8154,N_8023);
nor U8258 (N_8258,N_8005,N_8060);
nor U8259 (N_8259,N_8082,N_8002);
or U8260 (N_8260,N_8146,N_8072);
nor U8261 (N_8261,N_8157,N_8042);
nand U8262 (N_8262,N_8053,N_8155);
nor U8263 (N_8263,N_8010,N_8106);
or U8264 (N_8264,N_8066,N_8009);
xor U8265 (N_8265,N_8017,N_8098);
nor U8266 (N_8266,N_8019,N_8127);
nor U8267 (N_8267,N_8067,N_8035);
nand U8268 (N_8268,N_8138,N_8117);
and U8269 (N_8269,N_8110,N_8136);
and U8270 (N_8270,N_8075,N_8100);
and U8271 (N_8271,N_8143,N_8145);
or U8272 (N_8272,N_8154,N_8070);
or U8273 (N_8273,N_8035,N_8032);
nand U8274 (N_8274,N_8066,N_8059);
or U8275 (N_8275,N_8127,N_8002);
nand U8276 (N_8276,N_8117,N_8113);
nor U8277 (N_8277,N_8056,N_8076);
xor U8278 (N_8278,N_8137,N_8125);
or U8279 (N_8279,N_8037,N_8062);
nand U8280 (N_8280,N_8011,N_8009);
nand U8281 (N_8281,N_8075,N_8117);
nor U8282 (N_8282,N_8056,N_8057);
nand U8283 (N_8283,N_8042,N_8088);
nand U8284 (N_8284,N_8104,N_8074);
nor U8285 (N_8285,N_8073,N_8055);
nand U8286 (N_8286,N_8055,N_8087);
nor U8287 (N_8287,N_8111,N_8035);
nor U8288 (N_8288,N_8018,N_8081);
nor U8289 (N_8289,N_8062,N_8143);
nor U8290 (N_8290,N_8058,N_8048);
or U8291 (N_8291,N_8078,N_8032);
and U8292 (N_8292,N_8034,N_8121);
nor U8293 (N_8293,N_8020,N_8060);
and U8294 (N_8294,N_8150,N_8141);
nand U8295 (N_8295,N_8039,N_8044);
or U8296 (N_8296,N_8002,N_8134);
and U8297 (N_8297,N_8091,N_8039);
xor U8298 (N_8298,N_8158,N_8075);
and U8299 (N_8299,N_8141,N_8142);
and U8300 (N_8300,N_8158,N_8058);
and U8301 (N_8301,N_8075,N_8092);
or U8302 (N_8302,N_8119,N_8135);
nand U8303 (N_8303,N_8026,N_8094);
and U8304 (N_8304,N_8079,N_8093);
and U8305 (N_8305,N_8053,N_8149);
or U8306 (N_8306,N_8146,N_8101);
nand U8307 (N_8307,N_8040,N_8024);
or U8308 (N_8308,N_8021,N_8095);
nor U8309 (N_8309,N_8019,N_8035);
nand U8310 (N_8310,N_8146,N_8010);
or U8311 (N_8311,N_8050,N_8062);
or U8312 (N_8312,N_8103,N_8008);
and U8313 (N_8313,N_8107,N_8153);
nor U8314 (N_8314,N_8103,N_8114);
xnor U8315 (N_8315,N_8071,N_8085);
or U8316 (N_8316,N_8094,N_8078);
nor U8317 (N_8317,N_8106,N_8013);
xnor U8318 (N_8318,N_8025,N_8125);
nor U8319 (N_8319,N_8090,N_8103);
or U8320 (N_8320,N_8240,N_8317);
or U8321 (N_8321,N_8253,N_8191);
and U8322 (N_8322,N_8164,N_8293);
nand U8323 (N_8323,N_8308,N_8197);
nand U8324 (N_8324,N_8278,N_8224);
nor U8325 (N_8325,N_8319,N_8222);
or U8326 (N_8326,N_8177,N_8304);
nor U8327 (N_8327,N_8228,N_8289);
nand U8328 (N_8328,N_8246,N_8263);
and U8329 (N_8329,N_8239,N_8300);
or U8330 (N_8330,N_8165,N_8296);
nand U8331 (N_8331,N_8294,N_8290);
nor U8332 (N_8332,N_8242,N_8301);
and U8333 (N_8333,N_8201,N_8273);
nor U8334 (N_8334,N_8173,N_8217);
or U8335 (N_8335,N_8210,N_8299);
and U8336 (N_8336,N_8193,N_8272);
nor U8337 (N_8337,N_8176,N_8287);
nor U8338 (N_8338,N_8220,N_8248);
nor U8339 (N_8339,N_8254,N_8245);
xnor U8340 (N_8340,N_8232,N_8281);
nand U8341 (N_8341,N_8206,N_8305);
or U8342 (N_8342,N_8172,N_8169);
nor U8343 (N_8343,N_8227,N_8212);
and U8344 (N_8344,N_8204,N_8297);
nand U8345 (N_8345,N_8233,N_8184);
xnor U8346 (N_8346,N_8178,N_8261);
nor U8347 (N_8347,N_8282,N_8311);
xor U8348 (N_8348,N_8251,N_8194);
and U8349 (N_8349,N_8257,N_8270);
xnor U8350 (N_8350,N_8265,N_8259);
xor U8351 (N_8351,N_8185,N_8284);
nor U8352 (N_8352,N_8195,N_8247);
and U8353 (N_8353,N_8243,N_8260);
xor U8354 (N_8354,N_8252,N_8303);
nand U8355 (N_8355,N_8234,N_8288);
nor U8356 (N_8356,N_8198,N_8186);
nor U8357 (N_8357,N_8256,N_8269);
nand U8358 (N_8358,N_8192,N_8315);
or U8359 (N_8359,N_8309,N_8236);
nor U8360 (N_8360,N_8307,N_8238);
nand U8361 (N_8361,N_8189,N_8292);
nor U8362 (N_8362,N_8213,N_8205);
xnor U8363 (N_8363,N_8215,N_8310);
or U8364 (N_8364,N_8161,N_8221);
and U8365 (N_8365,N_8229,N_8218);
and U8366 (N_8366,N_8241,N_8313);
and U8367 (N_8367,N_8267,N_8237);
nor U8368 (N_8368,N_8188,N_8170);
nor U8369 (N_8369,N_8316,N_8182);
nand U8370 (N_8370,N_8314,N_8181);
nand U8371 (N_8371,N_8318,N_8271);
nor U8372 (N_8372,N_8255,N_8285);
and U8373 (N_8373,N_8283,N_8175);
xor U8374 (N_8374,N_8199,N_8268);
or U8375 (N_8375,N_8183,N_8200);
nor U8376 (N_8376,N_8280,N_8223);
and U8377 (N_8377,N_8209,N_8244);
nand U8378 (N_8378,N_8276,N_8264);
nor U8379 (N_8379,N_8230,N_8286);
nand U8380 (N_8380,N_8174,N_8166);
or U8381 (N_8381,N_8295,N_8277);
or U8382 (N_8382,N_8216,N_8211);
nor U8383 (N_8383,N_8235,N_8171);
and U8384 (N_8384,N_8214,N_8180);
nand U8385 (N_8385,N_8312,N_8306);
nor U8386 (N_8386,N_8266,N_8262);
nand U8387 (N_8387,N_8162,N_8179);
or U8388 (N_8388,N_8298,N_8160);
and U8389 (N_8389,N_8168,N_8208);
or U8390 (N_8390,N_8279,N_8291);
nor U8391 (N_8391,N_8258,N_8231);
and U8392 (N_8392,N_8203,N_8302);
or U8393 (N_8393,N_8190,N_8275);
and U8394 (N_8394,N_8219,N_8207);
or U8395 (N_8395,N_8163,N_8226);
and U8396 (N_8396,N_8250,N_8196);
nor U8397 (N_8397,N_8167,N_8274);
nor U8398 (N_8398,N_8249,N_8202);
or U8399 (N_8399,N_8225,N_8187);
or U8400 (N_8400,N_8181,N_8228);
and U8401 (N_8401,N_8267,N_8319);
nor U8402 (N_8402,N_8241,N_8300);
nor U8403 (N_8403,N_8248,N_8211);
and U8404 (N_8404,N_8168,N_8298);
nand U8405 (N_8405,N_8173,N_8304);
or U8406 (N_8406,N_8313,N_8169);
nand U8407 (N_8407,N_8178,N_8284);
or U8408 (N_8408,N_8237,N_8245);
or U8409 (N_8409,N_8239,N_8292);
or U8410 (N_8410,N_8313,N_8275);
and U8411 (N_8411,N_8310,N_8210);
nor U8412 (N_8412,N_8160,N_8213);
and U8413 (N_8413,N_8266,N_8250);
nor U8414 (N_8414,N_8186,N_8273);
or U8415 (N_8415,N_8216,N_8236);
nand U8416 (N_8416,N_8184,N_8217);
or U8417 (N_8417,N_8254,N_8207);
nor U8418 (N_8418,N_8251,N_8161);
nor U8419 (N_8419,N_8300,N_8200);
and U8420 (N_8420,N_8244,N_8161);
and U8421 (N_8421,N_8283,N_8245);
and U8422 (N_8422,N_8245,N_8313);
or U8423 (N_8423,N_8229,N_8274);
nor U8424 (N_8424,N_8301,N_8226);
and U8425 (N_8425,N_8277,N_8310);
or U8426 (N_8426,N_8260,N_8186);
xnor U8427 (N_8427,N_8281,N_8249);
or U8428 (N_8428,N_8301,N_8206);
nor U8429 (N_8429,N_8207,N_8248);
nand U8430 (N_8430,N_8298,N_8179);
nand U8431 (N_8431,N_8316,N_8279);
and U8432 (N_8432,N_8263,N_8228);
or U8433 (N_8433,N_8191,N_8182);
nand U8434 (N_8434,N_8266,N_8207);
nor U8435 (N_8435,N_8232,N_8276);
or U8436 (N_8436,N_8269,N_8204);
and U8437 (N_8437,N_8250,N_8309);
nand U8438 (N_8438,N_8224,N_8199);
or U8439 (N_8439,N_8233,N_8240);
nand U8440 (N_8440,N_8309,N_8195);
and U8441 (N_8441,N_8228,N_8234);
or U8442 (N_8442,N_8214,N_8252);
nand U8443 (N_8443,N_8266,N_8300);
or U8444 (N_8444,N_8222,N_8207);
and U8445 (N_8445,N_8205,N_8227);
nand U8446 (N_8446,N_8238,N_8197);
xor U8447 (N_8447,N_8246,N_8286);
nand U8448 (N_8448,N_8174,N_8203);
nand U8449 (N_8449,N_8210,N_8245);
nor U8450 (N_8450,N_8240,N_8209);
nand U8451 (N_8451,N_8279,N_8210);
or U8452 (N_8452,N_8198,N_8241);
or U8453 (N_8453,N_8275,N_8199);
nor U8454 (N_8454,N_8204,N_8208);
and U8455 (N_8455,N_8204,N_8237);
xnor U8456 (N_8456,N_8204,N_8264);
nor U8457 (N_8457,N_8270,N_8187);
and U8458 (N_8458,N_8266,N_8316);
or U8459 (N_8459,N_8198,N_8174);
nand U8460 (N_8460,N_8270,N_8164);
nor U8461 (N_8461,N_8212,N_8263);
nor U8462 (N_8462,N_8223,N_8267);
nor U8463 (N_8463,N_8252,N_8182);
xnor U8464 (N_8464,N_8233,N_8251);
nand U8465 (N_8465,N_8248,N_8206);
nand U8466 (N_8466,N_8231,N_8161);
nand U8467 (N_8467,N_8281,N_8186);
and U8468 (N_8468,N_8266,N_8236);
and U8469 (N_8469,N_8209,N_8313);
and U8470 (N_8470,N_8236,N_8286);
nand U8471 (N_8471,N_8219,N_8235);
nand U8472 (N_8472,N_8182,N_8160);
or U8473 (N_8473,N_8307,N_8181);
or U8474 (N_8474,N_8281,N_8228);
xnor U8475 (N_8475,N_8304,N_8169);
and U8476 (N_8476,N_8258,N_8298);
nand U8477 (N_8477,N_8275,N_8262);
nor U8478 (N_8478,N_8168,N_8314);
nand U8479 (N_8479,N_8291,N_8284);
and U8480 (N_8480,N_8358,N_8333);
or U8481 (N_8481,N_8321,N_8331);
and U8482 (N_8482,N_8478,N_8356);
and U8483 (N_8483,N_8441,N_8396);
or U8484 (N_8484,N_8459,N_8369);
and U8485 (N_8485,N_8407,N_8432);
nor U8486 (N_8486,N_8472,N_8352);
nand U8487 (N_8487,N_8389,N_8341);
and U8488 (N_8488,N_8421,N_8347);
nand U8489 (N_8489,N_8422,N_8397);
nand U8490 (N_8490,N_8391,N_8473);
nand U8491 (N_8491,N_8433,N_8360);
nor U8492 (N_8492,N_8332,N_8458);
nor U8493 (N_8493,N_8354,N_8345);
nor U8494 (N_8494,N_8336,N_8376);
nor U8495 (N_8495,N_8357,N_8320);
or U8496 (N_8496,N_8329,N_8443);
and U8497 (N_8497,N_8477,N_8334);
or U8498 (N_8498,N_8380,N_8339);
nor U8499 (N_8499,N_8465,N_8470);
nand U8500 (N_8500,N_8420,N_8335);
or U8501 (N_8501,N_8424,N_8383);
and U8502 (N_8502,N_8471,N_8476);
and U8503 (N_8503,N_8322,N_8330);
nor U8504 (N_8504,N_8463,N_8327);
or U8505 (N_8505,N_8323,N_8381);
and U8506 (N_8506,N_8403,N_8337);
nor U8507 (N_8507,N_8415,N_8457);
nor U8508 (N_8508,N_8361,N_8419);
and U8509 (N_8509,N_8435,N_8338);
or U8510 (N_8510,N_8417,N_8446);
nor U8511 (N_8511,N_8359,N_8467);
or U8512 (N_8512,N_8384,N_8449);
and U8513 (N_8513,N_8426,N_8429);
nand U8514 (N_8514,N_8448,N_8344);
or U8515 (N_8515,N_8427,N_8372);
nand U8516 (N_8516,N_8410,N_8442);
and U8517 (N_8517,N_8371,N_8438);
nand U8518 (N_8518,N_8366,N_8343);
nor U8519 (N_8519,N_8453,N_8405);
nand U8520 (N_8520,N_8423,N_8393);
nand U8521 (N_8521,N_8464,N_8439);
and U8522 (N_8522,N_8370,N_8466);
and U8523 (N_8523,N_8346,N_8411);
and U8524 (N_8524,N_8456,N_8428);
nor U8525 (N_8525,N_8474,N_8414);
nor U8526 (N_8526,N_8382,N_8388);
and U8527 (N_8527,N_8390,N_8402);
or U8528 (N_8528,N_8368,N_8454);
nand U8529 (N_8529,N_8349,N_8436);
nor U8530 (N_8530,N_8374,N_8412);
nor U8531 (N_8531,N_8434,N_8401);
nor U8532 (N_8532,N_8469,N_8462);
nor U8533 (N_8533,N_8406,N_8378);
nor U8534 (N_8534,N_8364,N_8395);
nor U8535 (N_8535,N_8425,N_8461);
or U8536 (N_8536,N_8387,N_8386);
nand U8537 (N_8537,N_8375,N_8479);
and U8538 (N_8538,N_8440,N_8418);
nand U8539 (N_8539,N_8394,N_8365);
and U8540 (N_8540,N_8409,N_8431);
or U8541 (N_8541,N_8398,N_8437);
and U8542 (N_8542,N_8362,N_8385);
and U8543 (N_8543,N_8416,N_8324);
or U8544 (N_8544,N_8326,N_8367);
nand U8545 (N_8545,N_8451,N_8377);
or U8546 (N_8546,N_8447,N_8400);
nor U8547 (N_8547,N_8430,N_8353);
and U8548 (N_8548,N_8404,N_8452);
nor U8549 (N_8549,N_8350,N_8399);
nor U8550 (N_8550,N_8325,N_8348);
nand U8551 (N_8551,N_8460,N_8328);
xnor U8552 (N_8552,N_8413,N_8455);
nor U8553 (N_8553,N_8408,N_8468);
xor U8554 (N_8554,N_8342,N_8379);
nor U8555 (N_8555,N_8392,N_8450);
nor U8556 (N_8556,N_8355,N_8363);
nor U8557 (N_8557,N_8340,N_8444);
xor U8558 (N_8558,N_8351,N_8445);
nand U8559 (N_8559,N_8373,N_8475);
or U8560 (N_8560,N_8363,N_8364);
and U8561 (N_8561,N_8360,N_8445);
nand U8562 (N_8562,N_8457,N_8465);
nor U8563 (N_8563,N_8333,N_8355);
nand U8564 (N_8564,N_8340,N_8441);
nor U8565 (N_8565,N_8387,N_8322);
or U8566 (N_8566,N_8379,N_8334);
nor U8567 (N_8567,N_8478,N_8375);
nor U8568 (N_8568,N_8420,N_8373);
or U8569 (N_8569,N_8472,N_8353);
xor U8570 (N_8570,N_8347,N_8431);
nor U8571 (N_8571,N_8430,N_8377);
or U8572 (N_8572,N_8470,N_8383);
nor U8573 (N_8573,N_8375,N_8433);
or U8574 (N_8574,N_8352,N_8431);
nand U8575 (N_8575,N_8444,N_8332);
nand U8576 (N_8576,N_8346,N_8336);
nand U8577 (N_8577,N_8323,N_8424);
nand U8578 (N_8578,N_8424,N_8433);
and U8579 (N_8579,N_8356,N_8391);
and U8580 (N_8580,N_8333,N_8339);
nor U8581 (N_8581,N_8383,N_8435);
nor U8582 (N_8582,N_8445,N_8424);
and U8583 (N_8583,N_8448,N_8321);
xnor U8584 (N_8584,N_8475,N_8429);
or U8585 (N_8585,N_8418,N_8420);
and U8586 (N_8586,N_8476,N_8470);
xnor U8587 (N_8587,N_8325,N_8327);
xnor U8588 (N_8588,N_8413,N_8380);
nor U8589 (N_8589,N_8375,N_8441);
and U8590 (N_8590,N_8475,N_8381);
and U8591 (N_8591,N_8442,N_8452);
or U8592 (N_8592,N_8478,N_8398);
or U8593 (N_8593,N_8395,N_8342);
and U8594 (N_8594,N_8420,N_8371);
nor U8595 (N_8595,N_8479,N_8438);
or U8596 (N_8596,N_8354,N_8392);
and U8597 (N_8597,N_8478,N_8376);
or U8598 (N_8598,N_8376,N_8433);
and U8599 (N_8599,N_8404,N_8461);
nand U8600 (N_8600,N_8351,N_8426);
or U8601 (N_8601,N_8414,N_8340);
xor U8602 (N_8602,N_8395,N_8386);
nor U8603 (N_8603,N_8363,N_8396);
nor U8604 (N_8604,N_8410,N_8321);
and U8605 (N_8605,N_8329,N_8336);
nand U8606 (N_8606,N_8404,N_8372);
or U8607 (N_8607,N_8367,N_8435);
nand U8608 (N_8608,N_8331,N_8468);
nand U8609 (N_8609,N_8478,N_8429);
xor U8610 (N_8610,N_8387,N_8412);
nor U8611 (N_8611,N_8345,N_8321);
and U8612 (N_8612,N_8418,N_8465);
nor U8613 (N_8613,N_8479,N_8345);
nor U8614 (N_8614,N_8344,N_8386);
xor U8615 (N_8615,N_8460,N_8437);
nor U8616 (N_8616,N_8327,N_8431);
and U8617 (N_8617,N_8414,N_8429);
nand U8618 (N_8618,N_8463,N_8479);
and U8619 (N_8619,N_8430,N_8370);
or U8620 (N_8620,N_8381,N_8479);
or U8621 (N_8621,N_8415,N_8417);
nand U8622 (N_8622,N_8382,N_8361);
or U8623 (N_8623,N_8409,N_8435);
and U8624 (N_8624,N_8329,N_8333);
and U8625 (N_8625,N_8378,N_8360);
or U8626 (N_8626,N_8396,N_8457);
xor U8627 (N_8627,N_8345,N_8477);
xnor U8628 (N_8628,N_8461,N_8375);
nand U8629 (N_8629,N_8357,N_8463);
nand U8630 (N_8630,N_8323,N_8394);
or U8631 (N_8631,N_8411,N_8351);
xor U8632 (N_8632,N_8414,N_8462);
nor U8633 (N_8633,N_8320,N_8442);
and U8634 (N_8634,N_8322,N_8460);
nor U8635 (N_8635,N_8467,N_8442);
or U8636 (N_8636,N_8460,N_8409);
nand U8637 (N_8637,N_8411,N_8443);
and U8638 (N_8638,N_8461,N_8395);
or U8639 (N_8639,N_8405,N_8449);
or U8640 (N_8640,N_8638,N_8591);
and U8641 (N_8641,N_8511,N_8583);
and U8642 (N_8642,N_8544,N_8553);
nor U8643 (N_8643,N_8513,N_8536);
or U8644 (N_8644,N_8589,N_8611);
nand U8645 (N_8645,N_8519,N_8526);
xor U8646 (N_8646,N_8559,N_8564);
and U8647 (N_8647,N_8541,N_8554);
nand U8648 (N_8648,N_8606,N_8576);
and U8649 (N_8649,N_8532,N_8524);
nor U8650 (N_8650,N_8579,N_8505);
and U8651 (N_8651,N_8530,N_8627);
nor U8652 (N_8652,N_8568,N_8499);
or U8653 (N_8653,N_8613,N_8497);
and U8654 (N_8654,N_8634,N_8484);
or U8655 (N_8655,N_8506,N_8514);
nand U8656 (N_8656,N_8535,N_8572);
nor U8657 (N_8657,N_8542,N_8560);
and U8658 (N_8658,N_8537,N_8493);
and U8659 (N_8659,N_8498,N_8561);
or U8660 (N_8660,N_8490,N_8639);
nand U8661 (N_8661,N_8573,N_8637);
xnor U8662 (N_8662,N_8528,N_8546);
and U8663 (N_8663,N_8616,N_8628);
and U8664 (N_8664,N_8584,N_8580);
and U8665 (N_8665,N_8509,N_8617);
and U8666 (N_8666,N_8630,N_8549);
nand U8667 (N_8667,N_8590,N_8539);
xor U8668 (N_8668,N_8598,N_8522);
nand U8669 (N_8669,N_8480,N_8512);
or U8670 (N_8670,N_8582,N_8609);
nor U8671 (N_8671,N_8552,N_8548);
xnor U8672 (N_8672,N_8501,N_8515);
nor U8673 (N_8673,N_8496,N_8614);
nor U8674 (N_8674,N_8504,N_8588);
nand U8675 (N_8675,N_8543,N_8605);
and U8676 (N_8676,N_8636,N_8608);
nor U8677 (N_8677,N_8551,N_8578);
and U8678 (N_8678,N_8594,N_8500);
nor U8679 (N_8679,N_8596,N_8487);
and U8680 (N_8680,N_8494,N_8565);
nor U8681 (N_8681,N_8557,N_8550);
nand U8682 (N_8682,N_8581,N_8622);
nand U8683 (N_8683,N_8600,N_8597);
nor U8684 (N_8684,N_8486,N_8489);
nand U8685 (N_8685,N_8629,N_8567);
and U8686 (N_8686,N_8623,N_8635);
nor U8687 (N_8687,N_8566,N_8619);
or U8688 (N_8688,N_8621,N_8492);
or U8689 (N_8689,N_8520,N_8604);
or U8690 (N_8690,N_8538,N_8618);
and U8691 (N_8691,N_8586,N_8563);
or U8692 (N_8692,N_8575,N_8488);
nand U8693 (N_8693,N_8593,N_8525);
or U8694 (N_8694,N_8610,N_8485);
and U8695 (N_8695,N_8602,N_8585);
or U8696 (N_8696,N_8508,N_8615);
nand U8697 (N_8697,N_8531,N_8607);
or U8698 (N_8698,N_8603,N_8633);
xnor U8699 (N_8699,N_8555,N_8592);
nor U8700 (N_8700,N_8481,N_8540);
nand U8701 (N_8701,N_8556,N_8545);
nor U8702 (N_8702,N_8495,N_8533);
xnor U8703 (N_8703,N_8507,N_8599);
or U8704 (N_8704,N_8569,N_8631);
nand U8705 (N_8705,N_8517,N_8595);
or U8706 (N_8706,N_8571,N_8518);
nor U8707 (N_8707,N_8626,N_8521);
or U8708 (N_8708,N_8577,N_8624);
and U8709 (N_8709,N_8570,N_8547);
nand U8710 (N_8710,N_8562,N_8558);
xor U8711 (N_8711,N_8510,N_8534);
and U8712 (N_8712,N_8502,N_8483);
or U8713 (N_8713,N_8527,N_8625);
or U8714 (N_8714,N_8523,N_8620);
nor U8715 (N_8715,N_8587,N_8503);
or U8716 (N_8716,N_8632,N_8491);
and U8717 (N_8717,N_8516,N_8601);
nor U8718 (N_8718,N_8482,N_8612);
or U8719 (N_8719,N_8529,N_8574);
or U8720 (N_8720,N_8565,N_8535);
or U8721 (N_8721,N_8569,N_8608);
nand U8722 (N_8722,N_8580,N_8541);
and U8723 (N_8723,N_8617,N_8597);
nand U8724 (N_8724,N_8611,N_8607);
or U8725 (N_8725,N_8586,N_8569);
and U8726 (N_8726,N_8571,N_8497);
or U8727 (N_8727,N_8503,N_8491);
xnor U8728 (N_8728,N_8569,N_8618);
nor U8729 (N_8729,N_8481,N_8578);
and U8730 (N_8730,N_8481,N_8548);
or U8731 (N_8731,N_8580,N_8536);
or U8732 (N_8732,N_8519,N_8550);
and U8733 (N_8733,N_8564,N_8524);
or U8734 (N_8734,N_8616,N_8506);
and U8735 (N_8735,N_8510,N_8558);
nor U8736 (N_8736,N_8617,N_8514);
or U8737 (N_8737,N_8605,N_8537);
nand U8738 (N_8738,N_8513,N_8490);
nand U8739 (N_8739,N_8535,N_8546);
and U8740 (N_8740,N_8513,N_8518);
nor U8741 (N_8741,N_8601,N_8612);
and U8742 (N_8742,N_8519,N_8498);
or U8743 (N_8743,N_8541,N_8602);
nand U8744 (N_8744,N_8579,N_8501);
nand U8745 (N_8745,N_8611,N_8610);
nor U8746 (N_8746,N_8594,N_8617);
nor U8747 (N_8747,N_8575,N_8566);
nand U8748 (N_8748,N_8489,N_8566);
xnor U8749 (N_8749,N_8517,N_8481);
and U8750 (N_8750,N_8628,N_8526);
or U8751 (N_8751,N_8570,N_8618);
nand U8752 (N_8752,N_8497,N_8530);
nor U8753 (N_8753,N_8571,N_8557);
or U8754 (N_8754,N_8515,N_8607);
or U8755 (N_8755,N_8483,N_8525);
nor U8756 (N_8756,N_8492,N_8584);
or U8757 (N_8757,N_8614,N_8622);
nor U8758 (N_8758,N_8590,N_8584);
and U8759 (N_8759,N_8602,N_8603);
or U8760 (N_8760,N_8637,N_8513);
nand U8761 (N_8761,N_8622,N_8506);
and U8762 (N_8762,N_8482,N_8503);
and U8763 (N_8763,N_8528,N_8638);
or U8764 (N_8764,N_8551,N_8572);
nor U8765 (N_8765,N_8505,N_8585);
nand U8766 (N_8766,N_8580,N_8506);
nor U8767 (N_8767,N_8607,N_8630);
or U8768 (N_8768,N_8601,N_8563);
nor U8769 (N_8769,N_8496,N_8559);
nand U8770 (N_8770,N_8608,N_8583);
nand U8771 (N_8771,N_8618,N_8562);
or U8772 (N_8772,N_8555,N_8604);
and U8773 (N_8773,N_8515,N_8563);
or U8774 (N_8774,N_8550,N_8634);
nor U8775 (N_8775,N_8480,N_8491);
nand U8776 (N_8776,N_8631,N_8517);
nor U8777 (N_8777,N_8560,N_8532);
nor U8778 (N_8778,N_8581,N_8557);
and U8779 (N_8779,N_8488,N_8506);
nor U8780 (N_8780,N_8541,N_8510);
or U8781 (N_8781,N_8523,N_8623);
and U8782 (N_8782,N_8583,N_8482);
xor U8783 (N_8783,N_8608,N_8502);
or U8784 (N_8784,N_8489,N_8508);
and U8785 (N_8785,N_8507,N_8555);
and U8786 (N_8786,N_8613,N_8636);
nor U8787 (N_8787,N_8592,N_8632);
nor U8788 (N_8788,N_8560,N_8581);
nor U8789 (N_8789,N_8597,N_8615);
and U8790 (N_8790,N_8515,N_8579);
nand U8791 (N_8791,N_8559,N_8527);
nand U8792 (N_8792,N_8534,N_8507);
nand U8793 (N_8793,N_8564,N_8555);
or U8794 (N_8794,N_8500,N_8536);
or U8795 (N_8795,N_8531,N_8609);
nor U8796 (N_8796,N_8520,N_8544);
nor U8797 (N_8797,N_8603,N_8595);
nand U8798 (N_8798,N_8550,N_8581);
nor U8799 (N_8799,N_8545,N_8523);
nand U8800 (N_8800,N_8743,N_8678);
nand U8801 (N_8801,N_8784,N_8796);
or U8802 (N_8802,N_8715,N_8696);
nand U8803 (N_8803,N_8730,N_8707);
or U8804 (N_8804,N_8684,N_8718);
or U8805 (N_8805,N_8733,N_8661);
nor U8806 (N_8806,N_8685,N_8657);
and U8807 (N_8807,N_8665,N_8735);
and U8808 (N_8808,N_8770,N_8689);
or U8809 (N_8809,N_8782,N_8656);
or U8810 (N_8810,N_8728,N_8680);
nor U8811 (N_8811,N_8671,N_8791);
and U8812 (N_8812,N_8788,N_8721);
nand U8813 (N_8813,N_8729,N_8754);
or U8814 (N_8814,N_8737,N_8642);
nand U8815 (N_8815,N_8768,N_8764);
and U8816 (N_8816,N_8759,N_8790);
nor U8817 (N_8817,N_8753,N_8792);
nand U8818 (N_8818,N_8644,N_8786);
nor U8819 (N_8819,N_8726,N_8663);
and U8820 (N_8820,N_8700,N_8652);
or U8821 (N_8821,N_8745,N_8758);
or U8822 (N_8822,N_8653,N_8709);
or U8823 (N_8823,N_8769,N_8761);
xor U8824 (N_8824,N_8668,N_8712);
or U8825 (N_8825,N_8698,N_8778);
nor U8826 (N_8826,N_8708,N_8767);
or U8827 (N_8827,N_8722,N_8738);
and U8828 (N_8828,N_8673,N_8748);
nor U8829 (N_8829,N_8724,N_8780);
or U8830 (N_8830,N_8752,N_8762);
xnor U8831 (N_8831,N_8777,N_8731);
nand U8832 (N_8832,N_8659,N_8691);
nor U8833 (N_8833,N_8772,N_8765);
nor U8834 (N_8834,N_8694,N_8719);
nor U8835 (N_8835,N_8740,N_8676);
xnor U8836 (N_8836,N_8785,N_8714);
nor U8837 (N_8837,N_8679,N_8697);
xor U8838 (N_8838,N_8686,N_8775);
nor U8839 (N_8839,N_8797,N_8674);
nor U8840 (N_8840,N_8682,N_8706);
or U8841 (N_8841,N_8749,N_8744);
or U8842 (N_8842,N_8732,N_8787);
or U8843 (N_8843,N_8757,N_8720);
or U8844 (N_8844,N_8773,N_8692);
nor U8845 (N_8845,N_8670,N_8660);
nand U8846 (N_8846,N_8646,N_8643);
and U8847 (N_8847,N_8739,N_8667);
nor U8848 (N_8848,N_8725,N_8746);
and U8849 (N_8849,N_8723,N_8742);
and U8850 (N_8850,N_8693,N_8675);
xor U8851 (N_8851,N_8771,N_8690);
xnor U8852 (N_8852,N_8799,N_8717);
nor U8853 (N_8853,N_8783,N_8766);
xor U8854 (N_8854,N_8755,N_8760);
nand U8855 (N_8855,N_8649,N_8640);
nor U8856 (N_8856,N_8713,N_8751);
and U8857 (N_8857,N_8798,N_8672);
nand U8858 (N_8858,N_8641,N_8664);
nand U8859 (N_8859,N_8650,N_8794);
nand U8860 (N_8860,N_8711,N_8704);
and U8861 (N_8861,N_8756,N_8716);
or U8862 (N_8862,N_8687,N_8747);
or U8863 (N_8863,N_8699,N_8795);
xor U8864 (N_8864,N_8793,N_8648);
or U8865 (N_8865,N_8734,N_8774);
nand U8866 (N_8866,N_8645,N_8781);
nand U8867 (N_8867,N_8702,N_8776);
or U8868 (N_8868,N_8677,N_8727);
or U8869 (N_8869,N_8763,N_8658);
and U8870 (N_8870,N_8695,N_8741);
xor U8871 (N_8871,N_8779,N_8750);
or U8872 (N_8872,N_8662,N_8666);
or U8873 (N_8873,N_8705,N_8647);
nor U8874 (N_8874,N_8651,N_8688);
or U8875 (N_8875,N_8654,N_8701);
nand U8876 (N_8876,N_8710,N_8736);
nand U8877 (N_8877,N_8789,N_8655);
and U8878 (N_8878,N_8703,N_8669);
nor U8879 (N_8879,N_8683,N_8681);
or U8880 (N_8880,N_8787,N_8665);
nor U8881 (N_8881,N_8674,N_8675);
and U8882 (N_8882,N_8741,N_8694);
nor U8883 (N_8883,N_8745,N_8670);
or U8884 (N_8884,N_8761,N_8731);
and U8885 (N_8885,N_8736,N_8715);
and U8886 (N_8886,N_8721,N_8640);
nor U8887 (N_8887,N_8785,N_8731);
xor U8888 (N_8888,N_8741,N_8792);
or U8889 (N_8889,N_8762,N_8793);
xnor U8890 (N_8890,N_8756,N_8745);
and U8891 (N_8891,N_8754,N_8721);
nand U8892 (N_8892,N_8686,N_8742);
xnor U8893 (N_8893,N_8673,N_8782);
xnor U8894 (N_8894,N_8769,N_8684);
or U8895 (N_8895,N_8793,N_8728);
and U8896 (N_8896,N_8779,N_8759);
or U8897 (N_8897,N_8715,N_8758);
nor U8898 (N_8898,N_8680,N_8780);
nor U8899 (N_8899,N_8785,N_8784);
or U8900 (N_8900,N_8734,N_8658);
or U8901 (N_8901,N_8717,N_8751);
and U8902 (N_8902,N_8683,N_8655);
or U8903 (N_8903,N_8656,N_8643);
nor U8904 (N_8904,N_8765,N_8761);
xor U8905 (N_8905,N_8640,N_8704);
or U8906 (N_8906,N_8757,N_8779);
or U8907 (N_8907,N_8745,N_8688);
nand U8908 (N_8908,N_8713,N_8680);
and U8909 (N_8909,N_8705,N_8750);
and U8910 (N_8910,N_8782,N_8722);
nor U8911 (N_8911,N_8703,N_8705);
nand U8912 (N_8912,N_8701,N_8780);
nand U8913 (N_8913,N_8717,N_8741);
xor U8914 (N_8914,N_8678,N_8776);
and U8915 (N_8915,N_8694,N_8658);
and U8916 (N_8916,N_8665,N_8717);
nor U8917 (N_8917,N_8784,N_8724);
or U8918 (N_8918,N_8750,N_8661);
or U8919 (N_8919,N_8746,N_8662);
and U8920 (N_8920,N_8774,N_8733);
xnor U8921 (N_8921,N_8641,N_8694);
nand U8922 (N_8922,N_8719,N_8764);
nand U8923 (N_8923,N_8667,N_8733);
nand U8924 (N_8924,N_8767,N_8741);
and U8925 (N_8925,N_8756,N_8784);
nand U8926 (N_8926,N_8754,N_8702);
and U8927 (N_8927,N_8674,N_8713);
nor U8928 (N_8928,N_8705,N_8663);
or U8929 (N_8929,N_8645,N_8785);
or U8930 (N_8930,N_8659,N_8727);
nand U8931 (N_8931,N_8677,N_8739);
and U8932 (N_8932,N_8705,N_8699);
and U8933 (N_8933,N_8657,N_8699);
and U8934 (N_8934,N_8643,N_8798);
or U8935 (N_8935,N_8674,N_8728);
xor U8936 (N_8936,N_8684,N_8661);
and U8937 (N_8937,N_8776,N_8723);
and U8938 (N_8938,N_8766,N_8650);
xor U8939 (N_8939,N_8641,N_8768);
nor U8940 (N_8940,N_8752,N_8655);
xor U8941 (N_8941,N_8703,N_8666);
nand U8942 (N_8942,N_8793,N_8714);
or U8943 (N_8943,N_8696,N_8706);
or U8944 (N_8944,N_8682,N_8677);
xnor U8945 (N_8945,N_8773,N_8687);
or U8946 (N_8946,N_8752,N_8765);
nor U8947 (N_8947,N_8754,N_8783);
or U8948 (N_8948,N_8772,N_8684);
nor U8949 (N_8949,N_8771,N_8731);
nand U8950 (N_8950,N_8750,N_8717);
and U8951 (N_8951,N_8713,N_8694);
nand U8952 (N_8952,N_8647,N_8764);
or U8953 (N_8953,N_8766,N_8716);
nand U8954 (N_8954,N_8752,N_8649);
or U8955 (N_8955,N_8774,N_8671);
nor U8956 (N_8956,N_8795,N_8731);
nor U8957 (N_8957,N_8673,N_8728);
and U8958 (N_8958,N_8674,N_8748);
nand U8959 (N_8959,N_8659,N_8796);
nor U8960 (N_8960,N_8959,N_8806);
or U8961 (N_8961,N_8833,N_8835);
nand U8962 (N_8962,N_8898,N_8818);
nand U8963 (N_8963,N_8927,N_8946);
or U8964 (N_8964,N_8951,N_8876);
nand U8965 (N_8965,N_8885,N_8873);
nand U8966 (N_8966,N_8883,N_8940);
nor U8967 (N_8967,N_8903,N_8936);
nor U8968 (N_8968,N_8801,N_8888);
nand U8969 (N_8969,N_8842,N_8813);
and U8970 (N_8970,N_8911,N_8919);
and U8971 (N_8971,N_8906,N_8934);
xnor U8972 (N_8972,N_8908,N_8923);
or U8973 (N_8973,N_8848,N_8823);
or U8974 (N_8974,N_8874,N_8808);
xor U8975 (N_8975,N_8939,N_8872);
nor U8976 (N_8976,N_8916,N_8831);
nand U8977 (N_8977,N_8922,N_8825);
nand U8978 (N_8978,N_8944,N_8953);
and U8979 (N_8979,N_8947,N_8847);
and U8980 (N_8980,N_8879,N_8851);
nor U8981 (N_8981,N_8859,N_8819);
nand U8982 (N_8982,N_8935,N_8932);
and U8983 (N_8983,N_8834,N_8810);
or U8984 (N_8984,N_8845,N_8817);
xor U8985 (N_8985,N_8832,N_8836);
nor U8986 (N_8986,N_8933,N_8804);
and U8987 (N_8987,N_8850,N_8956);
and U8988 (N_8988,N_8913,N_8802);
nor U8989 (N_8989,N_8899,N_8941);
nor U8990 (N_8990,N_8943,N_8849);
nand U8991 (N_8991,N_8928,N_8877);
or U8992 (N_8992,N_8867,N_8924);
nand U8993 (N_8993,N_8895,N_8920);
and U8994 (N_8994,N_8861,N_8829);
or U8995 (N_8995,N_8881,N_8875);
nor U8996 (N_8996,N_8826,N_8930);
nand U8997 (N_8997,N_8809,N_8958);
nor U8998 (N_8998,N_8840,N_8871);
xnor U8999 (N_8999,N_8917,N_8821);
and U9000 (N_9000,N_8815,N_8830);
or U9001 (N_9001,N_8907,N_8901);
xnor U9002 (N_9002,N_8870,N_8828);
xnor U9003 (N_9003,N_8905,N_8878);
or U9004 (N_9004,N_8814,N_8957);
and U9005 (N_9005,N_8889,N_8822);
nor U9006 (N_9006,N_8918,N_8909);
and U9007 (N_9007,N_8827,N_8904);
or U9008 (N_9008,N_8914,N_8915);
and U9009 (N_9009,N_8890,N_8893);
nand U9010 (N_9010,N_8884,N_8857);
or U9011 (N_9011,N_8816,N_8955);
nand U9012 (N_9012,N_8852,N_8843);
nand U9013 (N_9013,N_8805,N_8931);
xnor U9014 (N_9014,N_8950,N_8837);
and U9015 (N_9015,N_8948,N_8860);
nor U9016 (N_9016,N_8902,N_8812);
and U9017 (N_9017,N_8900,N_8938);
nor U9018 (N_9018,N_8844,N_8891);
and U9019 (N_9019,N_8866,N_8886);
nand U9020 (N_9020,N_8811,N_8942);
and U9021 (N_9021,N_8807,N_8862);
nor U9022 (N_9022,N_8869,N_8952);
nand U9023 (N_9023,N_8868,N_8863);
and U9024 (N_9024,N_8882,N_8838);
or U9025 (N_9025,N_8954,N_8864);
or U9026 (N_9026,N_8824,N_8839);
and U9027 (N_9027,N_8846,N_8820);
and U9028 (N_9028,N_8910,N_8926);
or U9029 (N_9029,N_8892,N_8803);
nor U9030 (N_9030,N_8937,N_8841);
or U9031 (N_9031,N_8925,N_8858);
and U9032 (N_9032,N_8897,N_8945);
nor U9033 (N_9033,N_8912,N_8887);
xnor U9034 (N_9034,N_8880,N_8896);
or U9035 (N_9035,N_8854,N_8853);
nand U9036 (N_9036,N_8894,N_8856);
or U9037 (N_9037,N_8929,N_8855);
and U9038 (N_9038,N_8865,N_8921);
nor U9039 (N_9039,N_8949,N_8800);
and U9040 (N_9040,N_8938,N_8876);
xor U9041 (N_9041,N_8878,N_8902);
and U9042 (N_9042,N_8889,N_8948);
nand U9043 (N_9043,N_8831,N_8837);
nor U9044 (N_9044,N_8952,N_8950);
or U9045 (N_9045,N_8864,N_8875);
and U9046 (N_9046,N_8956,N_8939);
nor U9047 (N_9047,N_8852,N_8875);
nor U9048 (N_9048,N_8880,N_8805);
or U9049 (N_9049,N_8870,N_8861);
xor U9050 (N_9050,N_8837,N_8955);
and U9051 (N_9051,N_8801,N_8924);
nand U9052 (N_9052,N_8880,N_8901);
and U9053 (N_9053,N_8828,N_8837);
and U9054 (N_9054,N_8832,N_8885);
nor U9055 (N_9055,N_8941,N_8868);
or U9056 (N_9056,N_8955,N_8833);
or U9057 (N_9057,N_8929,N_8924);
or U9058 (N_9058,N_8924,N_8847);
and U9059 (N_9059,N_8805,N_8845);
and U9060 (N_9060,N_8946,N_8938);
xor U9061 (N_9061,N_8924,N_8932);
and U9062 (N_9062,N_8855,N_8875);
and U9063 (N_9063,N_8917,N_8849);
nor U9064 (N_9064,N_8863,N_8917);
nand U9065 (N_9065,N_8873,N_8903);
nor U9066 (N_9066,N_8863,N_8840);
nor U9067 (N_9067,N_8872,N_8811);
and U9068 (N_9068,N_8824,N_8936);
and U9069 (N_9069,N_8813,N_8924);
and U9070 (N_9070,N_8927,N_8923);
and U9071 (N_9071,N_8938,N_8958);
nor U9072 (N_9072,N_8938,N_8853);
nand U9073 (N_9073,N_8870,N_8805);
nor U9074 (N_9074,N_8885,N_8934);
nand U9075 (N_9075,N_8898,N_8827);
or U9076 (N_9076,N_8835,N_8943);
or U9077 (N_9077,N_8878,N_8861);
and U9078 (N_9078,N_8884,N_8830);
or U9079 (N_9079,N_8930,N_8911);
or U9080 (N_9080,N_8888,N_8826);
and U9081 (N_9081,N_8812,N_8838);
or U9082 (N_9082,N_8959,N_8926);
or U9083 (N_9083,N_8943,N_8845);
xnor U9084 (N_9084,N_8849,N_8873);
and U9085 (N_9085,N_8881,N_8948);
or U9086 (N_9086,N_8903,N_8842);
and U9087 (N_9087,N_8915,N_8816);
xnor U9088 (N_9088,N_8880,N_8833);
nor U9089 (N_9089,N_8877,N_8954);
xor U9090 (N_9090,N_8893,N_8814);
nor U9091 (N_9091,N_8934,N_8889);
or U9092 (N_9092,N_8808,N_8938);
or U9093 (N_9093,N_8957,N_8901);
and U9094 (N_9094,N_8845,N_8816);
and U9095 (N_9095,N_8885,N_8926);
nand U9096 (N_9096,N_8836,N_8953);
nor U9097 (N_9097,N_8919,N_8861);
nor U9098 (N_9098,N_8841,N_8811);
or U9099 (N_9099,N_8801,N_8900);
nand U9100 (N_9100,N_8948,N_8854);
and U9101 (N_9101,N_8804,N_8856);
or U9102 (N_9102,N_8832,N_8877);
and U9103 (N_9103,N_8952,N_8919);
or U9104 (N_9104,N_8924,N_8862);
nand U9105 (N_9105,N_8947,N_8955);
and U9106 (N_9106,N_8831,N_8848);
xnor U9107 (N_9107,N_8856,N_8854);
and U9108 (N_9108,N_8942,N_8863);
or U9109 (N_9109,N_8832,N_8870);
nor U9110 (N_9110,N_8941,N_8940);
xnor U9111 (N_9111,N_8846,N_8807);
or U9112 (N_9112,N_8873,N_8914);
nor U9113 (N_9113,N_8807,N_8928);
xor U9114 (N_9114,N_8904,N_8916);
or U9115 (N_9115,N_8896,N_8865);
or U9116 (N_9116,N_8852,N_8921);
xor U9117 (N_9117,N_8861,N_8897);
nand U9118 (N_9118,N_8857,N_8851);
or U9119 (N_9119,N_8811,N_8883);
nand U9120 (N_9120,N_9119,N_8976);
nand U9121 (N_9121,N_9004,N_8965);
or U9122 (N_9122,N_9083,N_9063);
xnor U9123 (N_9123,N_9074,N_8991);
and U9124 (N_9124,N_9085,N_9017);
nor U9125 (N_9125,N_9094,N_9009);
or U9126 (N_9126,N_9064,N_9003);
and U9127 (N_9127,N_9087,N_9072);
nand U9128 (N_9128,N_9099,N_9026);
xor U9129 (N_9129,N_9065,N_9061);
or U9130 (N_9130,N_9024,N_9035);
nor U9131 (N_9131,N_8994,N_9034);
nand U9132 (N_9132,N_9092,N_9014);
nor U9133 (N_9133,N_9104,N_9047);
nor U9134 (N_9134,N_9098,N_8997);
nand U9135 (N_9135,N_9091,N_9013);
or U9136 (N_9136,N_9048,N_8970);
nand U9137 (N_9137,N_9078,N_9005);
nand U9138 (N_9138,N_9059,N_9033);
nand U9139 (N_9139,N_9050,N_8975);
or U9140 (N_9140,N_9067,N_8966);
nand U9141 (N_9141,N_9027,N_9023);
nor U9142 (N_9142,N_9012,N_8978);
and U9143 (N_9143,N_9053,N_8990);
nor U9144 (N_9144,N_8983,N_9028);
or U9145 (N_9145,N_9041,N_9022);
or U9146 (N_9146,N_9036,N_9062);
and U9147 (N_9147,N_9018,N_9114);
nor U9148 (N_9148,N_9032,N_8977);
and U9149 (N_9149,N_9040,N_9068);
and U9150 (N_9150,N_8973,N_9110);
nor U9151 (N_9151,N_9029,N_9102);
nor U9152 (N_9152,N_8963,N_8999);
nor U9153 (N_9153,N_9118,N_9069);
nor U9154 (N_9154,N_9019,N_9007);
or U9155 (N_9155,N_9039,N_9037);
nor U9156 (N_9156,N_8968,N_9051);
nor U9157 (N_9157,N_9093,N_8972);
and U9158 (N_9158,N_9105,N_8998);
or U9159 (N_9159,N_8981,N_9044);
and U9160 (N_9160,N_8988,N_9060);
nor U9161 (N_9161,N_9115,N_8960);
xnor U9162 (N_9162,N_9021,N_9077);
and U9163 (N_9163,N_9076,N_9080);
nor U9164 (N_9164,N_9000,N_9052);
or U9165 (N_9165,N_9073,N_8979);
or U9166 (N_9166,N_8986,N_9006);
or U9167 (N_9167,N_9016,N_9055);
nor U9168 (N_9168,N_9109,N_9046);
and U9169 (N_9169,N_9001,N_9108);
or U9170 (N_9170,N_9075,N_9057);
and U9171 (N_9171,N_8992,N_9038);
nand U9172 (N_9172,N_9031,N_8967);
nor U9173 (N_9173,N_9106,N_8980);
or U9174 (N_9174,N_9010,N_8993);
nand U9175 (N_9175,N_9112,N_9086);
and U9176 (N_9176,N_9043,N_9030);
nand U9177 (N_9177,N_9111,N_8962);
xor U9178 (N_9178,N_9071,N_9103);
xnor U9179 (N_9179,N_9095,N_8995);
and U9180 (N_9180,N_8987,N_9117);
nand U9181 (N_9181,N_8984,N_9042);
nand U9182 (N_9182,N_9020,N_9015);
nand U9183 (N_9183,N_8964,N_9049);
and U9184 (N_9184,N_8969,N_9008);
and U9185 (N_9185,N_9054,N_8982);
nor U9186 (N_9186,N_9070,N_8961);
xnor U9187 (N_9187,N_9089,N_8989);
nor U9188 (N_9188,N_9088,N_8971);
and U9189 (N_9189,N_9081,N_9082);
or U9190 (N_9190,N_9058,N_9025);
nor U9191 (N_9191,N_9100,N_9097);
and U9192 (N_9192,N_9045,N_8985);
or U9193 (N_9193,N_9002,N_9090);
nor U9194 (N_9194,N_8996,N_9113);
or U9195 (N_9195,N_9116,N_9011);
nand U9196 (N_9196,N_9101,N_9096);
xor U9197 (N_9197,N_9079,N_9056);
nand U9198 (N_9198,N_9066,N_8974);
and U9199 (N_9199,N_9107,N_9084);
nor U9200 (N_9200,N_9084,N_9051);
nor U9201 (N_9201,N_8995,N_9014);
xnor U9202 (N_9202,N_9021,N_9034);
xnor U9203 (N_9203,N_9066,N_9097);
or U9204 (N_9204,N_9078,N_8964);
and U9205 (N_9205,N_9075,N_8990);
nor U9206 (N_9206,N_9038,N_9095);
nor U9207 (N_9207,N_9109,N_8995);
nand U9208 (N_9208,N_8998,N_9053);
nor U9209 (N_9209,N_9104,N_9054);
nand U9210 (N_9210,N_8980,N_9043);
or U9211 (N_9211,N_9107,N_8978);
and U9212 (N_9212,N_8987,N_9015);
or U9213 (N_9213,N_9049,N_9099);
nor U9214 (N_9214,N_9083,N_9034);
nand U9215 (N_9215,N_9048,N_8997);
or U9216 (N_9216,N_8980,N_9099);
and U9217 (N_9217,N_9098,N_9106);
xnor U9218 (N_9218,N_9012,N_9058);
nor U9219 (N_9219,N_8963,N_9044);
or U9220 (N_9220,N_9081,N_9009);
xnor U9221 (N_9221,N_9102,N_8982);
nand U9222 (N_9222,N_9040,N_9060);
nand U9223 (N_9223,N_9029,N_9107);
and U9224 (N_9224,N_9016,N_9044);
xnor U9225 (N_9225,N_9058,N_9076);
or U9226 (N_9226,N_9036,N_9099);
nor U9227 (N_9227,N_9016,N_8982);
nand U9228 (N_9228,N_9093,N_8991);
and U9229 (N_9229,N_9063,N_9098);
and U9230 (N_9230,N_9004,N_9027);
or U9231 (N_9231,N_9037,N_8989);
and U9232 (N_9232,N_9018,N_8961);
and U9233 (N_9233,N_9071,N_9075);
or U9234 (N_9234,N_9090,N_9035);
nand U9235 (N_9235,N_8974,N_9059);
nor U9236 (N_9236,N_8991,N_9062);
nor U9237 (N_9237,N_9024,N_9089);
or U9238 (N_9238,N_8992,N_9092);
nand U9239 (N_9239,N_9060,N_9097);
and U9240 (N_9240,N_8960,N_8975);
nand U9241 (N_9241,N_8964,N_9037);
and U9242 (N_9242,N_8993,N_8975);
nor U9243 (N_9243,N_8978,N_8984);
nand U9244 (N_9244,N_9018,N_9087);
and U9245 (N_9245,N_9085,N_9079);
xor U9246 (N_9246,N_9111,N_9108);
nand U9247 (N_9247,N_9018,N_9092);
or U9248 (N_9248,N_9053,N_9064);
nand U9249 (N_9249,N_9104,N_9030);
nor U9250 (N_9250,N_9114,N_9020);
nand U9251 (N_9251,N_8991,N_9046);
and U9252 (N_9252,N_9119,N_9101);
xor U9253 (N_9253,N_9035,N_9057);
nor U9254 (N_9254,N_8975,N_9062);
nor U9255 (N_9255,N_9002,N_9104);
or U9256 (N_9256,N_9054,N_9112);
nand U9257 (N_9257,N_9052,N_8996);
nor U9258 (N_9258,N_8999,N_9043);
nand U9259 (N_9259,N_9084,N_9035);
nand U9260 (N_9260,N_9067,N_9044);
nor U9261 (N_9261,N_9081,N_9020);
nand U9262 (N_9262,N_9116,N_9039);
xor U9263 (N_9263,N_8982,N_9096);
xor U9264 (N_9264,N_9086,N_9027);
and U9265 (N_9265,N_9069,N_9051);
nand U9266 (N_9266,N_9046,N_8973);
nand U9267 (N_9267,N_9016,N_9008);
and U9268 (N_9268,N_8981,N_8985);
and U9269 (N_9269,N_9099,N_9111);
xnor U9270 (N_9270,N_9022,N_8962);
or U9271 (N_9271,N_9012,N_8994);
nand U9272 (N_9272,N_9030,N_9113);
nand U9273 (N_9273,N_8961,N_9026);
nand U9274 (N_9274,N_8978,N_9101);
and U9275 (N_9275,N_9007,N_8993);
or U9276 (N_9276,N_8985,N_9046);
nand U9277 (N_9277,N_8961,N_8993);
nand U9278 (N_9278,N_9011,N_8997);
nand U9279 (N_9279,N_9069,N_9015);
xnor U9280 (N_9280,N_9184,N_9270);
or U9281 (N_9281,N_9141,N_9228);
nor U9282 (N_9282,N_9159,N_9259);
and U9283 (N_9283,N_9220,N_9276);
and U9284 (N_9284,N_9191,N_9164);
nor U9285 (N_9285,N_9150,N_9193);
xor U9286 (N_9286,N_9267,N_9277);
nor U9287 (N_9287,N_9134,N_9173);
or U9288 (N_9288,N_9176,N_9133);
xnor U9289 (N_9289,N_9252,N_9246);
nand U9290 (N_9290,N_9204,N_9138);
and U9291 (N_9291,N_9123,N_9129);
nor U9292 (N_9292,N_9120,N_9236);
nor U9293 (N_9293,N_9131,N_9275);
nand U9294 (N_9294,N_9180,N_9253);
xnor U9295 (N_9295,N_9168,N_9222);
nand U9296 (N_9296,N_9249,N_9187);
and U9297 (N_9297,N_9240,N_9251);
or U9298 (N_9298,N_9254,N_9132);
or U9299 (N_9299,N_9231,N_9210);
nand U9300 (N_9300,N_9189,N_9219);
nor U9301 (N_9301,N_9188,N_9221);
and U9302 (N_9302,N_9271,N_9167);
and U9303 (N_9303,N_9166,N_9195);
and U9304 (N_9304,N_9146,N_9147);
and U9305 (N_9305,N_9160,N_9215);
or U9306 (N_9306,N_9234,N_9243);
xnor U9307 (N_9307,N_9199,N_9257);
nor U9308 (N_9308,N_9239,N_9128);
or U9309 (N_9309,N_9157,N_9190);
nor U9310 (N_9310,N_9121,N_9248);
and U9311 (N_9311,N_9196,N_9261);
nor U9312 (N_9312,N_9125,N_9126);
or U9313 (N_9313,N_9136,N_9181);
and U9314 (N_9314,N_9200,N_9237);
and U9315 (N_9315,N_9272,N_9172);
or U9316 (N_9316,N_9163,N_9124);
and U9317 (N_9317,N_9233,N_9211);
nand U9318 (N_9318,N_9244,N_9177);
or U9319 (N_9319,N_9192,N_9137);
nor U9320 (N_9320,N_9212,N_9202);
or U9321 (N_9321,N_9245,N_9214);
and U9322 (N_9322,N_9274,N_9151);
nor U9323 (N_9323,N_9207,N_9279);
nor U9324 (N_9324,N_9266,N_9135);
and U9325 (N_9325,N_9148,N_9127);
or U9326 (N_9326,N_9155,N_9232);
and U9327 (N_9327,N_9256,N_9226);
or U9328 (N_9328,N_9224,N_9158);
nand U9329 (N_9329,N_9258,N_9227);
and U9330 (N_9330,N_9186,N_9264);
xor U9331 (N_9331,N_9229,N_9153);
or U9332 (N_9332,N_9218,N_9242);
nor U9333 (N_9333,N_9169,N_9223);
xor U9334 (N_9334,N_9152,N_9241);
nor U9335 (N_9335,N_9262,N_9198);
or U9336 (N_9336,N_9206,N_9143);
and U9337 (N_9337,N_9268,N_9156);
xnor U9338 (N_9338,N_9260,N_9205);
and U9339 (N_9339,N_9144,N_9235);
nand U9340 (N_9340,N_9140,N_9273);
xor U9341 (N_9341,N_9209,N_9247);
or U9342 (N_9342,N_9255,N_9175);
nor U9343 (N_9343,N_9154,N_9183);
nor U9344 (N_9344,N_9197,N_9217);
and U9345 (N_9345,N_9225,N_9278);
nor U9346 (N_9346,N_9208,N_9178);
nand U9347 (N_9347,N_9216,N_9250);
nor U9348 (N_9348,N_9165,N_9142);
nand U9349 (N_9349,N_9149,N_9122);
nand U9350 (N_9350,N_9203,N_9230);
or U9351 (N_9351,N_9185,N_9265);
or U9352 (N_9352,N_9182,N_9170);
and U9353 (N_9353,N_9269,N_9238);
xnor U9354 (N_9354,N_9174,N_9213);
nor U9355 (N_9355,N_9162,N_9171);
or U9356 (N_9356,N_9201,N_9161);
nand U9357 (N_9357,N_9139,N_9145);
or U9358 (N_9358,N_9263,N_9194);
nand U9359 (N_9359,N_9130,N_9179);
or U9360 (N_9360,N_9177,N_9228);
or U9361 (N_9361,N_9231,N_9266);
and U9362 (N_9362,N_9263,N_9228);
nand U9363 (N_9363,N_9191,N_9204);
nand U9364 (N_9364,N_9252,N_9265);
nand U9365 (N_9365,N_9243,N_9210);
and U9366 (N_9366,N_9120,N_9194);
and U9367 (N_9367,N_9222,N_9125);
and U9368 (N_9368,N_9158,N_9149);
and U9369 (N_9369,N_9274,N_9244);
nor U9370 (N_9370,N_9227,N_9159);
xor U9371 (N_9371,N_9227,N_9238);
and U9372 (N_9372,N_9277,N_9204);
and U9373 (N_9373,N_9270,N_9254);
nor U9374 (N_9374,N_9140,N_9162);
and U9375 (N_9375,N_9214,N_9247);
xor U9376 (N_9376,N_9276,N_9124);
and U9377 (N_9377,N_9266,N_9236);
and U9378 (N_9378,N_9134,N_9123);
and U9379 (N_9379,N_9192,N_9218);
xor U9380 (N_9380,N_9194,N_9142);
or U9381 (N_9381,N_9122,N_9279);
nand U9382 (N_9382,N_9252,N_9247);
and U9383 (N_9383,N_9273,N_9242);
nor U9384 (N_9384,N_9231,N_9279);
and U9385 (N_9385,N_9252,N_9139);
nand U9386 (N_9386,N_9242,N_9134);
nand U9387 (N_9387,N_9206,N_9178);
nand U9388 (N_9388,N_9270,N_9152);
nand U9389 (N_9389,N_9253,N_9132);
nor U9390 (N_9390,N_9133,N_9121);
xor U9391 (N_9391,N_9133,N_9267);
nor U9392 (N_9392,N_9130,N_9164);
nor U9393 (N_9393,N_9189,N_9218);
nor U9394 (N_9394,N_9131,N_9174);
and U9395 (N_9395,N_9181,N_9133);
xor U9396 (N_9396,N_9269,N_9276);
xor U9397 (N_9397,N_9138,N_9146);
or U9398 (N_9398,N_9151,N_9271);
nor U9399 (N_9399,N_9192,N_9252);
or U9400 (N_9400,N_9261,N_9191);
nand U9401 (N_9401,N_9241,N_9227);
or U9402 (N_9402,N_9191,N_9165);
nand U9403 (N_9403,N_9256,N_9252);
nand U9404 (N_9404,N_9251,N_9163);
or U9405 (N_9405,N_9170,N_9211);
xor U9406 (N_9406,N_9244,N_9148);
or U9407 (N_9407,N_9239,N_9210);
or U9408 (N_9408,N_9214,N_9257);
nor U9409 (N_9409,N_9150,N_9206);
or U9410 (N_9410,N_9132,N_9194);
and U9411 (N_9411,N_9140,N_9124);
or U9412 (N_9412,N_9265,N_9276);
and U9413 (N_9413,N_9211,N_9190);
or U9414 (N_9414,N_9191,N_9170);
nor U9415 (N_9415,N_9234,N_9179);
nand U9416 (N_9416,N_9120,N_9260);
or U9417 (N_9417,N_9259,N_9215);
nand U9418 (N_9418,N_9209,N_9264);
nor U9419 (N_9419,N_9259,N_9235);
or U9420 (N_9420,N_9191,N_9161);
or U9421 (N_9421,N_9125,N_9156);
and U9422 (N_9422,N_9122,N_9262);
xor U9423 (N_9423,N_9197,N_9263);
xnor U9424 (N_9424,N_9154,N_9220);
or U9425 (N_9425,N_9241,N_9171);
or U9426 (N_9426,N_9224,N_9195);
or U9427 (N_9427,N_9248,N_9256);
and U9428 (N_9428,N_9264,N_9151);
nand U9429 (N_9429,N_9163,N_9150);
xor U9430 (N_9430,N_9152,N_9150);
or U9431 (N_9431,N_9251,N_9174);
or U9432 (N_9432,N_9151,N_9141);
and U9433 (N_9433,N_9156,N_9279);
and U9434 (N_9434,N_9202,N_9270);
xor U9435 (N_9435,N_9154,N_9215);
xnor U9436 (N_9436,N_9224,N_9263);
nor U9437 (N_9437,N_9220,N_9172);
or U9438 (N_9438,N_9132,N_9162);
nand U9439 (N_9439,N_9139,N_9233);
nand U9440 (N_9440,N_9339,N_9299);
or U9441 (N_9441,N_9414,N_9307);
and U9442 (N_9442,N_9431,N_9347);
and U9443 (N_9443,N_9311,N_9303);
nand U9444 (N_9444,N_9387,N_9429);
xor U9445 (N_9445,N_9306,N_9320);
nor U9446 (N_9446,N_9390,N_9432);
nor U9447 (N_9447,N_9365,N_9406);
or U9448 (N_9448,N_9329,N_9349);
nand U9449 (N_9449,N_9368,N_9425);
and U9450 (N_9450,N_9340,N_9395);
nor U9451 (N_9451,N_9435,N_9430);
and U9452 (N_9452,N_9384,N_9400);
nor U9453 (N_9453,N_9287,N_9391);
or U9454 (N_9454,N_9294,N_9379);
nor U9455 (N_9455,N_9316,N_9330);
nand U9456 (N_9456,N_9410,N_9351);
or U9457 (N_9457,N_9293,N_9312);
or U9458 (N_9458,N_9416,N_9439);
xnor U9459 (N_9459,N_9280,N_9381);
or U9460 (N_9460,N_9359,N_9282);
nand U9461 (N_9461,N_9413,N_9399);
nor U9462 (N_9462,N_9362,N_9319);
and U9463 (N_9463,N_9367,N_9314);
xnor U9464 (N_9464,N_9412,N_9385);
and U9465 (N_9465,N_9376,N_9427);
nor U9466 (N_9466,N_9315,N_9372);
nor U9467 (N_9467,N_9345,N_9296);
xor U9468 (N_9468,N_9428,N_9389);
and U9469 (N_9469,N_9334,N_9356);
or U9470 (N_9470,N_9378,N_9301);
nor U9471 (N_9471,N_9373,N_9404);
nor U9472 (N_9472,N_9408,N_9352);
nor U9473 (N_9473,N_9392,N_9289);
nor U9474 (N_9474,N_9417,N_9333);
nor U9475 (N_9475,N_9342,N_9292);
or U9476 (N_9476,N_9341,N_9353);
xnor U9477 (N_9477,N_9300,N_9302);
nor U9478 (N_9478,N_9360,N_9394);
and U9479 (N_9479,N_9371,N_9332);
nand U9480 (N_9480,N_9369,N_9322);
and U9481 (N_9481,N_9363,N_9323);
nand U9482 (N_9482,N_9426,N_9366);
or U9483 (N_9483,N_9398,N_9438);
nand U9484 (N_9484,N_9325,N_9423);
xor U9485 (N_9485,N_9421,N_9411);
xnor U9486 (N_9486,N_9328,N_9281);
nand U9487 (N_9487,N_9317,N_9326);
nand U9488 (N_9488,N_9375,N_9338);
and U9489 (N_9489,N_9324,N_9321);
nor U9490 (N_9490,N_9419,N_9437);
nand U9491 (N_9491,N_9364,N_9424);
nand U9492 (N_9492,N_9377,N_9386);
nand U9493 (N_9493,N_9388,N_9433);
nor U9494 (N_9494,N_9357,N_9361);
and U9495 (N_9495,N_9331,N_9290);
nor U9496 (N_9496,N_9397,N_9420);
or U9497 (N_9497,N_9284,N_9337);
and U9498 (N_9498,N_9374,N_9313);
and U9499 (N_9499,N_9310,N_9355);
and U9500 (N_9500,N_9396,N_9350);
or U9501 (N_9501,N_9436,N_9327);
xnor U9502 (N_9502,N_9415,N_9422);
or U9503 (N_9503,N_9407,N_9402);
nand U9504 (N_9504,N_9358,N_9295);
or U9505 (N_9505,N_9335,N_9297);
nor U9506 (N_9506,N_9285,N_9383);
nand U9507 (N_9507,N_9346,N_9336);
nor U9508 (N_9508,N_9403,N_9418);
and U9509 (N_9509,N_9298,N_9288);
and U9510 (N_9510,N_9309,N_9305);
or U9511 (N_9511,N_9434,N_9380);
and U9512 (N_9512,N_9405,N_9308);
nor U9513 (N_9513,N_9283,N_9401);
or U9514 (N_9514,N_9343,N_9354);
nor U9515 (N_9515,N_9286,N_9370);
or U9516 (N_9516,N_9393,N_9382);
nand U9517 (N_9517,N_9409,N_9318);
xor U9518 (N_9518,N_9344,N_9348);
nor U9519 (N_9519,N_9304,N_9291);
nand U9520 (N_9520,N_9379,N_9366);
nand U9521 (N_9521,N_9394,N_9289);
nor U9522 (N_9522,N_9352,N_9359);
or U9523 (N_9523,N_9420,N_9356);
or U9524 (N_9524,N_9369,N_9423);
and U9525 (N_9525,N_9381,N_9335);
or U9526 (N_9526,N_9412,N_9384);
nand U9527 (N_9527,N_9349,N_9295);
or U9528 (N_9528,N_9393,N_9311);
and U9529 (N_9529,N_9327,N_9386);
nand U9530 (N_9530,N_9421,N_9399);
or U9531 (N_9531,N_9383,N_9409);
nor U9532 (N_9532,N_9423,N_9342);
nor U9533 (N_9533,N_9395,N_9414);
nor U9534 (N_9534,N_9428,N_9366);
and U9535 (N_9535,N_9315,N_9439);
and U9536 (N_9536,N_9378,N_9374);
or U9537 (N_9537,N_9322,N_9357);
nand U9538 (N_9538,N_9428,N_9354);
nor U9539 (N_9539,N_9301,N_9310);
nand U9540 (N_9540,N_9296,N_9437);
nand U9541 (N_9541,N_9389,N_9414);
and U9542 (N_9542,N_9338,N_9430);
nand U9543 (N_9543,N_9283,N_9314);
nor U9544 (N_9544,N_9391,N_9288);
or U9545 (N_9545,N_9435,N_9346);
or U9546 (N_9546,N_9429,N_9307);
or U9547 (N_9547,N_9320,N_9395);
and U9548 (N_9548,N_9303,N_9408);
or U9549 (N_9549,N_9372,N_9388);
nor U9550 (N_9550,N_9290,N_9340);
or U9551 (N_9551,N_9355,N_9379);
and U9552 (N_9552,N_9318,N_9361);
or U9553 (N_9553,N_9287,N_9301);
or U9554 (N_9554,N_9280,N_9355);
nand U9555 (N_9555,N_9341,N_9334);
or U9556 (N_9556,N_9430,N_9339);
nor U9557 (N_9557,N_9340,N_9402);
nand U9558 (N_9558,N_9383,N_9323);
nor U9559 (N_9559,N_9407,N_9410);
or U9560 (N_9560,N_9300,N_9376);
nand U9561 (N_9561,N_9333,N_9394);
or U9562 (N_9562,N_9425,N_9350);
nand U9563 (N_9563,N_9326,N_9381);
or U9564 (N_9564,N_9332,N_9381);
and U9565 (N_9565,N_9390,N_9315);
nor U9566 (N_9566,N_9419,N_9408);
and U9567 (N_9567,N_9421,N_9320);
nand U9568 (N_9568,N_9346,N_9399);
and U9569 (N_9569,N_9362,N_9366);
nand U9570 (N_9570,N_9431,N_9342);
nand U9571 (N_9571,N_9372,N_9370);
nand U9572 (N_9572,N_9435,N_9321);
nand U9573 (N_9573,N_9331,N_9330);
or U9574 (N_9574,N_9283,N_9394);
nand U9575 (N_9575,N_9425,N_9347);
nor U9576 (N_9576,N_9329,N_9322);
nor U9577 (N_9577,N_9297,N_9324);
nor U9578 (N_9578,N_9314,N_9417);
nand U9579 (N_9579,N_9428,N_9285);
and U9580 (N_9580,N_9355,N_9343);
and U9581 (N_9581,N_9333,N_9316);
or U9582 (N_9582,N_9295,N_9297);
nor U9583 (N_9583,N_9432,N_9340);
or U9584 (N_9584,N_9410,N_9355);
xnor U9585 (N_9585,N_9380,N_9321);
nand U9586 (N_9586,N_9437,N_9422);
and U9587 (N_9587,N_9379,N_9427);
nor U9588 (N_9588,N_9370,N_9308);
and U9589 (N_9589,N_9393,N_9371);
or U9590 (N_9590,N_9322,N_9318);
and U9591 (N_9591,N_9394,N_9396);
and U9592 (N_9592,N_9355,N_9389);
nor U9593 (N_9593,N_9427,N_9331);
and U9594 (N_9594,N_9333,N_9314);
nand U9595 (N_9595,N_9386,N_9310);
or U9596 (N_9596,N_9291,N_9393);
and U9597 (N_9597,N_9325,N_9320);
and U9598 (N_9598,N_9427,N_9289);
or U9599 (N_9599,N_9416,N_9368);
or U9600 (N_9600,N_9587,N_9462);
nand U9601 (N_9601,N_9487,N_9517);
nor U9602 (N_9602,N_9473,N_9566);
and U9603 (N_9603,N_9533,N_9557);
or U9604 (N_9604,N_9539,N_9505);
nor U9605 (N_9605,N_9463,N_9497);
and U9606 (N_9606,N_9565,N_9447);
xnor U9607 (N_9607,N_9571,N_9537);
or U9608 (N_9608,N_9468,N_9454);
nor U9609 (N_9609,N_9522,N_9508);
and U9610 (N_9610,N_9547,N_9544);
nor U9611 (N_9611,N_9579,N_9569);
nor U9612 (N_9612,N_9501,N_9452);
nor U9613 (N_9613,N_9491,N_9582);
and U9614 (N_9614,N_9549,N_9532);
nor U9615 (N_9615,N_9531,N_9475);
nand U9616 (N_9616,N_9570,N_9445);
nor U9617 (N_9617,N_9558,N_9456);
nor U9618 (N_9618,N_9536,N_9583);
and U9619 (N_9619,N_9498,N_9513);
or U9620 (N_9620,N_9490,N_9478);
nand U9621 (N_9621,N_9576,N_9585);
or U9622 (N_9622,N_9519,N_9460);
nor U9623 (N_9623,N_9524,N_9559);
nand U9624 (N_9624,N_9514,N_9469);
nor U9625 (N_9625,N_9553,N_9472);
and U9626 (N_9626,N_9567,N_9546);
and U9627 (N_9627,N_9467,N_9485);
or U9628 (N_9628,N_9542,N_9563);
xnor U9629 (N_9629,N_9476,N_9444);
or U9630 (N_9630,N_9499,N_9525);
nor U9631 (N_9631,N_9595,N_9592);
and U9632 (N_9632,N_9550,N_9535);
or U9633 (N_9633,N_9593,N_9599);
and U9634 (N_9634,N_9481,N_9448);
nand U9635 (N_9635,N_9459,N_9528);
nor U9636 (N_9636,N_9594,N_9545);
nand U9637 (N_9637,N_9474,N_9502);
nand U9638 (N_9638,N_9560,N_9580);
and U9639 (N_9639,N_9457,N_9450);
nor U9640 (N_9640,N_9561,N_9596);
and U9641 (N_9641,N_9488,N_9584);
nor U9642 (N_9642,N_9458,N_9573);
xor U9643 (N_9643,N_9554,N_9495);
and U9644 (N_9644,N_9449,N_9480);
or U9645 (N_9645,N_9496,N_9464);
and U9646 (N_9646,N_9466,N_9470);
and U9647 (N_9647,N_9518,N_9515);
xor U9648 (N_9648,N_9512,N_9586);
xnor U9649 (N_9649,N_9574,N_9503);
xnor U9650 (N_9650,N_9581,N_9541);
and U9651 (N_9651,N_9465,N_9510);
nand U9652 (N_9652,N_9440,N_9572);
and U9653 (N_9653,N_9493,N_9556);
nand U9654 (N_9654,N_9461,N_9506);
and U9655 (N_9655,N_9504,N_9591);
or U9656 (N_9656,N_9527,N_9486);
and U9657 (N_9657,N_9520,N_9555);
and U9658 (N_9658,N_9455,N_9507);
nand U9659 (N_9659,N_9471,N_9441);
nor U9660 (N_9660,N_9552,N_9484);
nand U9661 (N_9661,N_9538,N_9516);
nor U9662 (N_9662,N_9530,N_9540);
nand U9663 (N_9663,N_9494,N_9575);
and U9664 (N_9664,N_9446,N_9551);
or U9665 (N_9665,N_9589,N_9523);
nand U9666 (N_9666,N_9489,N_9500);
or U9667 (N_9667,N_9492,N_9529);
nand U9668 (N_9668,N_9543,N_9598);
and U9669 (N_9669,N_9479,N_9451);
xnor U9670 (N_9670,N_9588,N_9477);
and U9671 (N_9671,N_9482,N_9442);
nor U9672 (N_9672,N_9597,N_9564);
nor U9673 (N_9673,N_9562,N_9511);
or U9674 (N_9674,N_9577,N_9526);
nand U9675 (N_9675,N_9590,N_9534);
nand U9676 (N_9676,N_9453,N_9443);
nor U9677 (N_9677,N_9509,N_9578);
or U9678 (N_9678,N_9568,N_9521);
nor U9679 (N_9679,N_9483,N_9548);
or U9680 (N_9680,N_9582,N_9471);
and U9681 (N_9681,N_9476,N_9578);
and U9682 (N_9682,N_9552,N_9504);
or U9683 (N_9683,N_9542,N_9546);
nor U9684 (N_9684,N_9559,N_9596);
or U9685 (N_9685,N_9556,N_9553);
nand U9686 (N_9686,N_9523,N_9461);
nor U9687 (N_9687,N_9470,N_9593);
or U9688 (N_9688,N_9462,N_9531);
or U9689 (N_9689,N_9571,N_9574);
and U9690 (N_9690,N_9505,N_9551);
nand U9691 (N_9691,N_9503,N_9463);
nand U9692 (N_9692,N_9556,N_9523);
and U9693 (N_9693,N_9490,N_9531);
or U9694 (N_9694,N_9575,N_9448);
xor U9695 (N_9695,N_9531,N_9557);
or U9696 (N_9696,N_9502,N_9446);
nor U9697 (N_9697,N_9510,N_9491);
nor U9698 (N_9698,N_9577,N_9544);
or U9699 (N_9699,N_9577,N_9585);
xnor U9700 (N_9700,N_9466,N_9555);
nand U9701 (N_9701,N_9448,N_9478);
nand U9702 (N_9702,N_9578,N_9555);
nand U9703 (N_9703,N_9559,N_9494);
or U9704 (N_9704,N_9585,N_9572);
nand U9705 (N_9705,N_9487,N_9528);
xor U9706 (N_9706,N_9591,N_9596);
or U9707 (N_9707,N_9450,N_9476);
or U9708 (N_9708,N_9519,N_9459);
nand U9709 (N_9709,N_9596,N_9461);
and U9710 (N_9710,N_9501,N_9514);
nand U9711 (N_9711,N_9553,N_9495);
nor U9712 (N_9712,N_9572,N_9478);
nor U9713 (N_9713,N_9462,N_9444);
xor U9714 (N_9714,N_9512,N_9505);
or U9715 (N_9715,N_9455,N_9501);
and U9716 (N_9716,N_9492,N_9454);
or U9717 (N_9717,N_9551,N_9444);
nor U9718 (N_9718,N_9541,N_9569);
nand U9719 (N_9719,N_9541,N_9550);
nor U9720 (N_9720,N_9467,N_9594);
xor U9721 (N_9721,N_9575,N_9499);
and U9722 (N_9722,N_9592,N_9487);
nor U9723 (N_9723,N_9456,N_9539);
or U9724 (N_9724,N_9526,N_9498);
xor U9725 (N_9725,N_9562,N_9513);
xnor U9726 (N_9726,N_9547,N_9451);
nor U9727 (N_9727,N_9550,N_9467);
and U9728 (N_9728,N_9548,N_9552);
and U9729 (N_9729,N_9441,N_9458);
or U9730 (N_9730,N_9519,N_9569);
or U9731 (N_9731,N_9489,N_9581);
or U9732 (N_9732,N_9453,N_9595);
and U9733 (N_9733,N_9490,N_9450);
nor U9734 (N_9734,N_9574,N_9584);
or U9735 (N_9735,N_9499,N_9479);
nand U9736 (N_9736,N_9524,N_9554);
nand U9737 (N_9737,N_9576,N_9441);
and U9738 (N_9738,N_9484,N_9553);
and U9739 (N_9739,N_9582,N_9585);
xnor U9740 (N_9740,N_9570,N_9496);
xor U9741 (N_9741,N_9475,N_9508);
nor U9742 (N_9742,N_9451,N_9513);
xnor U9743 (N_9743,N_9519,N_9587);
nor U9744 (N_9744,N_9582,N_9520);
and U9745 (N_9745,N_9465,N_9460);
and U9746 (N_9746,N_9457,N_9488);
nor U9747 (N_9747,N_9498,N_9587);
and U9748 (N_9748,N_9559,N_9501);
and U9749 (N_9749,N_9530,N_9458);
nand U9750 (N_9750,N_9506,N_9523);
and U9751 (N_9751,N_9553,N_9456);
xor U9752 (N_9752,N_9566,N_9492);
nand U9753 (N_9753,N_9478,N_9522);
and U9754 (N_9754,N_9555,N_9553);
or U9755 (N_9755,N_9593,N_9477);
and U9756 (N_9756,N_9499,N_9573);
and U9757 (N_9757,N_9486,N_9517);
xor U9758 (N_9758,N_9532,N_9452);
xnor U9759 (N_9759,N_9585,N_9454);
nand U9760 (N_9760,N_9677,N_9667);
and U9761 (N_9761,N_9687,N_9620);
and U9762 (N_9762,N_9695,N_9665);
nand U9763 (N_9763,N_9756,N_9745);
or U9764 (N_9764,N_9672,N_9607);
or U9765 (N_9765,N_9726,N_9635);
xnor U9766 (N_9766,N_9755,N_9746);
or U9767 (N_9767,N_9738,N_9713);
nor U9768 (N_9768,N_9628,N_9660);
nor U9769 (N_9769,N_9697,N_9643);
nor U9770 (N_9770,N_9706,N_9751);
or U9771 (N_9771,N_9669,N_9729);
or U9772 (N_9772,N_9601,N_9703);
and U9773 (N_9773,N_9685,N_9614);
and U9774 (N_9774,N_9615,N_9683);
nor U9775 (N_9775,N_9624,N_9630);
or U9776 (N_9776,N_9720,N_9722);
xnor U9777 (N_9777,N_9693,N_9647);
nor U9778 (N_9778,N_9639,N_9602);
nand U9779 (N_9779,N_9757,N_9719);
nor U9780 (N_9780,N_9725,N_9676);
nor U9781 (N_9781,N_9690,N_9734);
or U9782 (N_9782,N_9735,N_9705);
xnor U9783 (N_9783,N_9711,N_9600);
and U9784 (N_9784,N_9727,N_9623);
xor U9785 (N_9785,N_9750,N_9724);
or U9786 (N_9786,N_9721,N_9717);
nand U9787 (N_9787,N_9652,N_9758);
or U9788 (N_9788,N_9646,N_9655);
xnor U9789 (N_9789,N_9642,N_9648);
nor U9790 (N_9790,N_9694,N_9673);
nand U9791 (N_9791,N_9744,N_9638);
and U9792 (N_9792,N_9662,N_9731);
nand U9793 (N_9793,N_9653,N_9641);
nand U9794 (N_9794,N_9644,N_9736);
nor U9795 (N_9795,N_9686,N_9688);
and U9796 (N_9796,N_9730,N_9748);
or U9797 (N_9797,N_9710,N_9753);
and U9798 (N_9798,N_9664,N_9625);
nand U9799 (N_9799,N_9609,N_9743);
and U9800 (N_9800,N_9631,N_9671);
nor U9801 (N_9801,N_9627,N_9732);
and U9802 (N_9802,N_9741,N_9759);
nor U9803 (N_9803,N_9709,N_9696);
nor U9804 (N_9804,N_9700,N_9604);
or U9805 (N_9805,N_9659,N_9684);
or U9806 (N_9806,N_9714,N_9608);
nor U9807 (N_9807,N_9728,N_9613);
nand U9808 (N_9808,N_9610,N_9658);
xnor U9809 (N_9809,N_9712,N_9715);
or U9810 (N_9810,N_9621,N_9708);
nand U9811 (N_9811,N_9619,N_9702);
nand U9812 (N_9812,N_9618,N_9739);
or U9813 (N_9813,N_9689,N_9692);
nor U9814 (N_9814,N_9632,N_9645);
or U9815 (N_9815,N_9606,N_9723);
xor U9816 (N_9816,N_9707,N_9740);
xor U9817 (N_9817,N_9661,N_9651);
xnor U9818 (N_9818,N_9634,N_9636);
nand U9819 (N_9819,N_9611,N_9656);
or U9820 (N_9820,N_9640,N_9699);
nand U9821 (N_9821,N_9678,N_9650);
xor U9822 (N_9822,N_9612,N_9718);
nand U9823 (N_9823,N_9616,N_9637);
and U9824 (N_9824,N_9622,N_9754);
or U9825 (N_9825,N_9674,N_9679);
and U9826 (N_9826,N_9675,N_9704);
or U9827 (N_9827,N_9663,N_9749);
or U9828 (N_9828,N_9742,N_9654);
xor U9829 (N_9829,N_9698,N_9680);
and U9830 (N_9830,N_9605,N_9670);
nand U9831 (N_9831,N_9649,N_9716);
and U9832 (N_9832,N_9733,N_9629);
nor U9833 (N_9833,N_9668,N_9657);
nand U9834 (N_9834,N_9681,N_9752);
or U9835 (N_9835,N_9603,N_9633);
or U9836 (N_9836,N_9691,N_9666);
or U9837 (N_9837,N_9737,N_9747);
or U9838 (N_9838,N_9701,N_9626);
nand U9839 (N_9839,N_9617,N_9682);
and U9840 (N_9840,N_9753,N_9676);
nor U9841 (N_9841,N_9662,N_9739);
or U9842 (N_9842,N_9733,N_9623);
or U9843 (N_9843,N_9717,N_9680);
nand U9844 (N_9844,N_9603,N_9754);
nor U9845 (N_9845,N_9724,N_9700);
and U9846 (N_9846,N_9621,N_9731);
and U9847 (N_9847,N_9625,N_9611);
nand U9848 (N_9848,N_9657,N_9694);
nand U9849 (N_9849,N_9703,N_9704);
nand U9850 (N_9850,N_9654,N_9753);
xor U9851 (N_9851,N_9750,N_9748);
nand U9852 (N_9852,N_9748,N_9693);
and U9853 (N_9853,N_9625,N_9754);
and U9854 (N_9854,N_9725,N_9753);
nand U9855 (N_9855,N_9676,N_9708);
and U9856 (N_9856,N_9721,N_9660);
or U9857 (N_9857,N_9607,N_9754);
nand U9858 (N_9858,N_9645,N_9662);
nor U9859 (N_9859,N_9631,N_9668);
or U9860 (N_9860,N_9666,N_9746);
nand U9861 (N_9861,N_9678,N_9626);
or U9862 (N_9862,N_9652,N_9722);
and U9863 (N_9863,N_9651,N_9694);
xnor U9864 (N_9864,N_9690,N_9600);
nand U9865 (N_9865,N_9614,N_9670);
or U9866 (N_9866,N_9754,N_9651);
nor U9867 (N_9867,N_9708,N_9601);
and U9868 (N_9868,N_9693,N_9630);
and U9869 (N_9869,N_9658,N_9687);
and U9870 (N_9870,N_9628,N_9704);
or U9871 (N_9871,N_9717,N_9730);
nor U9872 (N_9872,N_9647,N_9726);
or U9873 (N_9873,N_9702,N_9698);
and U9874 (N_9874,N_9647,N_9678);
xnor U9875 (N_9875,N_9647,N_9759);
nor U9876 (N_9876,N_9701,N_9728);
and U9877 (N_9877,N_9687,N_9603);
and U9878 (N_9878,N_9600,N_9705);
nor U9879 (N_9879,N_9757,N_9645);
and U9880 (N_9880,N_9657,N_9759);
or U9881 (N_9881,N_9672,N_9679);
or U9882 (N_9882,N_9704,N_9706);
nor U9883 (N_9883,N_9745,N_9737);
nand U9884 (N_9884,N_9644,N_9632);
nor U9885 (N_9885,N_9742,N_9687);
and U9886 (N_9886,N_9680,N_9688);
xnor U9887 (N_9887,N_9641,N_9673);
xnor U9888 (N_9888,N_9713,N_9714);
or U9889 (N_9889,N_9643,N_9719);
nor U9890 (N_9890,N_9756,N_9656);
or U9891 (N_9891,N_9724,N_9630);
or U9892 (N_9892,N_9707,N_9709);
or U9893 (N_9893,N_9669,N_9656);
and U9894 (N_9894,N_9627,N_9625);
nand U9895 (N_9895,N_9663,N_9685);
nand U9896 (N_9896,N_9680,N_9676);
xor U9897 (N_9897,N_9722,N_9703);
or U9898 (N_9898,N_9633,N_9625);
and U9899 (N_9899,N_9615,N_9700);
nand U9900 (N_9900,N_9743,N_9624);
nor U9901 (N_9901,N_9638,N_9694);
nor U9902 (N_9902,N_9747,N_9686);
nor U9903 (N_9903,N_9706,N_9671);
or U9904 (N_9904,N_9699,N_9737);
nor U9905 (N_9905,N_9691,N_9645);
and U9906 (N_9906,N_9627,N_9633);
or U9907 (N_9907,N_9618,N_9651);
nor U9908 (N_9908,N_9759,N_9708);
nand U9909 (N_9909,N_9736,N_9727);
and U9910 (N_9910,N_9607,N_9634);
or U9911 (N_9911,N_9648,N_9655);
and U9912 (N_9912,N_9741,N_9636);
and U9913 (N_9913,N_9670,N_9674);
and U9914 (N_9914,N_9603,N_9642);
nor U9915 (N_9915,N_9687,N_9659);
xnor U9916 (N_9916,N_9633,N_9653);
or U9917 (N_9917,N_9727,N_9677);
and U9918 (N_9918,N_9698,N_9625);
nand U9919 (N_9919,N_9603,N_9667);
or U9920 (N_9920,N_9906,N_9802);
nor U9921 (N_9921,N_9790,N_9799);
nand U9922 (N_9922,N_9866,N_9893);
nand U9923 (N_9923,N_9841,N_9899);
xor U9924 (N_9924,N_9872,N_9821);
or U9925 (N_9925,N_9840,N_9912);
or U9926 (N_9926,N_9919,N_9856);
nand U9927 (N_9927,N_9855,N_9845);
or U9928 (N_9928,N_9878,N_9777);
nor U9929 (N_9929,N_9907,N_9886);
nand U9930 (N_9930,N_9787,N_9775);
nand U9931 (N_9931,N_9908,N_9896);
nand U9932 (N_9932,N_9911,N_9818);
nand U9933 (N_9933,N_9887,N_9763);
nand U9934 (N_9934,N_9891,N_9869);
nor U9935 (N_9935,N_9881,N_9794);
or U9936 (N_9936,N_9768,N_9898);
or U9937 (N_9937,N_9762,N_9765);
and U9938 (N_9938,N_9865,N_9864);
or U9939 (N_9939,N_9803,N_9825);
or U9940 (N_9940,N_9782,N_9903);
and U9941 (N_9941,N_9839,N_9834);
or U9942 (N_9942,N_9876,N_9889);
nand U9943 (N_9943,N_9905,N_9868);
and U9944 (N_9944,N_9867,N_9830);
nand U9945 (N_9945,N_9791,N_9861);
or U9946 (N_9946,N_9902,N_9792);
xor U9947 (N_9947,N_9811,N_9764);
xnor U9948 (N_9948,N_9852,N_9854);
nand U9949 (N_9949,N_9850,N_9847);
xnor U9950 (N_9950,N_9895,N_9831);
nor U9951 (N_9951,N_9822,N_9904);
nor U9952 (N_9952,N_9836,N_9781);
or U9953 (N_9953,N_9814,N_9800);
xor U9954 (N_9954,N_9877,N_9813);
xor U9955 (N_9955,N_9873,N_9807);
and U9956 (N_9956,N_9795,N_9892);
or U9957 (N_9957,N_9857,N_9772);
nand U9958 (N_9958,N_9819,N_9894);
and U9959 (N_9959,N_9833,N_9849);
or U9960 (N_9960,N_9914,N_9816);
nor U9961 (N_9961,N_9843,N_9897);
nand U9962 (N_9962,N_9917,N_9785);
nor U9963 (N_9963,N_9766,N_9880);
or U9964 (N_9964,N_9808,N_9783);
nand U9965 (N_9965,N_9801,N_9798);
or U9966 (N_9966,N_9796,N_9817);
nand U9967 (N_9967,N_9890,N_9835);
or U9968 (N_9968,N_9860,N_9773);
and U9969 (N_9969,N_9853,N_9885);
nand U9970 (N_9970,N_9884,N_9842);
nand U9971 (N_9971,N_9760,N_9793);
or U9972 (N_9972,N_9779,N_9915);
nor U9973 (N_9973,N_9870,N_9846);
and U9974 (N_9974,N_9810,N_9784);
and U9975 (N_9975,N_9909,N_9883);
nand U9976 (N_9976,N_9900,N_9875);
or U9977 (N_9977,N_9828,N_9851);
or U9978 (N_9978,N_9859,N_9809);
nand U9979 (N_9979,N_9832,N_9913);
or U9980 (N_9980,N_9826,N_9812);
or U9981 (N_9981,N_9901,N_9806);
xor U9982 (N_9982,N_9882,N_9879);
and U9983 (N_9983,N_9774,N_9804);
nor U9984 (N_9984,N_9888,N_9863);
and U9985 (N_9985,N_9776,N_9788);
xnor U9986 (N_9986,N_9862,N_9910);
nor U9987 (N_9987,N_9829,N_9871);
nor U9988 (N_9988,N_9838,N_9918);
and U9989 (N_9989,N_9797,N_9789);
nor U9990 (N_9990,N_9786,N_9805);
nor U9991 (N_9991,N_9761,N_9767);
nor U9992 (N_9992,N_9824,N_9827);
or U9993 (N_9993,N_9815,N_9820);
and U9994 (N_9994,N_9780,N_9844);
or U9995 (N_9995,N_9769,N_9837);
nor U9996 (N_9996,N_9771,N_9916);
nand U9997 (N_9997,N_9778,N_9770);
or U9998 (N_9998,N_9848,N_9858);
nand U9999 (N_9999,N_9823,N_9874);
nor U10000 (N_10000,N_9843,N_9900);
or U10001 (N_10001,N_9905,N_9852);
xnor U10002 (N_10002,N_9838,N_9817);
nand U10003 (N_10003,N_9881,N_9762);
nor U10004 (N_10004,N_9870,N_9827);
nor U10005 (N_10005,N_9892,N_9797);
xor U10006 (N_10006,N_9855,N_9910);
nor U10007 (N_10007,N_9834,N_9836);
nor U10008 (N_10008,N_9900,N_9822);
and U10009 (N_10009,N_9883,N_9904);
nor U10010 (N_10010,N_9831,N_9911);
or U10011 (N_10011,N_9812,N_9915);
nor U10012 (N_10012,N_9877,N_9887);
or U10013 (N_10013,N_9783,N_9802);
or U10014 (N_10014,N_9871,N_9890);
or U10015 (N_10015,N_9831,N_9883);
or U10016 (N_10016,N_9788,N_9914);
nor U10017 (N_10017,N_9838,N_9785);
xnor U10018 (N_10018,N_9767,N_9901);
nor U10019 (N_10019,N_9874,N_9883);
nand U10020 (N_10020,N_9816,N_9788);
and U10021 (N_10021,N_9882,N_9859);
or U10022 (N_10022,N_9761,N_9891);
xnor U10023 (N_10023,N_9776,N_9821);
or U10024 (N_10024,N_9867,N_9803);
nand U10025 (N_10025,N_9891,N_9786);
nand U10026 (N_10026,N_9790,N_9839);
nand U10027 (N_10027,N_9863,N_9892);
and U10028 (N_10028,N_9808,N_9768);
xor U10029 (N_10029,N_9778,N_9789);
and U10030 (N_10030,N_9771,N_9856);
nor U10031 (N_10031,N_9862,N_9888);
or U10032 (N_10032,N_9765,N_9794);
nor U10033 (N_10033,N_9802,N_9771);
and U10034 (N_10034,N_9795,N_9826);
nand U10035 (N_10035,N_9830,N_9908);
nor U10036 (N_10036,N_9862,N_9828);
nand U10037 (N_10037,N_9779,N_9858);
or U10038 (N_10038,N_9912,N_9872);
and U10039 (N_10039,N_9856,N_9914);
xnor U10040 (N_10040,N_9868,N_9906);
and U10041 (N_10041,N_9783,N_9827);
nand U10042 (N_10042,N_9874,N_9854);
nor U10043 (N_10043,N_9889,N_9856);
nor U10044 (N_10044,N_9852,N_9788);
nor U10045 (N_10045,N_9914,N_9785);
nor U10046 (N_10046,N_9783,N_9909);
or U10047 (N_10047,N_9812,N_9782);
nor U10048 (N_10048,N_9827,N_9848);
nor U10049 (N_10049,N_9818,N_9871);
nand U10050 (N_10050,N_9879,N_9813);
xnor U10051 (N_10051,N_9845,N_9792);
and U10052 (N_10052,N_9866,N_9777);
and U10053 (N_10053,N_9909,N_9885);
nand U10054 (N_10054,N_9806,N_9866);
xor U10055 (N_10055,N_9871,N_9808);
nand U10056 (N_10056,N_9849,N_9909);
and U10057 (N_10057,N_9856,N_9861);
xnor U10058 (N_10058,N_9902,N_9836);
and U10059 (N_10059,N_9835,N_9790);
and U10060 (N_10060,N_9851,N_9791);
nand U10061 (N_10061,N_9770,N_9839);
nor U10062 (N_10062,N_9914,N_9794);
nor U10063 (N_10063,N_9803,N_9864);
nor U10064 (N_10064,N_9911,N_9776);
xor U10065 (N_10065,N_9909,N_9769);
and U10066 (N_10066,N_9791,N_9792);
and U10067 (N_10067,N_9776,N_9877);
and U10068 (N_10068,N_9841,N_9763);
nor U10069 (N_10069,N_9777,N_9915);
nand U10070 (N_10070,N_9896,N_9816);
nor U10071 (N_10071,N_9778,N_9821);
and U10072 (N_10072,N_9804,N_9764);
or U10073 (N_10073,N_9907,N_9911);
nand U10074 (N_10074,N_9812,N_9900);
or U10075 (N_10075,N_9831,N_9809);
nor U10076 (N_10076,N_9884,N_9786);
nor U10077 (N_10077,N_9822,N_9858);
nor U10078 (N_10078,N_9787,N_9805);
and U10079 (N_10079,N_9804,N_9781);
or U10080 (N_10080,N_9952,N_10052);
and U10081 (N_10081,N_10022,N_10007);
nand U10082 (N_10082,N_10029,N_9939);
nand U10083 (N_10083,N_10048,N_10055);
nor U10084 (N_10084,N_10043,N_9936);
nor U10085 (N_10085,N_9924,N_10020);
nor U10086 (N_10086,N_10018,N_9962);
xor U10087 (N_10087,N_10074,N_10041);
and U10088 (N_10088,N_9956,N_9979);
nor U10089 (N_10089,N_10046,N_9923);
xnor U10090 (N_10090,N_10031,N_10069);
nand U10091 (N_10091,N_9934,N_10008);
and U10092 (N_10092,N_9955,N_9959);
and U10093 (N_10093,N_10001,N_10063);
nor U10094 (N_10094,N_9922,N_9988);
or U10095 (N_10095,N_9967,N_9976);
and U10096 (N_10096,N_10030,N_9926);
xnor U10097 (N_10097,N_9930,N_10045);
and U10098 (N_10098,N_9941,N_10054);
nand U10099 (N_10099,N_9965,N_9950);
nor U10100 (N_10100,N_9946,N_10059);
nand U10101 (N_10101,N_9945,N_9961);
nor U10102 (N_10102,N_10068,N_10076);
or U10103 (N_10103,N_9931,N_9929);
nor U10104 (N_10104,N_9994,N_9937);
and U10105 (N_10105,N_10067,N_10010);
nand U10106 (N_10106,N_10003,N_10002);
and U10107 (N_10107,N_9953,N_9987);
xor U10108 (N_10108,N_9932,N_10033);
nor U10109 (N_10109,N_9973,N_10072);
nor U10110 (N_10110,N_10075,N_9982);
nand U10111 (N_10111,N_10040,N_9984);
and U10112 (N_10112,N_10027,N_9938);
nor U10113 (N_10113,N_10026,N_9963);
nor U10114 (N_10114,N_9981,N_10050);
and U10115 (N_10115,N_10024,N_9998);
nand U10116 (N_10116,N_9943,N_9993);
nand U10117 (N_10117,N_10061,N_9971);
nand U10118 (N_10118,N_9978,N_10060);
xor U10119 (N_10119,N_10017,N_9989);
nor U10120 (N_10120,N_9999,N_9997);
nand U10121 (N_10121,N_10051,N_10032);
or U10122 (N_10122,N_9977,N_10047);
nand U10123 (N_10123,N_10070,N_10005);
or U10124 (N_10124,N_10023,N_9957);
nand U10125 (N_10125,N_9972,N_10057);
and U10126 (N_10126,N_10037,N_9940);
or U10127 (N_10127,N_9933,N_10073);
and U10128 (N_10128,N_10035,N_9928);
nor U10129 (N_10129,N_10078,N_10012);
and U10130 (N_10130,N_10066,N_10044);
or U10131 (N_10131,N_9975,N_9958);
and U10132 (N_10132,N_10025,N_9986);
nand U10133 (N_10133,N_9969,N_10011);
nand U10134 (N_10134,N_9985,N_10065);
or U10135 (N_10135,N_10056,N_10053);
xor U10136 (N_10136,N_10000,N_10016);
or U10137 (N_10137,N_10013,N_9935);
nand U10138 (N_10138,N_10042,N_9980);
or U10139 (N_10139,N_9947,N_10028);
and U10140 (N_10140,N_9983,N_10019);
xor U10141 (N_10141,N_9966,N_10014);
nor U10142 (N_10142,N_9920,N_9954);
and U10143 (N_10143,N_9996,N_9995);
or U10144 (N_10144,N_9951,N_10064);
and U10145 (N_10145,N_9944,N_10034);
or U10146 (N_10146,N_10062,N_9948);
or U10147 (N_10147,N_10038,N_9925);
nand U10148 (N_10148,N_9990,N_10036);
nand U10149 (N_10149,N_10015,N_10006);
nand U10150 (N_10150,N_10021,N_9991);
nand U10151 (N_10151,N_10009,N_9927);
nor U10152 (N_10152,N_10039,N_10071);
nand U10153 (N_10153,N_10058,N_9974);
nand U10154 (N_10154,N_9949,N_9921);
or U10155 (N_10155,N_9960,N_9964);
and U10156 (N_10156,N_9968,N_10079);
and U10157 (N_10157,N_10049,N_9970);
nand U10158 (N_10158,N_9942,N_10004);
nand U10159 (N_10159,N_10077,N_9992);
nor U10160 (N_10160,N_9941,N_10070);
or U10161 (N_10161,N_10061,N_9996);
nand U10162 (N_10162,N_9925,N_10042);
and U10163 (N_10163,N_10022,N_9984);
nand U10164 (N_10164,N_9981,N_10059);
and U10165 (N_10165,N_10060,N_9947);
and U10166 (N_10166,N_10041,N_10014);
and U10167 (N_10167,N_9976,N_9998);
or U10168 (N_10168,N_10009,N_10053);
nand U10169 (N_10169,N_9985,N_9937);
nor U10170 (N_10170,N_10006,N_10028);
and U10171 (N_10171,N_10073,N_10048);
xnor U10172 (N_10172,N_9998,N_10049);
xnor U10173 (N_10173,N_9957,N_10055);
xor U10174 (N_10174,N_10073,N_10075);
or U10175 (N_10175,N_9957,N_10078);
and U10176 (N_10176,N_9922,N_9941);
nand U10177 (N_10177,N_10030,N_9944);
or U10178 (N_10178,N_9967,N_10026);
and U10179 (N_10179,N_10039,N_10057);
or U10180 (N_10180,N_10004,N_10064);
nand U10181 (N_10181,N_9983,N_9930);
or U10182 (N_10182,N_9998,N_10068);
nand U10183 (N_10183,N_10074,N_9935);
xnor U10184 (N_10184,N_10036,N_9980);
nand U10185 (N_10185,N_10036,N_9939);
nor U10186 (N_10186,N_9967,N_9970);
or U10187 (N_10187,N_10059,N_10030);
or U10188 (N_10188,N_10064,N_10074);
or U10189 (N_10189,N_10035,N_9974);
nand U10190 (N_10190,N_10051,N_10062);
nor U10191 (N_10191,N_10061,N_10043);
or U10192 (N_10192,N_10011,N_10023);
nor U10193 (N_10193,N_9964,N_9971);
and U10194 (N_10194,N_10023,N_10064);
or U10195 (N_10195,N_9993,N_9992);
nor U10196 (N_10196,N_10073,N_10028);
xor U10197 (N_10197,N_9981,N_10007);
nand U10198 (N_10198,N_9936,N_10071);
nor U10199 (N_10199,N_9993,N_9989);
xor U10200 (N_10200,N_10037,N_9958);
or U10201 (N_10201,N_10038,N_10056);
nor U10202 (N_10202,N_9935,N_10040);
or U10203 (N_10203,N_9950,N_9985);
and U10204 (N_10204,N_10047,N_9920);
xor U10205 (N_10205,N_10008,N_10028);
nand U10206 (N_10206,N_9937,N_9925);
or U10207 (N_10207,N_10000,N_9927);
nand U10208 (N_10208,N_10040,N_9995);
nor U10209 (N_10209,N_9974,N_9971);
or U10210 (N_10210,N_10041,N_10006);
or U10211 (N_10211,N_9975,N_10057);
nor U10212 (N_10212,N_10003,N_10048);
nor U10213 (N_10213,N_9953,N_10067);
and U10214 (N_10214,N_9930,N_9989);
nand U10215 (N_10215,N_9929,N_9927);
nand U10216 (N_10216,N_9964,N_9940);
or U10217 (N_10217,N_10051,N_9995);
xor U10218 (N_10218,N_10036,N_9923);
and U10219 (N_10219,N_9978,N_10035);
nand U10220 (N_10220,N_9970,N_9956);
xor U10221 (N_10221,N_9988,N_9947);
and U10222 (N_10222,N_10040,N_10021);
xnor U10223 (N_10223,N_10060,N_9931);
or U10224 (N_10224,N_9941,N_9923);
nand U10225 (N_10225,N_9955,N_9947);
nor U10226 (N_10226,N_10028,N_9957);
and U10227 (N_10227,N_10058,N_9981);
or U10228 (N_10228,N_9925,N_10069);
nand U10229 (N_10229,N_9958,N_9972);
xnor U10230 (N_10230,N_9920,N_10065);
nor U10231 (N_10231,N_9981,N_9959);
or U10232 (N_10232,N_10045,N_9965);
nor U10233 (N_10233,N_9941,N_10028);
or U10234 (N_10234,N_9945,N_9951);
nor U10235 (N_10235,N_10028,N_9925);
or U10236 (N_10236,N_10039,N_9983);
or U10237 (N_10237,N_10059,N_9962);
nand U10238 (N_10238,N_10077,N_9969);
or U10239 (N_10239,N_9965,N_9985);
nor U10240 (N_10240,N_10176,N_10150);
and U10241 (N_10241,N_10123,N_10118);
and U10242 (N_10242,N_10195,N_10086);
or U10243 (N_10243,N_10156,N_10107);
nor U10244 (N_10244,N_10234,N_10143);
and U10245 (N_10245,N_10084,N_10166);
and U10246 (N_10246,N_10174,N_10230);
and U10247 (N_10247,N_10152,N_10220);
nor U10248 (N_10248,N_10211,N_10169);
nor U10249 (N_10249,N_10238,N_10111);
xnor U10250 (N_10250,N_10147,N_10205);
and U10251 (N_10251,N_10106,N_10089);
nor U10252 (N_10252,N_10170,N_10140);
nor U10253 (N_10253,N_10134,N_10225);
nand U10254 (N_10254,N_10215,N_10148);
nor U10255 (N_10255,N_10130,N_10110);
nor U10256 (N_10256,N_10221,N_10112);
or U10257 (N_10257,N_10132,N_10201);
nor U10258 (N_10258,N_10184,N_10232);
nor U10259 (N_10259,N_10109,N_10182);
or U10260 (N_10260,N_10159,N_10228);
xor U10261 (N_10261,N_10120,N_10083);
nor U10262 (N_10262,N_10196,N_10227);
and U10263 (N_10263,N_10124,N_10128);
and U10264 (N_10264,N_10210,N_10092);
and U10265 (N_10265,N_10108,N_10181);
nand U10266 (N_10266,N_10165,N_10142);
or U10267 (N_10267,N_10218,N_10131);
or U10268 (N_10268,N_10200,N_10186);
nand U10269 (N_10269,N_10236,N_10129);
or U10270 (N_10270,N_10100,N_10154);
nor U10271 (N_10271,N_10188,N_10093);
nand U10272 (N_10272,N_10204,N_10231);
nand U10273 (N_10273,N_10121,N_10105);
nor U10274 (N_10274,N_10117,N_10164);
nand U10275 (N_10275,N_10119,N_10217);
nand U10276 (N_10276,N_10209,N_10080);
or U10277 (N_10277,N_10149,N_10189);
nand U10278 (N_10278,N_10177,N_10167);
nor U10279 (N_10279,N_10222,N_10135);
or U10280 (N_10280,N_10082,N_10226);
nor U10281 (N_10281,N_10161,N_10155);
nand U10282 (N_10282,N_10157,N_10203);
nor U10283 (N_10283,N_10163,N_10187);
and U10284 (N_10284,N_10098,N_10099);
or U10285 (N_10285,N_10213,N_10104);
xnor U10286 (N_10286,N_10229,N_10202);
and U10287 (N_10287,N_10101,N_10237);
or U10288 (N_10288,N_10085,N_10239);
nor U10289 (N_10289,N_10212,N_10146);
and U10290 (N_10290,N_10206,N_10081);
and U10291 (N_10291,N_10125,N_10191);
or U10292 (N_10292,N_10168,N_10114);
nor U10293 (N_10293,N_10127,N_10162);
and U10294 (N_10294,N_10103,N_10095);
or U10295 (N_10295,N_10199,N_10190);
nand U10296 (N_10296,N_10116,N_10126);
nor U10297 (N_10297,N_10153,N_10096);
or U10298 (N_10298,N_10094,N_10198);
or U10299 (N_10299,N_10160,N_10113);
nor U10300 (N_10300,N_10219,N_10180);
nand U10301 (N_10301,N_10139,N_10138);
nor U10302 (N_10302,N_10090,N_10216);
nor U10303 (N_10303,N_10133,N_10102);
and U10304 (N_10304,N_10173,N_10194);
and U10305 (N_10305,N_10183,N_10208);
xnor U10306 (N_10306,N_10223,N_10207);
nor U10307 (N_10307,N_10087,N_10235);
nor U10308 (N_10308,N_10197,N_10178);
and U10309 (N_10309,N_10097,N_10144);
or U10310 (N_10310,N_10088,N_10171);
or U10311 (N_10311,N_10179,N_10233);
nand U10312 (N_10312,N_10145,N_10158);
nand U10313 (N_10313,N_10137,N_10192);
nor U10314 (N_10314,N_10175,N_10224);
nor U10315 (N_10315,N_10141,N_10136);
and U10316 (N_10316,N_10115,N_10091);
nand U10317 (N_10317,N_10185,N_10214);
or U10318 (N_10318,N_10122,N_10193);
nand U10319 (N_10319,N_10151,N_10172);
or U10320 (N_10320,N_10193,N_10156);
and U10321 (N_10321,N_10096,N_10137);
or U10322 (N_10322,N_10232,N_10105);
or U10323 (N_10323,N_10162,N_10081);
and U10324 (N_10324,N_10205,N_10143);
nor U10325 (N_10325,N_10189,N_10215);
nor U10326 (N_10326,N_10113,N_10211);
nor U10327 (N_10327,N_10168,N_10185);
or U10328 (N_10328,N_10153,N_10124);
and U10329 (N_10329,N_10115,N_10207);
xor U10330 (N_10330,N_10091,N_10165);
and U10331 (N_10331,N_10157,N_10146);
xnor U10332 (N_10332,N_10123,N_10149);
or U10333 (N_10333,N_10229,N_10232);
or U10334 (N_10334,N_10088,N_10209);
nand U10335 (N_10335,N_10126,N_10148);
nor U10336 (N_10336,N_10163,N_10156);
nor U10337 (N_10337,N_10080,N_10193);
and U10338 (N_10338,N_10152,N_10238);
or U10339 (N_10339,N_10166,N_10175);
nand U10340 (N_10340,N_10188,N_10200);
and U10341 (N_10341,N_10161,N_10146);
or U10342 (N_10342,N_10084,N_10151);
and U10343 (N_10343,N_10109,N_10161);
and U10344 (N_10344,N_10224,N_10235);
and U10345 (N_10345,N_10087,N_10112);
nand U10346 (N_10346,N_10114,N_10105);
nor U10347 (N_10347,N_10201,N_10173);
xnor U10348 (N_10348,N_10181,N_10137);
nor U10349 (N_10349,N_10190,N_10207);
and U10350 (N_10350,N_10091,N_10087);
and U10351 (N_10351,N_10084,N_10225);
and U10352 (N_10352,N_10081,N_10147);
nand U10353 (N_10353,N_10186,N_10220);
nand U10354 (N_10354,N_10148,N_10179);
nor U10355 (N_10355,N_10226,N_10171);
nor U10356 (N_10356,N_10134,N_10186);
nand U10357 (N_10357,N_10094,N_10197);
nor U10358 (N_10358,N_10194,N_10083);
and U10359 (N_10359,N_10101,N_10182);
or U10360 (N_10360,N_10108,N_10148);
and U10361 (N_10361,N_10131,N_10198);
or U10362 (N_10362,N_10149,N_10238);
or U10363 (N_10363,N_10140,N_10115);
nor U10364 (N_10364,N_10239,N_10237);
or U10365 (N_10365,N_10218,N_10088);
xnor U10366 (N_10366,N_10215,N_10199);
or U10367 (N_10367,N_10164,N_10123);
or U10368 (N_10368,N_10158,N_10206);
and U10369 (N_10369,N_10168,N_10189);
and U10370 (N_10370,N_10161,N_10207);
nand U10371 (N_10371,N_10110,N_10121);
or U10372 (N_10372,N_10236,N_10127);
or U10373 (N_10373,N_10220,N_10203);
nor U10374 (N_10374,N_10088,N_10119);
nand U10375 (N_10375,N_10163,N_10238);
and U10376 (N_10376,N_10154,N_10143);
nand U10377 (N_10377,N_10139,N_10231);
xor U10378 (N_10378,N_10175,N_10128);
nor U10379 (N_10379,N_10147,N_10145);
or U10380 (N_10380,N_10151,N_10205);
nand U10381 (N_10381,N_10200,N_10128);
nand U10382 (N_10382,N_10120,N_10091);
nand U10383 (N_10383,N_10204,N_10135);
xor U10384 (N_10384,N_10205,N_10119);
xor U10385 (N_10385,N_10138,N_10234);
nor U10386 (N_10386,N_10106,N_10146);
and U10387 (N_10387,N_10129,N_10119);
or U10388 (N_10388,N_10180,N_10088);
and U10389 (N_10389,N_10127,N_10188);
nor U10390 (N_10390,N_10192,N_10145);
nand U10391 (N_10391,N_10148,N_10167);
and U10392 (N_10392,N_10157,N_10115);
or U10393 (N_10393,N_10183,N_10081);
or U10394 (N_10394,N_10183,N_10239);
nand U10395 (N_10395,N_10177,N_10135);
nand U10396 (N_10396,N_10117,N_10217);
nor U10397 (N_10397,N_10107,N_10230);
and U10398 (N_10398,N_10178,N_10215);
nand U10399 (N_10399,N_10111,N_10233);
nor U10400 (N_10400,N_10334,N_10309);
or U10401 (N_10401,N_10249,N_10393);
or U10402 (N_10402,N_10272,N_10271);
and U10403 (N_10403,N_10348,N_10377);
nor U10404 (N_10404,N_10296,N_10277);
xor U10405 (N_10405,N_10283,N_10364);
or U10406 (N_10406,N_10269,N_10344);
and U10407 (N_10407,N_10371,N_10355);
nor U10408 (N_10408,N_10362,N_10304);
nand U10409 (N_10409,N_10307,N_10397);
nand U10410 (N_10410,N_10273,N_10335);
nand U10411 (N_10411,N_10342,N_10381);
and U10412 (N_10412,N_10246,N_10257);
nor U10413 (N_10413,N_10322,N_10294);
nor U10414 (N_10414,N_10350,N_10399);
nand U10415 (N_10415,N_10317,N_10326);
and U10416 (N_10416,N_10343,N_10345);
nor U10417 (N_10417,N_10265,N_10254);
or U10418 (N_10418,N_10298,N_10300);
nor U10419 (N_10419,N_10324,N_10332);
xor U10420 (N_10420,N_10285,N_10297);
nor U10421 (N_10421,N_10396,N_10242);
and U10422 (N_10422,N_10339,N_10276);
nor U10423 (N_10423,N_10386,N_10383);
and U10424 (N_10424,N_10320,N_10248);
and U10425 (N_10425,N_10284,N_10379);
and U10426 (N_10426,N_10394,N_10328);
or U10427 (N_10427,N_10329,N_10280);
nor U10428 (N_10428,N_10352,N_10250);
or U10429 (N_10429,N_10323,N_10252);
nand U10430 (N_10430,N_10353,N_10241);
and U10431 (N_10431,N_10245,N_10243);
or U10432 (N_10432,N_10366,N_10281);
and U10433 (N_10433,N_10368,N_10262);
nor U10434 (N_10434,N_10263,N_10389);
and U10435 (N_10435,N_10299,N_10319);
nand U10436 (N_10436,N_10259,N_10287);
nand U10437 (N_10437,N_10351,N_10361);
or U10438 (N_10438,N_10354,N_10346);
nor U10439 (N_10439,N_10260,N_10275);
or U10440 (N_10440,N_10376,N_10286);
xnor U10441 (N_10441,N_10356,N_10278);
nor U10442 (N_10442,N_10295,N_10388);
and U10443 (N_10443,N_10380,N_10244);
or U10444 (N_10444,N_10251,N_10369);
or U10445 (N_10445,N_10291,N_10292);
or U10446 (N_10446,N_10374,N_10310);
and U10447 (N_10447,N_10331,N_10256);
and U10448 (N_10448,N_10301,N_10311);
or U10449 (N_10449,N_10370,N_10274);
and U10450 (N_10450,N_10312,N_10279);
or U10451 (N_10451,N_10270,N_10395);
nor U10452 (N_10452,N_10303,N_10318);
nand U10453 (N_10453,N_10391,N_10340);
or U10454 (N_10454,N_10333,N_10282);
or U10455 (N_10455,N_10314,N_10373);
nor U10456 (N_10456,N_10372,N_10293);
and U10457 (N_10457,N_10253,N_10347);
nand U10458 (N_10458,N_10302,N_10336);
nand U10459 (N_10459,N_10316,N_10382);
nor U10460 (N_10460,N_10313,N_10367);
nand U10461 (N_10461,N_10358,N_10266);
and U10462 (N_10462,N_10267,N_10387);
nand U10463 (N_10463,N_10337,N_10357);
xor U10464 (N_10464,N_10365,N_10338);
or U10465 (N_10465,N_10385,N_10398);
nor U10466 (N_10466,N_10390,N_10268);
or U10467 (N_10467,N_10290,N_10325);
nand U10468 (N_10468,N_10264,N_10349);
and U10469 (N_10469,N_10392,N_10306);
or U10470 (N_10470,N_10247,N_10315);
and U10471 (N_10471,N_10305,N_10261);
and U10472 (N_10472,N_10341,N_10384);
nand U10473 (N_10473,N_10258,N_10308);
nand U10474 (N_10474,N_10360,N_10363);
xor U10475 (N_10475,N_10288,N_10378);
or U10476 (N_10476,N_10255,N_10327);
nand U10477 (N_10477,N_10359,N_10375);
or U10478 (N_10478,N_10321,N_10240);
nor U10479 (N_10479,N_10330,N_10289);
and U10480 (N_10480,N_10310,N_10318);
and U10481 (N_10481,N_10357,N_10331);
nand U10482 (N_10482,N_10373,N_10319);
nor U10483 (N_10483,N_10345,N_10346);
and U10484 (N_10484,N_10326,N_10294);
or U10485 (N_10485,N_10277,N_10264);
xnor U10486 (N_10486,N_10360,N_10377);
and U10487 (N_10487,N_10387,N_10294);
or U10488 (N_10488,N_10240,N_10361);
and U10489 (N_10489,N_10360,N_10274);
nor U10490 (N_10490,N_10276,N_10279);
xor U10491 (N_10491,N_10398,N_10311);
nor U10492 (N_10492,N_10309,N_10382);
nor U10493 (N_10493,N_10271,N_10313);
nand U10494 (N_10494,N_10254,N_10283);
or U10495 (N_10495,N_10349,N_10398);
or U10496 (N_10496,N_10339,N_10290);
nand U10497 (N_10497,N_10313,N_10244);
or U10498 (N_10498,N_10351,N_10284);
or U10499 (N_10499,N_10315,N_10316);
nand U10500 (N_10500,N_10294,N_10355);
nand U10501 (N_10501,N_10267,N_10343);
nor U10502 (N_10502,N_10250,N_10317);
nand U10503 (N_10503,N_10380,N_10302);
nor U10504 (N_10504,N_10382,N_10335);
nand U10505 (N_10505,N_10363,N_10303);
or U10506 (N_10506,N_10269,N_10370);
nand U10507 (N_10507,N_10243,N_10394);
or U10508 (N_10508,N_10309,N_10374);
nor U10509 (N_10509,N_10361,N_10312);
or U10510 (N_10510,N_10395,N_10264);
nor U10511 (N_10511,N_10398,N_10283);
and U10512 (N_10512,N_10314,N_10380);
nand U10513 (N_10513,N_10349,N_10240);
nor U10514 (N_10514,N_10282,N_10260);
nand U10515 (N_10515,N_10342,N_10396);
or U10516 (N_10516,N_10283,N_10292);
or U10517 (N_10517,N_10357,N_10380);
nand U10518 (N_10518,N_10283,N_10345);
and U10519 (N_10519,N_10348,N_10240);
and U10520 (N_10520,N_10332,N_10303);
or U10521 (N_10521,N_10329,N_10354);
nand U10522 (N_10522,N_10271,N_10379);
nor U10523 (N_10523,N_10330,N_10247);
nor U10524 (N_10524,N_10352,N_10310);
or U10525 (N_10525,N_10257,N_10278);
nor U10526 (N_10526,N_10317,N_10290);
nor U10527 (N_10527,N_10367,N_10282);
or U10528 (N_10528,N_10314,N_10355);
nor U10529 (N_10529,N_10259,N_10382);
and U10530 (N_10530,N_10393,N_10279);
nand U10531 (N_10531,N_10397,N_10385);
nor U10532 (N_10532,N_10382,N_10251);
nand U10533 (N_10533,N_10295,N_10393);
nor U10534 (N_10534,N_10377,N_10300);
nor U10535 (N_10535,N_10344,N_10333);
and U10536 (N_10536,N_10376,N_10396);
xnor U10537 (N_10537,N_10243,N_10314);
or U10538 (N_10538,N_10379,N_10380);
nand U10539 (N_10539,N_10370,N_10383);
or U10540 (N_10540,N_10383,N_10294);
or U10541 (N_10541,N_10349,N_10384);
nor U10542 (N_10542,N_10343,N_10285);
nor U10543 (N_10543,N_10372,N_10249);
nor U10544 (N_10544,N_10360,N_10388);
or U10545 (N_10545,N_10364,N_10356);
or U10546 (N_10546,N_10254,N_10271);
or U10547 (N_10547,N_10315,N_10309);
xnor U10548 (N_10548,N_10376,N_10254);
or U10549 (N_10549,N_10324,N_10354);
nor U10550 (N_10550,N_10304,N_10356);
nand U10551 (N_10551,N_10355,N_10318);
or U10552 (N_10552,N_10348,N_10291);
nor U10553 (N_10553,N_10307,N_10351);
nor U10554 (N_10554,N_10292,N_10347);
or U10555 (N_10555,N_10348,N_10271);
xnor U10556 (N_10556,N_10268,N_10396);
nor U10557 (N_10557,N_10259,N_10321);
and U10558 (N_10558,N_10361,N_10305);
or U10559 (N_10559,N_10300,N_10263);
or U10560 (N_10560,N_10552,N_10459);
or U10561 (N_10561,N_10431,N_10451);
and U10562 (N_10562,N_10524,N_10403);
nor U10563 (N_10563,N_10477,N_10468);
nand U10564 (N_10564,N_10549,N_10548);
or U10565 (N_10565,N_10519,N_10536);
or U10566 (N_10566,N_10454,N_10413);
nor U10567 (N_10567,N_10490,N_10506);
and U10568 (N_10568,N_10445,N_10415);
nor U10569 (N_10569,N_10491,N_10523);
or U10570 (N_10570,N_10407,N_10417);
xnor U10571 (N_10571,N_10492,N_10527);
or U10572 (N_10572,N_10432,N_10467);
or U10573 (N_10573,N_10481,N_10430);
or U10574 (N_10574,N_10483,N_10489);
xor U10575 (N_10575,N_10500,N_10525);
nor U10576 (N_10576,N_10473,N_10484);
and U10577 (N_10577,N_10505,N_10482);
or U10578 (N_10578,N_10550,N_10528);
and U10579 (N_10579,N_10486,N_10558);
or U10580 (N_10580,N_10410,N_10555);
xnor U10581 (N_10581,N_10520,N_10557);
and U10582 (N_10582,N_10400,N_10539);
nand U10583 (N_10583,N_10531,N_10499);
nand U10584 (N_10584,N_10414,N_10426);
and U10585 (N_10585,N_10479,N_10416);
or U10586 (N_10586,N_10406,N_10502);
nor U10587 (N_10587,N_10534,N_10465);
nor U10588 (N_10588,N_10433,N_10504);
and U10589 (N_10589,N_10423,N_10553);
and U10590 (N_10590,N_10480,N_10463);
xor U10591 (N_10591,N_10441,N_10515);
and U10592 (N_10592,N_10556,N_10434);
and U10593 (N_10593,N_10478,N_10530);
or U10594 (N_10594,N_10538,N_10509);
or U10595 (N_10595,N_10476,N_10475);
xnor U10596 (N_10596,N_10455,N_10438);
or U10597 (N_10597,N_10472,N_10452);
xnor U10598 (N_10598,N_10450,N_10429);
or U10599 (N_10599,N_10424,N_10469);
xor U10600 (N_10600,N_10512,N_10510);
nand U10601 (N_10601,N_10507,N_10453);
nor U10602 (N_10602,N_10526,N_10404);
nor U10603 (N_10603,N_10488,N_10543);
nor U10604 (N_10604,N_10495,N_10487);
nor U10605 (N_10605,N_10447,N_10464);
nor U10606 (N_10606,N_10551,N_10440);
and U10607 (N_10607,N_10401,N_10462);
xor U10608 (N_10608,N_10419,N_10474);
xnor U10609 (N_10609,N_10540,N_10402);
nor U10610 (N_10610,N_10533,N_10493);
xnor U10611 (N_10611,N_10498,N_10521);
xor U10612 (N_10612,N_10466,N_10442);
and U10613 (N_10613,N_10443,N_10503);
nand U10614 (N_10614,N_10514,N_10448);
and U10615 (N_10615,N_10541,N_10529);
xnor U10616 (N_10616,N_10411,N_10508);
nor U10617 (N_10617,N_10449,N_10532);
and U10618 (N_10618,N_10554,N_10516);
nand U10619 (N_10619,N_10436,N_10412);
or U10620 (N_10620,N_10439,N_10518);
nor U10621 (N_10621,N_10457,N_10546);
or U10622 (N_10622,N_10458,N_10460);
nor U10623 (N_10623,N_10544,N_10405);
nor U10624 (N_10624,N_10427,N_10409);
and U10625 (N_10625,N_10537,N_10559);
xor U10626 (N_10626,N_10496,N_10535);
and U10627 (N_10627,N_10418,N_10420);
nor U10628 (N_10628,N_10522,N_10485);
or U10629 (N_10629,N_10497,N_10408);
or U10630 (N_10630,N_10435,N_10446);
nor U10631 (N_10631,N_10421,N_10461);
and U10632 (N_10632,N_10444,N_10517);
and U10633 (N_10633,N_10542,N_10425);
nor U10634 (N_10634,N_10456,N_10437);
nor U10635 (N_10635,N_10471,N_10547);
and U10636 (N_10636,N_10545,N_10511);
and U10637 (N_10637,N_10428,N_10501);
or U10638 (N_10638,N_10513,N_10470);
nor U10639 (N_10639,N_10494,N_10422);
nor U10640 (N_10640,N_10461,N_10499);
nor U10641 (N_10641,N_10530,N_10454);
or U10642 (N_10642,N_10524,N_10484);
nor U10643 (N_10643,N_10410,N_10543);
nor U10644 (N_10644,N_10473,N_10425);
and U10645 (N_10645,N_10518,N_10550);
nor U10646 (N_10646,N_10552,N_10479);
xor U10647 (N_10647,N_10439,N_10537);
nor U10648 (N_10648,N_10457,N_10466);
and U10649 (N_10649,N_10500,N_10406);
or U10650 (N_10650,N_10468,N_10403);
or U10651 (N_10651,N_10421,N_10458);
and U10652 (N_10652,N_10461,N_10542);
nand U10653 (N_10653,N_10463,N_10484);
xor U10654 (N_10654,N_10430,N_10402);
nand U10655 (N_10655,N_10481,N_10469);
or U10656 (N_10656,N_10507,N_10504);
xor U10657 (N_10657,N_10423,N_10467);
nor U10658 (N_10658,N_10459,N_10533);
and U10659 (N_10659,N_10430,N_10426);
nand U10660 (N_10660,N_10473,N_10469);
or U10661 (N_10661,N_10466,N_10521);
nand U10662 (N_10662,N_10506,N_10539);
nand U10663 (N_10663,N_10557,N_10411);
nand U10664 (N_10664,N_10461,N_10549);
nand U10665 (N_10665,N_10469,N_10408);
nor U10666 (N_10666,N_10553,N_10509);
nor U10667 (N_10667,N_10412,N_10417);
and U10668 (N_10668,N_10467,N_10447);
xnor U10669 (N_10669,N_10449,N_10521);
nor U10670 (N_10670,N_10511,N_10550);
or U10671 (N_10671,N_10429,N_10523);
nand U10672 (N_10672,N_10518,N_10551);
nor U10673 (N_10673,N_10511,N_10441);
nor U10674 (N_10674,N_10473,N_10531);
or U10675 (N_10675,N_10422,N_10411);
or U10676 (N_10676,N_10493,N_10480);
nor U10677 (N_10677,N_10449,N_10482);
and U10678 (N_10678,N_10532,N_10416);
nor U10679 (N_10679,N_10434,N_10521);
and U10680 (N_10680,N_10559,N_10517);
nor U10681 (N_10681,N_10503,N_10404);
or U10682 (N_10682,N_10542,N_10409);
nand U10683 (N_10683,N_10404,N_10517);
and U10684 (N_10684,N_10455,N_10539);
and U10685 (N_10685,N_10490,N_10487);
nor U10686 (N_10686,N_10476,N_10491);
nor U10687 (N_10687,N_10514,N_10493);
nand U10688 (N_10688,N_10432,N_10492);
nand U10689 (N_10689,N_10559,N_10413);
nor U10690 (N_10690,N_10538,N_10427);
nand U10691 (N_10691,N_10426,N_10555);
and U10692 (N_10692,N_10498,N_10427);
nand U10693 (N_10693,N_10459,N_10411);
nor U10694 (N_10694,N_10544,N_10407);
and U10695 (N_10695,N_10460,N_10416);
and U10696 (N_10696,N_10445,N_10462);
and U10697 (N_10697,N_10457,N_10489);
or U10698 (N_10698,N_10550,N_10414);
and U10699 (N_10699,N_10475,N_10531);
xor U10700 (N_10700,N_10409,N_10557);
nand U10701 (N_10701,N_10407,N_10428);
and U10702 (N_10702,N_10556,N_10441);
and U10703 (N_10703,N_10428,N_10468);
xor U10704 (N_10704,N_10519,N_10522);
or U10705 (N_10705,N_10430,N_10446);
nand U10706 (N_10706,N_10493,N_10465);
or U10707 (N_10707,N_10510,N_10506);
and U10708 (N_10708,N_10474,N_10403);
or U10709 (N_10709,N_10465,N_10503);
and U10710 (N_10710,N_10521,N_10463);
nor U10711 (N_10711,N_10531,N_10543);
nor U10712 (N_10712,N_10419,N_10426);
and U10713 (N_10713,N_10412,N_10408);
xor U10714 (N_10714,N_10538,N_10466);
and U10715 (N_10715,N_10543,N_10552);
nand U10716 (N_10716,N_10470,N_10415);
nor U10717 (N_10717,N_10557,N_10533);
xor U10718 (N_10718,N_10518,N_10474);
nand U10719 (N_10719,N_10439,N_10432);
nand U10720 (N_10720,N_10712,N_10566);
or U10721 (N_10721,N_10628,N_10694);
or U10722 (N_10722,N_10666,N_10684);
nor U10723 (N_10723,N_10565,N_10676);
xnor U10724 (N_10724,N_10618,N_10713);
nand U10725 (N_10725,N_10603,N_10562);
or U10726 (N_10726,N_10589,N_10681);
or U10727 (N_10727,N_10653,N_10682);
xnor U10728 (N_10728,N_10576,N_10658);
nor U10729 (N_10729,N_10607,N_10572);
xor U10730 (N_10730,N_10637,N_10641);
nand U10731 (N_10731,N_10668,N_10595);
and U10732 (N_10732,N_10616,N_10627);
nor U10733 (N_10733,N_10649,N_10591);
and U10734 (N_10734,N_10669,N_10645);
or U10735 (N_10735,N_10609,N_10575);
or U10736 (N_10736,N_10635,N_10652);
or U10737 (N_10737,N_10673,N_10708);
nor U10738 (N_10738,N_10655,N_10568);
nor U10739 (N_10739,N_10710,N_10581);
xor U10740 (N_10740,N_10711,N_10640);
and U10741 (N_10741,N_10593,N_10683);
nand U10742 (N_10742,N_10570,N_10588);
nand U10743 (N_10743,N_10672,N_10714);
nand U10744 (N_10744,N_10717,N_10642);
nand U10745 (N_10745,N_10650,N_10602);
nand U10746 (N_10746,N_10661,N_10662);
nor U10747 (N_10747,N_10692,N_10634);
and U10748 (N_10748,N_10585,N_10571);
or U10749 (N_10749,N_10630,N_10660);
or U10750 (N_10750,N_10698,N_10719);
nand U10751 (N_10751,N_10690,N_10622);
xnor U10752 (N_10752,N_10646,N_10590);
nand U10753 (N_10753,N_10617,N_10689);
xnor U10754 (N_10754,N_10716,N_10677);
xnor U10755 (N_10755,N_10573,N_10612);
or U10756 (N_10756,N_10619,N_10706);
and U10757 (N_10757,N_10586,N_10671);
nand U10758 (N_10758,N_10623,N_10648);
or U10759 (N_10759,N_10624,N_10691);
nand U10760 (N_10760,N_10701,N_10674);
and U10761 (N_10761,N_10569,N_10608);
xnor U10762 (N_10762,N_10643,N_10625);
and U10763 (N_10763,N_10577,N_10582);
and U10764 (N_10764,N_10705,N_10580);
nor U10765 (N_10765,N_10564,N_10615);
or U10766 (N_10766,N_10584,N_10563);
nor U10767 (N_10767,N_10620,N_10610);
nand U10768 (N_10768,N_10656,N_10667);
nor U10769 (N_10769,N_10700,N_10699);
nor U10770 (N_10770,N_10665,N_10695);
nor U10771 (N_10771,N_10604,N_10594);
xor U10772 (N_10772,N_10574,N_10614);
nand U10773 (N_10773,N_10583,N_10709);
nand U10774 (N_10774,N_10696,N_10632);
xor U10775 (N_10775,N_10678,N_10629);
or U10776 (N_10776,N_10657,N_10679);
xnor U10777 (N_10777,N_10647,N_10664);
and U10778 (N_10778,N_10636,N_10686);
or U10779 (N_10779,N_10707,N_10626);
or U10780 (N_10780,N_10680,N_10613);
or U10781 (N_10781,N_10561,N_10702);
nor U10782 (N_10782,N_10688,N_10644);
nand U10783 (N_10783,N_10601,N_10715);
and U10784 (N_10784,N_10654,N_10685);
and U10785 (N_10785,N_10651,N_10639);
and U10786 (N_10786,N_10663,N_10600);
xnor U10787 (N_10787,N_10704,N_10599);
and U10788 (N_10788,N_10638,N_10592);
or U10789 (N_10789,N_10597,N_10560);
or U10790 (N_10790,N_10697,N_10578);
nor U10791 (N_10791,N_10587,N_10703);
nand U10792 (N_10792,N_10633,N_10631);
and U10793 (N_10793,N_10605,N_10670);
or U10794 (N_10794,N_10611,N_10579);
and U10795 (N_10795,N_10598,N_10675);
or U10796 (N_10796,N_10606,N_10596);
xor U10797 (N_10797,N_10659,N_10718);
nor U10798 (N_10798,N_10693,N_10621);
xnor U10799 (N_10799,N_10687,N_10567);
nand U10800 (N_10800,N_10625,N_10713);
and U10801 (N_10801,N_10592,N_10637);
and U10802 (N_10802,N_10598,N_10619);
xnor U10803 (N_10803,N_10590,N_10683);
or U10804 (N_10804,N_10673,N_10693);
nor U10805 (N_10805,N_10709,N_10654);
nor U10806 (N_10806,N_10690,N_10638);
nor U10807 (N_10807,N_10619,N_10689);
nand U10808 (N_10808,N_10655,N_10603);
or U10809 (N_10809,N_10674,N_10715);
nor U10810 (N_10810,N_10620,N_10570);
nor U10811 (N_10811,N_10682,N_10595);
and U10812 (N_10812,N_10683,N_10611);
and U10813 (N_10813,N_10660,N_10686);
xnor U10814 (N_10814,N_10584,N_10560);
and U10815 (N_10815,N_10579,N_10637);
or U10816 (N_10816,N_10623,N_10636);
nor U10817 (N_10817,N_10666,N_10614);
nor U10818 (N_10818,N_10698,N_10645);
nor U10819 (N_10819,N_10630,N_10602);
nand U10820 (N_10820,N_10608,N_10641);
or U10821 (N_10821,N_10576,N_10683);
and U10822 (N_10822,N_10632,N_10637);
or U10823 (N_10823,N_10690,N_10706);
nand U10824 (N_10824,N_10617,N_10706);
nand U10825 (N_10825,N_10625,N_10615);
and U10826 (N_10826,N_10560,N_10644);
or U10827 (N_10827,N_10594,N_10576);
nor U10828 (N_10828,N_10651,N_10674);
nand U10829 (N_10829,N_10585,N_10614);
nand U10830 (N_10830,N_10580,N_10579);
and U10831 (N_10831,N_10659,N_10578);
or U10832 (N_10832,N_10710,N_10642);
xor U10833 (N_10833,N_10708,N_10629);
and U10834 (N_10834,N_10608,N_10665);
nand U10835 (N_10835,N_10612,N_10643);
xnor U10836 (N_10836,N_10591,N_10695);
nor U10837 (N_10837,N_10645,N_10670);
nor U10838 (N_10838,N_10593,N_10715);
and U10839 (N_10839,N_10710,N_10668);
xor U10840 (N_10840,N_10688,N_10713);
and U10841 (N_10841,N_10711,N_10612);
xor U10842 (N_10842,N_10634,N_10595);
nand U10843 (N_10843,N_10693,N_10614);
or U10844 (N_10844,N_10588,N_10665);
nor U10845 (N_10845,N_10705,N_10601);
and U10846 (N_10846,N_10701,N_10715);
nor U10847 (N_10847,N_10600,N_10578);
nor U10848 (N_10848,N_10634,N_10646);
xnor U10849 (N_10849,N_10568,N_10570);
nand U10850 (N_10850,N_10625,N_10578);
and U10851 (N_10851,N_10648,N_10717);
and U10852 (N_10852,N_10624,N_10636);
nor U10853 (N_10853,N_10621,N_10610);
and U10854 (N_10854,N_10616,N_10688);
nor U10855 (N_10855,N_10590,N_10638);
or U10856 (N_10856,N_10656,N_10682);
nor U10857 (N_10857,N_10571,N_10586);
nor U10858 (N_10858,N_10640,N_10587);
and U10859 (N_10859,N_10716,N_10578);
nand U10860 (N_10860,N_10580,N_10707);
or U10861 (N_10861,N_10590,N_10701);
nor U10862 (N_10862,N_10632,N_10650);
nor U10863 (N_10863,N_10614,N_10641);
nand U10864 (N_10864,N_10689,N_10717);
nand U10865 (N_10865,N_10682,N_10707);
xor U10866 (N_10866,N_10585,N_10625);
nor U10867 (N_10867,N_10575,N_10576);
or U10868 (N_10868,N_10715,N_10696);
nand U10869 (N_10869,N_10647,N_10644);
or U10870 (N_10870,N_10649,N_10700);
nor U10871 (N_10871,N_10610,N_10582);
and U10872 (N_10872,N_10597,N_10702);
and U10873 (N_10873,N_10664,N_10689);
nor U10874 (N_10874,N_10651,N_10598);
and U10875 (N_10875,N_10711,N_10693);
nand U10876 (N_10876,N_10686,N_10583);
or U10877 (N_10877,N_10702,N_10622);
or U10878 (N_10878,N_10605,N_10620);
nand U10879 (N_10879,N_10696,N_10708);
nand U10880 (N_10880,N_10789,N_10748);
or U10881 (N_10881,N_10795,N_10786);
or U10882 (N_10882,N_10756,N_10858);
or U10883 (N_10883,N_10741,N_10827);
nand U10884 (N_10884,N_10726,N_10792);
and U10885 (N_10885,N_10796,N_10768);
nor U10886 (N_10886,N_10875,N_10830);
xnor U10887 (N_10887,N_10806,N_10820);
nand U10888 (N_10888,N_10769,N_10738);
or U10889 (N_10889,N_10735,N_10841);
nand U10890 (N_10890,N_10753,N_10800);
nor U10891 (N_10891,N_10851,N_10823);
or U10892 (N_10892,N_10817,N_10736);
xnor U10893 (N_10893,N_10864,N_10863);
and U10894 (N_10894,N_10879,N_10764);
nand U10895 (N_10895,N_10754,N_10816);
nand U10896 (N_10896,N_10788,N_10731);
nand U10897 (N_10897,N_10846,N_10771);
and U10898 (N_10898,N_10834,N_10844);
nand U10899 (N_10899,N_10782,N_10773);
or U10900 (N_10900,N_10856,N_10824);
or U10901 (N_10901,N_10868,N_10776);
nand U10902 (N_10902,N_10751,N_10848);
and U10903 (N_10903,N_10758,N_10843);
or U10904 (N_10904,N_10798,N_10878);
nor U10905 (N_10905,N_10759,N_10766);
and U10906 (N_10906,N_10752,N_10873);
nor U10907 (N_10907,N_10742,N_10732);
nand U10908 (N_10908,N_10737,N_10745);
nand U10909 (N_10909,N_10826,N_10859);
and U10910 (N_10910,N_10870,N_10877);
xor U10911 (N_10911,N_10832,N_10866);
or U10912 (N_10912,N_10803,N_10727);
nand U10913 (N_10913,N_10770,N_10867);
or U10914 (N_10914,N_10833,N_10805);
or U10915 (N_10915,N_10860,N_10744);
and U10916 (N_10916,N_10779,N_10787);
nor U10917 (N_10917,N_10849,N_10855);
nand U10918 (N_10918,N_10755,N_10743);
nor U10919 (N_10919,N_10857,N_10840);
nand U10920 (N_10920,N_10750,N_10847);
nand U10921 (N_10921,N_10739,N_10845);
and U10922 (N_10922,N_10872,N_10740);
and U10923 (N_10923,N_10876,N_10865);
xor U10924 (N_10924,N_10821,N_10777);
nor U10925 (N_10925,N_10825,N_10730);
nand U10926 (N_10926,N_10813,N_10874);
and U10927 (N_10927,N_10775,N_10853);
or U10928 (N_10928,N_10762,N_10774);
and U10929 (N_10929,N_10838,N_10810);
and U10930 (N_10930,N_10828,N_10837);
or U10931 (N_10931,N_10807,N_10746);
or U10932 (N_10932,N_10729,N_10862);
xor U10933 (N_10933,N_10794,N_10811);
or U10934 (N_10934,N_10780,N_10812);
nor U10935 (N_10935,N_10869,N_10818);
nand U10936 (N_10936,N_10835,N_10808);
and U10937 (N_10937,N_10815,N_10733);
nand U10938 (N_10938,N_10802,N_10871);
nor U10939 (N_10939,N_10783,N_10722);
nand U10940 (N_10940,N_10852,N_10724);
nor U10941 (N_10941,N_10854,N_10861);
nor U10942 (N_10942,N_10829,N_10822);
nor U10943 (N_10943,N_10772,N_10781);
nand U10944 (N_10944,N_10831,N_10778);
nand U10945 (N_10945,N_10749,N_10793);
nor U10946 (N_10946,N_10842,N_10723);
or U10947 (N_10947,N_10801,N_10767);
nor U10948 (N_10948,N_10765,N_10760);
xor U10949 (N_10949,N_10757,N_10799);
nand U10950 (N_10950,N_10734,N_10809);
or U10951 (N_10951,N_10814,N_10784);
nor U10952 (N_10952,N_10790,N_10804);
nand U10953 (N_10953,N_10728,N_10720);
nor U10954 (N_10954,N_10839,N_10725);
and U10955 (N_10955,N_10797,N_10791);
xnor U10956 (N_10956,N_10785,N_10819);
and U10957 (N_10957,N_10836,N_10850);
nand U10958 (N_10958,N_10763,N_10721);
nand U10959 (N_10959,N_10747,N_10761);
nor U10960 (N_10960,N_10875,N_10824);
and U10961 (N_10961,N_10740,N_10786);
and U10962 (N_10962,N_10770,N_10777);
and U10963 (N_10963,N_10720,N_10730);
nor U10964 (N_10964,N_10833,N_10871);
nand U10965 (N_10965,N_10791,N_10775);
nor U10966 (N_10966,N_10721,N_10756);
or U10967 (N_10967,N_10838,N_10765);
or U10968 (N_10968,N_10829,N_10854);
and U10969 (N_10969,N_10779,N_10760);
nor U10970 (N_10970,N_10830,N_10739);
nand U10971 (N_10971,N_10813,N_10799);
and U10972 (N_10972,N_10839,N_10770);
and U10973 (N_10973,N_10817,N_10797);
nor U10974 (N_10974,N_10830,N_10755);
xnor U10975 (N_10975,N_10812,N_10817);
nand U10976 (N_10976,N_10832,N_10777);
or U10977 (N_10977,N_10830,N_10860);
and U10978 (N_10978,N_10801,N_10784);
nand U10979 (N_10979,N_10790,N_10827);
nor U10980 (N_10980,N_10732,N_10806);
and U10981 (N_10981,N_10722,N_10864);
nor U10982 (N_10982,N_10852,N_10865);
nor U10983 (N_10983,N_10736,N_10735);
and U10984 (N_10984,N_10774,N_10721);
nand U10985 (N_10985,N_10778,N_10850);
or U10986 (N_10986,N_10751,N_10765);
nor U10987 (N_10987,N_10798,N_10752);
nand U10988 (N_10988,N_10831,N_10731);
and U10989 (N_10989,N_10855,N_10859);
xnor U10990 (N_10990,N_10765,N_10844);
nand U10991 (N_10991,N_10753,N_10814);
nand U10992 (N_10992,N_10876,N_10766);
or U10993 (N_10993,N_10862,N_10836);
nand U10994 (N_10994,N_10796,N_10870);
nor U10995 (N_10995,N_10739,N_10843);
xnor U10996 (N_10996,N_10844,N_10774);
xor U10997 (N_10997,N_10727,N_10842);
and U10998 (N_10998,N_10859,N_10770);
and U10999 (N_10999,N_10850,N_10748);
nor U11000 (N_11000,N_10876,N_10866);
xnor U11001 (N_11001,N_10862,N_10828);
and U11002 (N_11002,N_10811,N_10805);
nand U11003 (N_11003,N_10828,N_10750);
nand U11004 (N_11004,N_10857,N_10795);
xnor U11005 (N_11005,N_10739,N_10847);
nand U11006 (N_11006,N_10876,N_10757);
or U11007 (N_11007,N_10740,N_10783);
and U11008 (N_11008,N_10809,N_10798);
or U11009 (N_11009,N_10734,N_10755);
and U11010 (N_11010,N_10860,N_10865);
or U11011 (N_11011,N_10829,N_10743);
nor U11012 (N_11012,N_10807,N_10814);
nand U11013 (N_11013,N_10721,N_10855);
and U11014 (N_11014,N_10745,N_10739);
nor U11015 (N_11015,N_10786,N_10758);
and U11016 (N_11016,N_10845,N_10867);
or U11017 (N_11017,N_10873,N_10877);
and U11018 (N_11018,N_10855,N_10866);
nor U11019 (N_11019,N_10874,N_10754);
or U11020 (N_11020,N_10771,N_10811);
xor U11021 (N_11021,N_10844,N_10787);
and U11022 (N_11022,N_10872,N_10844);
xor U11023 (N_11023,N_10815,N_10775);
nor U11024 (N_11024,N_10738,N_10774);
nand U11025 (N_11025,N_10793,N_10837);
or U11026 (N_11026,N_10727,N_10854);
or U11027 (N_11027,N_10797,N_10798);
or U11028 (N_11028,N_10871,N_10869);
or U11029 (N_11029,N_10871,N_10768);
nand U11030 (N_11030,N_10862,N_10873);
xor U11031 (N_11031,N_10836,N_10746);
or U11032 (N_11032,N_10788,N_10767);
and U11033 (N_11033,N_10774,N_10773);
or U11034 (N_11034,N_10770,N_10822);
nand U11035 (N_11035,N_10858,N_10765);
or U11036 (N_11036,N_10872,N_10785);
and U11037 (N_11037,N_10821,N_10878);
nand U11038 (N_11038,N_10848,N_10856);
nand U11039 (N_11039,N_10744,N_10787);
nor U11040 (N_11040,N_10886,N_10943);
nor U11041 (N_11041,N_11037,N_11007);
xor U11042 (N_11042,N_11015,N_10930);
or U11043 (N_11043,N_11019,N_10908);
xnor U11044 (N_11044,N_10948,N_10912);
nor U11045 (N_11045,N_10974,N_10905);
nand U11046 (N_11046,N_10911,N_11016);
nand U11047 (N_11047,N_10904,N_10919);
or U11048 (N_11048,N_10967,N_10979);
nand U11049 (N_11049,N_11029,N_10944);
nor U11050 (N_11050,N_10927,N_10994);
and U11051 (N_11051,N_10946,N_10906);
nand U11052 (N_11052,N_11023,N_10881);
nand U11053 (N_11053,N_10907,N_10986);
or U11054 (N_11054,N_10988,N_10902);
or U11055 (N_11055,N_10952,N_11002);
nor U11056 (N_11056,N_10966,N_11039);
nor U11057 (N_11057,N_10933,N_10897);
nand U11058 (N_11058,N_10982,N_11008);
xor U11059 (N_11059,N_10955,N_11024);
and U11060 (N_11060,N_11011,N_10909);
nand U11061 (N_11061,N_11004,N_10889);
or U11062 (N_11062,N_10996,N_10899);
nor U11063 (N_11063,N_10903,N_11014);
and U11064 (N_11064,N_10938,N_10926);
nand U11065 (N_11065,N_11001,N_10925);
or U11066 (N_11066,N_10950,N_10900);
and U11067 (N_11067,N_10995,N_10997);
or U11068 (N_11068,N_10956,N_10949);
nor U11069 (N_11069,N_10880,N_11010);
and U11070 (N_11070,N_10921,N_10983);
nor U11071 (N_11071,N_10892,N_10971);
nor U11072 (N_11072,N_11031,N_10954);
and U11073 (N_11073,N_10989,N_10984);
xnor U11074 (N_11074,N_10951,N_10940);
and U11075 (N_11075,N_11005,N_11038);
nor U11076 (N_11076,N_10991,N_10969);
nand U11077 (N_11077,N_10962,N_10923);
xor U11078 (N_11078,N_10960,N_10913);
nor U11079 (N_11079,N_11032,N_10890);
xnor U11080 (N_11080,N_11027,N_10882);
nand U11081 (N_11081,N_11034,N_10910);
and U11082 (N_11082,N_10980,N_11003);
or U11083 (N_11083,N_10916,N_10887);
nor U11084 (N_11084,N_10959,N_10895);
nor U11085 (N_11085,N_10885,N_10993);
or U11086 (N_11086,N_10939,N_10884);
xnor U11087 (N_11087,N_10936,N_11026);
nor U11088 (N_11088,N_10981,N_10898);
nand U11089 (N_11089,N_10888,N_10924);
and U11090 (N_11090,N_10914,N_11006);
and U11091 (N_11091,N_11021,N_10953);
or U11092 (N_11092,N_10992,N_11013);
nand U11093 (N_11093,N_10945,N_10891);
or U11094 (N_11094,N_10934,N_10965);
and U11095 (N_11095,N_10917,N_10999);
or U11096 (N_11096,N_10915,N_10932);
or U11097 (N_11097,N_11030,N_10947);
and U11098 (N_11098,N_11033,N_10928);
xor U11099 (N_11099,N_10970,N_10973);
xnor U11100 (N_11100,N_11036,N_11000);
or U11101 (N_11101,N_11028,N_10963);
nand U11102 (N_11102,N_11018,N_10896);
nor U11103 (N_11103,N_10918,N_10931);
nand U11104 (N_11104,N_10964,N_10893);
and U11105 (N_11105,N_10883,N_10920);
nor U11106 (N_11106,N_10942,N_11012);
or U11107 (N_11107,N_11025,N_10978);
and U11108 (N_11108,N_10990,N_10975);
and U11109 (N_11109,N_11017,N_10941);
nand U11110 (N_11110,N_10968,N_10998);
nor U11111 (N_11111,N_10977,N_11009);
and U11112 (N_11112,N_10922,N_10976);
or U11113 (N_11113,N_11020,N_10901);
xor U11114 (N_11114,N_10894,N_10987);
nor U11115 (N_11115,N_11022,N_10972);
nand U11116 (N_11116,N_11035,N_10957);
nand U11117 (N_11117,N_10929,N_10937);
nor U11118 (N_11118,N_10985,N_10961);
nor U11119 (N_11119,N_10958,N_10935);
nor U11120 (N_11120,N_10982,N_10998);
nor U11121 (N_11121,N_10898,N_11029);
nor U11122 (N_11122,N_10943,N_10985);
xnor U11123 (N_11123,N_10895,N_11015);
or U11124 (N_11124,N_11013,N_10990);
nand U11125 (N_11125,N_10992,N_10978);
nand U11126 (N_11126,N_11015,N_10973);
nor U11127 (N_11127,N_10950,N_10889);
nor U11128 (N_11128,N_11022,N_10982);
or U11129 (N_11129,N_11022,N_10913);
nor U11130 (N_11130,N_10905,N_10933);
or U11131 (N_11131,N_10940,N_10903);
xor U11132 (N_11132,N_10997,N_11004);
nor U11133 (N_11133,N_10992,N_10915);
or U11134 (N_11134,N_10909,N_10981);
nand U11135 (N_11135,N_10882,N_10924);
nand U11136 (N_11136,N_10915,N_11038);
nand U11137 (N_11137,N_10999,N_11005);
or U11138 (N_11138,N_10949,N_10986);
or U11139 (N_11139,N_10939,N_11001);
and U11140 (N_11140,N_10941,N_10926);
and U11141 (N_11141,N_10896,N_10937);
nor U11142 (N_11142,N_10956,N_10998);
and U11143 (N_11143,N_10892,N_10998);
nand U11144 (N_11144,N_11010,N_10885);
nand U11145 (N_11145,N_10923,N_11006);
and U11146 (N_11146,N_10996,N_10917);
nand U11147 (N_11147,N_11032,N_10966);
or U11148 (N_11148,N_11002,N_11037);
and U11149 (N_11149,N_10916,N_10937);
and U11150 (N_11150,N_10923,N_11039);
nor U11151 (N_11151,N_10956,N_10882);
nor U11152 (N_11152,N_10925,N_10940);
and U11153 (N_11153,N_10975,N_11007);
or U11154 (N_11154,N_10951,N_10900);
or U11155 (N_11155,N_10955,N_10900);
or U11156 (N_11156,N_10971,N_10905);
nor U11157 (N_11157,N_10970,N_10934);
or U11158 (N_11158,N_10943,N_10962);
or U11159 (N_11159,N_10926,N_11025);
nand U11160 (N_11160,N_10987,N_10891);
nor U11161 (N_11161,N_11038,N_10993);
nand U11162 (N_11162,N_10942,N_10896);
nor U11163 (N_11163,N_11038,N_10935);
and U11164 (N_11164,N_10916,N_11031);
xor U11165 (N_11165,N_10947,N_10968);
nand U11166 (N_11166,N_10917,N_10931);
xnor U11167 (N_11167,N_10979,N_10999);
xor U11168 (N_11168,N_10977,N_10924);
or U11169 (N_11169,N_10897,N_10917);
nand U11170 (N_11170,N_10880,N_10928);
nor U11171 (N_11171,N_11016,N_10898);
nor U11172 (N_11172,N_10932,N_11001);
or U11173 (N_11173,N_10988,N_10938);
nand U11174 (N_11174,N_10905,N_10932);
nor U11175 (N_11175,N_10943,N_11006);
and U11176 (N_11176,N_11028,N_10899);
and U11177 (N_11177,N_10962,N_10958);
or U11178 (N_11178,N_10919,N_10950);
or U11179 (N_11179,N_10903,N_11029);
nor U11180 (N_11180,N_10977,N_10893);
nand U11181 (N_11181,N_10886,N_10934);
nand U11182 (N_11182,N_11028,N_10897);
nand U11183 (N_11183,N_10887,N_11028);
and U11184 (N_11184,N_11017,N_10993);
or U11185 (N_11185,N_11024,N_10910);
and U11186 (N_11186,N_10999,N_10944);
and U11187 (N_11187,N_10964,N_10913);
and U11188 (N_11188,N_10907,N_10922);
or U11189 (N_11189,N_11029,N_10900);
nor U11190 (N_11190,N_10884,N_11033);
or U11191 (N_11191,N_10967,N_11019);
or U11192 (N_11192,N_11018,N_11015);
and U11193 (N_11193,N_11030,N_10979);
nand U11194 (N_11194,N_11006,N_10935);
and U11195 (N_11195,N_10892,N_11010);
and U11196 (N_11196,N_11005,N_10994);
nor U11197 (N_11197,N_10893,N_10887);
xnor U11198 (N_11198,N_10948,N_10926);
or U11199 (N_11199,N_10886,N_10905);
nor U11200 (N_11200,N_11178,N_11127);
or U11201 (N_11201,N_11074,N_11107);
or U11202 (N_11202,N_11045,N_11181);
or U11203 (N_11203,N_11059,N_11190);
xnor U11204 (N_11204,N_11093,N_11097);
or U11205 (N_11205,N_11069,N_11122);
nand U11206 (N_11206,N_11194,N_11163);
nor U11207 (N_11207,N_11049,N_11102);
nor U11208 (N_11208,N_11174,N_11098);
nand U11209 (N_11209,N_11100,N_11119);
nor U11210 (N_11210,N_11165,N_11058);
or U11211 (N_11211,N_11084,N_11179);
and U11212 (N_11212,N_11070,N_11088);
nor U11213 (N_11213,N_11180,N_11167);
nor U11214 (N_11214,N_11053,N_11048);
or U11215 (N_11215,N_11054,N_11162);
nand U11216 (N_11216,N_11067,N_11061);
and U11217 (N_11217,N_11136,N_11113);
nor U11218 (N_11218,N_11157,N_11191);
xnor U11219 (N_11219,N_11099,N_11160);
and U11220 (N_11220,N_11164,N_11175);
and U11221 (N_11221,N_11080,N_11065);
nor U11222 (N_11222,N_11135,N_11144);
and U11223 (N_11223,N_11117,N_11166);
and U11224 (N_11224,N_11124,N_11103);
and U11225 (N_11225,N_11159,N_11083);
and U11226 (N_11226,N_11156,N_11130);
nand U11227 (N_11227,N_11114,N_11056);
and U11228 (N_11228,N_11057,N_11068);
and U11229 (N_11229,N_11043,N_11185);
or U11230 (N_11230,N_11055,N_11063);
xor U11231 (N_11231,N_11052,N_11125);
and U11232 (N_11232,N_11196,N_11089);
nand U11233 (N_11233,N_11044,N_11077);
or U11234 (N_11234,N_11096,N_11133);
xor U11235 (N_11235,N_11072,N_11198);
and U11236 (N_11236,N_11140,N_11050);
nand U11237 (N_11237,N_11071,N_11172);
nor U11238 (N_11238,N_11195,N_11118);
nor U11239 (N_11239,N_11076,N_11197);
nor U11240 (N_11240,N_11108,N_11115);
nand U11241 (N_11241,N_11109,N_11128);
and U11242 (N_11242,N_11078,N_11134);
nand U11243 (N_11243,N_11051,N_11106);
nand U11244 (N_11244,N_11142,N_11101);
nand U11245 (N_11245,N_11139,N_11146);
nand U11246 (N_11246,N_11092,N_11090);
xnor U11247 (N_11247,N_11062,N_11105);
nand U11248 (N_11248,N_11155,N_11189);
nand U11249 (N_11249,N_11170,N_11132);
nand U11250 (N_11250,N_11147,N_11186);
xor U11251 (N_11251,N_11150,N_11040);
or U11252 (N_11252,N_11041,N_11199);
and U11253 (N_11253,N_11183,N_11046);
xnor U11254 (N_11254,N_11129,N_11066);
xnor U11255 (N_11255,N_11060,N_11104);
nand U11256 (N_11256,N_11047,N_11131);
or U11257 (N_11257,N_11171,N_11094);
nor U11258 (N_11258,N_11082,N_11042);
nor U11259 (N_11259,N_11192,N_11177);
and U11260 (N_11260,N_11075,N_11095);
nor U11261 (N_11261,N_11079,N_11087);
and U11262 (N_11262,N_11111,N_11158);
nand U11263 (N_11263,N_11154,N_11112);
nor U11264 (N_11264,N_11148,N_11184);
nand U11265 (N_11265,N_11152,N_11188);
xnor U11266 (N_11266,N_11081,N_11138);
nor U11267 (N_11267,N_11143,N_11169);
nand U11268 (N_11268,N_11121,N_11126);
and U11269 (N_11269,N_11073,N_11182);
nand U11270 (N_11270,N_11110,N_11137);
or U11271 (N_11271,N_11153,N_11161);
or U11272 (N_11272,N_11168,N_11085);
or U11273 (N_11273,N_11123,N_11091);
xor U11274 (N_11274,N_11187,N_11120);
nand U11275 (N_11275,N_11173,N_11116);
or U11276 (N_11276,N_11176,N_11086);
and U11277 (N_11277,N_11193,N_11151);
nand U11278 (N_11278,N_11145,N_11141);
or U11279 (N_11279,N_11064,N_11149);
or U11280 (N_11280,N_11140,N_11060);
nor U11281 (N_11281,N_11121,N_11155);
xnor U11282 (N_11282,N_11139,N_11064);
nor U11283 (N_11283,N_11043,N_11110);
or U11284 (N_11284,N_11184,N_11194);
nand U11285 (N_11285,N_11149,N_11110);
and U11286 (N_11286,N_11091,N_11147);
xor U11287 (N_11287,N_11104,N_11041);
xor U11288 (N_11288,N_11157,N_11118);
or U11289 (N_11289,N_11195,N_11064);
nor U11290 (N_11290,N_11044,N_11165);
nand U11291 (N_11291,N_11180,N_11099);
nand U11292 (N_11292,N_11045,N_11040);
nand U11293 (N_11293,N_11073,N_11084);
nor U11294 (N_11294,N_11114,N_11167);
nand U11295 (N_11295,N_11183,N_11061);
and U11296 (N_11296,N_11164,N_11134);
and U11297 (N_11297,N_11070,N_11074);
and U11298 (N_11298,N_11158,N_11057);
xor U11299 (N_11299,N_11064,N_11191);
and U11300 (N_11300,N_11136,N_11092);
nor U11301 (N_11301,N_11052,N_11152);
or U11302 (N_11302,N_11085,N_11182);
nand U11303 (N_11303,N_11146,N_11162);
or U11304 (N_11304,N_11183,N_11137);
or U11305 (N_11305,N_11157,N_11135);
or U11306 (N_11306,N_11116,N_11080);
nand U11307 (N_11307,N_11060,N_11198);
or U11308 (N_11308,N_11164,N_11111);
nor U11309 (N_11309,N_11070,N_11188);
and U11310 (N_11310,N_11149,N_11152);
nand U11311 (N_11311,N_11063,N_11118);
nand U11312 (N_11312,N_11086,N_11080);
nor U11313 (N_11313,N_11096,N_11139);
nor U11314 (N_11314,N_11060,N_11092);
or U11315 (N_11315,N_11148,N_11107);
or U11316 (N_11316,N_11199,N_11196);
or U11317 (N_11317,N_11191,N_11101);
xnor U11318 (N_11318,N_11162,N_11147);
and U11319 (N_11319,N_11097,N_11042);
and U11320 (N_11320,N_11180,N_11129);
nand U11321 (N_11321,N_11153,N_11125);
or U11322 (N_11322,N_11167,N_11178);
nand U11323 (N_11323,N_11132,N_11081);
nor U11324 (N_11324,N_11152,N_11060);
nand U11325 (N_11325,N_11064,N_11174);
nor U11326 (N_11326,N_11102,N_11098);
xor U11327 (N_11327,N_11194,N_11041);
nand U11328 (N_11328,N_11177,N_11155);
nand U11329 (N_11329,N_11072,N_11090);
or U11330 (N_11330,N_11068,N_11111);
xnor U11331 (N_11331,N_11068,N_11186);
nand U11332 (N_11332,N_11090,N_11121);
and U11333 (N_11333,N_11183,N_11053);
nor U11334 (N_11334,N_11050,N_11059);
and U11335 (N_11335,N_11192,N_11135);
or U11336 (N_11336,N_11144,N_11054);
nand U11337 (N_11337,N_11098,N_11139);
or U11338 (N_11338,N_11165,N_11158);
xnor U11339 (N_11339,N_11069,N_11046);
or U11340 (N_11340,N_11151,N_11132);
nand U11341 (N_11341,N_11101,N_11181);
and U11342 (N_11342,N_11083,N_11170);
and U11343 (N_11343,N_11049,N_11166);
nand U11344 (N_11344,N_11055,N_11162);
xor U11345 (N_11345,N_11157,N_11148);
or U11346 (N_11346,N_11069,N_11143);
nor U11347 (N_11347,N_11047,N_11184);
and U11348 (N_11348,N_11065,N_11041);
or U11349 (N_11349,N_11044,N_11116);
xnor U11350 (N_11350,N_11045,N_11055);
nor U11351 (N_11351,N_11057,N_11069);
or U11352 (N_11352,N_11062,N_11125);
nand U11353 (N_11353,N_11060,N_11159);
and U11354 (N_11354,N_11142,N_11116);
nor U11355 (N_11355,N_11072,N_11061);
nor U11356 (N_11356,N_11051,N_11056);
nand U11357 (N_11357,N_11093,N_11175);
and U11358 (N_11358,N_11078,N_11104);
or U11359 (N_11359,N_11067,N_11197);
nor U11360 (N_11360,N_11300,N_11331);
and U11361 (N_11361,N_11260,N_11201);
nand U11362 (N_11362,N_11269,N_11295);
and U11363 (N_11363,N_11253,N_11222);
and U11364 (N_11364,N_11213,N_11327);
nand U11365 (N_11365,N_11348,N_11310);
and U11366 (N_11366,N_11350,N_11321);
or U11367 (N_11367,N_11209,N_11204);
nor U11368 (N_11368,N_11234,N_11254);
or U11369 (N_11369,N_11340,N_11257);
or U11370 (N_11370,N_11330,N_11336);
nor U11371 (N_11371,N_11338,N_11273);
nor U11372 (N_11372,N_11217,N_11276);
or U11373 (N_11373,N_11332,N_11233);
xnor U11374 (N_11374,N_11344,N_11214);
nor U11375 (N_11375,N_11322,N_11270);
and U11376 (N_11376,N_11262,N_11268);
nor U11377 (N_11377,N_11290,N_11335);
nor U11378 (N_11378,N_11207,N_11337);
and U11379 (N_11379,N_11285,N_11242);
or U11380 (N_11380,N_11248,N_11232);
or U11381 (N_11381,N_11317,N_11357);
or U11382 (N_11382,N_11249,N_11216);
and U11383 (N_11383,N_11224,N_11354);
or U11384 (N_11384,N_11309,N_11359);
or U11385 (N_11385,N_11297,N_11293);
nand U11386 (N_11386,N_11333,N_11305);
nor U11387 (N_11387,N_11349,N_11205);
nand U11388 (N_11388,N_11200,N_11229);
and U11389 (N_11389,N_11313,N_11334);
nand U11390 (N_11390,N_11246,N_11311);
nand U11391 (N_11391,N_11235,N_11281);
or U11392 (N_11392,N_11292,N_11241);
or U11393 (N_11393,N_11264,N_11343);
nor U11394 (N_11394,N_11221,N_11261);
or U11395 (N_11395,N_11303,N_11324);
xor U11396 (N_11396,N_11284,N_11206);
or U11397 (N_11397,N_11315,N_11286);
nor U11398 (N_11398,N_11208,N_11223);
nor U11399 (N_11399,N_11237,N_11228);
xor U11400 (N_11400,N_11271,N_11258);
or U11401 (N_11401,N_11203,N_11266);
nor U11402 (N_11402,N_11318,N_11298);
xor U11403 (N_11403,N_11277,N_11226);
nand U11404 (N_11404,N_11274,N_11304);
nand U11405 (N_11405,N_11215,N_11356);
or U11406 (N_11406,N_11263,N_11265);
and U11407 (N_11407,N_11329,N_11325);
nor U11408 (N_11408,N_11220,N_11296);
nand U11409 (N_11409,N_11339,N_11251);
or U11410 (N_11410,N_11212,N_11308);
nand U11411 (N_11411,N_11288,N_11211);
or U11412 (N_11412,N_11275,N_11245);
and U11413 (N_11413,N_11231,N_11283);
or U11414 (N_11414,N_11239,N_11236);
xor U11415 (N_11415,N_11289,N_11219);
nor U11416 (N_11416,N_11225,N_11238);
or U11417 (N_11417,N_11341,N_11287);
xnor U11418 (N_11418,N_11279,N_11358);
nand U11419 (N_11419,N_11243,N_11347);
xor U11420 (N_11420,N_11355,N_11328);
or U11421 (N_11421,N_11272,N_11345);
xor U11422 (N_11422,N_11250,N_11316);
or U11423 (N_11423,N_11259,N_11247);
xnor U11424 (N_11424,N_11291,N_11326);
nand U11425 (N_11425,N_11306,N_11218);
nor U11426 (N_11426,N_11319,N_11210);
xnor U11427 (N_11427,N_11352,N_11267);
nand U11428 (N_11428,N_11312,N_11353);
nand U11429 (N_11429,N_11320,N_11301);
or U11430 (N_11430,N_11323,N_11346);
and U11431 (N_11431,N_11227,N_11302);
nor U11432 (N_11432,N_11282,N_11314);
nand U11433 (N_11433,N_11230,N_11278);
nor U11434 (N_11434,N_11202,N_11256);
nand U11435 (N_11435,N_11342,N_11294);
nor U11436 (N_11436,N_11280,N_11244);
and U11437 (N_11437,N_11240,N_11252);
nand U11438 (N_11438,N_11351,N_11255);
and U11439 (N_11439,N_11307,N_11299);
and U11440 (N_11440,N_11355,N_11236);
or U11441 (N_11441,N_11347,N_11228);
or U11442 (N_11442,N_11211,N_11297);
or U11443 (N_11443,N_11235,N_11234);
nand U11444 (N_11444,N_11205,N_11296);
or U11445 (N_11445,N_11328,N_11271);
nand U11446 (N_11446,N_11275,N_11299);
and U11447 (N_11447,N_11323,N_11295);
or U11448 (N_11448,N_11239,N_11216);
xor U11449 (N_11449,N_11220,N_11257);
or U11450 (N_11450,N_11336,N_11354);
xor U11451 (N_11451,N_11214,N_11216);
and U11452 (N_11452,N_11275,N_11322);
nand U11453 (N_11453,N_11282,N_11236);
nand U11454 (N_11454,N_11239,N_11232);
or U11455 (N_11455,N_11231,N_11334);
nand U11456 (N_11456,N_11247,N_11236);
nand U11457 (N_11457,N_11286,N_11204);
xnor U11458 (N_11458,N_11341,N_11257);
xor U11459 (N_11459,N_11309,N_11305);
nor U11460 (N_11460,N_11281,N_11302);
or U11461 (N_11461,N_11287,N_11328);
or U11462 (N_11462,N_11354,N_11257);
or U11463 (N_11463,N_11300,N_11334);
xor U11464 (N_11464,N_11343,N_11218);
nand U11465 (N_11465,N_11231,N_11307);
or U11466 (N_11466,N_11294,N_11290);
nor U11467 (N_11467,N_11268,N_11204);
and U11468 (N_11468,N_11327,N_11218);
nand U11469 (N_11469,N_11277,N_11208);
nor U11470 (N_11470,N_11257,N_11351);
or U11471 (N_11471,N_11301,N_11227);
nor U11472 (N_11472,N_11221,N_11342);
nand U11473 (N_11473,N_11326,N_11202);
nand U11474 (N_11474,N_11277,N_11261);
or U11475 (N_11475,N_11247,N_11346);
nor U11476 (N_11476,N_11332,N_11331);
nor U11477 (N_11477,N_11234,N_11296);
or U11478 (N_11478,N_11320,N_11324);
or U11479 (N_11479,N_11232,N_11230);
nand U11480 (N_11480,N_11285,N_11209);
or U11481 (N_11481,N_11247,N_11204);
xor U11482 (N_11482,N_11313,N_11321);
nand U11483 (N_11483,N_11292,N_11281);
xor U11484 (N_11484,N_11313,N_11246);
and U11485 (N_11485,N_11343,N_11233);
or U11486 (N_11486,N_11209,N_11279);
xnor U11487 (N_11487,N_11280,N_11205);
xor U11488 (N_11488,N_11255,N_11304);
nand U11489 (N_11489,N_11257,N_11269);
and U11490 (N_11490,N_11356,N_11307);
or U11491 (N_11491,N_11316,N_11315);
nand U11492 (N_11492,N_11317,N_11208);
nand U11493 (N_11493,N_11210,N_11229);
or U11494 (N_11494,N_11294,N_11201);
or U11495 (N_11495,N_11339,N_11202);
nor U11496 (N_11496,N_11328,N_11278);
and U11497 (N_11497,N_11359,N_11338);
and U11498 (N_11498,N_11282,N_11267);
nand U11499 (N_11499,N_11315,N_11232);
nand U11500 (N_11500,N_11262,N_11263);
or U11501 (N_11501,N_11262,N_11318);
nand U11502 (N_11502,N_11334,N_11296);
and U11503 (N_11503,N_11328,N_11347);
xnor U11504 (N_11504,N_11328,N_11303);
xnor U11505 (N_11505,N_11321,N_11311);
nor U11506 (N_11506,N_11202,N_11320);
or U11507 (N_11507,N_11288,N_11216);
nor U11508 (N_11508,N_11324,N_11340);
nand U11509 (N_11509,N_11286,N_11331);
xnor U11510 (N_11510,N_11244,N_11290);
nand U11511 (N_11511,N_11358,N_11212);
and U11512 (N_11512,N_11201,N_11303);
nor U11513 (N_11513,N_11207,N_11287);
and U11514 (N_11514,N_11328,N_11317);
nor U11515 (N_11515,N_11344,N_11209);
xnor U11516 (N_11516,N_11266,N_11342);
and U11517 (N_11517,N_11233,N_11315);
nor U11518 (N_11518,N_11309,N_11276);
or U11519 (N_11519,N_11359,N_11211);
and U11520 (N_11520,N_11393,N_11517);
and U11521 (N_11521,N_11409,N_11515);
or U11522 (N_11522,N_11400,N_11480);
xor U11523 (N_11523,N_11428,N_11443);
or U11524 (N_11524,N_11383,N_11495);
and U11525 (N_11525,N_11473,N_11445);
and U11526 (N_11526,N_11377,N_11469);
and U11527 (N_11527,N_11430,N_11474);
nor U11528 (N_11528,N_11432,N_11508);
or U11529 (N_11529,N_11494,N_11498);
or U11530 (N_11530,N_11361,N_11388);
nand U11531 (N_11531,N_11437,N_11424);
nand U11532 (N_11532,N_11435,N_11419);
nor U11533 (N_11533,N_11425,N_11512);
and U11534 (N_11534,N_11470,N_11457);
or U11535 (N_11535,N_11399,N_11458);
or U11536 (N_11536,N_11504,N_11387);
nor U11537 (N_11537,N_11362,N_11496);
and U11538 (N_11538,N_11446,N_11472);
xnor U11539 (N_11539,N_11415,N_11374);
nor U11540 (N_11540,N_11366,N_11444);
nand U11541 (N_11541,N_11367,N_11489);
and U11542 (N_11542,N_11396,N_11441);
and U11543 (N_11543,N_11509,N_11394);
nor U11544 (N_11544,N_11418,N_11410);
nand U11545 (N_11545,N_11483,N_11385);
and U11546 (N_11546,N_11365,N_11510);
nand U11547 (N_11547,N_11384,N_11406);
nor U11548 (N_11548,N_11392,N_11461);
nor U11549 (N_11549,N_11395,N_11481);
nor U11550 (N_11550,N_11364,N_11370);
or U11551 (N_11551,N_11466,N_11513);
nor U11552 (N_11552,N_11368,N_11511);
and U11553 (N_11553,N_11401,N_11405);
or U11554 (N_11554,N_11417,N_11454);
and U11555 (N_11555,N_11493,N_11500);
nand U11556 (N_11556,N_11372,N_11397);
or U11557 (N_11557,N_11439,N_11423);
nand U11558 (N_11558,N_11412,N_11416);
and U11559 (N_11559,N_11478,N_11440);
or U11560 (N_11560,N_11518,N_11468);
nand U11561 (N_11561,N_11452,N_11465);
or U11562 (N_11562,N_11507,N_11413);
and U11563 (N_11563,N_11476,N_11408);
nand U11564 (N_11564,N_11464,N_11485);
nor U11565 (N_11565,N_11502,N_11456);
or U11566 (N_11566,N_11363,N_11360);
xnor U11567 (N_11567,N_11514,N_11450);
nand U11568 (N_11568,N_11404,N_11421);
xor U11569 (N_11569,N_11488,N_11375);
nor U11570 (N_11570,N_11453,N_11422);
nor U11571 (N_11571,N_11433,N_11369);
xnor U11572 (N_11572,N_11391,N_11390);
nand U11573 (N_11573,N_11497,N_11492);
nand U11574 (N_11574,N_11462,N_11379);
or U11575 (N_11575,N_11447,N_11477);
and U11576 (N_11576,N_11484,N_11482);
nand U11577 (N_11577,N_11519,N_11427);
nor U11578 (N_11578,N_11503,N_11426);
xor U11579 (N_11579,N_11436,N_11438);
xor U11580 (N_11580,N_11455,N_11491);
nand U11581 (N_11581,N_11380,N_11506);
or U11582 (N_11582,N_11449,N_11486);
nor U11583 (N_11583,N_11402,N_11411);
xnor U11584 (N_11584,N_11448,N_11442);
nand U11585 (N_11585,N_11463,N_11516);
and U11586 (N_11586,N_11451,N_11487);
xor U11587 (N_11587,N_11414,N_11371);
or U11588 (N_11588,N_11389,N_11467);
xor U11589 (N_11589,N_11460,N_11471);
or U11590 (N_11590,N_11475,N_11501);
xor U11591 (N_11591,N_11403,N_11382);
and U11592 (N_11592,N_11505,N_11420);
and U11593 (N_11593,N_11376,N_11434);
and U11594 (N_11594,N_11407,N_11429);
xor U11595 (N_11595,N_11381,N_11459);
nor U11596 (N_11596,N_11378,N_11490);
nand U11597 (N_11597,N_11386,N_11499);
nand U11598 (N_11598,N_11479,N_11398);
and U11599 (N_11599,N_11373,N_11431);
xnor U11600 (N_11600,N_11432,N_11392);
or U11601 (N_11601,N_11401,N_11373);
nand U11602 (N_11602,N_11364,N_11504);
and U11603 (N_11603,N_11367,N_11426);
nand U11604 (N_11604,N_11497,N_11503);
xor U11605 (N_11605,N_11452,N_11468);
or U11606 (N_11606,N_11421,N_11392);
nor U11607 (N_11607,N_11377,N_11376);
or U11608 (N_11608,N_11365,N_11505);
nand U11609 (N_11609,N_11383,N_11502);
xnor U11610 (N_11610,N_11434,N_11444);
nor U11611 (N_11611,N_11505,N_11461);
and U11612 (N_11612,N_11404,N_11484);
nor U11613 (N_11613,N_11437,N_11390);
nand U11614 (N_11614,N_11430,N_11379);
nor U11615 (N_11615,N_11452,N_11517);
nand U11616 (N_11616,N_11459,N_11437);
or U11617 (N_11617,N_11445,N_11511);
and U11618 (N_11618,N_11385,N_11501);
or U11619 (N_11619,N_11482,N_11432);
nor U11620 (N_11620,N_11511,N_11420);
xor U11621 (N_11621,N_11380,N_11419);
nor U11622 (N_11622,N_11472,N_11512);
nand U11623 (N_11623,N_11415,N_11393);
or U11624 (N_11624,N_11447,N_11435);
nor U11625 (N_11625,N_11448,N_11374);
or U11626 (N_11626,N_11462,N_11360);
nand U11627 (N_11627,N_11414,N_11368);
xnor U11628 (N_11628,N_11416,N_11361);
and U11629 (N_11629,N_11498,N_11518);
xor U11630 (N_11630,N_11415,N_11398);
or U11631 (N_11631,N_11455,N_11503);
or U11632 (N_11632,N_11461,N_11437);
nor U11633 (N_11633,N_11360,N_11474);
and U11634 (N_11634,N_11438,N_11394);
or U11635 (N_11635,N_11445,N_11368);
and U11636 (N_11636,N_11372,N_11366);
or U11637 (N_11637,N_11431,N_11368);
or U11638 (N_11638,N_11481,N_11375);
or U11639 (N_11639,N_11481,N_11486);
nor U11640 (N_11640,N_11419,N_11492);
nand U11641 (N_11641,N_11460,N_11378);
or U11642 (N_11642,N_11421,N_11361);
and U11643 (N_11643,N_11490,N_11462);
xnor U11644 (N_11644,N_11380,N_11502);
nand U11645 (N_11645,N_11469,N_11398);
or U11646 (N_11646,N_11377,N_11420);
and U11647 (N_11647,N_11477,N_11496);
xnor U11648 (N_11648,N_11422,N_11417);
nor U11649 (N_11649,N_11395,N_11401);
nor U11650 (N_11650,N_11401,N_11463);
nor U11651 (N_11651,N_11376,N_11362);
nor U11652 (N_11652,N_11474,N_11516);
nand U11653 (N_11653,N_11503,N_11454);
or U11654 (N_11654,N_11366,N_11410);
nand U11655 (N_11655,N_11484,N_11435);
and U11656 (N_11656,N_11449,N_11465);
and U11657 (N_11657,N_11366,N_11464);
or U11658 (N_11658,N_11381,N_11376);
nor U11659 (N_11659,N_11497,N_11474);
and U11660 (N_11660,N_11426,N_11446);
xor U11661 (N_11661,N_11494,N_11403);
nand U11662 (N_11662,N_11509,N_11488);
or U11663 (N_11663,N_11475,N_11496);
xor U11664 (N_11664,N_11493,N_11409);
nor U11665 (N_11665,N_11389,N_11455);
nand U11666 (N_11666,N_11461,N_11509);
or U11667 (N_11667,N_11496,N_11429);
nor U11668 (N_11668,N_11400,N_11391);
and U11669 (N_11669,N_11425,N_11498);
or U11670 (N_11670,N_11459,N_11424);
nand U11671 (N_11671,N_11437,N_11402);
and U11672 (N_11672,N_11518,N_11466);
and U11673 (N_11673,N_11459,N_11404);
and U11674 (N_11674,N_11419,N_11485);
nor U11675 (N_11675,N_11367,N_11401);
xor U11676 (N_11676,N_11499,N_11382);
nor U11677 (N_11677,N_11382,N_11444);
nand U11678 (N_11678,N_11429,N_11501);
and U11679 (N_11679,N_11416,N_11446);
nor U11680 (N_11680,N_11562,N_11663);
nand U11681 (N_11681,N_11563,N_11661);
nand U11682 (N_11682,N_11605,N_11664);
and U11683 (N_11683,N_11676,N_11523);
nand U11684 (N_11684,N_11608,N_11577);
or U11685 (N_11685,N_11620,N_11611);
or U11686 (N_11686,N_11542,N_11596);
nor U11687 (N_11687,N_11649,N_11555);
and U11688 (N_11688,N_11547,N_11591);
and U11689 (N_11689,N_11554,N_11616);
and U11690 (N_11690,N_11597,N_11643);
nor U11691 (N_11691,N_11646,N_11625);
nand U11692 (N_11692,N_11668,N_11535);
xor U11693 (N_11693,N_11536,N_11581);
nor U11694 (N_11694,N_11524,N_11594);
nor U11695 (N_11695,N_11624,N_11585);
nand U11696 (N_11696,N_11635,N_11565);
nor U11697 (N_11697,N_11614,N_11607);
or U11698 (N_11698,N_11595,N_11651);
nand U11699 (N_11699,N_11539,N_11604);
or U11700 (N_11700,N_11574,N_11618);
and U11701 (N_11701,N_11546,N_11582);
xor U11702 (N_11702,N_11670,N_11675);
xnor U11703 (N_11703,N_11568,N_11576);
nand U11704 (N_11704,N_11601,N_11575);
and U11705 (N_11705,N_11525,N_11650);
nor U11706 (N_11706,N_11619,N_11590);
and U11707 (N_11707,N_11677,N_11580);
xnor U11708 (N_11708,N_11659,N_11667);
and U11709 (N_11709,N_11522,N_11612);
and U11710 (N_11710,N_11660,N_11615);
nand U11711 (N_11711,N_11630,N_11537);
nor U11712 (N_11712,N_11672,N_11598);
and U11713 (N_11713,N_11533,N_11556);
and U11714 (N_11714,N_11665,N_11566);
and U11715 (N_11715,N_11636,N_11527);
nand U11716 (N_11716,N_11540,N_11632);
nand U11717 (N_11717,N_11586,N_11674);
and U11718 (N_11718,N_11617,N_11606);
nand U11719 (N_11719,N_11633,N_11631);
and U11720 (N_11720,N_11629,N_11645);
xor U11721 (N_11721,N_11571,N_11623);
and U11722 (N_11722,N_11621,N_11573);
or U11723 (N_11723,N_11641,N_11553);
and U11724 (N_11724,N_11609,N_11521);
xnor U11725 (N_11725,N_11543,N_11678);
and U11726 (N_11726,N_11648,N_11671);
or U11727 (N_11727,N_11587,N_11529);
nand U11728 (N_11728,N_11532,N_11579);
nand U11729 (N_11729,N_11558,N_11541);
nor U11730 (N_11730,N_11679,N_11530);
or U11731 (N_11731,N_11600,N_11572);
nor U11732 (N_11732,N_11610,N_11531);
nor U11733 (N_11733,N_11602,N_11640);
nand U11734 (N_11734,N_11652,N_11569);
or U11735 (N_11735,N_11528,N_11526);
nand U11736 (N_11736,N_11638,N_11538);
nor U11737 (N_11737,N_11545,N_11657);
nand U11738 (N_11738,N_11551,N_11626);
nor U11739 (N_11739,N_11666,N_11662);
or U11740 (N_11740,N_11628,N_11642);
or U11741 (N_11741,N_11550,N_11658);
xor U11742 (N_11742,N_11639,N_11549);
and U11743 (N_11743,N_11655,N_11588);
and U11744 (N_11744,N_11561,N_11634);
xor U11745 (N_11745,N_11560,N_11564);
or U11746 (N_11746,N_11603,N_11599);
or U11747 (N_11747,N_11654,N_11559);
and U11748 (N_11748,N_11544,N_11589);
nand U11749 (N_11749,N_11592,N_11593);
and U11750 (N_11750,N_11583,N_11584);
nand U11751 (N_11751,N_11557,N_11534);
and U11752 (N_11752,N_11653,N_11578);
nand U11753 (N_11753,N_11637,N_11552);
nor U11754 (N_11754,N_11673,N_11622);
nor U11755 (N_11755,N_11669,N_11647);
or U11756 (N_11756,N_11570,N_11644);
nor U11757 (N_11757,N_11520,N_11627);
xor U11758 (N_11758,N_11656,N_11613);
nand U11759 (N_11759,N_11567,N_11548);
nor U11760 (N_11760,N_11665,N_11634);
or U11761 (N_11761,N_11634,N_11607);
nor U11762 (N_11762,N_11525,N_11653);
and U11763 (N_11763,N_11616,N_11572);
nand U11764 (N_11764,N_11552,N_11596);
or U11765 (N_11765,N_11673,N_11581);
xor U11766 (N_11766,N_11663,N_11667);
nor U11767 (N_11767,N_11624,N_11630);
or U11768 (N_11768,N_11584,N_11577);
or U11769 (N_11769,N_11599,N_11658);
nand U11770 (N_11770,N_11558,N_11632);
xnor U11771 (N_11771,N_11638,N_11596);
nand U11772 (N_11772,N_11598,N_11593);
nand U11773 (N_11773,N_11619,N_11645);
nand U11774 (N_11774,N_11605,N_11550);
or U11775 (N_11775,N_11650,N_11543);
nand U11776 (N_11776,N_11637,N_11622);
or U11777 (N_11777,N_11641,N_11534);
nor U11778 (N_11778,N_11608,N_11547);
or U11779 (N_11779,N_11545,N_11559);
or U11780 (N_11780,N_11620,N_11621);
nand U11781 (N_11781,N_11669,N_11664);
nand U11782 (N_11782,N_11555,N_11630);
nor U11783 (N_11783,N_11570,N_11582);
nor U11784 (N_11784,N_11591,N_11654);
and U11785 (N_11785,N_11609,N_11643);
nor U11786 (N_11786,N_11659,N_11603);
nor U11787 (N_11787,N_11531,N_11671);
nand U11788 (N_11788,N_11604,N_11662);
nand U11789 (N_11789,N_11636,N_11535);
and U11790 (N_11790,N_11529,N_11635);
and U11791 (N_11791,N_11663,N_11607);
or U11792 (N_11792,N_11551,N_11641);
nor U11793 (N_11793,N_11607,N_11553);
and U11794 (N_11794,N_11575,N_11524);
nand U11795 (N_11795,N_11563,N_11621);
nor U11796 (N_11796,N_11666,N_11621);
nor U11797 (N_11797,N_11600,N_11664);
nand U11798 (N_11798,N_11549,N_11612);
and U11799 (N_11799,N_11598,N_11654);
or U11800 (N_11800,N_11586,N_11676);
and U11801 (N_11801,N_11641,N_11608);
and U11802 (N_11802,N_11594,N_11674);
or U11803 (N_11803,N_11592,N_11658);
and U11804 (N_11804,N_11620,N_11609);
nand U11805 (N_11805,N_11651,N_11552);
and U11806 (N_11806,N_11564,N_11676);
or U11807 (N_11807,N_11673,N_11604);
nor U11808 (N_11808,N_11593,N_11605);
nand U11809 (N_11809,N_11599,N_11544);
and U11810 (N_11810,N_11604,N_11558);
and U11811 (N_11811,N_11523,N_11565);
nor U11812 (N_11812,N_11574,N_11632);
nand U11813 (N_11813,N_11631,N_11637);
and U11814 (N_11814,N_11623,N_11558);
nor U11815 (N_11815,N_11614,N_11538);
nand U11816 (N_11816,N_11543,N_11608);
nor U11817 (N_11817,N_11534,N_11649);
nor U11818 (N_11818,N_11578,N_11599);
nor U11819 (N_11819,N_11527,N_11547);
or U11820 (N_11820,N_11655,N_11657);
nand U11821 (N_11821,N_11539,N_11568);
nand U11822 (N_11822,N_11528,N_11543);
xnor U11823 (N_11823,N_11669,N_11637);
nor U11824 (N_11824,N_11543,N_11545);
or U11825 (N_11825,N_11622,N_11649);
or U11826 (N_11826,N_11521,N_11673);
nand U11827 (N_11827,N_11603,N_11527);
or U11828 (N_11828,N_11570,N_11621);
nand U11829 (N_11829,N_11624,N_11669);
or U11830 (N_11830,N_11527,N_11561);
nor U11831 (N_11831,N_11668,N_11583);
nor U11832 (N_11832,N_11601,N_11537);
and U11833 (N_11833,N_11522,N_11672);
or U11834 (N_11834,N_11581,N_11583);
and U11835 (N_11835,N_11660,N_11572);
nand U11836 (N_11836,N_11625,N_11583);
and U11837 (N_11837,N_11558,N_11675);
nand U11838 (N_11838,N_11588,N_11604);
or U11839 (N_11839,N_11571,N_11598);
or U11840 (N_11840,N_11750,N_11809);
or U11841 (N_11841,N_11740,N_11710);
xnor U11842 (N_11842,N_11813,N_11702);
or U11843 (N_11843,N_11807,N_11780);
and U11844 (N_11844,N_11788,N_11776);
nand U11845 (N_11845,N_11681,N_11821);
xor U11846 (N_11846,N_11798,N_11783);
or U11847 (N_11847,N_11696,N_11730);
xor U11848 (N_11848,N_11699,N_11722);
and U11849 (N_11849,N_11820,N_11723);
nor U11850 (N_11850,N_11727,N_11773);
or U11851 (N_11851,N_11705,N_11703);
nor U11852 (N_11852,N_11759,N_11801);
nand U11853 (N_11853,N_11683,N_11735);
nor U11854 (N_11854,N_11717,N_11767);
nand U11855 (N_11855,N_11824,N_11778);
nand U11856 (N_11856,N_11785,N_11802);
nor U11857 (N_11857,N_11694,N_11770);
nand U11858 (N_11858,N_11834,N_11704);
nand U11859 (N_11859,N_11713,N_11764);
or U11860 (N_11860,N_11791,N_11836);
nand U11861 (N_11861,N_11760,N_11706);
and U11862 (N_11862,N_11823,N_11726);
or U11863 (N_11863,N_11810,N_11765);
xnor U11864 (N_11864,N_11736,N_11769);
and U11865 (N_11865,N_11757,N_11800);
or U11866 (N_11866,N_11748,N_11733);
xor U11867 (N_11867,N_11805,N_11701);
or U11868 (N_11868,N_11732,N_11734);
or U11869 (N_11869,N_11691,N_11728);
nor U11870 (N_11870,N_11711,N_11777);
or U11871 (N_11871,N_11793,N_11754);
or U11872 (N_11872,N_11761,N_11787);
xor U11873 (N_11873,N_11827,N_11781);
nor U11874 (N_11874,N_11689,N_11693);
nor U11875 (N_11875,N_11816,N_11811);
or U11876 (N_11876,N_11737,N_11774);
and U11877 (N_11877,N_11687,N_11818);
or U11878 (N_11878,N_11690,N_11839);
nor U11879 (N_11879,N_11744,N_11747);
or U11880 (N_11880,N_11753,N_11775);
nand U11881 (N_11881,N_11692,N_11831);
or U11882 (N_11882,N_11719,N_11804);
and U11883 (N_11883,N_11822,N_11790);
nand U11884 (N_11884,N_11731,N_11738);
xnor U11885 (N_11885,N_11797,N_11712);
or U11886 (N_11886,N_11743,N_11806);
nand U11887 (N_11887,N_11838,N_11799);
xor U11888 (N_11888,N_11718,N_11755);
xnor U11889 (N_11889,N_11794,N_11763);
and U11890 (N_11890,N_11795,N_11758);
nor U11891 (N_11891,N_11784,N_11762);
and U11892 (N_11892,N_11749,N_11720);
nand U11893 (N_11893,N_11779,N_11782);
nand U11894 (N_11894,N_11746,N_11721);
xor U11895 (N_11895,N_11826,N_11830);
xnor U11896 (N_11896,N_11837,N_11808);
nor U11897 (N_11897,N_11829,N_11825);
and U11898 (N_11898,N_11698,N_11686);
or U11899 (N_11899,N_11715,N_11796);
nor U11900 (N_11900,N_11803,N_11814);
nor U11901 (N_11901,N_11697,N_11771);
nand U11902 (N_11902,N_11684,N_11708);
nor U11903 (N_11903,N_11819,N_11709);
or U11904 (N_11904,N_11741,N_11768);
and U11905 (N_11905,N_11786,N_11828);
or U11906 (N_11906,N_11685,N_11739);
or U11907 (N_11907,N_11792,N_11729);
xor U11908 (N_11908,N_11833,N_11766);
or U11909 (N_11909,N_11832,N_11745);
nor U11910 (N_11910,N_11695,N_11815);
and U11911 (N_11911,N_11751,N_11714);
or U11912 (N_11912,N_11812,N_11817);
nor U11913 (N_11913,N_11688,N_11789);
and U11914 (N_11914,N_11680,N_11716);
nand U11915 (N_11915,N_11835,N_11772);
xnor U11916 (N_11916,N_11752,N_11707);
xor U11917 (N_11917,N_11742,N_11682);
xnor U11918 (N_11918,N_11756,N_11724);
or U11919 (N_11919,N_11725,N_11700);
nand U11920 (N_11920,N_11759,N_11732);
or U11921 (N_11921,N_11717,N_11822);
nor U11922 (N_11922,N_11752,N_11700);
nand U11923 (N_11923,N_11728,N_11789);
or U11924 (N_11924,N_11832,N_11827);
nand U11925 (N_11925,N_11767,N_11782);
nor U11926 (N_11926,N_11742,N_11805);
or U11927 (N_11927,N_11725,N_11769);
and U11928 (N_11928,N_11811,N_11684);
and U11929 (N_11929,N_11831,N_11720);
or U11930 (N_11930,N_11837,N_11704);
nand U11931 (N_11931,N_11813,N_11680);
nand U11932 (N_11932,N_11734,N_11690);
nand U11933 (N_11933,N_11776,N_11700);
or U11934 (N_11934,N_11687,N_11777);
and U11935 (N_11935,N_11822,N_11796);
and U11936 (N_11936,N_11815,N_11684);
or U11937 (N_11937,N_11808,N_11818);
and U11938 (N_11938,N_11821,N_11709);
nor U11939 (N_11939,N_11820,N_11761);
xor U11940 (N_11940,N_11744,N_11746);
and U11941 (N_11941,N_11719,N_11750);
nor U11942 (N_11942,N_11787,N_11767);
and U11943 (N_11943,N_11689,N_11831);
nand U11944 (N_11944,N_11760,N_11782);
and U11945 (N_11945,N_11720,N_11695);
and U11946 (N_11946,N_11756,N_11723);
or U11947 (N_11947,N_11803,N_11737);
nor U11948 (N_11948,N_11803,N_11712);
nor U11949 (N_11949,N_11711,N_11739);
and U11950 (N_11950,N_11831,N_11694);
nor U11951 (N_11951,N_11737,N_11816);
nor U11952 (N_11952,N_11799,N_11701);
nand U11953 (N_11953,N_11681,N_11788);
and U11954 (N_11954,N_11788,N_11695);
or U11955 (N_11955,N_11793,N_11837);
xnor U11956 (N_11956,N_11822,N_11768);
xor U11957 (N_11957,N_11730,N_11682);
nor U11958 (N_11958,N_11738,N_11720);
or U11959 (N_11959,N_11709,N_11686);
and U11960 (N_11960,N_11823,N_11813);
nand U11961 (N_11961,N_11713,N_11754);
nor U11962 (N_11962,N_11753,N_11723);
xor U11963 (N_11963,N_11738,N_11766);
nor U11964 (N_11964,N_11723,N_11744);
or U11965 (N_11965,N_11807,N_11822);
and U11966 (N_11966,N_11778,N_11691);
nor U11967 (N_11967,N_11791,N_11818);
and U11968 (N_11968,N_11726,N_11754);
nor U11969 (N_11969,N_11708,N_11779);
nor U11970 (N_11970,N_11803,N_11688);
nor U11971 (N_11971,N_11835,N_11764);
or U11972 (N_11972,N_11836,N_11837);
nor U11973 (N_11973,N_11710,N_11806);
or U11974 (N_11974,N_11691,N_11697);
and U11975 (N_11975,N_11741,N_11709);
and U11976 (N_11976,N_11784,N_11716);
and U11977 (N_11977,N_11794,N_11739);
and U11978 (N_11978,N_11829,N_11746);
nand U11979 (N_11979,N_11708,N_11816);
nand U11980 (N_11980,N_11802,N_11814);
nor U11981 (N_11981,N_11813,N_11689);
nand U11982 (N_11982,N_11743,N_11776);
and U11983 (N_11983,N_11703,N_11759);
nor U11984 (N_11984,N_11741,N_11773);
and U11985 (N_11985,N_11682,N_11739);
and U11986 (N_11986,N_11754,N_11685);
nor U11987 (N_11987,N_11781,N_11685);
nor U11988 (N_11988,N_11810,N_11685);
and U11989 (N_11989,N_11791,N_11802);
and U11990 (N_11990,N_11681,N_11703);
nor U11991 (N_11991,N_11788,N_11796);
and U11992 (N_11992,N_11827,N_11784);
nor U11993 (N_11993,N_11816,N_11832);
or U11994 (N_11994,N_11748,N_11737);
nor U11995 (N_11995,N_11779,N_11772);
nor U11996 (N_11996,N_11828,N_11741);
and U11997 (N_11997,N_11818,N_11825);
nor U11998 (N_11998,N_11708,N_11811);
nor U11999 (N_11999,N_11814,N_11692);
nand U12000 (N_12000,N_11994,N_11982);
or U12001 (N_12001,N_11962,N_11853);
nand U12002 (N_12002,N_11913,N_11972);
xnor U12003 (N_12003,N_11965,N_11996);
or U12004 (N_12004,N_11867,N_11969);
or U12005 (N_12005,N_11874,N_11984);
and U12006 (N_12006,N_11882,N_11912);
nor U12007 (N_12007,N_11904,N_11907);
nand U12008 (N_12008,N_11918,N_11959);
nor U12009 (N_12009,N_11983,N_11860);
nor U12010 (N_12010,N_11850,N_11910);
or U12011 (N_12011,N_11854,N_11875);
xor U12012 (N_12012,N_11990,N_11968);
and U12013 (N_12013,N_11845,N_11976);
xnor U12014 (N_12014,N_11942,N_11946);
and U12015 (N_12015,N_11920,N_11840);
or U12016 (N_12016,N_11916,N_11967);
and U12017 (N_12017,N_11985,N_11899);
nand U12018 (N_12018,N_11950,N_11883);
or U12019 (N_12019,N_11973,N_11865);
xor U12020 (N_12020,N_11940,N_11851);
or U12021 (N_12021,N_11905,N_11914);
nand U12022 (N_12022,N_11919,N_11892);
nor U12023 (N_12023,N_11992,N_11862);
nand U12024 (N_12024,N_11906,N_11869);
nor U12025 (N_12025,N_11885,N_11980);
nor U12026 (N_12026,N_11966,N_11929);
or U12027 (N_12027,N_11847,N_11997);
or U12028 (N_12028,N_11975,N_11931);
or U12029 (N_12029,N_11995,N_11872);
nand U12030 (N_12030,N_11936,N_11954);
and U12031 (N_12031,N_11897,N_11871);
and U12032 (N_12032,N_11844,N_11999);
xnor U12033 (N_12033,N_11848,N_11998);
nand U12034 (N_12034,N_11970,N_11981);
nand U12035 (N_12035,N_11925,N_11900);
nand U12036 (N_12036,N_11974,N_11879);
nor U12037 (N_12037,N_11941,N_11877);
and U12038 (N_12038,N_11961,N_11955);
and U12039 (N_12039,N_11988,N_11934);
and U12040 (N_12040,N_11891,N_11949);
nand U12041 (N_12041,N_11911,N_11889);
xnor U12042 (N_12042,N_11932,N_11937);
or U12043 (N_12043,N_11846,N_11873);
nand U12044 (N_12044,N_11902,N_11922);
xor U12045 (N_12045,N_11855,N_11939);
nand U12046 (N_12046,N_11858,N_11887);
and U12047 (N_12047,N_11886,N_11948);
xor U12048 (N_12048,N_11977,N_11963);
nand U12049 (N_12049,N_11868,N_11933);
nand U12050 (N_12050,N_11958,N_11993);
nor U12051 (N_12051,N_11987,N_11951);
nor U12052 (N_12052,N_11866,N_11878);
nand U12053 (N_12053,N_11927,N_11895);
or U12054 (N_12054,N_11896,N_11928);
or U12055 (N_12055,N_11903,N_11861);
nand U12056 (N_12056,N_11971,N_11841);
and U12057 (N_12057,N_11870,N_11842);
nor U12058 (N_12058,N_11864,N_11978);
nand U12059 (N_12059,N_11947,N_11849);
nand U12060 (N_12060,N_11888,N_11893);
and U12061 (N_12061,N_11857,N_11930);
and U12062 (N_12062,N_11923,N_11952);
nor U12063 (N_12063,N_11956,N_11859);
nor U12064 (N_12064,N_11960,N_11880);
or U12065 (N_12065,N_11915,N_11979);
nand U12066 (N_12066,N_11964,N_11890);
nand U12067 (N_12067,N_11943,N_11991);
and U12068 (N_12068,N_11852,N_11945);
nand U12069 (N_12069,N_11909,N_11924);
or U12070 (N_12070,N_11957,N_11898);
and U12071 (N_12071,N_11944,N_11926);
or U12072 (N_12072,N_11881,N_11938);
nor U12073 (N_12073,N_11856,N_11901);
or U12074 (N_12074,N_11894,N_11908);
and U12075 (N_12075,N_11986,N_11917);
and U12076 (N_12076,N_11843,N_11921);
nand U12077 (N_12077,N_11863,N_11989);
xor U12078 (N_12078,N_11953,N_11884);
or U12079 (N_12079,N_11935,N_11876);
or U12080 (N_12080,N_11975,N_11951);
and U12081 (N_12081,N_11901,N_11926);
nor U12082 (N_12082,N_11854,N_11963);
nor U12083 (N_12083,N_11866,N_11873);
and U12084 (N_12084,N_11910,N_11980);
and U12085 (N_12085,N_11931,N_11870);
xnor U12086 (N_12086,N_11996,N_11941);
nor U12087 (N_12087,N_11844,N_11908);
nor U12088 (N_12088,N_11965,N_11840);
nor U12089 (N_12089,N_11872,N_11844);
nand U12090 (N_12090,N_11942,N_11963);
or U12091 (N_12091,N_11998,N_11874);
or U12092 (N_12092,N_11867,N_11863);
nor U12093 (N_12093,N_11914,N_11853);
nand U12094 (N_12094,N_11952,N_11964);
or U12095 (N_12095,N_11922,N_11982);
and U12096 (N_12096,N_11949,N_11970);
or U12097 (N_12097,N_11963,N_11904);
nand U12098 (N_12098,N_11867,N_11849);
and U12099 (N_12099,N_11897,N_11863);
and U12100 (N_12100,N_11866,N_11999);
and U12101 (N_12101,N_11937,N_11910);
nand U12102 (N_12102,N_11898,N_11965);
nor U12103 (N_12103,N_11923,N_11956);
nor U12104 (N_12104,N_11951,N_11874);
nand U12105 (N_12105,N_11919,N_11887);
nand U12106 (N_12106,N_11936,N_11876);
and U12107 (N_12107,N_11990,N_11991);
nor U12108 (N_12108,N_11992,N_11852);
xor U12109 (N_12109,N_11975,N_11867);
and U12110 (N_12110,N_11874,N_11938);
nor U12111 (N_12111,N_11906,N_11927);
or U12112 (N_12112,N_11886,N_11943);
nor U12113 (N_12113,N_11934,N_11948);
or U12114 (N_12114,N_11980,N_11929);
nor U12115 (N_12115,N_11844,N_11897);
xor U12116 (N_12116,N_11914,N_11899);
nor U12117 (N_12117,N_11856,N_11963);
and U12118 (N_12118,N_11965,N_11970);
xor U12119 (N_12119,N_11960,N_11924);
and U12120 (N_12120,N_11894,N_11910);
nor U12121 (N_12121,N_11964,N_11872);
nor U12122 (N_12122,N_11885,N_11934);
nand U12123 (N_12123,N_11843,N_11953);
xor U12124 (N_12124,N_11938,N_11994);
nand U12125 (N_12125,N_11952,N_11876);
nor U12126 (N_12126,N_11955,N_11929);
nor U12127 (N_12127,N_11858,N_11982);
nand U12128 (N_12128,N_11945,N_11919);
nand U12129 (N_12129,N_11971,N_11892);
nand U12130 (N_12130,N_11879,N_11936);
nor U12131 (N_12131,N_11846,N_11928);
nor U12132 (N_12132,N_11929,N_11945);
xnor U12133 (N_12133,N_11861,N_11945);
xnor U12134 (N_12134,N_11958,N_11970);
and U12135 (N_12135,N_11920,N_11995);
and U12136 (N_12136,N_11977,N_11895);
xor U12137 (N_12137,N_11870,N_11928);
nor U12138 (N_12138,N_11984,N_11948);
and U12139 (N_12139,N_11949,N_11956);
nand U12140 (N_12140,N_11905,N_11930);
nand U12141 (N_12141,N_11935,N_11954);
xnor U12142 (N_12142,N_11907,N_11858);
nand U12143 (N_12143,N_11893,N_11986);
nand U12144 (N_12144,N_11909,N_11963);
nand U12145 (N_12145,N_11946,N_11987);
nor U12146 (N_12146,N_11986,N_11843);
nor U12147 (N_12147,N_11997,N_11965);
and U12148 (N_12148,N_11925,N_11849);
nand U12149 (N_12149,N_11992,N_11929);
nand U12150 (N_12150,N_11843,N_11987);
nand U12151 (N_12151,N_11939,N_11918);
nor U12152 (N_12152,N_11858,N_11880);
xnor U12153 (N_12153,N_11897,N_11850);
or U12154 (N_12154,N_11910,N_11930);
or U12155 (N_12155,N_11872,N_11877);
and U12156 (N_12156,N_11961,N_11907);
or U12157 (N_12157,N_11878,N_11912);
xnor U12158 (N_12158,N_11885,N_11971);
and U12159 (N_12159,N_11873,N_11955);
nand U12160 (N_12160,N_12076,N_12003);
nand U12161 (N_12161,N_12033,N_12029);
nor U12162 (N_12162,N_12116,N_12074);
or U12163 (N_12163,N_12068,N_12053);
nor U12164 (N_12164,N_12137,N_12042);
nor U12165 (N_12165,N_12037,N_12150);
and U12166 (N_12166,N_12096,N_12084);
nand U12167 (N_12167,N_12009,N_12103);
and U12168 (N_12168,N_12107,N_12129);
xnor U12169 (N_12169,N_12145,N_12088);
nor U12170 (N_12170,N_12006,N_12122);
and U12171 (N_12171,N_12044,N_12092);
and U12172 (N_12172,N_12140,N_12026);
and U12173 (N_12173,N_12035,N_12020);
nor U12174 (N_12174,N_12011,N_12014);
nand U12175 (N_12175,N_12108,N_12104);
xor U12176 (N_12176,N_12133,N_12059);
or U12177 (N_12177,N_12034,N_12111);
or U12178 (N_12178,N_12078,N_12019);
and U12179 (N_12179,N_12017,N_12113);
nand U12180 (N_12180,N_12063,N_12132);
and U12181 (N_12181,N_12115,N_12032);
nand U12182 (N_12182,N_12021,N_12156);
or U12183 (N_12183,N_12093,N_12075);
nor U12184 (N_12184,N_12036,N_12117);
or U12185 (N_12185,N_12131,N_12030);
and U12186 (N_12186,N_12031,N_12008);
nand U12187 (N_12187,N_12046,N_12040);
and U12188 (N_12188,N_12056,N_12127);
and U12189 (N_12189,N_12016,N_12083);
and U12190 (N_12190,N_12055,N_12144);
nand U12191 (N_12191,N_12043,N_12070);
or U12192 (N_12192,N_12018,N_12024);
or U12193 (N_12193,N_12000,N_12005);
nand U12194 (N_12194,N_12012,N_12062);
nor U12195 (N_12195,N_12001,N_12110);
nor U12196 (N_12196,N_12154,N_12126);
nor U12197 (N_12197,N_12146,N_12155);
and U12198 (N_12198,N_12085,N_12128);
and U12199 (N_12199,N_12086,N_12069);
xor U12200 (N_12200,N_12039,N_12067);
and U12201 (N_12201,N_12023,N_12151);
xor U12202 (N_12202,N_12058,N_12010);
and U12203 (N_12203,N_12118,N_12123);
nor U12204 (N_12204,N_12106,N_12091);
nor U12205 (N_12205,N_12130,N_12098);
nand U12206 (N_12206,N_12095,N_12027);
nand U12207 (N_12207,N_12090,N_12089);
and U12208 (N_12208,N_12071,N_12072);
or U12209 (N_12209,N_12054,N_12013);
or U12210 (N_12210,N_12094,N_12120);
nor U12211 (N_12211,N_12048,N_12143);
nand U12212 (N_12212,N_12050,N_12077);
nand U12213 (N_12213,N_12052,N_12147);
nor U12214 (N_12214,N_12105,N_12124);
xor U12215 (N_12215,N_12057,N_12139);
nand U12216 (N_12216,N_12136,N_12041);
and U12217 (N_12217,N_12004,N_12060);
and U12218 (N_12218,N_12081,N_12022);
or U12219 (N_12219,N_12102,N_12134);
xor U12220 (N_12220,N_12049,N_12101);
and U12221 (N_12221,N_12114,N_12073);
or U12222 (N_12222,N_12159,N_12007);
xor U12223 (N_12223,N_12065,N_12080);
nor U12224 (N_12224,N_12135,N_12015);
nand U12225 (N_12225,N_12121,N_12153);
and U12226 (N_12226,N_12138,N_12141);
xor U12227 (N_12227,N_12125,N_12087);
nor U12228 (N_12228,N_12158,N_12079);
and U12229 (N_12229,N_12038,N_12002);
nand U12230 (N_12230,N_12119,N_12142);
or U12231 (N_12231,N_12157,N_12099);
and U12232 (N_12232,N_12100,N_12082);
nand U12233 (N_12233,N_12028,N_12061);
or U12234 (N_12234,N_12148,N_12097);
xnor U12235 (N_12235,N_12064,N_12066);
nor U12236 (N_12236,N_12109,N_12025);
nor U12237 (N_12237,N_12045,N_12051);
and U12238 (N_12238,N_12112,N_12152);
and U12239 (N_12239,N_12149,N_12047);
xnor U12240 (N_12240,N_12134,N_12049);
xnor U12241 (N_12241,N_12114,N_12021);
nand U12242 (N_12242,N_12073,N_12153);
or U12243 (N_12243,N_12024,N_12133);
xor U12244 (N_12244,N_12122,N_12133);
and U12245 (N_12245,N_12119,N_12032);
nand U12246 (N_12246,N_12152,N_12049);
xor U12247 (N_12247,N_12084,N_12132);
and U12248 (N_12248,N_12104,N_12039);
and U12249 (N_12249,N_12116,N_12146);
or U12250 (N_12250,N_12064,N_12010);
nand U12251 (N_12251,N_12155,N_12005);
nand U12252 (N_12252,N_12137,N_12097);
nor U12253 (N_12253,N_12083,N_12154);
nand U12254 (N_12254,N_12098,N_12009);
xnor U12255 (N_12255,N_12010,N_12040);
or U12256 (N_12256,N_12131,N_12015);
or U12257 (N_12257,N_12009,N_12068);
nand U12258 (N_12258,N_12019,N_12143);
and U12259 (N_12259,N_12025,N_12111);
nor U12260 (N_12260,N_12061,N_12122);
xnor U12261 (N_12261,N_12089,N_12026);
or U12262 (N_12262,N_12041,N_12073);
xor U12263 (N_12263,N_12159,N_12096);
nor U12264 (N_12264,N_12023,N_12019);
nand U12265 (N_12265,N_12148,N_12081);
nor U12266 (N_12266,N_12041,N_12103);
and U12267 (N_12267,N_12155,N_12082);
or U12268 (N_12268,N_12059,N_12069);
nor U12269 (N_12269,N_12079,N_12097);
nor U12270 (N_12270,N_12001,N_12123);
and U12271 (N_12271,N_12022,N_12016);
or U12272 (N_12272,N_12144,N_12026);
xnor U12273 (N_12273,N_12159,N_12100);
xor U12274 (N_12274,N_12114,N_12069);
or U12275 (N_12275,N_12102,N_12094);
nor U12276 (N_12276,N_12079,N_12022);
nand U12277 (N_12277,N_12037,N_12109);
nand U12278 (N_12278,N_12053,N_12144);
nand U12279 (N_12279,N_12147,N_12019);
nor U12280 (N_12280,N_12140,N_12098);
or U12281 (N_12281,N_12132,N_12099);
nand U12282 (N_12282,N_12013,N_12061);
and U12283 (N_12283,N_12020,N_12011);
or U12284 (N_12284,N_12040,N_12117);
nor U12285 (N_12285,N_12117,N_12011);
nor U12286 (N_12286,N_12100,N_12024);
xnor U12287 (N_12287,N_12084,N_12110);
xnor U12288 (N_12288,N_12110,N_12011);
nand U12289 (N_12289,N_12062,N_12131);
and U12290 (N_12290,N_12071,N_12113);
nor U12291 (N_12291,N_12088,N_12058);
and U12292 (N_12292,N_12037,N_12107);
nor U12293 (N_12293,N_12102,N_12041);
nand U12294 (N_12294,N_12103,N_12072);
and U12295 (N_12295,N_12097,N_12003);
nand U12296 (N_12296,N_12090,N_12074);
xnor U12297 (N_12297,N_12150,N_12118);
xnor U12298 (N_12298,N_12100,N_12143);
nor U12299 (N_12299,N_12039,N_12055);
and U12300 (N_12300,N_12098,N_12049);
or U12301 (N_12301,N_12097,N_12157);
xor U12302 (N_12302,N_12105,N_12012);
nand U12303 (N_12303,N_12089,N_12000);
and U12304 (N_12304,N_12025,N_12151);
nand U12305 (N_12305,N_12056,N_12148);
and U12306 (N_12306,N_12056,N_12109);
nor U12307 (N_12307,N_12143,N_12149);
nand U12308 (N_12308,N_12108,N_12111);
and U12309 (N_12309,N_12137,N_12039);
and U12310 (N_12310,N_12118,N_12080);
or U12311 (N_12311,N_12095,N_12096);
or U12312 (N_12312,N_12021,N_12005);
nor U12313 (N_12313,N_12156,N_12157);
nor U12314 (N_12314,N_12058,N_12089);
nor U12315 (N_12315,N_12021,N_12080);
nand U12316 (N_12316,N_12053,N_12135);
and U12317 (N_12317,N_12010,N_12015);
or U12318 (N_12318,N_12012,N_12116);
and U12319 (N_12319,N_12119,N_12103);
xor U12320 (N_12320,N_12280,N_12235);
nand U12321 (N_12321,N_12170,N_12186);
nand U12322 (N_12322,N_12289,N_12259);
and U12323 (N_12323,N_12251,N_12305);
and U12324 (N_12324,N_12246,N_12188);
or U12325 (N_12325,N_12316,N_12231);
and U12326 (N_12326,N_12213,N_12228);
and U12327 (N_12327,N_12211,N_12203);
nor U12328 (N_12328,N_12274,N_12223);
xor U12329 (N_12329,N_12266,N_12192);
nand U12330 (N_12330,N_12303,N_12297);
nand U12331 (N_12331,N_12205,N_12284);
nand U12332 (N_12332,N_12288,N_12194);
and U12333 (N_12333,N_12279,N_12262);
nand U12334 (N_12334,N_12299,N_12168);
and U12335 (N_12335,N_12193,N_12254);
xnor U12336 (N_12336,N_12237,N_12209);
and U12337 (N_12337,N_12199,N_12277);
or U12338 (N_12338,N_12177,N_12278);
nor U12339 (N_12339,N_12224,N_12230);
or U12340 (N_12340,N_12196,N_12314);
and U12341 (N_12341,N_12302,N_12304);
nor U12342 (N_12342,N_12260,N_12214);
or U12343 (N_12343,N_12182,N_12232);
and U12344 (N_12344,N_12239,N_12269);
nand U12345 (N_12345,N_12309,N_12187);
nand U12346 (N_12346,N_12291,N_12276);
and U12347 (N_12347,N_12225,N_12184);
or U12348 (N_12348,N_12272,N_12238);
or U12349 (N_12349,N_12243,N_12295);
or U12350 (N_12350,N_12172,N_12226);
nor U12351 (N_12351,N_12261,N_12307);
and U12352 (N_12352,N_12267,N_12294);
or U12353 (N_12353,N_12317,N_12221);
or U12354 (N_12354,N_12311,N_12210);
nor U12355 (N_12355,N_12256,N_12169);
or U12356 (N_12356,N_12215,N_12200);
and U12357 (N_12357,N_12174,N_12175);
or U12358 (N_12358,N_12318,N_12282);
xor U12359 (N_12359,N_12176,N_12292);
and U12360 (N_12360,N_12202,N_12298);
nand U12361 (N_12361,N_12189,N_12219);
nor U12362 (N_12362,N_12300,N_12207);
nor U12363 (N_12363,N_12160,N_12178);
and U12364 (N_12364,N_12296,N_12248);
or U12365 (N_12365,N_12183,N_12240);
xor U12366 (N_12366,N_12212,N_12287);
or U12367 (N_12367,N_12171,N_12281);
nand U12368 (N_12368,N_12252,N_12283);
nor U12369 (N_12369,N_12217,N_12181);
or U12370 (N_12370,N_12244,N_12161);
and U12371 (N_12371,N_12249,N_12185);
nand U12372 (N_12372,N_12312,N_12180);
and U12373 (N_12373,N_12164,N_12308);
nor U12374 (N_12374,N_12250,N_12285);
nand U12375 (N_12375,N_12229,N_12273);
xor U12376 (N_12376,N_12247,N_12198);
nor U12377 (N_12377,N_12204,N_12220);
nand U12378 (N_12378,N_12216,N_12234);
or U12379 (N_12379,N_12264,N_12222);
and U12380 (N_12380,N_12319,N_12242);
nor U12381 (N_12381,N_12241,N_12227);
nor U12382 (N_12382,N_12286,N_12268);
and U12383 (N_12383,N_12313,N_12271);
or U12384 (N_12384,N_12253,N_12290);
xor U12385 (N_12385,N_12167,N_12245);
or U12386 (N_12386,N_12306,N_12315);
xnor U12387 (N_12387,N_12270,N_12265);
nand U12388 (N_12388,N_12206,N_12191);
nor U12389 (N_12389,N_12310,N_12195);
and U12390 (N_12390,N_12218,N_12263);
and U12391 (N_12391,N_12190,N_12257);
and U12392 (N_12392,N_12173,N_12208);
and U12393 (N_12393,N_12275,N_12166);
xnor U12394 (N_12394,N_12255,N_12301);
and U12395 (N_12395,N_12258,N_12165);
nor U12396 (N_12396,N_12162,N_12293);
nand U12397 (N_12397,N_12179,N_12236);
nor U12398 (N_12398,N_12197,N_12201);
or U12399 (N_12399,N_12233,N_12163);
xnor U12400 (N_12400,N_12228,N_12198);
and U12401 (N_12401,N_12299,N_12203);
and U12402 (N_12402,N_12298,N_12187);
nor U12403 (N_12403,N_12318,N_12237);
nand U12404 (N_12404,N_12303,N_12216);
nor U12405 (N_12405,N_12254,N_12192);
xor U12406 (N_12406,N_12315,N_12204);
or U12407 (N_12407,N_12319,N_12257);
nor U12408 (N_12408,N_12265,N_12241);
and U12409 (N_12409,N_12256,N_12186);
nand U12410 (N_12410,N_12247,N_12194);
nand U12411 (N_12411,N_12223,N_12194);
or U12412 (N_12412,N_12255,N_12311);
or U12413 (N_12413,N_12246,N_12273);
or U12414 (N_12414,N_12167,N_12220);
or U12415 (N_12415,N_12178,N_12230);
nand U12416 (N_12416,N_12279,N_12283);
nand U12417 (N_12417,N_12226,N_12297);
nor U12418 (N_12418,N_12246,N_12182);
nor U12419 (N_12419,N_12278,N_12289);
or U12420 (N_12420,N_12266,N_12230);
and U12421 (N_12421,N_12220,N_12309);
and U12422 (N_12422,N_12247,N_12161);
or U12423 (N_12423,N_12194,N_12269);
nand U12424 (N_12424,N_12244,N_12218);
or U12425 (N_12425,N_12250,N_12209);
nand U12426 (N_12426,N_12225,N_12318);
xor U12427 (N_12427,N_12295,N_12240);
nor U12428 (N_12428,N_12300,N_12304);
and U12429 (N_12429,N_12208,N_12244);
and U12430 (N_12430,N_12285,N_12181);
and U12431 (N_12431,N_12194,N_12234);
and U12432 (N_12432,N_12160,N_12314);
or U12433 (N_12433,N_12182,N_12257);
xnor U12434 (N_12434,N_12234,N_12302);
and U12435 (N_12435,N_12170,N_12253);
nand U12436 (N_12436,N_12206,N_12265);
xnor U12437 (N_12437,N_12160,N_12251);
nand U12438 (N_12438,N_12305,N_12191);
nand U12439 (N_12439,N_12279,N_12212);
nand U12440 (N_12440,N_12175,N_12258);
or U12441 (N_12441,N_12187,N_12211);
or U12442 (N_12442,N_12234,N_12161);
nand U12443 (N_12443,N_12223,N_12260);
or U12444 (N_12444,N_12309,N_12231);
nor U12445 (N_12445,N_12260,N_12246);
xnor U12446 (N_12446,N_12209,N_12254);
nor U12447 (N_12447,N_12217,N_12301);
or U12448 (N_12448,N_12189,N_12192);
nand U12449 (N_12449,N_12236,N_12213);
xnor U12450 (N_12450,N_12209,N_12257);
xor U12451 (N_12451,N_12290,N_12285);
and U12452 (N_12452,N_12257,N_12174);
nor U12453 (N_12453,N_12299,N_12298);
nand U12454 (N_12454,N_12230,N_12240);
or U12455 (N_12455,N_12189,N_12247);
and U12456 (N_12456,N_12207,N_12269);
and U12457 (N_12457,N_12170,N_12200);
or U12458 (N_12458,N_12170,N_12256);
nand U12459 (N_12459,N_12284,N_12237);
nand U12460 (N_12460,N_12240,N_12190);
or U12461 (N_12461,N_12286,N_12302);
or U12462 (N_12462,N_12267,N_12273);
and U12463 (N_12463,N_12304,N_12197);
or U12464 (N_12464,N_12260,N_12161);
or U12465 (N_12465,N_12264,N_12258);
and U12466 (N_12466,N_12169,N_12191);
nor U12467 (N_12467,N_12164,N_12254);
xor U12468 (N_12468,N_12277,N_12270);
nor U12469 (N_12469,N_12241,N_12275);
or U12470 (N_12470,N_12163,N_12224);
nand U12471 (N_12471,N_12260,N_12295);
or U12472 (N_12472,N_12249,N_12258);
nor U12473 (N_12473,N_12253,N_12283);
and U12474 (N_12474,N_12290,N_12210);
and U12475 (N_12475,N_12207,N_12306);
or U12476 (N_12476,N_12305,N_12176);
or U12477 (N_12477,N_12196,N_12222);
and U12478 (N_12478,N_12222,N_12249);
and U12479 (N_12479,N_12268,N_12244);
and U12480 (N_12480,N_12440,N_12417);
nor U12481 (N_12481,N_12355,N_12374);
and U12482 (N_12482,N_12358,N_12363);
and U12483 (N_12483,N_12323,N_12470);
or U12484 (N_12484,N_12424,N_12407);
nor U12485 (N_12485,N_12438,N_12341);
or U12486 (N_12486,N_12437,N_12330);
nand U12487 (N_12487,N_12385,N_12446);
nand U12488 (N_12488,N_12473,N_12428);
and U12489 (N_12489,N_12445,N_12423);
xor U12490 (N_12490,N_12328,N_12351);
or U12491 (N_12491,N_12463,N_12395);
xnor U12492 (N_12492,N_12436,N_12321);
and U12493 (N_12493,N_12462,N_12370);
nor U12494 (N_12494,N_12337,N_12468);
or U12495 (N_12495,N_12379,N_12455);
or U12496 (N_12496,N_12465,N_12454);
or U12497 (N_12497,N_12430,N_12368);
nand U12498 (N_12498,N_12360,N_12466);
or U12499 (N_12499,N_12434,N_12441);
or U12500 (N_12500,N_12479,N_12467);
and U12501 (N_12501,N_12435,N_12366);
and U12502 (N_12502,N_12406,N_12426);
nand U12503 (N_12503,N_12329,N_12415);
or U12504 (N_12504,N_12353,N_12452);
nor U12505 (N_12505,N_12384,N_12344);
and U12506 (N_12506,N_12460,N_12387);
nand U12507 (N_12507,N_12361,N_12420);
nand U12508 (N_12508,N_12472,N_12369);
and U12509 (N_12509,N_12410,N_12331);
nand U12510 (N_12510,N_12442,N_12380);
nor U12511 (N_12511,N_12346,N_12421);
nor U12512 (N_12512,N_12354,N_12414);
or U12513 (N_12513,N_12377,N_12401);
and U12514 (N_12514,N_12429,N_12388);
nand U12515 (N_12515,N_12413,N_12398);
or U12516 (N_12516,N_12332,N_12396);
and U12517 (N_12517,N_12411,N_12419);
and U12518 (N_12518,N_12362,N_12327);
or U12519 (N_12519,N_12456,N_12427);
nand U12520 (N_12520,N_12399,N_12433);
and U12521 (N_12521,N_12412,N_12340);
nand U12522 (N_12522,N_12403,N_12322);
and U12523 (N_12523,N_12345,N_12432);
and U12524 (N_12524,N_12390,N_12339);
and U12525 (N_12525,N_12409,N_12402);
and U12526 (N_12526,N_12357,N_12349);
and U12527 (N_12527,N_12444,N_12431);
nand U12528 (N_12528,N_12451,N_12335);
nor U12529 (N_12529,N_12373,N_12375);
nor U12530 (N_12530,N_12453,N_12422);
nand U12531 (N_12531,N_12459,N_12394);
and U12532 (N_12532,N_12382,N_12383);
and U12533 (N_12533,N_12461,N_12334);
nor U12534 (N_12534,N_12464,N_12400);
or U12535 (N_12535,N_12405,N_12338);
and U12536 (N_12536,N_12449,N_12478);
or U12537 (N_12537,N_12347,N_12381);
nor U12538 (N_12538,N_12386,N_12475);
xor U12539 (N_12539,N_12352,N_12367);
nand U12540 (N_12540,N_12350,N_12364);
or U12541 (N_12541,N_12378,N_12356);
xor U12542 (N_12542,N_12450,N_12458);
nor U12543 (N_12543,N_12448,N_12443);
nand U12544 (N_12544,N_12389,N_12457);
or U12545 (N_12545,N_12359,N_12320);
nand U12546 (N_12546,N_12324,N_12325);
nor U12547 (N_12547,N_12333,N_12474);
nor U12548 (N_12548,N_12343,N_12477);
and U12549 (N_12549,N_12348,N_12404);
and U12550 (N_12550,N_12476,N_12342);
nor U12551 (N_12551,N_12416,N_12392);
nand U12552 (N_12552,N_12439,N_12336);
or U12553 (N_12553,N_12471,N_12393);
nor U12554 (N_12554,N_12447,N_12425);
nand U12555 (N_12555,N_12469,N_12326);
and U12556 (N_12556,N_12372,N_12391);
or U12557 (N_12557,N_12408,N_12365);
nand U12558 (N_12558,N_12371,N_12418);
and U12559 (N_12559,N_12397,N_12376);
or U12560 (N_12560,N_12330,N_12353);
nand U12561 (N_12561,N_12451,N_12467);
and U12562 (N_12562,N_12333,N_12388);
xor U12563 (N_12563,N_12342,N_12401);
xor U12564 (N_12564,N_12437,N_12349);
nor U12565 (N_12565,N_12325,N_12472);
and U12566 (N_12566,N_12456,N_12428);
nand U12567 (N_12567,N_12384,N_12458);
and U12568 (N_12568,N_12445,N_12378);
and U12569 (N_12569,N_12326,N_12394);
and U12570 (N_12570,N_12408,N_12355);
or U12571 (N_12571,N_12425,N_12329);
nand U12572 (N_12572,N_12411,N_12472);
or U12573 (N_12573,N_12417,N_12328);
and U12574 (N_12574,N_12396,N_12361);
xnor U12575 (N_12575,N_12407,N_12354);
or U12576 (N_12576,N_12369,N_12412);
and U12577 (N_12577,N_12377,N_12448);
or U12578 (N_12578,N_12430,N_12400);
nand U12579 (N_12579,N_12440,N_12394);
nor U12580 (N_12580,N_12454,N_12416);
nand U12581 (N_12581,N_12347,N_12389);
and U12582 (N_12582,N_12380,N_12422);
nand U12583 (N_12583,N_12450,N_12420);
nor U12584 (N_12584,N_12385,N_12381);
nor U12585 (N_12585,N_12386,N_12403);
nand U12586 (N_12586,N_12333,N_12352);
nor U12587 (N_12587,N_12390,N_12360);
nor U12588 (N_12588,N_12445,N_12405);
nand U12589 (N_12589,N_12466,N_12454);
nand U12590 (N_12590,N_12382,N_12420);
and U12591 (N_12591,N_12435,N_12389);
nand U12592 (N_12592,N_12322,N_12396);
or U12593 (N_12593,N_12366,N_12474);
nand U12594 (N_12594,N_12380,N_12448);
nor U12595 (N_12595,N_12417,N_12477);
nand U12596 (N_12596,N_12402,N_12364);
and U12597 (N_12597,N_12411,N_12360);
and U12598 (N_12598,N_12390,N_12473);
and U12599 (N_12599,N_12460,N_12351);
xor U12600 (N_12600,N_12397,N_12331);
or U12601 (N_12601,N_12368,N_12390);
or U12602 (N_12602,N_12472,N_12384);
nor U12603 (N_12603,N_12413,N_12353);
and U12604 (N_12604,N_12325,N_12403);
or U12605 (N_12605,N_12330,N_12426);
nand U12606 (N_12606,N_12462,N_12393);
and U12607 (N_12607,N_12419,N_12322);
or U12608 (N_12608,N_12449,N_12358);
nor U12609 (N_12609,N_12398,N_12455);
nand U12610 (N_12610,N_12445,N_12404);
or U12611 (N_12611,N_12414,N_12368);
or U12612 (N_12612,N_12431,N_12454);
nor U12613 (N_12613,N_12361,N_12462);
nor U12614 (N_12614,N_12322,N_12442);
nand U12615 (N_12615,N_12320,N_12470);
nor U12616 (N_12616,N_12425,N_12407);
nor U12617 (N_12617,N_12324,N_12371);
nand U12618 (N_12618,N_12376,N_12464);
nor U12619 (N_12619,N_12348,N_12464);
and U12620 (N_12620,N_12333,N_12431);
and U12621 (N_12621,N_12435,N_12356);
nand U12622 (N_12622,N_12425,N_12324);
nor U12623 (N_12623,N_12432,N_12477);
nand U12624 (N_12624,N_12335,N_12339);
nor U12625 (N_12625,N_12427,N_12434);
xnor U12626 (N_12626,N_12367,N_12473);
nand U12627 (N_12627,N_12360,N_12443);
or U12628 (N_12628,N_12474,N_12414);
nor U12629 (N_12629,N_12391,N_12478);
and U12630 (N_12630,N_12458,N_12324);
nand U12631 (N_12631,N_12363,N_12382);
or U12632 (N_12632,N_12433,N_12342);
nand U12633 (N_12633,N_12432,N_12361);
or U12634 (N_12634,N_12356,N_12369);
or U12635 (N_12635,N_12408,N_12374);
or U12636 (N_12636,N_12373,N_12394);
nand U12637 (N_12637,N_12437,N_12320);
or U12638 (N_12638,N_12337,N_12424);
nand U12639 (N_12639,N_12460,N_12446);
nand U12640 (N_12640,N_12625,N_12564);
or U12641 (N_12641,N_12582,N_12493);
or U12642 (N_12642,N_12523,N_12511);
nand U12643 (N_12643,N_12487,N_12506);
nor U12644 (N_12644,N_12518,N_12588);
or U12645 (N_12645,N_12578,N_12531);
or U12646 (N_12646,N_12555,N_12623);
nor U12647 (N_12647,N_12502,N_12596);
and U12648 (N_12648,N_12522,N_12554);
nand U12649 (N_12649,N_12601,N_12496);
or U12650 (N_12650,N_12509,N_12587);
and U12651 (N_12651,N_12558,N_12635);
nand U12652 (N_12652,N_12499,N_12530);
and U12653 (N_12653,N_12593,N_12600);
nor U12654 (N_12654,N_12566,N_12544);
xor U12655 (N_12655,N_12565,N_12581);
nand U12656 (N_12656,N_12569,N_12637);
or U12657 (N_12657,N_12512,N_12494);
or U12658 (N_12658,N_12547,N_12500);
or U12659 (N_12659,N_12561,N_12548);
xor U12660 (N_12660,N_12606,N_12480);
and U12661 (N_12661,N_12485,N_12598);
or U12662 (N_12662,N_12612,N_12560);
or U12663 (N_12663,N_12498,N_12534);
or U12664 (N_12664,N_12605,N_12627);
and U12665 (N_12665,N_12621,N_12615);
xor U12666 (N_12666,N_12573,N_12639);
or U12667 (N_12667,N_12527,N_12538);
or U12668 (N_12668,N_12504,N_12495);
nand U12669 (N_12669,N_12526,N_12489);
or U12670 (N_12670,N_12630,N_12619);
xor U12671 (N_12671,N_12599,N_12628);
and U12672 (N_12672,N_12568,N_12611);
nor U12673 (N_12673,N_12481,N_12546);
nand U12674 (N_12674,N_12556,N_12629);
or U12675 (N_12675,N_12550,N_12505);
nor U12676 (N_12676,N_12603,N_12559);
or U12677 (N_12677,N_12540,N_12492);
nor U12678 (N_12678,N_12545,N_12516);
or U12679 (N_12679,N_12508,N_12549);
nor U12680 (N_12680,N_12631,N_12490);
nand U12681 (N_12681,N_12577,N_12608);
nand U12682 (N_12682,N_12486,N_12517);
nor U12683 (N_12683,N_12622,N_12562);
and U12684 (N_12684,N_12563,N_12616);
xor U12685 (N_12685,N_12579,N_12594);
nand U12686 (N_12686,N_12503,N_12589);
and U12687 (N_12687,N_12586,N_12535);
nor U12688 (N_12688,N_12521,N_12542);
nand U12689 (N_12689,N_12497,N_12541);
nand U12690 (N_12690,N_12515,N_12519);
nor U12691 (N_12691,N_12525,N_12624);
or U12692 (N_12692,N_12570,N_12610);
or U12693 (N_12693,N_12482,N_12529);
nor U12694 (N_12694,N_12626,N_12617);
xnor U12695 (N_12695,N_12543,N_12632);
nand U12696 (N_12696,N_12636,N_12507);
xnor U12697 (N_12697,N_12583,N_12613);
and U12698 (N_12698,N_12510,N_12597);
nand U12699 (N_12699,N_12491,N_12533);
or U12700 (N_12700,N_12591,N_12614);
nand U12701 (N_12701,N_12572,N_12576);
nor U12702 (N_12702,N_12585,N_12484);
xnor U12703 (N_12703,N_12537,N_12607);
nor U12704 (N_12704,N_12575,N_12618);
nand U12705 (N_12705,N_12553,N_12580);
nor U12706 (N_12706,N_12514,N_12551);
nand U12707 (N_12707,N_12528,N_12604);
xor U12708 (N_12708,N_12501,N_12488);
and U12709 (N_12709,N_12524,N_12634);
or U12710 (N_12710,N_12638,N_12557);
and U12711 (N_12711,N_12567,N_12536);
nand U12712 (N_12712,N_12552,N_12609);
and U12713 (N_12713,N_12483,N_12571);
or U12714 (N_12714,N_12633,N_12620);
and U12715 (N_12715,N_12532,N_12590);
and U12716 (N_12716,N_12513,N_12574);
and U12717 (N_12717,N_12592,N_12539);
nor U12718 (N_12718,N_12584,N_12520);
and U12719 (N_12719,N_12602,N_12595);
nor U12720 (N_12720,N_12553,N_12617);
or U12721 (N_12721,N_12546,N_12562);
nand U12722 (N_12722,N_12487,N_12545);
or U12723 (N_12723,N_12613,N_12557);
nor U12724 (N_12724,N_12580,N_12503);
nand U12725 (N_12725,N_12489,N_12504);
nor U12726 (N_12726,N_12490,N_12506);
and U12727 (N_12727,N_12590,N_12568);
and U12728 (N_12728,N_12614,N_12570);
and U12729 (N_12729,N_12608,N_12541);
or U12730 (N_12730,N_12622,N_12599);
and U12731 (N_12731,N_12622,N_12616);
nor U12732 (N_12732,N_12530,N_12558);
nand U12733 (N_12733,N_12633,N_12503);
or U12734 (N_12734,N_12482,N_12567);
nand U12735 (N_12735,N_12566,N_12639);
nand U12736 (N_12736,N_12549,N_12481);
or U12737 (N_12737,N_12523,N_12486);
or U12738 (N_12738,N_12552,N_12511);
and U12739 (N_12739,N_12574,N_12491);
nand U12740 (N_12740,N_12530,N_12579);
xor U12741 (N_12741,N_12591,N_12572);
or U12742 (N_12742,N_12580,N_12601);
nand U12743 (N_12743,N_12615,N_12529);
or U12744 (N_12744,N_12525,N_12563);
or U12745 (N_12745,N_12556,N_12545);
nor U12746 (N_12746,N_12609,N_12508);
and U12747 (N_12747,N_12499,N_12489);
nand U12748 (N_12748,N_12584,N_12511);
xnor U12749 (N_12749,N_12633,N_12506);
and U12750 (N_12750,N_12600,N_12615);
nand U12751 (N_12751,N_12480,N_12591);
nand U12752 (N_12752,N_12521,N_12493);
nand U12753 (N_12753,N_12536,N_12621);
nor U12754 (N_12754,N_12571,N_12625);
nand U12755 (N_12755,N_12586,N_12557);
nor U12756 (N_12756,N_12557,N_12560);
nand U12757 (N_12757,N_12537,N_12550);
or U12758 (N_12758,N_12622,N_12582);
and U12759 (N_12759,N_12548,N_12583);
or U12760 (N_12760,N_12626,N_12576);
nand U12761 (N_12761,N_12506,N_12616);
and U12762 (N_12762,N_12521,N_12599);
or U12763 (N_12763,N_12622,N_12628);
or U12764 (N_12764,N_12610,N_12558);
nand U12765 (N_12765,N_12615,N_12499);
nor U12766 (N_12766,N_12619,N_12485);
nor U12767 (N_12767,N_12493,N_12630);
nand U12768 (N_12768,N_12575,N_12485);
and U12769 (N_12769,N_12628,N_12550);
and U12770 (N_12770,N_12548,N_12482);
nand U12771 (N_12771,N_12562,N_12506);
nand U12772 (N_12772,N_12523,N_12490);
xnor U12773 (N_12773,N_12582,N_12593);
nand U12774 (N_12774,N_12483,N_12524);
xnor U12775 (N_12775,N_12506,N_12572);
or U12776 (N_12776,N_12546,N_12605);
nor U12777 (N_12777,N_12635,N_12516);
xor U12778 (N_12778,N_12553,N_12593);
or U12779 (N_12779,N_12570,N_12488);
nand U12780 (N_12780,N_12618,N_12500);
xnor U12781 (N_12781,N_12516,N_12576);
nor U12782 (N_12782,N_12609,N_12625);
nor U12783 (N_12783,N_12526,N_12545);
nand U12784 (N_12784,N_12634,N_12541);
or U12785 (N_12785,N_12609,N_12530);
and U12786 (N_12786,N_12587,N_12605);
and U12787 (N_12787,N_12564,N_12480);
or U12788 (N_12788,N_12598,N_12561);
or U12789 (N_12789,N_12605,N_12547);
or U12790 (N_12790,N_12634,N_12572);
and U12791 (N_12791,N_12626,N_12526);
and U12792 (N_12792,N_12491,N_12629);
and U12793 (N_12793,N_12558,N_12508);
and U12794 (N_12794,N_12594,N_12535);
and U12795 (N_12795,N_12567,N_12487);
nand U12796 (N_12796,N_12508,N_12525);
and U12797 (N_12797,N_12549,N_12621);
nand U12798 (N_12798,N_12579,N_12627);
nor U12799 (N_12799,N_12516,N_12515);
or U12800 (N_12800,N_12672,N_12642);
nand U12801 (N_12801,N_12754,N_12742);
and U12802 (N_12802,N_12755,N_12778);
or U12803 (N_12803,N_12699,N_12690);
and U12804 (N_12804,N_12676,N_12779);
nor U12805 (N_12805,N_12700,N_12715);
and U12806 (N_12806,N_12711,N_12654);
and U12807 (N_12807,N_12725,N_12780);
nand U12808 (N_12808,N_12692,N_12798);
nor U12809 (N_12809,N_12763,N_12720);
nor U12810 (N_12810,N_12752,N_12669);
and U12811 (N_12811,N_12760,N_12777);
xor U12812 (N_12812,N_12773,N_12658);
nor U12813 (N_12813,N_12783,N_12774);
nand U12814 (N_12814,N_12791,N_12750);
nor U12815 (N_12815,N_12686,N_12721);
nand U12816 (N_12816,N_12650,N_12747);
nor U12817 (N_12817,N_12709,N_12651);
nand U12818 (N_12818,N_12681,N_12697);
and U12819 (N_12819,N_12683,N_12731);
and U12820 (N_12820,N_12652,N_12768);
nor U12821 (N_12821,N_12741,N_12667);
nand U12822 (N_12822,N_12703,N_12740);
and U12823 (N_12823,N_12761,N_12786);
or U12824 (N_12824,N_12756,N_12706);
or U12825 (N_12825,N_12648,N_12765);
nor U12826 (N_12826,N_12653,N_12674);
and U12827 (N_12827,N_12730,N_12663);
nand U12828 (N_12828,N_12641,N_12746);
nand U12829 (N_12829,N_12657,N_12766);
or U12830 (N_12830,N_12794,N_12705);
or U12831 (N_12831,N_12718,N_12767);
or U12832 (N_12832,N_12696,N_12724);
nor U12833 (N_12833,N_12701,N_12691);
nand U12834 (N_12834,N_12726,N_12735);
nand U12835 (N_12835,N_12675,N_12781);
nand U12836 (N_12836,N_12789,N_12790);
and U12837 (N_12837,N_12797,N_12795);
nand U12838 (N_12838,N_12733,N_12769);
or U12839 (N_12839,N_12748,N_12719);
nand U12840 (N_12840,N_12728,N_12785);
or U12841 (N_12841,N_12714,N_12753);
xnor U12842 (N_12842,N_12784,N_12670);
or U12843 (N_12843,N_12661,N_12684);
xor U12844 (N_12844,N_12673,N_12775);
xor U12845 (N_12845,N_12799,N_12680);
xor U12846 (N_12846,N_12757,N_12682);
xnor U12847 (N_12847,N_12782,N_12723);
or U12848 (N_12848,N_12665,N_12713);
nand U12849 (N_12849,N_12722,N_12685);
and U12850 (N_12850,N_12727,N_12646);
nor U12851 (N_12851,N_12655,N_12737);
nand U12852 (N_12852,N_12668,N_12770);
nor U12853 (N_12853,N_12698,N_12643);
and U12854 (N_12854,N_12688,N_12732);
or U12855 (N_12855,N_12678,N_12716);
or U12856 (N_12856,N_12751,N_12745);
xor U12857 (N_12857,N_12644,N_12762);
xor U12858 (N_12858,N_12744,N_12677);
and U12859 (N_12859,N_12645,N_12792);
or U12860 (N_12860,N_12659,N_12796);
nor U12861 (N_12861,N_12787,N_12708);
nand U12862 (N_12862,N_12759,N_12647);
nand U12863 (N_12863,N_12793,N_12649);
or U12864 (N_12864,N_12666,N_12749);
and U12865 (N_12865,N_12771,N_12640);
or U12866 (N_12866,N_12734,N_12662);
nand U12867 (N_12867,N_12656,N_12689);
nor U12868 (N_12868,N_12671,N_12660);
and U12869 (N_12869,N_12772,N_12687);
or U12870 (N_12870,N_12736,N_12764);
nor U12871 (N_12871,N_12788,N_12717);
and U12872 (N_12872,N_12729,N_12758);
or U12873 (N_12873,N_12738,N_12776);
and U12874 (N_12874,N_12694,N_12679);
nand U12875 (N_12875,N_12702,N_12704);
xnor U12876 (N_12876,N_12707,N_12739);
nor U12877 (N_12877,N_12664,N_12710);
xnor U12878 (N_12878,N_12695,N_12693);
and U12879 (N_12879,N_12743,N_12712);
nand U12880 (N_12880,N_12762,N_12689);
and U12881 (N_12881,N_12775,N_12716);
and U12882 (N_12882,N_12728,N_12739);
and U12883 (N_12883,N_12709,N_12724);
and U12884 (N_12884,N_12660,N_12679);
nor U12885 (N_12885,N_12731,N_12753);
nor U12886 (N_12886,N_12791,N_12690);
nor U12887 (N_12887,N_12767,N_12654);
nor U12888 (N_12888,N_12745,N_12773);
nand U12889 (N_12889,N_12666,N_12705);
xnor U12890 (N_12890,N_12748,N_12791);
or U12891 (N_12891,N_12714,N_12698);
and U12892 (N_12892,N_12779,N_12711);
nor U12893 (N_12893,N_12653,N_12748);
nor U12894 (N_12894,N_12767,N_12761);
nand U12895 (N_12895,N_12765,N_12740);
nand U12896 (N_12896,N_12682,N_12794);
nor U12897 (N_12897,N_12766,N_12753);
or U12898 (N_12898,N_12651,N_12734);
nand U12899 (N_12899,N_12776,N_12700);
or U12900 (N_12900,N_12786,N_12661);
and U12901 (N_12901,N_12732,N_12693);
nor U12902 (N_12902,N_12755,N_12762);
and U12903 (N_12903,N_12759,N_12728);
and U12904 (N_12904,N_12782,N_12668);
nand U12905 (N_12905,N_12702,N_12780);
and U12906 (N_12906,N_12646,N_12693);
and U12907 (N_12907,N_12693,N_12734);
and U12908 (N_12908,N_12790,N_12666);
and U12909 (N_12909,N_12705,N_12715);
and U12910 (N_12910,N_12647,N_12732);
nand U12911 (N_12911,N_12658,N_12795);
and U12912 (N_12912,N_12715,N_12780);
nor U12913 (N_12913,N_12731,N_12668);
or U12914 (N_12914,N_12649,N_12644);
nor U12915 (N_12915,N_12663,N_12769);
and U12916 (N_12916,N_12721,N_12687);
nor U12917 (N_12917,N_12647,N_12651);
and U12918 (N_12918,N_12746,N_12716);
or U12919 (N_12919,N_12734,N_12785);
or U12920 (N_12920,N_12744,N_12752);
or U12921 (N_12921,N_12716,N_12698);
nand U12922 (N_12922,N_12763,N_12775);
nor U12923 (N_12923,N_12699,N_12722);
and U12924 (N_12924,N_12667,N_12662);
xnor U12925 (N_12925,N_12712,N_12655);
nor U12926 (N_12926,N_12709,N_12646);
nand U12927 (N_12927,N_12770,N_12711);
or U12928 (N_12928,N_12644,N_12774);
and U12929 (N_12929,N_12737,N_12681);
xnor U12930 (N_12930,N_12742,N_12664);
xnor U12931 (N_12931,N_12713,N_12709);
nor U12932 (N_12932,N_12693,N_12684);
and U12933 (N_12933,N_12783,N_12737);
nand U12934 (N_12934,N_12742,N_12640);
and U12935 (N_12935,N_12730,N_12702);
nand U12936 (N_12936,N_12682,N_12777);
nor U12937 (N_12937,N_12721,N_12706);
or U12938 (N_12938,N_12764,N_12756);
or U12939 (N_12939,N_12796,N_12693);
nor U12940 (N_12940,N_12640,N_12719);
nor U12941 (N_12941,N_12720,N_12781);
nand U12942 (N_12942,N_12734,N_12640);
nand U12943 (N_12943,N_12784,N_12695);
xnor U12944 (N_12944,N_12741,N_12709);
or U12945 (N_12945,N_12649,N_12650);
nor U12946 (N_12946,N_12738,N_12782);
nand U12947 (N_12947,N_12789,N_12648);
and U12948 (N_12948,N_12673,N_12756);
or U12949 (N_12949,N_12671,N_12740);
or U12950 (N_12950,N_12764,N_12726);
xor U12951 (N_12951,N_12762,N_12749);
and U12952 (N_12952,N_12671,N_12776);
or U12953 (N_12953,N_12736,N_12713);
nand U12954 (N_12954,N_12727,N_12678);
or U12955 (N_12955,N_12737,N_12756);
nand U12956 (N_12956,N_12708,N_12755);
and U12957 (N_12957,N_12742,N_12734);
nand U12958 (N_12958,N_12797,N_12746);
and U12959 (N_12959,N_12725,N_12686);
nand U12960 (N_12960,N_12924,N_12958);
nor U12961 (N_12961,N_12847,N_12835);
and U12962 (N_12962,N_12834,N_12807);
or U12963 (N_12963,N_12817,N_12816);
nor U12964 (N_12964,N_12903,N_12808);
or U12965 (N_12965,N_12805,N_12802);
or U12966 (N_12966,N_12803,N_12896);
nand U12967 (N_12967,N_12891,N_12933);
nor U12968 (N_12968,N_12894,N_12844);
nand U12969 (N_12969,N_12836,N_12826);
and U12970 (N_12970,N_12957,N_12830);
nor U12971 (N_12971,N_12854,N_12810);
and U12972 (N_12972,N_12814,N_12956);
or U12973 (N_12973,N_12880,N_12948);
and U12974 (N_12974,N_12918,N_12823);
nand U12975 (N_12975,N_12881,N_12926);
or U12976 (N_12976,N_12865,N_12825);
and U12977 (N_12977,N_12876,N_12801);
and U12978 (N_12978,N_12867,N_12829);
nand U12979 (N_12979,N_12886,N_12889);
and U12980 (N_12980,N_12959,N_12846);
nor U12981 (N_12981,N_12811,N_12890);
nand U12982 (N_12982,N_12954,N_12947);
nand U12983 (N_12983,N_12800,N_12900);
xor U12984 (N_12984,N_12925,N_12913);
or U12985 (N_12985,N_12938,N_12906);
nand U12986 (N_12986,N_12872,N_12914);
or U12987 (N_12987,N_12868,N_12871);
nor U12988 (N_12988,N_12859,N_12923);
nor U12989 (N_12989,N_12833,N_12927);
nor U12990 (N_12990,N_12937,N_12822);
xor U12991 (N_12991,N_12873,N_12951);
nor U12992 (N_12992,N_12892,N_12949);
and U12993 (N_12993,N_12911,N_12853);
or U12994 (N_12994,N_12922,N_12841);
or U12995 (N_12995,N_12824,N_12862);
and U12996 (N_12996,N_12955,N_12942);
and U12997 (N_12997,N_12929,N_12866);
nor U12998 (N_12998,N_12931,N_12883);
nor U12999 (N_12999,N_12946,N_12898);
nor U13000 (N_13000,N_12904,N_12818);
or U13001 (N_13001,N_12843,N_12910);
xor U13002 (N_13002,N_12950,N_12884);
and U13003 (N_13003,N_12945,N_12920);
or U13004 (N_13004,N_12857,N_12934);
or U13005 (N_13005,N_12917,N_12899);
or U13006 (N_13006,N_12940,N_12909);
or U13007 (N_13007,N_12928,N_12902);
xor U13008 (N_13008,N_12935,N_12901);
or U13009 (N_13009,N_12921,N_12821);
and U13010 (N_13010,N_12815,N_12893);
or U13011 (N_13011,N_12839,N_12840);
xnor U13012 (N_13012,N_12885,N_12813);
and U13013 (N_13013,N_12887,N_12837);
or U13014 (N_13014,N_12919,N_12855);
xnor U13015 (N_13015,N_12888,N_12877);
and U13016 (N_13016,N_12863,N_12941);
nor U13017 (N_13017,N_12895,N_12870);
or U13018 (N_13018,N_12882,N_12842);
or U13019 (N_13019,N_12932,N_12809);
or U13020 (N_13020,N_12930,N_12806);
nand U13021 (N_13021,N_12861,N_12907);
nor U13022 (N_13022,N_12804,N_12812);
or U13023 (N_13023,N_12878,N_12875);
xnor U13024 (N_13024,N_12905,N_12915);
xor U13025 (N_13025,N_12831,N_12845);
nor U13026 (N_13026,N_12916,N_12912);
nand U13027 (N_13027,N_12851,N_12943);
and U13028 (N_13028,N_12832,N_12827);
and U13029 (N_13029,N_12953,N_12828);
xnor U13030 (N_13030,N_12864,N_12897);
and U13031 (N_13031,N_12944,N_12849);
and U13032 (N_13032,N_12848,N_12838);
xor U13033 (N_13033,N_12850,N_12939);
nor U13034 (N_13034,N_12820,N_12936);
nand U13035 (N_13035,N_12869,N_12879);
or U13036 (N_13036,N_12874,N_12858);
nor U13037 (N_13037,N_12856,N_12819);
and U13038 (N_13038,N_12852,N_12952);
nand U13039 (N_13039,N_12860,N_12908);
nor U13040 (N_13040,N_12954,N_12910);
and U13041 (N_13041,N_12934,N_12927);
nor U13042 (N_13042,N_12924,N_12800);
or U13043 (N_13043,N_12825,N_12843);
nor U13044 (N_13044,N_12805,N_12912);
and U13045 (N_13045,N_12938,N_12957);
nor U13046 (N_13046,N_12933,N_12929);
nand U13047 (N_13047,N_12832,N_12812);
or U13048 (N_13048,N_12941,N_12920);
nor U13049 (N_13049,N_12806,N_12953);
nand U13050 (N_13050,N_12802,N_12863);
nor U13051 (N_13051,N_12906,N_12871);
and U13052 (N_13052,N_12884,N_12838);
nand U13053 (N_13053,N_12845,N_12916);
or U13054 (N_13054,N_12862,N_12926);
nand U13055 (N_13055,N_12812,N_12959);
nand U13056 (N_13056,N_12956,N_12930);
nand U13057 (N_13057,N_12869,N_12880);
nor U13058 (N_13058,N_12948,N_12812);
and U13059 (N_13059,N_12832,N_12903);
and U13060 (N_13060,N_12872,N_12958);
nand U13061 (N_13061,N_12855,N_12869);
and U13062 (N_13062,N_12833,N_12818);
and U13063 (N_13063,N_12837,N_12814);
nand U13064 (N_13064,N_12866,N_12898);
and U13065 (N_13065,N_12936,N_12826);
and U13066 (N_13066,N_12803,N_12943);
xor U13067 (N_13067,N_12858,N_12828);
xnor U13068 (N_13068,N_12816,N_12929);
or U13069 (N_13069,N_12917,N_12829);
nor U13070 (N_13070,N_12912,N_12841);
and U13071 (N_13071,N_12935,N_12905);
or U13072 (N_13072,N_12872,N_12878);
nor U13073 (N_13073,N_12954,N_12847);
and U13074 (N_13074,N_12852,N_12841);
nand U13075 (N_13075,N_12912,N_12930);
nand U13076 (N_13076,N_12924,N_12941);
or U13077 (N_13077,N_12955,N_12891);
nor U13078 (N_13078,N_12884,N_12859);
nor U13079 (N_13079,N_12866,N_12952);
and U13080 (N_13080,N_12927,N_12933);
or U13081 (N_13081,N_12939,N_12803);
nand U13082 (N_13082,N_12830,N_12896);
or U13083 (N_13083,N_12869,N_12843);
and U13084 (N_13084,N_12805,N_12857);
or U13085 (N_13085,N_12834,N_12921);
xnor U13086 (N_13086,N_12899,N_12876);
nand U13087 (N_13087,N_12946,N_12913);
and U13088 (N_13088,N_12902,N_12831);
and U13089 (N_13089,N_12815,N_12919);
or U13090 (N_13090,N_12891,N_12894);
and U13091 (N_13091,N_12908,N_12907);
nor U13092 (N_13092,N_12946,N_12856);
nor U13093 (N_13093,N_12804,N_12871);
and U13094 (N_13094,N_12913,N_12849);
or U13095 (N_13095,N_12839,N_12954);
nand U13096 (N_13096,N_12958,N_12863);
and U13097 (N_13097,N_12927,N_12873);
and U13098 (N_13098,N_12835,N_12809);
and U13099 (N_13099,N_12902,N_12812);
or U13100 (N_13100,N_12825,N_12820);
and U13101 (N_13101,N_12840,N_12913);
nor U13102 (N_13102,N_12903,N_12846);
or U13103 (N_13103,N_12908,N_12811);
nand U13104 (N_13104,N_12917,N_12914);
nand U13105 (N_13105,N_12821,N_12827);
xor U13106 (N_13106,N_12942,N_12937);
and U13107 (N_13107,N_12954,N_12823);
nor U13108 (N_13108,N_12813,N_12912);
nand U13109 (N_13109,N_12942,N_12834);
nand U13110 (N_13110,N_12938,N_12864);
xnor U13111 (N_13111,N_12820,N_12959);
and U13112 (N_13112,N_12915,N_12808);
nor U13113 (N_13113,N_12819,N_12823);
and U13114 (N_13114,N_12870,N_12930);
nor U13115 (N_13115,N_12812,N_12843);
nor U13116 (N_13116,N_12934,N_12816);
or U13117 (N_13117,N_12897,N_12934);
and U13118 (N_13118,N_12936,N_12814);
or U13119 (N_13119,N_12829,N_12828);
nor U13120 (N_13120,N_13026,N_13016);
or U13121 (N_13121,N_13104,N_13032);
or U13122 (N_13122,N_13017,N_13007);
and U13123 (N_13123,N_12967,N_13079);
nand U13124 (N_13124,N_12971,N_12984);
nor U13125 (N_13125,N_13115,N_13041);
nand U13126 (N_13126,N_13036,N_13097);
nand U13127 (N_13127,N_13069,N_13024);
or U13128 (N_13128,N_12965,N_13072);
and U13129 (N_13129,N_12983,N_13002);
and U13130 (N_13130,N_13020,N_13076);
or U13131 (N_13131,N_13015,N_13114);
nand U13132 (N_13132,N_13109,N_13038);
nand U13133 (N_13133,N_13084,N_12975);
nand U13134 (N_13134,N_13006,N_12998);
nor U13135 (N_13135,N_13062,N_13110);
or U13136 (N_13136,N_13000,N_13093);
or U13137 (N_13137,N_13005,N_13112);
nand U13138 (N_13138,N_12990,N_12961);
and U13139 (N_13139,N_13111,N_13094);
xor U13140 (N_13140,N_12994,N_13012);
and U13141 (N_13141,N_13008,N_13119);
xnor U13142 (N_13142,N_13004,N_12968);
and U13143 (N_13143,N_13025,N_13075);
nor U13144 (N_13144,N_13064,N_13113);
nand U13145 (N_13145,N_13107,N_13023);
nand U13146 (N_13146,N_13116,N_12986);
and U13147 (N_13147,N_13080,N_13105);
nor U13148 (N_13148,N_13053,N_12963);
or U13149 (N_13149,N_12966,N_13083);
nor U13150 (N_13150,N_13092,N_13051);
and U13151 (N_13151,N_12969,N_13046);
and U13152 (N_13152,N_13056,N_13034);
nor U13153 (N_13153,N_13001,N_12985);
and U13154 (N_13154,N_12979,N_13065);
or U13155 (N_13155,N_13085,N_13045);
or U13156 (N_13156,N_12995,N_12973);
or U13157 (N_13157,N_12997,N_13013);
and U13158 (N_13158,N_12996,N_12992);
nor U13159 (N_13159,N_12981,N_13058);
and U13160 (N_13160,N_13074,N_13066);
nor U13161 (N_13161,N_12980,N_12962);
xnor U13162 (N_13162,N_13052,N_13088);
nor U13163 (N_13163,N_13049,N_12964);
nand U13164 (N_13164,N_13060,N_13003);
or U13165 (N_13165,N_12960,N_13068);
nand U13166 (N_13166,N_13082,N_13090);
nand U13167 (N_13167,N_13081,N_12970);
or U13168 (N_13168,N_13108,N_13054);
nor U13169 (N_13169,N_12972,N_13102);
nor U13170 (N_13170,N_13101,N_12991);
nor U13171 (N_13171,N_13030,N_13091);
and U13172 (N_13172,N_13103,N_13044);
nand U13173 (N_13173,N_13061,N_13028);
nor U13174 (N_13174,N_13063,N_13048);
and U13175 (N_13175,N_13106,N_13118);
and U13176 (N_13176,N_13098,N_13100);
nor U13177 (N_13177,N_13037,N_12974);
and U13178 (N_13178,N_12978,N_13099);
or U13179 (N_13179,N_13011,N_13042);
nor U13180 (N_13180,N_13014,N_12977);
nand U13181 (N_13181,N_13087,N_13067);
and U13182 (N_13182,N_13033,N_13071);
and U13183 (N_13183,N_13021,N_13095);
nor U13184 (N_13184,N_13050,N_13055);
and U13185 (N_13185,N_12988,N_12999);
nand U13186 (N_13186,N_13078,N_13031);
nor U13187 (N_13187,N_13086,N_12982);
nor U13188 (N_13188,N_13027,N_12989);
or U13189 (N_13189,N_13089,N_12993);
nand U13190 (N_13190,N_13070,N_13010);
xnor U13191 (N_13191,N_13035,N_12987);
xor U13192 (N_13192,N_13019,N_13040);
and U13193 (N_13193,N_13073,N_13029);
nand U13194 (N_13194,N_13022,N_12976);
or U13195 (N_13195,N_13043,N_13018);
nor U13196 (N_13196,N_13059,N_13039);
nand U13197 (N_13197,N_13057,N_13047);
nand U13198 (N_13198,N_13077,N_13096);
and U13199 (N_13199,N_13009,N_13117);
and U13200 (N_13200,N_13091,N_13005);
nor U13201 (N_13201,N_12978,N_13050);
and U13202 (N_13202,N_13059,N_13082);
nor U13203 (N_13203,N_13003,N_12992);
nand U13204 (N_13204,N_13091,N_12993);
or U13205 (N_13205,N_13110,N_13065);
nand U13206 (N_13206,N_13097,N_12990);
or U13207 (N_13207,N_12993,N_13111);
or U13208 (N_13208,N_13013,N_13112);
and U13209 (N_13209,N_13087,N_13106);
or U13210 (N_13210,N_12965,N_12961);
nand U13211 (N_13211,N_13077,N_13057);
and U13212 (N_13212,N_12993,N_12976);
or U13213 (N_13213,N_13033,N_13038);
and U13214 (N_13214,N_13004,N_13107);
nor U13215 (N_13215,N_13072,N_12962);
nor U13216 (N_13216,N_12987,N_12963);
xnor U13217 (N_13217,N_13038,N_12978);
xor U13218 (N_13218,N_13057,N_13021);
nand U13219 (N_13219,N_13012,N_13110);
xor U13220 (N_13220,N_12980,N_12961);
or U13221 (N_13221,N_13091,N_13089);
nand U13222 (N_13222,N_12975,N_13080);
and U13223 (N_13223,N_13089,N_13027);
nor U13224 (N_13224,N_13115,N_13042);
and U13225 (N_13225,N_13105,N_13088);
nand U13226 (N_13226,N_12963,N_13101);
and U13227 (N_13227,N_13067,N_13042);
nor U13228 (N_13228,N_13106,N_12985);
nor U13229 (N_13229,N_13003,N_13104);
nor U13230 (N_13230,N_12979,N_13075);
nor U13231 (N_13231,N_12992,N_13008);
nand U13232 (N_13232,N_12986,N_13102);
nand U13233 (N_13233,N_12987,N_12964);
nand U13234 (N_13234,N_13039,N_13008);
and U13235 (N_13235,N_13081,N_13095);
and U13236 (N_13236,N_13110,N_13073);
nand U13237 (N_13237,N_12985,N_13116);
and U13238 (N_13238,N_13119,N_13017);
or U13239 (N_13239,N_13010,N_13092);
nor U13240 (N_13240,N_13119,N_13068);
xor U13241 (N_13241,N_13079,N_13052);
nor U13242 (N_13242,N_13101,N_13005);
nand U13243 (N_13243,N_13027,N_12966);
nor U13244 (N_13244,N_12960,N_13059);
nor U13245 (N_13245,N_13100,N_13079);
or U13246 (N_13246,N_13004,N_13016);
nand U13247 (N_13247,N_13112,N_13019);
and U13248 (N_13248,N_13074,N_13025);
nand U13249 (N_13249,N_13072,N_12970);
nor U13250 (N_13250,N_13047,N_13050);
or U13251 (N_13251,N_13011,N_12987);
nand U13252 (N_13252,N_13072,N_12995);
and U13253 (N_13253,N_13050,N_13084);
or U13254 (N_13254,N_13117,N_13045);
xor U13255 (N_13255,N_12995,N_12984);
nor U13256 (N_13256,N_13040,N_12983);
nor U13257 (N_13257,N_13076,N_13099);
xor U13258 (N_13258,N_13078,N_13020);
or U13259 (N_13259,N_13008,N_13052);
nor U13260 (N_13260,N_13057,N_13030);
nor U13261 (N_13261,N_12994,N_13089);
and U13262 (N_13262,N_13001,N_13050);
or U13263 (N_13263,N_13023,N_13056);
and U13264 (N_13264,N_13101,N_13090);
and U13265 (N_13265,N_13012,N_12981);
or U13266 (N_13266,N_13021,N_13025);
nand U13267 (N_13267,N_13063,N_13014);
nand U13268 (N_13268,N_13093,N_13099);
nor U13269 (N_13269,N_13014,N_12975);
nand U13270 (N_13270,N_13056,N_13097);
xor U13271 (N_13271,N_12987,N_12983);
nor U13272 (N_13272,N_12961,N_12962);
nor U13273 (N_13273,N_12990,N_13017);
xor U13274 (N_13274,N_12993,N_13015);
nand U13275 (N_13275,N_12980,N_13053);
xnor U13276 (N_13276,N_13114,N_12994);
nor U13277 (N_13277,N_13075,N_13005);
or U13278 (N_13278,N_13045,N_13114);
xnor U13279 (N_13279,N_13100,N_13057);
and U13280 (N_13280,N_13255,N_13202);
nor U13281 (N_13281,N_13271,N_13264);
and U13282 (N_13282,N_13241,N_13142);
or U13283 (N_13283,N_13262,N_13183);
or U13284 (N_13284,N_13199,N_13127);
nand U13285 (N_13285,N_13191,N_13216);
or U13286 (N_13286,N_13238,N_13252);
nor U13287 (N_13287,N_13133,N_13215);
or U13288 (N_13288,N_13151,N_13134);
and U13289 (N_13289,N_13177,N_13175);
and U13290 (N_13290,N_13274,N_13196);
nand U13291 (N_13291,N_13254,N_13146);
nand U13292 (N_13292,N_13275,N_13123);
nand U13293 (N_13293,N_13176,N_13157);
and U13294 (N_13294,N_13145,N_13223);
or U13295 (N_13295,N_13237,N_13180);
nand U13296 (N_13296,N_13273,N_13167);
nand U13297 (N_13297,N_13149,N_13169);
xnor U13298 (N_13298,N_13267,N_13230);
and U13299 (N_13299,N_13235,N_13265);
nand U13300 (N_13300,N_13179,N_13189);
or U13301 (N_13301,N_13239,N_13144);
nor U13302 (N_13302,N_13270,N_13168);
or U13303 (N_13303,N_13227,N_13212);
and U13304 (N_13304,N_13170,N_13128);
or U13305 (N_13305,N_13186,N_13135);
and U13306 (N_13306,N_13259,N_13185);
nor U13307 (N_13307,N_13165,N_13210);
and U13308 (N_13308,N_13250,N_13206);
or U13309 (N_13309,N_13207,N_13173);
and U13310 (N_13310,N_13218,N_13159);
or U13311 (N_13311,N_13171,N_13193);
nor U13312 (N_13312,N_13122,N_13152);
or U13313 (N_13313,N_13174,N_13263);
or U13314 (N_13314,N_13163,N_13245);
nor U13315 (N_13315,N_13147,N_13164);
nand U13316 (N_13316,N_13233,N_13221);
and U13317 (N_13317,N_13234,N_13125);
nor U13318 (N_13318,N_13261,N_13187);
and U13319 (N_13319,N_13132,N_13139);
nand U13320 (N_13320,N_13258,N_13197);
nand U13321 (N_13321,N_13278,N_13160);
and U13322 (N_13322,N_13126,N_13143);
nand U13323 (N_13323,N_13224,N_13182);
nand U13324 (N_13324,N_13242,N_13244);
or U13325 (N_13325,N_13148,N_13236);
nor U13326 (N_13326,N_13153,N_13194);
xor U13327 (N_13327,N_13130,N_13256);
or U13328 (N_13328,N_13124,N_13154);
and U13329 (N_13329,N_13162,N_13257);
nor U13330 (N_13330,N_13172,N_13226);
and U13331 (N_13331,N_13214,N_13120);
and U13332 (N_13332,N_13203,N_13141);
and U13333 (N_13333,N_13243,N_13181);
nor U13334 (N_13334,N_13136,N_13155);
nor U13335 (N_13335,N_13200,N_13208);
nand U13336 (N_13336,N_13232,N_13268);
nor U13337 (N_13337,N_13272,N_13138);
nor U13338 (N_13338,N_13231,N_13129);
or U13339 (N_13339,N_13166,N_13260);
nand U13340 (N_13340,N_13240,N_13229);
nor U13341 (N_13341,N_13251,N_13211);
and U13342 (N_13342,N_13201,N_13178);
nor U13343 (N_13343,N_13195,N_13269);
or U13344 (N_13344,N_13192,N_13198);
or U13345 (N_13345,N_13140,N_13277);
nor U13346 (N_13346,N_13161,N_13222);
xnor U13347 (N_13347,N_13188,N_13248);
nor U13348 (N_13348,N_13158,N_13246);
and U13349 (N_13349,N_13220,N_13131);
and U13350 (N_13350,N_13279,N_13213);
or U13351 (N_13351,N_13121,N_13156);
xor U13352 (N_13352,N_13228,N_13266);
xor U13353 (N_13353,N_13190,N_13209);
nor U13354 (N_13354,N_13150,N_13276);
xnor U13355 (N_13355,N_13217,N_13249);
nor U13356 (N_13356,N_13184,N_13204);
xnor U13357 (N_13357,N_13219,N_13225);
nor U13358 (N_13358,N_13253,N_13247);
nor U13359 (N_13359,N_13137,N_13205);
nand U13360 (N_13360,N_13268,N_13209);
or U13361 (N_13361,N_13227,N_13189);
xor U13362 (N_13362,N_13149,N_13136);
and U13363 (N_13363,N_13172,N_13123);
and U13364 (N_13364,N_13239,N_13161);
or U13365 (N_13365,N_13129,N_13222);
nand U13366 (N_13366,N_13268,N_13182);
nand U13367 (N_13367,N_13150,N_13254);
and U13368 (N_13368,N_13137,N_13183);
or U13369 (N_13369,N_13264,N_13127);
and U13370 (N_13370,N_13184,N_13207);
xor U13371 (N_13371,N_13212,N_13151);
nor U13372 (N_13372,N_13146,N_13213);
and U13373 (N_13373,N_13212,N_13268);
xnor U13374 (N_13374,N_13146,N_13257);
nand U13375 (N_13375,N_13215,N_13200);
and U13376 (N_13376,N_13226,N_13230);
nor U13377 (N_13377,N_13209,N_13146);
or U13378 (N_13378,N_13268,N_13145);
nor U13379 (N_13379,N_13188,N_13232);
nor U13380 (N_13380,N_13127,N_13187);
or U13381 (N_13381,N_13232,N_13263);
or U13382 (N_13382,N_13234,N_13204);
and U13383 (N_13383,N_13277,N_13270);
nor U13384 (N_13384,N_13210,N_13204);
nand U13385 (N_13385,N_13156,N_13209);
xor U13386 (N_13386,N_13170,N_13277);
or U13387 (N_13387,N_13205,N_13167);
and U13388 (N_13388,N_13141,N_13222);
nand U13389 (N_13389,N_13276,N_13271);
nor U13390 (N_13390,N_13272,N_13150);
or U13391 (N_13391,N_13246,N_13213);
or U13392 (N_13392,N_13190,N_13174);
nand U13393 (N_13393,N_13276,N_13279);
or U13394 (N_13394,N_13181,N_13186);
or U13395 (N_13395,N_13184,N_13160);
nand U13396 (N_13396,N_13156,N_13266);
nor U13397 (N_13397,N_13208,N_13178);
or U13398 (N_13398,N_13163,N_13165);
or U13399 (N_13399,N_13274,N_13143);
or U13400 (N_13400,N_13233,N_13262);
and U13401 (N_13401,N_13125,N_13207);
and U13402 (N_13402,N_13185,N_13155);
or U13403 (N_13403,N_13133,N_13137);
nand U13404 (N_13404,N_13233,N_13216);
and U13405 (N_13405,N_13237,N_13204);
nand U13406 (N_13406,N_13260,N_13214);
and U13407 (N_13407,N_13215,N_13142);
nand U13408 (N_13408,N_13229,N_13275);
nand U13409 (N_13409,N_13223,N_13206);
or U13410 (N_13410,N_13156,N_13260);
nor U13411 (N_13411,N_13225,N_13275);
xnor U13412 (N_13412,N_13199,N_13164);
and U13413 (N_13413,N_13219,N_13166);
and U13414 (N_13414,N_13165,N_13164);
xnor U13415 (N_13415,N_13258,N_13240);
xor U13416 (N_13416,N_13260,N_13160);
nor U13417 (N_13417,N_13183,N_13249);
xor U13418 (N_13418,N_13155,N_13276);
and U13419 (N_13419,N_13224,N_13147);
and U13420 (N_13420,N_13240,N_13255);
or U13421 (N_13421,N_13138,N_13253);
nand U13422 (N_13422,N_13156,N_13120);
and U13423 (N_13423,N_13275,N_13189);
nor U13424 (N_13424,N_13191,N_13183);
nor U13425 (N_13425,N_13254,N_13214);
xor U13426 (N_13426,N_13243,N_13188);
and U13427 (N_13427,N_13270,N_13164);
nor U13428 (N_13428,N_13191,N_13224);
or U13429 (N_13429,N_13177,N_13187);
nor U13430 (N_13430,N_13273,N_13262);
nor U13431 (N_13431,N_13206,N_13222);
and U13432 (N_13432,N_13232,N_13246);
nor U13433 (N_13433,N_13174,N_13233);
nand U13434 (N_13434,N_13217,N_13232);
or U13435 (N_13435,N_13174,N_13254);
or U13436 (N_13436,N_13220,N_13185);
and U13437 (N_13437,N_13184,N_13153);
and U13438 (N_13438,N_13141,N_13187);
nand U13439 (N_13439,N_13276,N_13194);
or U13440 (N_13440,N_13383,N_13398);
or U13441 (N_13441,N_13282,N_13433);
or U13442 (N_13442,N_13329,N_13407);
and U13443 (N_13443,N_13333,N_13375);
nor U13444 (N_13444,N_13369,N_13303);
nor U13445 (N_13445,N_13411,N_13323);
or U13446 (N_13446,N_13405,N_13352);
and U13447 (N_13447,N_13318,N_13364);
xnor U13448 (N_13448,N_13335,N_13334);
nor U13449 (N_13449,N_13302,N_13362);
nor U13450 (N_13450,N_13416,N_13321);
nor U13451 (N_13451,N_13366,N_13434);
and U13452 (N_13452,N_13314,N_13382);
nand U13453 (N_13453,N_13377,N_13308);
xnor U13454 (N_13454,N_13388,N_13307);
nor U13455 (N_13455,N_13344,N_13389);
and U13456 (N_13456,N_13378,N_13316);
nand U13457 (N_13457,N_13292,N_13370);
or U13458 (N_13458,N_13418,N_13356);
or U13459 (N_13459,N_13349,N_13331);
nor U13460 (N_13460,N_13410,N_13409);
and U13461 (N_13461,N_13320,N_13286);
and U13462 (N_13462,N_13295,N_13431);
or U13463 (N_13463,N_13430,N_13357);
nor U13464 (N_13464,N_13404,N_13290);
or U13465 (N_13465,N_13327,N_13392);
or U13466 (N_13466,N_13422,N_13421);
nand U13467 (N_13467,N_13428,N_13293);
and U13468 (N_13468,N_13435,N_13285);
and U13469 (N_13469,N_13399,N_13347);
nor U13470 (N_13470,N_13312,N_13313);
nand U13471 (N_13471,N_13351,N_13337);
nor U13472 (N_13472,N_13380,N_13424);
and U13473 (N_13473,N_13339,N_13374);
nand U13474 (N_13474,N_13400,N_13301);
nor U13475 (N_13475,N_13420,N_13324);
xnor U13476 (N_13476,N_13358,N_13336);
and U13477 (N_13477,N_13319,N_13298);
nand U13478 (N_13478,N_13294,N_13414);
or U13479 (N_13479,N_13417,N_13376);
nand U13480 (N_13480,N_13309,N_13340);
nor U13481 (N_13481,N_13311,N_13300);
and U13482 (N_13482,N_13345,N_13342);
nor U13483 (N_13483,N_13287,N_13426);
nand U13484 (N_13484,N_13401,N_13284);
or U13485 (N_13485,N_13281,N_13332);
and U13486 (N_13486,N_13427,N_13338);
or U13487 (N_13487,N_13305,N_13363);
and U13488 (N_13488,N_13304,N_13341);
nand U13489 (N_13489,N_13436,N_13406);
nand U13490 (N_13490,N_13432,N_13346);
nor U13491 (N_13491,N_13322,N_13385);
nor U13492 (N_13492,N_13423,N_13361);
and U13493 (N_13493,N_13368,N_13354);
or U13494 (N_13494,N_13429,N_13289);
and U13495 (N_13495,N_13373,N_13437);
and U13496 (N_13496,N_13412,N_13330);
and U13497 (N_13497,N_13360,N_13381);
nand U13498 (N_13498,N_13390,N_13291);
xor U13499 (N_13499,N_13413,N_13365);
nor U13500 (N_13500,N_13283,N_13394);
nand U13501 (N_13501,N_13350,N_13325);
and U13502 (N_13502,N_13419,N_13396);
nor U13503 (N_13503,N_13379,N_13372);
nand U13504 (N_13504,N_13297,N_13403);
nand U13505 (N_13505,N_13408,N_13326);
or U13506 (N_13506,N_13402,N_13353);
nand U13507 (N_13507,N_13425,N_13355);
or U13508 (N_13508,N_13393,N_13359);
nand U13509 (N_13509,N_13310,N_13367);
nor U13510 (N_13510,N_13306,N_13391);
xnor U13511 (N_13511,N_13317,N_13386);
nor U13512 (N_13512,N_13299,N_13328);
or U13513 (N_13513,N_13315,N_13387);
xnor U13514 (N_13514,N_13371,N_13384);
and U13515 (N_13515,N_13288,N_13296);
or U13516 (N_13516,N_13343,N_13395);
nand U13517 (N_13517,N_13397,N_13348);
nor U13518 (N_13518,N_13439,N_13415);
xor U13519 (N_13519,N_13280,N_13438);
xor U13520 (N_13520,N_13407,N_13310);
nand U13521 (N_13521,N_13337,N_13354);
and U13522 (N_13522,N_13341,N_13372);
or U13523 (N_13523,N_13358,N_13339);
or U13524 (N_13524,N_13434,N_13344);
nand U13525 (N_13525,N_13308,N_13412);
or U13526 (N_13526,N_13305,N_13437);
xor U13527 (N_13527,N_13297,N_13335);
xnor U13528 (N_13528,N_13412,N_13341);
or U13529 (N_13529,N_13433,N_13325);
nand U13530 (N_13530,N_13412,N_13404);
and U13531 (N_13531,N_13300,N_13381);
nor U13532 (N_13532,N_13283,N_13380);
nand U13533 (N_13533,N_13396,N_13386);
nor U13534 (N_13534,N_13295,N_13331);
or U13535 (N_13535,N_13438,N_13314);
and U13536 (N_13536,N_13405,N_13325);
and U13537 (N_13537,N_13350,N_13368);
nand U13538 (N_13538,N_13290,N_13396);
or U13539 (N_13539,N_13381,N_13415);
nor U13540 (N_13540,N_13307,N_13397);
or U13541 (N_13541,N_13356,N_13344);
nand U13542 (N_13542,N_13360,N_13344);
or U13543 (N_13543,N_13436,N_13318);
xor U13544 (N_13544,N_13407,N_13332);
xnor U13545 (N_13545,N_13361,N_13326);
nand U13546 (N_13546,N_13323,N_13417);
or U13547 (N_13547,N_13359,N_13310);
nand U13548 (N_13548,N_13418,N_13387);
and U13549 (N_13549,N_13370,N_13351);
or U13550 (N_13550,N_13422,N_13321);
xor U13551 (N_13551,N_13432,N_13291);
and U13552 (N_13552,N_13403,N_13322);
nor U13553 (N_13553,N_13431,N_13426);
or U13554 (N_13554,N_13416,N_13382);
nand U13555 (N_13555,N_13309,N_13322);
nand U13556 (N_13556,N_13332,N_13385);
nand U13557 (N_13557,N_13349,N_13313);
or U13558 (N_13558,N_13292,N_13385);
nand U13559 (N_13559,N_13378,N_13435);
or U13560 (N_13560,N_13330,N_13426);
or U13561 (N_13561,N_13339,N_13331);
or U13562 (N_13562,N_13437,N_13343);
nor U13563 (N_13563,N_13354,N_13403);
nor U13564 (N_13564,N_13422,N_13328);
xnor U13565 (N_13565,N_13423,N_13315);
xnor U13566 (N_13566,N_13385,N_13423);
or U13567 (N_13567,N_13407,N_13437);
nand U13568 (N_13568,N_13305,N_13311);
nand U13569 (N_13569,N_13336,N_13414);
nand U13570 (N_13570,N_13395,N_13424);
nor U13571 (N_13571,N_13368,N_13359);
nand U13572 (N_13572,N_13348,N_13396);
xnor U13573 (N_13573,N_13348,N_13333);
nand U13574 (N_13574,N_13361,N_13374);
nand U13575 (N_13575,N_13313,N_13314);
nand U13576 (N_13576,N_13365,N_13307);
or U13577 (N_13577,N_13320,N_13398);
nand U13578 (N_13578,N_13318,N_13386);
nor U13579 (N_13579,N_13334,N_13435);
or U13580 (N_13580,N_13332,N_13356);
nand U13581 (N_13581,N_13409,N_13355);
nor U13582 (N_13582,N_13390,N_13394);
or U13583 (N_13583,N_13409,N_13343);
nand U13584 (N_13584,N_13324,N_13332);
nor U13585 (N_13585,N_13423,N_13348);
nor U13586 (N_13586,N_13326,N_13402);
nand U13587 (N_13587,N_13340,N_13369);
nand U13588 (N_13588,N_13369,N_13307);
nor U13589 (N_13589,N_13379,N_13354);
and U13590 (N_13590,N_13381,N_13328);
nand U13591 (N_13591,N_13404,N_13352);
nand U13592 (N_13592,N_13303,N_13332);
or U13593 (N_13593,N_13398,N_13433);
nor U13594 (N_13594,N_13364,N_13391);
nor U13595 (N_13595,N_13346,N_13332);
or U13596 (N_13596,N_13390,N_13389);
nor U13597 (N_13597,N_13302,N_13417);
xnor U13598 (N_13598,N_13323,N_13416);
nand U13599 (N_13599,N_13369,N_13321);
and U13600 (N_13600,N_13570,N_13545);
nor U13601 (N_13601,N_13521,N_13448);
or U13602 (N_13602,N_13532,N_13515);
or U13603 (N_13603,N_13556,N_13476);
nor U13604 (N_13604,N_13487,N_13473);
and U13605 (N_13605,N_13488,N_13577);
or U13606 (N_13606,N_13441,N_13548);
or U13607 (N_13607,N_13454,N_13520);
and U13608 (N_13608,N_13466,N_13581);
or U13609 (N_13609,N_13584,N_13455);
or U13610 (N_13610,N_13541,N_13568);
and U13611 (N_13611,N_13567,N_13503);
and U13612 (N_13612,N_13586,N_13537);
or U13613 (N_13613,N_13543,N_13500);
nand U13614 (N_13614,N_13526,N_13593);
and U13615 (N_13615,N_13524,N_13599);
and U13616 (N_13616,N_13549,N_13538);
nor U13617 (N_13617,N_13546,N_13533);
nor U13618 (N_13618,N_13573,N_13480);
nor U13619 (N_13619,N_13459,N_13507);
nor U13620 (N_13620,N_13542,N_13529);
and U13621 (N_13621,N_13453,N_13519);
xor U13622 (N_13622,N_13514,N_13564);
or U13623 (N_13623,N_13562,N_13484);
nand U13624 (N_13624,N_13591,N_13475);
and U13625 (N_13625,N_13540,N_13592);
nand U13626 (N_13626,N_13569,N_13530);
xor U13627 (N_13627,N_13497,N_13518);
nand U13628 (N_13628,N_13580,N_13494);
nor U13629 (N_13629,N_13486,N_13464);
and U13630 (N_13630,N_13574,N_13485);
nor U13631 (N_13631,N_13547,N_13445);
or U13632 (N_13632,N_13481,N_13536);
nand U13633 (N_13633,N_13516,N_13510);
and U13634 (N_13634,N_13463,N_13531);
nand U13635 (N_13635,N_13506,N_13499);
or U13636 (N_13636,N_13490,N_13550);
and U13637 (N_13637,N_13469,N_13461);
nor U13638 (N_13638,N_13496,N_13451);
and U13639 (N_13639,N_13509,N_13582);
and U13640 (N_13640,N_13458,N_13470);
or U13641 (N_13641,N_13444,N_13528);
nor U13642 (N_13642,N_13495,N_13557);
and U13643 (N_13643,N_13452,N_13501);
or U13644 (N_13644,N_13561,N_13551);
xnor U13645 (N_13645,N_13560,N_13576);
or U13646 (N_13646,N_13527,N_13525);
or U13647 (N_13647,N_13544,N_13558);
and U13648 (N_13648,N_13447,N_13585);
or U13649 (N_13649,N_13523,N_13565);
or U13650 (N_13650,N_13478,N_13589);
and U13651 (N_13651,N_13552,N_13502);
and U13652 (N_13652,N_13512,N_13498);
nor U13653 (N_13653,N_13443,N_13553);
and U13654 (N_13654,N_13493,N_13467);
or U13655 (N_13655,N_13554,N_13457);
or U13656 (N_13656,N_13472,N_13471);
and U13657 (N_13657,N_13555,N_13559);
xnor U13658 (N_13658,N_13578,N_13479);
nand U13659 (N_13659,N_13442,N_13579);
nand U13660 (N_13660,N_13513,N_13590);
or U13661 (N_13661,N_13460,N_13504);
nand U13662 (N_13662,N_13598,N_13508);
nor U13663 (N_13663,N_13440,N_13597);
nand U13664 (N_13664,N_13572,N_13587);
nor U13665 (N_13665,N_13595,N_13456);
nor U13666 (N_13666,N_13534,N_13449);
nand U13667 (N_13667,N_13575,N_13511);
and U13668 (N_13668,N_13596,N_13462);
and U13669 (N_13669,N_13468,N_13492);
nor U13670 (N_13670,N_13489,N_13539);
or U13671 (N_13671,N_13588,N_13491);
nor U13672 (N_13672,N_13477,N_13522);
or U13673 (N_13673,N_13450,N_13482);
and U13674 (N_13674,N_13474,N_13465);
or U13675 (N_13675,N_13535,N_13517);
nand U13676 (N_13676,N_13563,N_13446);
nand U13677 (N_13677,N_13566,N_13571);
nand U13678 (N_13678,N_13583,N_13594);
and U13679 (N_13679,N_13505,N_13483);
nand U13680 (N_13680,N_13545,N_13450);
nor U13681 (N_13681,N_13579,N_13516);
nand U13682 (N_13682,N_13598,N_13586);
nand U13683 (N_13683,N_13505,N_13472);
nor U13684 (N_13684,N_13523,N_13479);
nor U13685 (N_13685,N_13477,N_13580);
nand U13686 (N_13686,N_13444,N_13540);
or U13687 (N_13687,N_13522,N_13517);
nand U13688 (N_13688,N_13552,N_13495);
xor U13689 (N_13689,N_13455,N_13568);
and U13690 (N_13690,N_13548,N_13539);
nand U13691 (N_13691,N_13564,N_13522);
and U13692 (N_13692,N_13581,N_13583);
or U13693 (N_13693,N_13577,N_13565);
or U13694 (N_13694,N_13599,N_13550);
nor U13695 (N_13695,N_13490,N_13464);
nor U13696 (N_13696,N_13451,N_13552);
or U13697 (N_13697,N_13491,N_13461);
and U13698 (N_13698,N_13521,N_13490);
and U13699 (N_13699,N_13462,N_13461);
nand U13700 (N_13700,N_13472,N_13460);
nand U13701 (N_13701,N_13475,N_13569);
and U13702 (N_13702,N_13494,N_13564);
or U13703 (N_13703,N_13499,N_13559);
nand U13704 (N_13704,N_13542,N_13513);
or U13705 (N_13705,N_13440,N_13491);
and U13706 (N_13706,N_13523,N_13489);
nor U13707 (N_13707,N_13551,N_13553);
and U13708 (N_13708,N_13557,N_13442);
or U13709 (N_13709,N_13452,N_13548);
nor U13710 (N_13710,N_13442,N_13587);
and U13711 (N_13711,N_13554,N_13591);
nand U13712 (N_13712,N_13590,N_13546);
and U13713 (N_13713,N_13511,N_13542);
and U13714 (N_13714,N_13568,N_13504);
or U13715 (N_13715,N_13556,N_13497);
nor U13716 (N_13716,N_13593,N_13567);
or U13717 (N_13717,N_13581,N_13482);
nor U13718 (N_13718,N_13462,N_13510);
nand U13719 (N_13719,N_13482,N_13559);
xor U13720 (N_13720,N_13483,N_13521);
nor U13721 (N_13721,N_13579,N_13576);
nor U13722 (N_13722,N_13459,N_13516);
or U13723 (N_13723,N_13457,N_13485);
nor U13724 (N_13724,N_13552,N_13487);
and U13725 (N_13725,N_13503,N_13491);
or U13726 (N_13726,N_13490,N_13461);
and U13727 (N_13727,N_13563,N_13482);
and U13728 (N_13728,N_13483,N_13500);
and U13729 (N_13729,N_13591,N_13582);
nor U13730 (N_13730,N_13471,N_13461);
nor U13731 (N_13731,N_13440,N_13566);
or U13732 (N_13732,N_13441,N_13559);
and U13733 (N_13733,N_13546,N_13489);
nor U13734 (N_13734,N_13592,N_13475);
or U13735 (N_13735,N_13447,N_13535);
and U13736 (N_13736,N_13597,N_13565);
nor U13737 (N_13737,N_13502,N_13581);
or U13738 (N_13738,N_13598,N_13542);
and U13739 (N_13739,N_13550,N_13508);
or U13740 (N_13740,N_13558,N_13443);
nand U13741 (N_13741,N_13497,N_13583);
xor U13742 (N_13742,N_13530,N_13511);
nand U13743 (N_13743,N_13579,N_13510);
xnor U13744 (N_13744,N_13529,N_13448);
or U13745 (N_13745,N_13518,N_13457);
nor U13746 (N_13746,N_13523,N_13500);
nand U13747 (N_13747,N_13462,N_13491);
or U13748 (N_13748,N_13442,N_13565);
xnor U13749 (N_13749,N_13445,N_13552);
or U13750 (N_13750,N_13575,N_13480);
or U13751 (N_13751,N_13536,N_13512);
and U13752 (N_13752,N_13462,N_13509);
nand U13753 (N_13753,N_13586,N_13592);
and U13754 (N_13754,N_13540,N_13557);
nand U13755 (N_13755,N_13535,N_13564);
nand U13756 (N_13756,N_13457,N_13530);
and U13757 (N_13757,N_13589,N_13542);
nand U13758 (N_13758,N_13468,N_13597);
nand U13759 (N_13759,N_13442,N_13572);
nand U13760 (N_13760,N_13604,N_13642);
nor U13761 (N_13761,N_13721,N_13671);
or U13762 (N_13762,N_13683,N_13648);
nor U13763 (N_13763,N_13757,N_13708);
xor U13764 (N_13764,N_13653,N_13700);
nor U13765 (N_13765,N_13675,N_13670);
or U13766 (N_13766,N_13691,N_13698);
nor U13767 (N_13767,N_13684,N_13631);
nand U13768 (N_13768,N_13661,N_13738);
and U13769 (N_13769,N_13749,N_13693);
nor U13770 (N_13770,N_13742,N_13727);
nor U13771 (N_13771,N_13603,N_13645);
xnor U13772 (N_13772,N_13623,N_13625);
nor U13773 (N_13773,N_13696,N_13743);
and U13774 (N_13774,N_13664,N_13643);
nor U13775 (N_13775,N_13620,N_13614);
xnor U13776 (N_13776,N_13687,N_13607);
xor U13777 (N_13777,N_13739,N_13612);
xor U13778 (N_13778,N_13730,N_13712);
and U13779 (N_13779,N_13688,N_13704);
or U13780 (N_13780,N_13679,N_13735);
nor U13781 (N_13781,N_13690,N_13650);
and U13782 (N_13782,N_13723,N_13674);
xnor U13783 (N_13783,N_13668,N_13699);
nand U13784 (N_13784,N_13647,N_13662);
nor U13785 (N_13785,N_13710,N_13740);
or U13786 (N_13786,N_13616,N_13628);
and U13787 (N_13787,N_13666,N_13750);
and U13788 (N_13788,N_13609,N_13720);
nor U13789 (N_13789,N_13618,N_13641);
nor U13790 (N_13790,N_13639,N_13713);
nor U13791 (N_13791,N_13747,N_13619);
nand U13792 (N_13792,N_13706,N_13644);
nor U13793 (N_13793,N_13621,N_13652);
nand U13794 (N_13794,N_13629,N_13633);
nor U13795 (N_13795,N_13694,N_13680);
nor U13796 (N_13796,N_13686,N_13718);
xnor U13797 (N_13797,N_13677,N_13728);
nor U13798 (N_13798,N_13663,N_13709);
and U13799 (N_13799,N_13703,N_13751);
nor U13800 (N_13800,N_13654,N_13719);
nand U13801 (N_13801,N_13759,N_13657);
nand U13802 (N_13802,N_13758,N_13660);
nand U13803 (N_13803,N_13689,N_13697);
nand U13804 (N_13804,N_13729,N_13608);
nand U13805 (N_13805,N_13613,N_13756);
and U13806 (N_13806,N_13717,N_13725);
or U13807 (N_13807,N_13655,N_13702);
and U13808 (N_13808,N_13611,N_13673);
nand U13809 (N_13809,N_13715,N_13634);
and U13810 (N_13810,N_13748,N_13617);
or U13811 (N_13811,N_13640,N_13755);
and U13812 (N_13812,N_13605,N_13737);
nand U13813 (N_13813,N_13632,N_13732);
nor U13814 (N_13814,N_13635,N_13745);
and U13815 (N_13815,N_13736,N_13746);
nand U13816 (N_13816,N_13602,N_13622);
and U13817 (N_13817,N_13624,N_13658);
and U13818 (N_13818,N_13659,N_13733);
nor U13819 (N_13819,N_13754,N_13726);
xnor U13820 (N_13820,N_13667,N_13716);
xnor U13821 (N_13821,N_13741,N_13665);
nor U13822 (N_13822,N_13627,N_13734);
and U13823 (N_13823,N_13707,N_13711);
nand U13824 (N_13824,N_13606,N_13681);
and U13825 (N_13825,N_13601,N_13637);
nor U13826 (N_13826,N_13600,N_13646);
nand U13827 (N_13827,N_13669,N_13744);
nand U13828 (N_13828,N_13731,N_13610);
nand U13829 (N_13829,N_13676,N_13638);
nor U13830 (N_13830,N_13753,N_13695);
nand U13831 (N_13831,N_13651,N_13626);
or U13832 (N_13832,N_13722,N_13649);
nor U13833 (N_13833,N_13752,N_13630);
and U13834 (N_13834,N_13705,N_13615);
or U13835 (N_13835,N_13656,N_13682);
nor U13836 (N_13836,N_13636,N_13714);
nor U13837 (N_13837,N_13672,N_13701);
nor U13838 (N_13838,N_13724,N_13692);
nor U13839 (N_13839,N_13678,N_13685);
nand U13840 (N_13840,N_13680,N_13633);
nand U13841 (N_13841,N_13718,N_13654);
nand U13842 (N_13842,N_13754,N_13731);
and U13843 (N_13843,N_13714,N_13618);
or U13844 (N_13844,N_13614,N_13626);
or U13845 (N_13845,N_13646,N_13650);
xnor U13846 (N_13846,N_13687,N_13638);
nand U13847 (N_13847,N_13746,N_13678);
or U13848 (N_13848,N_13676,N_13733);
nand U13849 (N_13849,N_13673,N_13633);
xor U13850 (N_13850,N_13687,N_13647);
and U13851 (N_13851,N_13683,N_13643);
xnor U13852 (N_13852,N_13642,N_13738);
nor U13853 (N_13853,N_13641,N_13670);
or U13854 (N_13854,N_13612,N_13688);
nor U13855 (N_13855,N_13692,N_13713);
xor U13856 (N_13856,N_13652,N_13649);
xor U13857 (N_13857,N_13620,N_13659);
or U13858 (N_13858,N_13688,N_13750);
or U13859 (N_13859,N_13622,N_13705);
and U13860 (N_13860,N_13650,N_13720);
and U13861 (N_13861,N_13656,N_13614);
nor U13862 (N_13862,N_13692,N_13638);
nand U13863 (N_13863,N_13720,N_13718);
or U13864 (N_13864,N_13660,N_13609);
and U13865 (N_13865,N_13747,N_13622);
xnor U13866 (N_13866,N_13651,N_13607);
and U13867 (N_13867,N_13661,N_13633);
and U13868 (N_13868,N_13616,N_13727);
or U13869 (N_13869,N_13757,N_13647);
nand U13870 (N_13870,N_13653,N_13749);
or U13871 (N_13871,N_13621,N_13618);
nand U13872 (N_13872,N_13729,N_13710);
nor U13873 (N_13873,N_13692,N_13723);
nand U13874 (N_13874,N_13685,N_13670);
nor U13875 (N_13875,N_13746,N_13733);
and U13876 (N_13876,N_13742,N_13676);
or U13877 (N_13877,N_13734,N_13724);
or U13878 (N_13878,N_13694,N_13725);
and U13879 (N_13879,N_13730,N_13638);
xnor U13880 (N_13880,N_13750,N_13680);
and U13881 (N_13881,N_13607,N_13639);
nand U13882 (N_13882,N_13754,N_13643);
or U13883 (N_13883,N_13722,N_13732);
nor U13884 (N_13884,N_13669,N_13682);
nor U13885 (N_13885,N_13719,N_13692);
nand U13886 (N_13886,N_13672,N_13614);
or U13887 (N_13887,N_13688,N_13657);
xnor U13888 (N_13888,N_13688,N_13739);
nor U13889 (N_13889,N_13725,N_13640);
and U13890 (N_13890,N_13697,N_13661);
nor U13891 (N_13891,N_13674,N_13678);
nand U13892 (N_13892,N_13633,N_13711);
and U13893 (N_13893,N_13612,N_13715);
and U13894 (N_13894,N_13610,N_13688);
and U13895 (N_13895,N_13648,N_13642);
and U13896 (N_13896,N_13714,N_13655);
nor U13897 (N_13897,N_13720,N_13757);
nor U13898 (N_13898,N_13610,N_13652);
nand U13899 (N_13899,N_13661,N_13651);
nor U13900 (N_13900,N_13681,N_13711);
nor U13901 (N_13901,N_13662,N_13741);
and U13902 (N_13902,N_13754,N_13752);
nand U13903 (N_13903,N_13694,N_13670);
and U13904 (N_13904,N_13739,N_13613);
and U13905 (N_13905,N_13663,N_13704);
nor U13906 (N_13906,N_13663,N_13745);
nor U13907 (N_13907,N_13670,N_13754);
or U13908 (N_13908,N_13612,N_13722);
nand U13909 (N_13909,N_13752,N_13623);
nand U13910 (N_13910,N_13688,N_13743);
xnor U13911 (N_13911,N_13627,N_13675);
nor U13912 (N_13912,N_13752,N_13632);
nand U13913 (N_13913,N_13653,N_13614);
nand U13914 (N_13914,N_13665,N_13755);
or U13915 (N_13915,N_13679,N_13643);
and U13916 (N_13916,N_13634,N_13757);
and U13917 (N_13917,N_13679,N_13710);
nand U13918 (N_13918,N_13690,N_13695);
and U13919 (N_13919,N_13616,N_13697);
and U13920 (N_13920,N_13881,N_13858);
nand U13921 (N_13921,N_13868,N_13894);
nor U13922 (N_13922,N_13760,N_13834);
nor U13923 (N_13923,N_13790,N_13896);
nand U13924 (N_13924,N_13844,N_13827);
nor U13925 (N_13925,N_13783,N_13825);
and U13926 (N_13926,N_13883,N_13802);
and U13927 (N_13927,N_13807,N_13835);
nor U13928 (N_13928,N_13900,N_13848);
or U13929 (N_13929,N_13773,N_13917);
or U13930 (N_13930,N_13888,N_13795);
nand U13931 (N_13931,N_13903,N_13838);
or U13932 (N_13932,N_13822,N_13837);
or U13933 (N_13933,N_13819,N_13856);
nor U13934 (N_13934,N_13804,N_13919);
or U13935 (N_13935,N_13855,N_13885);
nor U13936 (N_13936,N_13869,N_13864);
or U13937 (N_13937,N_13785,N_13808);
nor U13938 (N_13938,N_13777,N_13876);
or U13939 (N_13939,N_13873,N_13870);
nand U13940 (N_13940,N_13763,N_13867);
xnor U13941 (N_13941,N_13779,N_13782);
and U13942 (N_13942,N_13914,N_13781);
nand U13943 (N_13943,N_13910,N_13771);
xnor U13944 (N_13944,N_13872,N_13915);
nor U13945 (N_13945,N_13798,N_13886);
or U13946 (N_13946,N_13843,N_13850);
nand U13947 (N_13947,N_13817,N_13871);
nand U13948 (N_13948,N_13810,N_13898);
nand U13949 (N_13949,N_13764,N_13895);
nand U13950 (N_13950,N_13788,N_13826);
xor U13951 (N_13951,N_13778,N_13828);
nor U13952 (N_13952,N_13904,N_13774);
nor U13953 (N_13953,N_13768,N_13784);
or U13954 (N_13954,N_13813,N_13880);
xor U13955 (N_13955,N_13776,N_13918);
nand U13956 (N_13956,N_13812,N_13860);
nor U13957 (N_13957,N_13824,N_13849);
xnor U13958 (N_13958,N_13806,N_13770);
or U13959 (N_13959,N_13799,N_13841);
nor U13960 (N_13960,N_13775,N_13809);
nor U13961 (N_13961,N_13890,N_13874);
nand U13962 (N_13962,N_13793,N_13911);
nor U13963 (N_13963,N_13803,N_13852);
or U13964 (N_13964,N_13907,N_13905);
and U13965 (N_13965,N_13893,N_13839);
or U13966 (N_13966,N_13902,N_13866);
or U13967 (N_13967,N_13859,N_13832);
and U13968 (N_13968,N_13851,N_13830);
or U13969 (N_13969,N_13865,N_13792);
and U13970 (N_13970,N_13801,N_13916);
nand U13971 (N_13971,N_13897,N_13796);
or U13972 (N_13972,N_13891,N_13889);
xnor U13973 (N_13973,N_13805,N_13829);
or U13974 (N_13974,N_13908,N_13786);
and U13975 (N_13975,N_13845,N_13901);
or U13976 (N_13976,N_13913,N_13846);
nor U13977 (N_13977,N_13840,N_13854);
and U13978 (N_13978,N_13791,N_13899);
nor U13979 (N_13979,N_13761,N_13857);
nor U13980 (N_13980,N_13831,N_13780);
xor U13981 (N_13981,N_13818,N_13877);
nor U13982 (N_13982,N_13789,N_13765);
and U13983 (N_13983,N_13882,N_13875);
or U13984 (N_13984,N_13794,N_13912);
or U13985 (N_13985,N_13847,N_13762);
nor U13986 (N_13986,N_13909,N_13816);
nand U13987 (N_13987,N_13820,N_13892);
or U13988 (N_13988,N_13766,N_13878);
or U13989 (N_13989,N_13769,N_13821);
nand U13990 (N_13990,N_13823,N_13767);
xor U13991 (N_13991,N_13842,N_13884);
xnor U13992 (N_13992,N_13862,N_13787);
nand U13993 (N_13993,N_13853,N_13797);
and U13994 (N_13994,N_13833,N_13879);
nor U13995 (N_13995,N_13815,N_13814);
xnor U13996 (N_13996,N_13836,N_13800);
and U13997 (N_13997,N_13811,N_13863);
and U13998 (N_13998,N_13772,N_13887);
or U13999 (N_13999,N_13906,N_13861);
or U14000 (N_14000,N_13770,N_13871);
nor U14001 (N_14001,N_13838,N_13833);
nor U14002 (N_14002,N_13906,N_13763);
nand U14003 (N_14003,N_13767,N_13820);
nand U14004 (N_14004,N_13901,N_13867);
nor U14005 (N_14005,N_13778,N_13894);
nand U14006 (N_14006,N_13860,N_13881);
and U14007 (N_14007,N_13789,N_13884);
or U14008 (N_14008,N_13797,N_13907);
and U14009 (N_14009,N_13852,N_13918);
nand U14010 (N_14010,N_13792,N_13838);
nor U14011 (N_14011,N_13810,N_13829);
nor U14012 (N_14012,N_13903,N_13795);
or U14013 (N_14013,N_13905,N_13813);
nor U14014 (N_14014,N_13809,N_13807);
nand U14015 (N_14015,N_13847,N_13761);
nor U14016 (N_14016,N_13858,N_13821);
nor U14017 (N_14017,N_13843,N_13888);
nor U14018 (N_14018,N_13777,N_13781);
or U14019 (N_14019,N_13867,N_13780);
and U14020 (N_14020,N_13903,N_13818);
nor U14021 (N_14021,N_13901,N_13789);
nand U14022 (N_14022,N_13846,N_13890);
or U14023 (N_14023,N_13875,N_13891);
nor U14024 (N_14024,N_13773,N_13901);
and U14025 (N_14025,N_13863,N_13898);
xnor U14026 (N_14026,N_13810,N_13841);
nor U14027 (N_14027,N_13792,N_13804);
or U14028 (N_14028,N_13874,N_13918);
nor U14029 (N_14029,N_13814,N_13792);
nor U14030 (N_14030,N_13844,N_13847);
nor U14031 (N_14031,N_13907,N_13829);
and U14032 (N_14032,N_13809,N_13835);
nor U14033 (N_14033,N_13833,N_13826);
or U14034 (N_14034,N_13884,N_13791);
nand U14035 (N_14035,N_13886,N_13832);
and U14036 (N_14036,N_13869,N_13906);
nor U14037 (N_14037,N_13849,N_13797);
nand U14038 (N_14038,N_13861,N_13880);
or U14039 (N_14039,N_13858,N_13901);
or U14040 (N_14040,N_13897,N_13882);
nand U14041 (N_14041,N_13775,N_13862);
nand U14042 (N_14042,N_13898,N_13837);
nor U14043 (N_14043,N_13811,N_13784);
nor U14044 (N_14044,N_13840,N_13784);
nor U14045 (N_14045,N_13913,N_13777);
nand U14046 (N_14046,N_13763,N_13783);
or U14047 (N_14047,N_13761,N_13870);
and U14048 (N_14048,N_13773,N_13823);
xnor U14049 (N_14049,N_13805,N_13843);
xor U14050 (N_14050,N_13876,N_13872);
nand U14051 (N_14051,N_13865,N_13894);
nand U14052 (N_14052,N_13876,N_13766);
and U14053 (N_14053,N_13875,N_13797);
or U14054 (N_14054,N_13770,N_13856);
nand U14055 (N_14055,N_13854,N_13904);
and U14056 (N_14056,N_13766,N_13790);
xnor U14057 (N_14057,N_13801,N_13777);
nor U14058 (N_14058,N_13819,N_13886);
nor U14059 (N_14059,N_13839,N_13917);
and U14060 (N_14060,N_13831,N_13889);
nor U14061 (N_14061,N_13775,N_13915);
nand U14062 (N_14062,N_13839,N_13765);
nor U14063 (N_14063,N_13871,N_13891);
and U14064 (N_14064,N_13794,N_13760);
nand U14065 (N_14065,N_13853,N_13793);
nand U14066 (N_14066,N_13881,N_13800);
nor U14067 (N_14067,N_13824,N_13806);
or U14068 (N_14068,N_13777,N_13818);
and U14069 (N_14069,N_13848,N_13855);
nand U14070 (N_14070,N_13804,N_13764);
and U14071 (N_14071,N_13895,N_13826);
nand U14072 (N_14072,N_13760,N_13805);
nor U14073 (N_14073,N_13862,N_13883);
and U14074 (N_14074,N_13913,N_13827);
nand U14075 (N_14075,N_13886,N_13773);
and U14076 (N_14076,N_13886,N_13849);
or U14077 (N_14077,N_13815,N_13834);
or U14078 (N_14078,N_13873,N_13871);
nor U14079 (N_14079,N_13828,N_13780);
or U14080 (N_14080,N_13973,N_14001);
nor U14081 (N_14081,N_14067,N_13967);
xnor U14082 (N_14082,N_14039,N_14061);
or U14083 (N_14083,N_14075,N_13995);
nand U14084 (N_14084,N_13956,N_13935);
and U14085 (N_14085,N_13978,N_14033);
and U14086 (N_14086,N_14032,N_14019);
nor U14087 (N_14087,N_13955,N_13997);
nor U14088 (N_14088,N_13941,N_13939);
nand U14089 (N_14089,N_14022,N_13996);
or U14090 (N_14090,N_14028,N_13976);
and U14091 (N_14091,N_14008,N_14047);
or U14092 (N_14092,N_13975,N_14025);
nand U14093 (N_14093,N_14042,N_14002);
nand U14094 (N_14094,N_13954,N_13926);
xnor U14095 (N_14095,N_13933,N_13940);
xor U14096 (N_14096,N_14030,N_13928);
nor U14097 (N_14097,N_13957,N_13922);
nor U14098 (N_14098,N_13920,N_13979);
nor U14099 (N_14099,N_14050,N_13929);
and U14100 (N_14100,N_14053,N_13931);
or U14101 (N_14101,N_14045,N_13945);
or U14102 (N_14102,N_14064,N_13977);
nand U14103 (N_14103,N_13943,N_14043);
or U14104 (N_14104,N_13934,N_13924);
and U14105 (N_14105,N_14077,N_14011);
nor U14106 (N_14106,N_13970,N_13993);
or U14107 (N_14107,N_14069,N_14010);
xnor U14108 (N_14108,N_13998,N_13982);
and U14109 (N_14109,N_13966,N_14057);
and U14110 (N_14110,N_14079,N_13927);
or U14111 (N_14111,N_13938,N_13988);
or U14112 (N_14112,N_14056,N_14015);
or U14113 (N_14113,N_14020,N_14065);
nand U14114 (N_14114,N_14071,N_14044);
nand U14115 (N_14115,N_13950,N_14023);
nor U14116 (N_14116,N_13930,N_14016);
nand U14117 (N_14117,N_13974,N_14068);
and U14118 (N_14118,N_13961,N_14070);
and U14119 (N_14119,N_14006,N_14024);
nor U14120 (N_14120,N_14021,N_13948);
nand U14121 (N_14121,N_14040,N_14049);
or U14122 (N_14122,N_13963,N_13983);
and U14123 (N_14123,N_13944,N_14013);
nor U14124 (N_14124,N_13968,N_14038);
xnor U14125 (N_14125,N_13984,N_13999);
and U14126 (N_14126,N_14005,N_13972);
nand U14127 (N_14127,N_14052,N_13942);
and U14128 (N_14128,N_14012,N_14007);
nand U14129 (N_14129,N_13921,N_14014);
nor U14130 (N_14130,N_13962,N_14074);
nand U14131 (N_14131,N_14063,N_14073);
nor U14132 (N_14132,N_13965,N_13986);
and U14133 (N_14133,N_14059,N_13992);
and U14134 (N_14134,N_13925,N_13994);
or U14135 (N_14135,N_13987,N_13923);
nor U14136 (N_14136,N_13951,N_13952);
nor U14137 (N_14137,N_13932,N_13969);
and U14138 (N_14138,N_14041,N_13960);
xnor U14139 (N_14139,N_13947,N_14035);
or U14140 (N_14140,N_14036,N_14055);
or U14141 (N_14141,N_14051,N_13991);
or U14142 (N_14142,N_14031,N_13964);
and U14143 (N_14143,N_14078,N_14060);
and U14144 (N_14144,N_14029,N_13989);
nor U14145 (N_14145,N_14018,N_14054);
nand U14146 (N_14146,N_13980,N_13981);
nor U14147 (N_14147,N_14076,N_13959);
nand U14148 (N_14148,N_14066,N_13946);
nor U14149 (N_14149,N_13937,N_13936);
and U14150 (N_14150,N_14058,N_14004);
nor U14151 (N_14151,N_14000,N_14037);
or U14152 (N_14152,N_14003,N_13958);
nand U14153 (N_14153,N_13990,N_14017);
and U14154 (N_14154,N_13985,N_14062);
nand U14155 (N_14155,N_13953,N_14009);
nor U14156 (N_14156,N_14027,N_14034);
xnor U14157 (N_14157,N_14072,N_14046);
and U14158 (N_14158,N_13949,N_13971);
and U14159 (N_14159,N_14048,N_14026);
and U14160 (N_14160,N_13979,N_14076);
nand U14161 (N_14161,N_14030,N_13971);
nand U14162 (N_14162,N_13942,N_13943);
nand U14163 (N_14163,N_14042,N_14056);
xnor U14164 (N_14164,N_13936,N_14000);
nand U14165 (N_14165,N_13988,N_13943);
or U14166 (N_14166,N_13946,N_13958);
nand U14167 (N_14167,N_14009,N_14067);
and U14168 (N_14168,N_14026,N_14047);
and U14169 (N_14169,N_14024,N_14023);
nor U14170 (N_14170,N_14027,N_13976);
xor U14171 (N_14171,N_13989,N_13981);
nand U14172 (N_14172,N_13986,N_14071);
nand U14173 (N_14173,N_13974,N_13963);
and U14174 (N_14174,N_14009,N_13925);
xnor U14175 (N_14175,N_13949,N_13942);
and U14176 (N_14176,N_14077,N_14056);
or U14177 (N_14177,N_13968,N_13949);
nor U14178 (N_14178,N_14028,N_13984);
nor U14179 (N_14179,N_13977,N_13958);
and U14180 (N_14180,N_13971,N_14042);
or U14181 (N_14181,N_13956,N_13940);
xnor U14182 (N_14182,N_14028,N_14034);
and U14183 (N_14183,N_13924,N_14008);
nand U14184 (N_14184,N_13971,N_14036);
or U14185 (N_14185,N_13984,N_14074);
and U14186 (N_14186,N_14008,N_13928);
or U14187 (N_14187,N_14079,N_13980);
or U14188 (N_14188,N_14070,N_14069);
nand U14189 (N_14189,N_14026,N_13955);
nand U14190 (N_14190,N_13946,N_13999);
and U14191 (N_14191,N_13996,N_14055);
or U14192 (N_14192,N_14074,N_13937);
or U14193 (N_14193,N_13981,N_14060);
nor U14194 (N_14194,N_14059,N_14048);
or U14195 (N_14195,N_14005,N_14016);
nor U14196 (N_14196,N_14015,N_14005);
and U14197 (N_14197,N_13990,N_13969);
nand U14198 (N_14198,N_13990,N_14003);
nor U14199 (N_14199,N_14024,N_14059);
and U14200 (N_14200,N_13949,N_13933);
or U14201 (N_14201,N_13950,N_13971);
or U14202 (N_14202,N_14042,N_13953);
nor U14203 (N_14203,N_13928,N_14053);
or U14204 (N_14204,N_13966,N_13998);
nor U14205 (N_14205,N_14039,N_13932);
and U14206 (N_14206,N_14006,N_14079);
and U14207 (N_14207,N_13965,N_13952);
nand U14208 (N_14208,N_14066,N_13997);
and U14209 (N_14209,N_13940,N_13960);
nand U14210 (N_14210,N_13988,N_13960);
xnor U14211 (N_14211,N_14025,N_13941);
nor U14212 (N_14212,N_13920,N_14027);
or U14213 (N_14213,N_14050,N_13973);
and U14214 (N_14214,N_13998,N_14020);
and U14215 (N_14215,N_14070,N_14047);
nor U14216 (N_14216,N_14052,N_13947);
and U14217 (N_14217,N_14045,N_14054);
nor U14218 (N_14218,N_14075,N_13992);
xnor U14219 (N_14219,N_13980,N_14031);
and U14220 (N_14220,N_14053,N_13987);
or U14221 (N_14221,N_14075,N_14051);
nor U14222 (N_14222,N_13966,N_14051);
nor U14223 (N_14223,N_14041,N_13945);
or U14224 (N_14224,N_14031,N_14034);
nand U14225 (N_14225,N_14059,N_13923);
nand U14226 (N_14226,N_14001,N_13928);
nor U14227 (N_14227,N_13921,N_13969);
nand U14228 (N_14228,N_14021,N_14035);
and U14229 (N_14229,N_13986,N_13970);
or U14230 (N_14230,N_13929,N_13948);
nor U14231 (N_14231,N_14051,N_13983);
nor U14232 (N_14232,N_14071,N_13924);
nor U14233 (N_14233,N_14039,N_13967);
and U14234 (N_14234,N_14076,N_14012);
and U14235 (N_14235,N_14038,N_13930);
and U14236 (N_14236,N_14058,N_13942);
or U14237 (N_14237,N_14027,N_13955);
nand U14238 (N_14238,N_13946,N_14002);
nor U14239 (N_14239,N_14053,N_13994);
or U14240 (N_14240,N_14099,N_14114);
or U14241 (N_14241,N_14132,N_14133);
nor U14242 (N_14242,N_14234,N_14188);
and U14243 (N_14243,N_14212,N_14210);
or U14244 (N_14244,N_14211,N_14093);
or U14245 (N_14245,N_14191,N_14120);
nor U14246 (N_14246,N_14083,N_14235);
or U14247 (N_14247,N_14228,N_14229);
and U14248 (N_14248,N_14080,N_14180);
nand U14249 (N_14249,N_14115,N_14110);
or U14250 (N_14250,N_14166,N_14217);
or U14251 (N_14251,N_14122,N_14109);
nor U14252 (N_14252,N_14124,N_14091);
and U14253 (N_14253,N_14206,N_14128);
or U14254 (N_14254,N_14216,N_14161);
nand U14255 (N_14255,N_14183,N_14088);
nor U14256 (N_14256,N_14104,N_14208);
or U14257 (N_14257,N_14193,N_14189);
and U14258 (N_14258,N_14136,N_14200);
nor U14259 (N_14259,N_14102,N_14186);
and U14260 (N_14260,N_14084,N_14129);
or U14261 (N_14261,N_14181,N_14225);
nand U14262 (N_14262,N_14201,N_14097);
and U14263 (N_14263,N_14160,N_14231);
nand U14264 (N_14264,N_14095,N_14236);
nand U14265 (N_14265,N_14121,N_14087);
and U14266 (N_14266,N_14101,N_14146);
and U14267 (N_14267,N_14155,N_14209);
and U14268 (N_14268,N_14195,N_14187);
xor U14269 (N_14269,N_14177,N_14105);
and U14270 (N_14270,N_14222,N_14164);
nand U14271 (N_14271,N_14113,N_14142);
nor U14272 (N_14272,N_14118,N_14194);
xor U14273 (N_14273,N_14130,N_14226);
nor U14274 (N_14274,N_14163,N_14223);
nor U14275 (N_14275,N_14117,N_14131);
or U14276 (N_14276,N_14185,N_14112);
nor U14277 (N_14277,N_14148,N_14137);
nor U14278 (N_14278,N_14135,N_14227);
nor U14279 (N_14279,N_14141,N_14179);
and U14280 (N_14280,N_14139,N_14103);
or U14281 (N_14281,N_14202,N_14150);
xnor U14282 (N_14282,N_14224,N_14213);
nand U14283 (N_14283,N_14143,N_14138);
or U14284 (N_14284,N_14196,N_14108);
xnor U14285 (N_14285,N_14230,N_14147);
nor U14286 (N_14286,N_14172,N_14081);
or U14287 (N_14287,N_14198,N_14096);
nor U14288 (N_14288,N_14158,N_14111);
or U14289 (N_14289,N_14218,N_14145);
nor U14290 (N_14290,N_14197,N_14127);
nor U14291 (N_14291,N_14219,N_14089);
and U14292 (N_14292,N_14221,N_14184);
or U14293 (N_14293,N_14144,N_14214);
nand U14294 (N_14294,N_14165,N_14207);
nor U14295 (N_14295,N_14159,N_14171);
or U14296 (N_14296,N_14192,N_14232);
and U14297 (N_14297,N_14205,N_14125);
nand U14298 (N_14298,N_14178,N_14156);
nor U14299 (N_14299,N_14215,N_14094);
and U14300 (N_14300,N_14123,N_14170);
and U14301 (N_14301,N_14092,N_14152);
nor U14302 (N_14302,N_14149,N_14106);
nand U14303 (N_14303,N_14220,N_14140);
or U14304 (N_14304,N_14175,N_14176);
or U14305 (N_14305,N_14134,N_14237);
and U14306 (N_14306,N_14174,N_14154);
xor U14307 (N_14307,N_14190,N_14169);
nor U14308 (N_14308,N_14238,N_14119);
and U14309 (N_14309,N_14167,N_14233);
or U14310 (N_14310,N_14173,N_14157);
or U14311 (N_14311,N_14082,N_14098);
nor U14312 (N_14312,N_14168,N_14203);
and U14313 (N_14313,N_14086,N_14239);
xnor U14314 (N_14314,N_14100,N_14153);
and U14315 (N_14315,N_14090,N_14085);
nor U14316 (N_14316,N_14182,N_14116);
and U14317 (N_14317,N_14199,N_14204);
and U14318 (N_14318,N_14126,N_14151);
nand U14319 (N_14319,N_14107,N_14162);
nand U14320 (N_14320,N_14228,N_14162);
nor U14321 (N_14321,N_14227,N_14158);
or U14322 (N_14322,N_14097,N_14220);
or U14323 (N_14323,N_14230,N_14084);
and U14324 (N_14324,N_14081,N_14190);
nor U14325 (N_14325,N_14119,N_14165);
or U14326 (N_14326,N_14223,N_14098);
or U14327 (N_14327,N_14216,N_14094);
nand U14328 (N_14328,N_14120,N_14132);
xnor U14329 (N_14329,N_14233,N_14200);
or U14330 (N_14330,N_14235,N_14196);
nor U14331 (N_14331,N_14092,N_14210);
and U14332 (N_14332,N_14127,N_14205);
or U14333 (N_14333,N_14217,N_14196);
and U14334 (N_14334,N_14232,N_14128);
nand U14335 (N_14335,N_14148,N_14133);
or U14336 (N_14336,N_14202,N_14089);
nand U14337 (N_14337,N_14138,N_14183);
nor U14338 (N_14338,N_14184,N_14113);
or U14339 (N_14339,N_14170,N_14190);
nand U14340 (N_14340,N_14117,N_14110);
xor U14341 (N_14341,N_14085,N_14111);
and U14342 (N_14342,N_14137,N_14083);
or U14343 (N_14343,N_14126,N_14160);
or U14344 (N_14344,N_14222,N_14167);
or U14345 (N_14345,N_14168,N_14109);
xnor U14346 (N_14346,N_14152,N_14086);
and U14347 (N_14347,N_14164,N_14205);
nand U14348 (N_14348,N_14213,N_14223);
nor U14349 (N_14349,N_14195,N_14204);
or U14350 (N_14350,N_14197,N_14114);
xor U14351 (N_14351,N_14221,N_14201);
and U14352 (N_14352,N_14219,N_14184);
and U14353 (N_14353,N_14230,N_14236);
and U14354 (N_14354,N_14205,N_14144);
and U14355 (N_14355,N_14221,N_14130);
nor U14356 (N_14356,N_14101,N_14091);
or U14357 (N_14357,N_14213,N_14116);
nand U14358 (N_14358,N_14233,N_14219);
nor U14359 (N_14359,N_14141,N_14231);
xor U14360 (N_14360,N_14104,N_14092);
nor U14361 (N_14361,N_14134,N_14110);
nand U14362 (N_14362,N_14148,N_14239);
nand U14363 (N_14363,N_14149,N_14221);
xor U14364 (N_14364,N_14113,N_14126);
nand U14365 (N_14365,N_14153,N_14182);
nand U14366 (N_14366,N_14081,N_14136);
nand U14367 (N_14367,N_14146,N_14214);
nand U14368 (N_14368,N_14180,N_14191);
nand U14369 (N_14369,N_14189,N_14204);
nand U14370 (N_14370,N_14094,N_14135);
and U14371 (N_14371,N_14234,N_14181);
and U14372 (N_14372,N_14165,N_14184);
and U14373 (N_14373,N_14238,N_14202);
nand U14374 (N_14374,N_14144,N_14218);
nor U14375 (N_14375,N_14147,N_14098);
nor U14376 (N_14376,N_14176,N_14089);
nand U14377 (N_14377,N_14093,N_14121);
and U14378 (N_14378,N_14129,N_14182);
or U14379 (N_14379,N_14153,N_14186);
xor U14380 (N_14380,N_14195,N_14160);
nor U14381 (N_14381,N_14235,N_14177);
nor U14382 (N_14382,N_14112,N_14211);
and U14383 (N_14383,N_14210,N_14098);
nor U14384 (N_14384,N_14161,N_14152);
or U14385 (N_14385,N_14089,N_14099);
and U14386 (N_14386,N_14197,N_14112);
and U14387 (N_14387,N_14182,N_14188);
and U14388 (N_14388,N_14225,N_14116);
nand U14389 (N_14389,N_14200,N_14236);
xor U14390 (N_14390,N_14117,N_14175);
nand U14391 (N_14391,N_14228,N_14130);
and U14392 (N_14392,N_14156,N_14098);
and U14393 (N_14393,N_14099,N_14086);
or U14394 (N_14394,N_14216,N_14206);
nor U14395 (N_14395,N_14125,N_14209);
and U14396 (N_14396,N_14122,N_14100);
nor U14397 (N_14397,N_14134,N_14188);
nor U14398 (N_14398,N_14174,N_14196);
or U14399 (N_14399,N_14174,N_14161);
and U14400 (N_14400,N_14288,N_14255);
nor U14401 (N_14401,N_14281,N_14343);
xnor U14402 (N_14402,N_14269,N_14349);
or U14403 (N_14403,N_14322,N_14378);
or U14404 (N_14404,N_14248,N_14310);
xnor U14405 (N_14405,N_14274,N_14266);
nor U14406 (N_14406,N_14348,N_14240);
or U14407 (N_14407,N_14361,N_14357);
nand U14408 (N_14408,N_14370,N_14331);
and U14409 (N_14409,N_14321,N_14333);
nand U14410 (N_14410,N_14366,N_14352);
nor U14411 (N_14411,N_14272,N_14347);
or U14412 (N_14412,N_14392,N_14271);
nor U14413 (N_14413,N_14390,N_14258);
nand U14414 (N_14414,N_14249,N_14290);
nand U14415 (N_14415,N_14386,N_14345);
nor U14416 (N_14416,N_14243,N_14393);
and U14417 (N_14417,N_14245,N_14324);
nand U14418 (N_14418,N_14277,N_14354);
nand U14419 (N_14419,N_14388,N_14346);
or U14420 (N_14420,N_14338,N_14325);
and U14421 (N_14421,N_14267,N_14292);
nor U14422 (N_14422,N_14261,N_14329);
or U14423 (N_14423,N_14336,N_14244);
and U14424 (N_14424,N_14306,N_14323);
and U14425 (N_14425,N_14313,N_14379);
nor U14426 (N_14426,N_14256,N_14394);
nand U14427 (N_14427,N_14314,N_14356);
xnor U14428 (N_14428,N_14257,N_14295);
nor U14429 (N_14429,N_14280,N_14254);
nor U14430 (N_14430,N_14263,N_14307);
or U14431 (N_14431,N_14376,N_14387);
xor U14432 (N_14432,N_14369,N_14320);
and U14433 (N_14433,N_14341,N_14300);
or U14434 (N_14434,N_14368,N_14304);
or U14435 (N_14435,N_14298,N_14260);
and U14436 (N_14436,N_14303,N_14279);
and U14437 (N_14437,N_14342,N_14296);
and U14438 (N_14438,N_14326,N_14318);
and U14439 (N_14439,N_14287,N_14293);
and U14440 (N_14440,N_14363,N_14332);
nand U14441 (N_14441,N_14252,N_14382);
or U14442 (N_14442,N_14283,N_14268);
nor U14443 (N_14443,N_14284,N_14377);
nand U14444 (N_14444,N_14355,N_14374);
nor U14445 (N_14445,N_14353,N_14397);
or U14446 (N_14446,N_14334,N_14286);
or U14447 (N_14447,N_14315,N_14251);
nand U14448 (N_14448,N_14285,N_14399);
and U14449 (N_14449,N_14259,N_14308);
or U14450 (N_14450,N_14351,N_14389);
and U14451 (N_14451,N_14241,N_14309);
or U14452 (N_14452,N_14301,N_14305);
or U14453 (N_14453,N_14311,N_14270);
nand U14454 (N_14454,N_14302,N_14330);
nand U14455 (N_14455,N_14364,N_14278);
or U14456 (N_14456,N_14319,N_14265);
nor U14457 (N_14457,N_14391,N_14340);
nor U14458 (N_14458,N_14297,N_14350);
and U14459 (N_14459,N_14246,N_14395);
and U14460 (N_14460,N_14328,N_14396);
and U14461 (N_14461,N_14381,N_14335);
or U14462 (N_14462,N_14299,N_14275);
xor U14463 (N_14463,N_14375,N_14282);
or U14464 (N_14464,N_14262,N_14373);
and U14465 (N_14465,N_14276,N_14383);
nor U14466 (N_14466,N_14253,N_14371);
nor U14467 (N_14467,N_14344,N_14264);
xnor U14468 (N_14468,N_14273,N_14362);
nor U14469 (N_14469,N_14337,N_14247);
and U14470 (N_14470,N_14385,N_14380);
nor U14471 (N_14471,N_14360,N_14372);
nor U14472 (N_14472,N_14398,N_14250);
nand U14473 (N_14473,N_14358,N_14289);
and U14474 (N_14474,N_14291,N_14359);
and U14475 (N_14475,N_14294,N_14367);
or U14476 (N_14476,N_14317,N_14316);
and U14477 (N_14477,N_14384,N_14365);
nand U14478 (N_14478,N_14312,N_14327);
nand U14479 (N_14479,N_14339,N_14242);
or U14480 (N_14480,N_14361,N_14349);
or U14481 (N_14481,N_14383,N_14344);
and U14482 (N_14482,N_14243,N_14312);
xnor U14483 (N_14483,N_14336,N_14391);
or U14484 (N_14484,N_14290,N_14314);
xnor U14485 (N_14485,N_14306,N_14396);
and U14486 (N_14486,N_14308,N_14375);
nand U14487 (N_14487,N_14381,N_14328);
and U14488 (N_14488,N_14348,N_14247);
and U14489 (N_14489,N_14328,N_14310);
nor U14490 (N_14490,N_14360,N_14314);
nand U14491 (N_14491,N_14261,N_14270);
nand U14492 (N_14492,N_14319,N_14363);
nor U14493 (N_14493,N_14255,N_14365);
and U14494 (N_14494,N_14292,N_14379);
or U14495 (N_14495,N_14287,N_14244);
nand U14496 (N_14496,N_14335,N_14333);
or U14497 (N_14497,N_14329,N_14370);
or U14498 (N_14498,N_14268,N_14394);
nor U14499 (N_14499,N_14265,N_14303);
xor U14500 (N_14500,N_14296,N_14331);
xor U14501 (N_14501,N_14346,N_14326);
and U14502 (N_14502,N_14317,N_14356);
or U14503 (N_14503,N_14382,N_14354);
xor U14504 (N_14504,N_14263,N_14372);
nor U14505 (N_14505,N_14326,N_14241);
nand U14506 (N_14506,N_14302,N_14345);
or U14507 (N_14507,N_14303,N_14393);
and U14508 (N_14508,N_14372,N_14306);
or U14509 (N_14509,N_14304,N_14339);
nor U14510 (N_14510,N_14285,N_14396);
or U14511 (N_14511,N_14294,N_14336);
nand U14512 (N_14512,N_14378,N_14269);
nor U14513 (N_14513,N_14273,N_14335);
or U14514 (N_14514,N_14376,N_14311);
nor U14515 (N_14515,N_14392,N_14373);
and U14516 (N_14516,N_14248,N_14343);
and U14517 (N_14517,N_14396,N_14304);
or U14518 (N_14518,N_14269,N_14331);
or U14519 (N_14519,N_14381,N_14259);
or U14520 (N_14520,N_14342,N_14373);
nand U14521 (N_14521,N_14383,N_14251);
nand U14522 (N_14522,N_14354,N_14289);
and U14523 (N_14523,N_14370,N_14245);
nand U14524 (N_14524,N_14372,N_14270);
or U14525 (N_14525,N_14358,N_14260);
and U14526 (N_14526,N_14248,N_14363);
nor U14527 (N_14527,N_14330,N_14326);
or U14528 (N_14528,N_14250,N_14260);
and U14529 (N_14529,N_14323,N_14273);
and U14530 (N_14530,N_14303,N_14390);
nor U14531 (N_14531,N_14361,N_14392);
nand U14532 (N_14532,N_14242,N_14283);
nand U14533 (N_14533,N_14354,N_14285);
and U14534 (N_14534,N_14390,N_14345);
or U14535 (N_14535,N_14378,N_14279);
and U14536 (N_14536,N_14339,N_14299);
and U14537 (N_14537,N_14371,N_14381);
xnor U14538 (N_14538,N_14356,N_14399);
and U14539 (N_14539,N_14387,N_14265);
and U14540 (N_14540,N_14337,N_14273);
nor U14541 (N_14541,N_14247,N_14289);
or U14542 (N_14542,N_14383,N_14380);
nor U14543 (N_14543,N_14281,N_14263);
nand U14544 (N_14544,N_14360,N_14384);
xnor U14545 (N_14545,N_14297,N_14275);
or U14546 (N_14546,N_14344,N_14319);
or U14547 (N_14547,N_14382,N_14284);
and U14548 (N_14548,N_14252,N_14399);
nor U14549 (N_14549,N_14393,N_14375);
nor U14550 (N_14550,N_14295,N_14266);
nor U14551 (N_14551,N_14370,N_14278);
nand U14552 (N_14552,N_14283,N_14293);
and U14553 (N_14553,N_14246,N_14381);
and U14554 (N_14554,N_14251,N_14356);
and U14555 (N_14555,N_14299,N_14365);
nor U14556 (N_14556,N_14273,N_14294);
nand U14557 (N_14557,N_14329,N_14349);
nor U14558 (N_14558,N_14299,N_14327);
or U14559 (N_14559,N_14274,N_14329);
nand U14560 (N_14560,N_14521,N_14460);
and U14561 (N_14561,N_14443,N_14523);
or U14562 (N_14562,N_14499,N_14458);
and U14563 (N_14563,N_14452,N_14545);
and U14564 (N_14564,N_14505,N_14532);
nor U14565 (N_14565,N_14535,N_14534);
xor U14566 (N_14566,N_14528,N_14542);
and U14567 (N_14567,N_14529,N_14412);
nand U14568 (N_14568,N_14502,N_14557);
or U14569 (N_14569,N_14513,N_14536);
or U14570 (N_14570,N_14453,N_14544);
or U14571 (N_14571,N_14509,N_14449);
nand U14572 (N_14572,N_14501,N_14402);
nor U14573 (N_14573,N_14457,N_14437);
and U14574 (N_14574,N_14445,N_14484);
nand U14575 (N_14575,N_14434,N_14508);
or U14576 (N_14576,N_14472,N_14483);
nand U14577 (N_14577,N_14500,N_14405);
and U14578 (N_14578,N_14419,N_14427);
nand U14579 (N_14579,N_14487,N_14423);
and U14580 (N_14580,N_14467,N_14474);
and U14581 (N_14581,N_14476,N_14498);
or U14582 (N_14582,N_14488,N_14516);
nor U14583 (N_14583,N_14441,N_14432);
nor U14584 (N_14584,N_14514,N_14520);
or U14585 (N_14585,N_14456,N_14485);
nor U14586 (N_14586,N_14494,N_14446);
or U14587 (N_14587,N_14539,N_14430);
and U14588 (N_14588,N_14531,N_14400);
and U14589 (N_14589,N_14482,N_14504);
nand U14590 (N_14590,N_14537,N_14438);
nor U14591 (N_14591,N_14550,N_14552);
xnor U14592 (N_14592,N_14489,N_14454);
or U14593 (N_14593,N_14543,N_14463);
or U14594 (N_14594,N_14462,N_14480);
nor U14595 (N_14595,N_14433,N_14422);
xor U14596 (N_14596,N_14473,N_14519);
or U14597 (N_14597,N_14426,N_14556);
nor U14598 (N_14598,N_14415,N_14541);
and U14599 (N_14599,N_14451,N_14470);
nand U14600 (N_14600,N_14479,N_14435);
and U14601 (N_14601,N_14421,N_14406);
nand U14602 (N_14602,N_14459,N_14478);
and U14603 (N_14603,N_14526,N_14404);
xor U14604 (N_14604,N_14510,N_14407);
nand U14605 (N_14605,N_14424,N_14503);
and U14606 (N_14606,N_14558,N_14481);
nor U14607 (N_14607,N_14471,N_14538);
and U14608 (N_14608,N_14429,N_14469);
and U14609 (N_14609,N_14492,N_14408);
nand U14610 (N_14610,N_14515,N_14448);
nor U14611 (N_14611,N_14468,N_14506);
and U14612 (N_14612,N_14547,N_14512);
xor U14613 (N_14613,N_14403,N_14530);
or U14614 (N_14614,N_14475,N_14546);
xnor U14615 (N_14615,N_14522,N_14559);
and U14616 (N_14616,N_14466,N_14409);
nand U14617 (N_14617,N_14401,N_14525);
nand U14618 (N_14618,N_14431,N_14518);
and U14619 (N_14619,N_14414,N_14551);
or U14620 (N_14620,N_14533,N_14436);
and U14621 (N_14621,N_14495,N_14548);
nand U14622 (N_14622,N_14486,N_14418);
nand U14623 (N_14623,N_14410,N_14553);
nand U14624 (N_14624,N_14540,N_14496);
and U14625 (N_14625,N_14493,N_14417);
xor U14626 (N_14626,N_14442,N_14461);
nand U14627 (N_14627,N_14511,N_14444);
nand U14628 (N_14628,N_14425,N_14450);
or U14629 (N_14629,N_14411,N_14555);
or U14630 (N_14630,N_14439,N_14420);
or U14631 (N_14631,N_14549,N_14464);
nor U14632 (N_14632,N_14527,N_14413);
nor U14633 (N_14633,N_14416,N_14517);
and U14634 (N_14634,N_14428,N_14524);
nand U14635 (N_14635,N_14447,N_14490);
or U14636 (N_14636,N_14507,N_14440);
nand U14637 (N_14637,N_14554,N_14455);
nor U14638 (N_14638,N_14477,N_14491);
and U14639 (N_14639,N_14465,N_14497);
nand U14640 (N_14640,N_14537,N_14501);
or U14641 (N_14641,N_14444,N_14401);
or U14642 (N_14642,N_14479,N_14472);
nand U14643 (N_14643,N_14485,N_14449);
or U14644 (N_14644,N_14401,N_14493);
and U14645 (N_14645,N_14429,N_14535);
nand U14646 (N_14646,N_14548,N_14529);
and U14647 (N_14647,N_14455,N_14419);
xor U14648 (N_14648,N_14534,N_14528);
and U14649 (N_14649,N_14435,N_14547);
nand U14650 (N_14650,N_14415,N_14467);
nand U14651 (N_14651,N_14430,N_14449);
or U14652 (N_14652,N_14557,N_14436);
and U14653 (N_14653,N_14492,N_14450);
nand U14654 (N_14654,N_14405,N_14525);
and U14655 (N_14655,N_14429,N_14533);
nor U14656 (N_14656,N_14408,N_14406);
or U14657 (N_14657,N_14494,N_14506);
and U14658 (N_14658,N_14402,N_14484);
or U14659 (N_14659,N_14492,N_14521);
or U14660 (N_14660,N_14416,N_14549);
nand U14661 (N_14661,N_14447,N_14541);
nor U14662 (N_14662,N_14524,N_14544);
nor U14663 (N_14663,N_14415,N_14443);
nand U14664 (N_14664,N_14514,N_14551);
nor U14665 (N_14665,N_14532,N_14512);
and U14666 (N_14666,N_14488,N_14509);
or U14667 (N_14667,N_14438,N_14476);
nor U14668 (N_14668,N_14432,N_14507);
or U14669 (N_14669,N_14471,N_14422);
nor U14670 (N_14670,N_14415,N_14421);
nor U14671 (N_14671,N_14425,N_14502);
and U14672 (N_14672,N_14518,N_14528);
or U14673 (N_14673,N_14506,N_14493);
and U14674 (N_14674,N_14508,N_14458);
nor U14675 (N_14675,N_14519,N_14466);
nor U14676 (N_14676,N_14467,N_14456);
nand U14677 (N_14677,N_14479,N_14436);
nor U14678 (N_14678,N_14512,N_14440);
or U14679 (N_14679,N_14557,N_14524);
nor U14680 (N_14680,N_14521,N_14430);
and U14681 (N_14681,N_14446,N_14465);
nand U14682 (N_14682,N_14486,N_14419);
and U14683 (N_14683,N_14441,N_14470);
nand U14684 (N_14684,N_14504,N_14471);
nor U14685 (N_14685,N_14545,N_14411);
and U14686 (N_14686,N_14517,N_14508);
or U14687 (N_14687,N_14515,N_14419);
or U14688 (N_14688,N_14521,N_14507);
and U14689 (N_14689,N_14419,N_14489);
or U14690 (N_14690,N_14410,N_14445);
or U14691 (N_14691,N_14459,N_14450);
or U14692 (N_14692,N_14406,N_14542);
nand U14693 (N_14693,N_14520,N_14543);
or U14694 (N_14694,N_14428,N_14439);
or U14695 (N_14695,N_14497,N_14425);
and U14696 (N_14696,N_14542,N_14400);
nor U14697 (N_14697,N_14484,N_14490);
nor U14698 (N_14698,N_14462,N_14509);
nand U14699 (N_14699,N_14411,N_14488);
nand U14700 (N_14700,N_14500,N_14481);
or U14701 (N_14701,N_14434,N_14406);
nor U14702 (N_14702,N_14495,N_14407);
nor U14703 (N_14703,N_14448,N_14442);
nand U14704 (N_14704,N_14554,N_14404);
or U14705 (N_14705,N_14488,N_14416);
or U14706 (N_14706,N_14453,N_14508);
and U14707 (N_14707,N_14537,N_14538);
or U14708 (N_14708,N_14538,N_14452);
or U14709 (N_14709,N_14545,N_14546);
nor U14710 (N_14710,N_14440,N_14461);
nand U14711 (N_14711,N_14408,N_14491);
and U14712 (N_14712,N_14445,N_14466);
nand U14713 (N_14713,N_14418,N_14458);
nand U14714 (N_14714,N_14461,N_14528);
or U14715 (N_14715,N_14480,N_14402);
and U14716 (N_14716,N_14530,N_14486);
nor U14717 (N_14717,N_14491,N_14466);
and U14718 (N_14718,N_14443,N_14496);
nor U14719 (N_14719,N_14406,N_14471);
or U14720 (N_14720,N_14643,N_14605);
nand U14721 (N_14721,N_14612,N_14593);
and U14722 (N_14722,N_14604,N_14599);
or U14723 (N_14723,N_14716,N_14675);
nor U14724 (N_14724,N_14568,N_14573);
and U14725 (N_14725,N_14715,N_14674);
and U14726 (N_14726,N_14641,N_14653);
xor U14727 (N_14727,N_14694,N_14669);
and U14728 (N_14728,N_14637,N_14642);
or U14729 (N_14729,N_14592,N_14651);
and U14730 (N_14730,N_14560,N_14665);
and U14731 (N_14731,N_14691,N_14611);
or U14732 (N_14732,N_14705,N_14634);
and U14733 (N_14733,N_14577,N_14613);
xnor U14734 (N_14734,N_14630,N_14590);
or U14735 (N_14735,N_14704,N_14627);
nand U14736 (N_14736,N_14618,N_14662);
or U14737 (N_14737,N_14644,N_14718);
nand U14738 (N_14738,N_14672,N_14615);
or U14739 (N_14739,N_14636,N_14580);
and U14740 (N_14740,N_14701,N_14633);
nand U14741 (N_14741,N_14579,N_14688);
nand U14742 (N_14742,N_14714,N_14671);
nand U14743 (N_14743,N_14683,N_14578);
nand U14744 (N_14744,N_14706,N_14631);
and U14745 (N_14745,N_14622,N_14713);
or U14746 (N_14746,N_14689,N_14658);
nand U14747 (N_14747,N_14610,N_14598);
and U14748 (N_14748,N_14565,N_14571);
and U14749 (N_14749,N_14673,N_14616);
nor U14750 (N_14750,N_14574,N_14586);
and U14751 (N_14751,N_14697,N_14623);
or U14752 (N_14752,N_14566,N_14679);
and U14753 (N_14753,N_14703,N_14680);
nor U14754 (N_14754,N_14695,N_14717);
or U14755 (N_14755,N_14626,N_14561);
and U14756 (N_14756,N_14617,N_14588);
and U14757 (N_14757,N_14666,N_14692);
nor U14758 (N_14758,N_14620,N_14681);
and U14759 (N_14759,N_14629,N_14583);
nor U14760 (N_14760,N_14656,N_14660);
nand U14761 (N_14761,N_14589,N_14597);
and U14762 (N_14762,N_14664,N_14621);
nor U14763 (N_14763,N_14647,N_14602);
and U14764 (N_14764,N_14670,N_14607);
xor U14765 (N_14765,N_14606,N_14575);
nor U14766 (N_14766,N_14668,N_14709);
nor U14767 (N_14767,N_14564,N_14603);
and U14768 (N_14768,N_14649,N_14609);
or U14769 (N_14769,N_14572,N_14682);
or U14770 (N_14770,N_14663,N_14594);
and U14771 (N_14771,N_14570,N_14652);
or U14772 (N_14772,N_14567,N_14576);
or U14773 (N_14773,N_14707,N_14700);
or U14774 (N_14774,N_14678,N_14661);
nor U14775 (N_14775,N_14614,N_14711);
and U14776 (N_14776,N_14632,N_14650);
nor U14777 (N_14777,N_14685,N_14708);
and U14778 (N_14778,N_14693,N_14712);
nand U14779 (N_14779,N_14676,N_14646);
xnor U14780 (N_14780,N_14625,N_14667);
nand U14781 (N_14781,N_14619,N_14659);
xnor U14782 (N_14782,N_14563,N_14690);
or U14783 (N_14783,N_14645,N_14624);
and U14784 (N_14784,N_14595,N_14696);
nand U14785 (N_14785,N_14596,N_14687);
xnor U14786 (N_14786,N_14686,N_14698);
and U14787 (N_14787,N_14585,N_14677);
or U14788 (N_14788,N_14638,N_14581);
and U14789 (N_14789,N_14719,N_14657);
nand U14790 (N_14790,N_14639,N_14702);
nand U14791 (N_14791,N_14640,N_14654);
and U14792 (N_14792,N_14601,N_14655);
nor U14793 (N_14793,N_14587,N_14608);
nand U14794 (N_14794,N_14569,N_14684);
or U14795 (N_14795,N_14699,N_14710);
nor U14796 (N_14796,N_14584,N_14635);
nor U14797 (N_14797,N_14591,N_14600);
and U14798 (N_14798,N_14628,N_14562);
nor U14799 (N_14799,N_14648,N_14582);
or U14800 (N_14800,N_14708,N_14700);
or U14801 (N_14801,N_14579,N_14641);
or U14802 (N_14802,N_14585,N_14709);
nor U14803 (N_14803,N_14709,N_14567);
and U14804 (N_14804,N_14617,N_14655);
and U14805 (N_14805,N_14595,N_14705);
nand U14806 (N_14806,N_14659,N_14575);
or U14807 (N_14807,N_14655,N_14660);
or U14808 (N_14808,N_14622,N_14647);
or U14809 (N_14809,N_14676,N_14711);
nand U14810 (N_14810,N_14690,N_14638);
nor U14811 (N_14811,N_14592,N_14695);
nand U14812 (N_14812,N_14632,N_14718);
nor U14813 (N_14813,N_14588,N_14614);
nor U14814 (N_14814,N_14572,N_14625);
nor U14815 (N_14815,N_14596,N_14656);
and U14816 (N_14816,N_14599,N_14696);
and U14817 (N_14817,N_14622,N_14641);
and U14818 (N_14818,N_14580,N_14592);
and U14819 (N_14819,N_14696,N_14606);
nor U14820 (N_14820,N_14709,N_14660);
nand U14821 (N_14821,N_14590,N_14699);
nor U14822 (N_14822,N_14620,N_14580);
xnor U14823 (N_14823,N_14697,N_14663);
and U14824 (N_14824,N_14626,N_14678);
nand U14825 (N_14825,N_14595,N_14564);
and U14826 (N_14826,N_14623,N_14667);
nand U14827 (N_14827,N_14566,N_14578);
and U14828 (N_14828,N_14629,N_14571);
nand U14829 (N_14829,N_14701,N_14719);
and U14830 (N_14830,N_14666,N_14605);
or U14831 (N_14831,N_14714,N_14712);
nand U14832 (N_14832,N_14673,N_14605);
xnor U14833 (N_14833,N_14629,N_14606);
or U14834 (N_14834,N_14618,N_14598);
or U14835 (N_14835,N_14635,N_14670);
or U14836 (N_14836,N_14641,N_14639);
and U14837 (N_14837,N_14708,N_14631);
nor U14838 (N_14838,N_14604,N_14657);
or U14839 (N_14839,N_14653,N_14583);
nor U14840 (N_14840,N_14611,N_14655);
xor U14841 (N_14841,N_14578,N_14606);
xor U14842 (N_14842,N_14686,N_14653);
or U14843 (N_14843,N_14588,N_14714);
and U14844 (N_14844,N_14659,N_14579);
and U14845 (N_14845,N_14619,N_14585);
or U14846 (N_14846,N_14670,N_14611);
nor U14847 (N_14847,N_14639,N_14671);
nand U14848 (N_14848,N_14625,N_14613);
nand U14849 (N_14849,N_14659,N_14635);
or U14850 (N_14850,N_14703,N_14607);
and U14851 (N_14851,N_14614,N_14594);
and U14852 (N_14852,N_14687,N_14671);
or U14853 (N_14853,N_14704,N_14679);
or U14854 (N_14854,N_14660,N_14614);
nor U14855 (N_14855,N_14607,N_14652);
nor U14856 (N_14856,N_14617,N_14717);
nand U14857 (N_14857,N_14605,N_14658);
or U14858 (N_14858,N_14589,N_14669);
nand U14859 (N_14859,N_14640,N_14580);
nor U14860 (N_14860,N_14670,N_14655);
nand U14861 (N_14861,N_14612,N_14706);
or U14862 (N_14862,N_14683,N_14700);
xnor U14863 (N_14863,N_14635,N_14574);
nand U14864 (N_14864,N_14672,N_14574);
nand U14865 (N_14865,N_14671,N_14708);
and U14866 (N_14866,N_14687,N_14633);
xor U14867 (N_14867,N_14618,N_14565);
or U14868 (N_14868,N_14662,N_14569);
or U14869 (N_14869,N_14638,N_14575);
nor U14870 (N_14870,N_14662,N_14690);
and U14871 (N_14871,N_14671,N_14665);
nand U14872 (N_14872,N_14644,N_14575);
nand U14873 (N_14873,N_14603,N_14677);
nor U14874 (N_14874,N_14693,N_14704);
and U14875 (N_14875,N_14673,N_14628);
or U14876 (N_14876,N_14716,N_14605);
xor U14877 (N_14877,N_14705,N_14652);
nand U14878 (N_14878,N_14594,N_14622);
nand U14879 (N_14879,N_14662,N_14597);
and U14880 (N_14880,N_14783,N_14798);
xnor U14881 (N_14881,N_14831,N_14846);
nor U14882 (N_14882,N_14727,N_14812);
nor U14883 (N_14883,N_14757,N_14816);
or U14884 (N_14884,N_14860,N_14748);
xnor U14885 (N_14885,N_14852,N_14740);
nor U14886 (N_14886,N_14723,N_14797);
and U14887 (N_14887,N_14870,N_14743);
nor U14888 (N_14888,N_14747,N_14828);
nand U14889 (N_14889,N_14874,N_14806);
and U14890 (N_14890,N_14833,N_14842);
nand U14891 (N_14891,N_14856,N_14792);
and U14892 (N_14892,N_14779,N_14753);
or U14893 (N_14893,N_14760,N_14859);
xnor U14894 (N_14894,N_14867,N_14830);
nand U14895 (N_14895,N_14780,N_14786);
nor U14896 (N_14896,N_14729,N_14868);
or U14897 (N_14897,N_14844,N_14721);
nor U14898 (N_14898,N_14835,N_14843);
nor U14899 (N_14899,N_14756,N_14829);
nor U14900 (N_14900,N_14725,N_14858);
nand U14901 (N_14901,N_14773,N_14742);
nand U14902 (N_14902,N_14788,N_14827);
xor U14903 (N_14903,N_14872,N_14839);
nand U14904 (N_14904,N_14876,N_14750);
nor U14905 (N_14905,N_14738,N_14803);
nand U14906 (N_14906,N_14777,N_14814);
and U14907 (N_14907,N_14820,N_14764);
and U14908 (N_14908,N_14815,N_14735);
and U14909 (N_14909,N_14782,N_14720);
nor U14910 (N_14910,N_14857,N_14771);
and U14911 (N_14911,N_14873,N_14763);
nor U14912 (N_14912,N_14849,N_14799);
xnor U14913 (N_14913,N_14871,N_14751);
and U14914 (N_14914,N_14734,N_14730);
and U14915 (N_14915,N_14801,N_14838);
nor U14916 (N_14916,N_14732,N_14879);
and U14917 (N_14917,N_14746,N_14855);
nand U14918 (N_14918,N_14778,N_14877);
nand U14919 (N_14919,N_14791,N_14767);
nor U14920 (N_14920,N_14776,N_14808);
and U14921 (N_14921,N_14749,N_14759);
or U14922 (N_14922,N_14768,N_14845);
or U14923 (N_14923,N_14739,N_14802);
nand U14924 (N_14924,N_14818,N_14728);
nand U14925 (N_14925,N_14863,N_14869);
and U14926 (N_14926,N_14726,N_14854);
nor U14927 (N_14927,N_14832,N_14787);
nor U14928 (N_14928,N_14847,N_14841);
and U14929 (N_14929,N_14737,N_14761);
nand U14930 (N_14930,N_14813,N_14796);
and U14931 (N_14931,N_14795,N_14772);
nor U14932 (N_14932,N_14781,N_14823);
and U14933 (N_14933,N_14800,N_14836);
nand U14934 (N_14934,N_14853,N_14811);
and U14935 (N_14935,N_14875,N_14789);
and U14936 (N_14936,N_14784,N_14826);
or U14937 (N_14937,N_14804,N_14821);
nand U14938 (N_14938,N_14790,N_14724);
or U14939 (N_14939,N_14822,N_14765);
nand U14940 (N_14940,N_14834,N_14805);
xor U14941 (N_14941,N_14766,N_14736);
or U14942 (N_14942,N_14762,N_14851);
nand U14943 (N_14943,N_14819,N_14840);
nand U14944 (N_14944,N_14770,N_14848);
and U14945 (N_14945,N_14774,N_14878);
nand U14946 (N_14946,N_14862,N_14810);
or U14947 (N_14947,N_14745,N_14741);
or U14948 (N_14948,N_14755,N_14793);
nor U14949 (N_14949,N_14837,N_14733);
nand U14950 (N_14950,N_14817,N_14850);
and U14951 (N_14951,N_14825,N_14866);
xnor U14952 (N_14952,N_14785,N_14731);
xnor U14953 (N_14953,N_14754,N_14861);
or U14954 (N_14954,N_14824,N_14794);
xor U14955 (N_14955,N_14744,N_14809);
nor U14956 (N_14956,N_14775,N_14722);
and U14957 (N_14957,N_14758,N_14864);
nor U14958 (N_14958,N_14769,N_14752);
nor U14959 (N_14959,N_14807,N_14865);
nor U14960 (N_14960,N_14724,N_14812);
nor U14961 (N_14961,N_14874,N_14795);
nor U14962 (N_14962,N_14781,N_14806);
and U14963 (N_14963,N_14833,N_14788);
xor U14964 (N_14964,N_14749,N_14724);
or U14965 (N_14965,N_14857,N_14875);
and U14966 (N_14966,N_14872,N_14758);
and U14967 (N_14967,N_14805,N_14796);
nor U14968 (N_14968,N_14842,N_14772);
nand U14969 (N_14969,N_14802,N_14805);
and U14970 (N_14970,N_14730,N_14807);
and U14971 (N_14971,N_14805,N_14824);
nand U14972 (N_14972,N_14781,N_14770);
nor U14973 (N_14973,N_14843,N_14792);
nor U14974 (N_14974,N_14819,N_14795);
and U14975 (N_14975,N_14791,N_14806);
nor U14976 (N_14976,N_14807,N_14863);
and U14977 (N_14977,N_14845,N_14757);
nor U14978 (N_14978,N_14724,N_14727);
or U14979 (N_14979,N_14743,N_14777);
nor U14980 (N_14980,N_14792,N_14777);
or U14981 (N_14981,N_14770,N_14788);
nand U14982 (N_14982,N_14798,N_14732);
and U14983 (N_14983,N_14771,N_14784);
nand U14984 (N_14984,N_14764,N_14731);
nand U14985 (N_14985,N_14788,N_14723);
xor U14986 (N_14986,N_14852,N_14810);
nor U14987 (N_14987,N_14839,N_14821);
nand U14988 (N_14988,N_14813,N_14762);
nand U14989 (N_14989,N_14748,N_14773);
or U14990 (N_14990,N_14870,N_14876);
nor U14991 (N_14991,N_14833,N_14729);
and U14992 (N_14992,N_14723,N_14757);
and U14993 (N_14993,N_14822,N_14825);
nor U14994 (N_14994,N_14836,N_14792);
nand U14995 (N_14995,N_14761,N_14768);
nand U14996 (N_14996,N_14792,N_14796);
nand U14997 (N_14997,N_14769,N_14726);
or U14998 (N_14998,N_14743,N_14742);
or U14999 (N_14999,N_14783,N_14849);
and U15000 (N_15000,N_14825,N_14878);
nor U15001 (N_15001,N_14763,N_14784);
or U15002 (N_15002,N_14742,N_14828);
xor U15003 (N_15003,N_14848,N_14856);
nor U15004 (N_15004,N_14814,N_14870);
nor U15005 (N_15005,N_14829,N_14750);
nor U15006 (N_15006,N_14732,N_14834);
xnor U15007 (N_15007,N_14836,N_14758);
and U15008 (N_15008,N_14755,N_14817);
nor U15009 (N_15009,N_14849,N_14755);
and U15010 (N_15010,N_14851,N_14799);
nor U15011 (N_15011,N_14856,N_14832);
or U15012 (N_15012,N_14861,N_14732);
xor U15013 (N_15013,N_14790,N_14862);
nor U15014 (N_15014,N_14773,N_14765);
nand U15015 (N_15015,N_14836,N_14817);
nor U15016 (N_15016,N_14861,N_14866);
nor U15017 (N_15017,N_14774,N_14830);
nand U15018 (N_15018,N_14790,N_14750);
and U15019 (N_15019,N_14819,N_14810);
nand U15020 (N_15020,N_14747,N_14726);
nor U15021 (N_15021,N_14778,N_14745);
nor U15022 (N_15022,N_14744,N_14724);
nor U15023 (N_15023,N_14777,N_14854);
nor U15024 (N_15024,N_14750,N_14837);
or U15025 (N_15025,N_14777,N_14839);
nor U15026 (N_15026,N_14721,N_14789);
xnor U15027 (N_15027,N_14789,N_14742);
or U15028 (N_15028,N_14775,N_14721);
nor U15029 (N_15029,N_14776,N_14826);
xnor U15030 (N_15030,N_14741,N_14772);
and U15031 (N_15031,N_14785,N_14752);
xnor U15032 (N_15032,N_14858,N_14748);
or U15033 (N_15033,N_14831,N_14814);
nor U15034 (N_15034,N_14735,N_14813);
nor U15035 (N_15035,N_14780,N_14865);
or U15036 (N_15036,N_14733,N_14824);
or U15037 (N_15037,N_14831,N_14819);
and U15038 (N_15038,N_14850,N_14779);
nor U15039 (N_15039,N_14837,N_14785);
xor U15040 (N_15040,N_14976,N_14972);
and U15041 (N_15041,N_14945,N_14881);
or U15042 (N_15042,N_14990,N_15012);
nand U15043 (N_15043,N_15015,N_14906);
xnor U15044 (N_15044,N_14911,N_14934);
nand U15045 (N_15045,N_14890,N_14901);
nor U15046 (N_15046,N_14917,N_14919);
and U15047 (N_15047,N_14998,N_14929);
and U15048 (N_15048,N_14896,N_14984);
nand U15049 (N_15049,N_15008,N_14883);
xor U15050 (N_15050,N_14925,N_14921);
nand U15051 (N_15051,N_15025,N_15013);
or U15052 (N_15052,N_14918,N_14992);
and U15053 (N_15053,N_14980,N_14951);
nand U15054 (N_15054,N_15034,N_14915);
nor U15055 (N_15055,N_15022,N_14965);
nor U15056 (N_15056,N_14958,N_14986);
nand U15057 (N_15057,N_14898,N_14916);
or U15058 (N_15058,N_14999,N_15016);
nor U15059 (N_15059,N_14904,N_14982);
nor U15060 (N_15060,N_15023,N_14910);
or U15061 (N_15061,N_14959,N_15027);
nor U15062 (N_15062,N_14997,N_14897);
nand U15063 (N_15063,N_15039,N_14985);
nor U15064 (N_15064,N_14969,N_14987);
or U15065 (N_15065,N_14935,N_15010);
nand U15066 (N_15066,N_14975,N_15038);
and U15067 (N_15067,N_14961,N_14970);
or U15068 (N_15068,N_14948,N_14944);
nand U15069 (N_15069,N_14887,N_14939);
and U15070 (N_15070,N_15019,N_15018);
and U15071 (N_15071,N_15029,N_14950);
nand U15072 (N_15072,N_14991,N_14905);
xor U15073 (N_15073,N_14930,N_15000);
or U15074 (N_15074,N_15017,N_14893);
nor U15075 (N_15075,N_14967,N_14962);
and U15076 (N_15076,N_14912,N_14947);
nor U15077 (N_15077,N_14920,N_14968);
or U15078 (N_15078,N_14889,N_14954);
or U15079 (N_15079,N_14971,N_14914);
and U15080 (N_15080,N_14931,N_14907);
and U15081 (N_15081,N_14891,N_14978);
nor U15082 (N_15082,N_14994,N_14946);
and U15083 (N_15083,N_14894,N_15028);
nor U15084 (N_15084,N_14952,N_14928);
nand U15085 (N_15085,N_14923,N_14996);
or U15086 (N_15086,N_15036,N_14979);
or U15087 (N_15087,N_14993,N_15031);
or U15088 (N_15088,N_15021,N_14989);
nand U15089 (N_15089,N_14988,N_14909);
nand U15090 (N_15090,N_14942,N_14956);
nand U15091 (N_15091,N_14977,N_14941);
nor U15092 (N_15092,N_15003,N_14936);
or U15093 (N_15093,N_14922,N_15009);
nor U15094 (N_15094,N_15006,N_14964);
or U15095 (N_15095,N_14913,N_14940);
and U15096 (N_15096,N_15001,N_14886);
and U15097 (N_15097,N_15007,N_14949);
and U15098 (N_15098,N_15035,N_14927);
nor U15099 (N_15099,N_14995,N_15011);
and U15100 (N_15100,N_14938,N_14908);
nand U15101 (N_15101,N_14888,N_15014);
nand U15102 (N_15102,N_14884,N_15004);
and U15103 (N_15103,N_14963,N_15024);
or U15104 (N_15104,N_14882,N_14902);
xor U15105 (N_15105,N_14957,N_14899);
or U15106 (N_15106,N_14953,N_14937);
or U15107 (N_15107,N_14892,N_14983);
or U15108 (N_15108,N_14900,N_14880);
xor U15109 (N_15109,N_14885,N_14960);
xor U15110 (N_15110,N_14966,N_14924);
or U15111 (N_15111,N_14974,N_14973);
xnor U15112 (N_15112,N_14895,N_14981);
nand U15113 (N_15113,N_14933,N_15026);
xnor U15114 (N_15114,N_15033,N_15005);
nor U15115 (N_15115,N_15002,N_14903);
nor U15116 (N_15116,N_15020,N_14926);
nand U15117 (N_15117,N_14955,N_15032);
or U15118 (N_15118,N_14943,N_15030);
nor U15119 (N_15119,N_14932,N_15037);
or U15120 (N_15120,N_14982,N_14941);
nor U15121 (N_15121,N_14899,N_14985);
nand U15122 (N_15122,N_14937,N_14940);
nor U15123 (N_15123,N_14981,N_14925);
nand U15124 (N_15124,N_15016,N_14920);
nand U15125 (N_15125,N_14905,N_14889);
nand U15126 (N_15126,N_15021,N_14894);
nand U15127 (N_15127,N_14923,N_14917);
or U15128 (N_15128,N_15034,N_14888);
and U15129 (N_15129,N_14986,N_14991);
xnor U15130 (N_15130,N_14888,N_14921);
nand U15131 (N_15131,N_14942,N_14989);
and U15132 (N_15132,N_14989,N_15018);
xnor U15133 (N_15133,N_15031,N_14880);
nand U15134 (N_15134,N_14992,N_15038);
or U15135 (N_15135,N_14919,N_14988);
nor U15136 (N_15136,N_14969,N_14947);
and U15137 (N_15137,N_14890,N_14957);
and U15138 (N_15138,N_14973,N_14951);
nand U15139 (N_15139,N_15021,N_15018);
xor U15140 (N_15140,N_14941,N_14901);
nand U15141 (N_15141,N_14977,N_14954);
nand U15142 (N_15142,N_14894,N_14932);
nor U15143 (N_15143,N_14924,N_14897);
nor U15144 (N_15144,N_14951,N_14917);
nor U15145 (N_15145,N_15013,N_14961);
xnor U15146 (N_15146,N_14997,N_14928);
nand U15147 (N_15147,N_14946,N_15018);
nand U15148 (N_15148,N_14936,N_14924);
nand U15149 (N_15149,N_14893,N_14948);
and U15150 (N_15150,N_14884,N_15012);
and U15151 (N_15151,N_14945,N_14978);
or U15152 (N_15152,N_14911,N_14981);
xor U15153 (N_15153,N_14968,N_14888);
nor U15154 (N_15154,N_14937,N_14954);
or U15155 (N_15155,N_15030,N_15039);
nor U15156 (N_15156,N_14925,N_15027);
and U15157 (N_15157,N_14972,N_14981);
nand U15158 (N_15158,N_14974,N_14936);
and U15159 (N_15159,N_14941,N_14935);
and U15160 (N_15160,N_14894,N_14897);
nor U15161 (N_15161,N_14963,N_15028);
or U15162 (N_15162,N_14987,N_14935);
or U15163 (N_15163,N_14932,N_14984);
and U15164 (N_15164,N_15016,N_14980);
and U15165 (N_15165,N_14896,N_14951);
and U15166 (N_15166,N_14987,N_14887);
nor U15167 (N_15167,N_14904,N_14935);
and U15168 (N_15168,N_15002,N_14949);
nand U15169 (N_15169,N_14923,N_14970);
and U15170 (N_15170,N_14890,N_15006);
or U15171 (N_15171,N_14945,N_14916);
nand U15172 (N_15172,N_14954,N_15038);
nand U15173 (N_15173,N_14978,N_15034);
or U15174 (N_15174,N_15035,N_15029);
or U15175 (N_15175,N_14891,N_14968);
and U15176 (N_15176,N_15001,N_14933);
nand U15177 (N_15177,N_15008,N_15027);
nand U15178 (N_15178,N_14906,N_15014);
nor U15179 (N_15179,N_15030,N_14918);
xnor U15180 (N_15180,N_14964,N_14954);
and U15181 (N_15181,N_14978,N_14972);
nor U15182 (N_15182,N_14979,N_14988);
xor U15183 (N_15183,N_15021,N_14991);
xor U15184 (N_15184,N_15006,N_14950);
or U15185 (N_15185,N_14986,N_14982);
and U15186 (N_15186,N_14965,N_14911);
and U15187 (N_15187,N_14891,N_14952);
and U15188 (N_15188,N_14965,N_15031);
xnor U15189 (N_15189,N_14914,N_14987);
and U15190 (N_15190,N_14893,N_15023);
xnor U15191 (N_15191,N_14923,N_14989);
or U15192 (N_15192,N_14977,N_14945);
nor U15193 (N_15193,N_15036,N_14930);
nor U15194 (N_15194,N_14944,N_15016);
xor U15195 (N_15195,N_14973,N_14910);
nand U15196 (N_15196,N_14890,N_15033);
and U15197 (N_15197,N_14956,N_15000);
and U15198 (N_15198,N_14886,N_15034);
nor U15199 (N_15199,N_15025,N_14907);
xnor U15200 (N_15200,N_15139,N_15122);
xor U15201 (N_15201,N_15047,N_15156);
and U15202 (N_15202,N_15130,N_15099);
nand U15203 (N_15203,N_15044,N_15090);
nand U15204 (N_15204,N_15068,N_15094);
nor U15205 (N_15205,N_15129,N_15097);
nor U15206 (N_15206,N_15197,N_15081);
nand U15207 (N_15207,N_15144,N_15134);
nor U15208 (N_15208,N_15184,N_15092);
nand U15209 (N_15209,N_15112,N_15138);
and U15210 (N_15210,N_15157,N_15182);
or U15211 (N_15211,N_15113,N_15128);
nand U15212 (N_15212,N_15075,N_15196);
nor U15213 (N_15213,N_15066,N_15072);
nand U15214 (N_15214,N_15082,N_15093);
nor U15215 (N_15215,N_15199,N_15193);
nor U15216 (N_15216,N_15104,N_15187);
nor U15217 (N_15217,N_15162,N_15150);
nor U15218 (N_15218,N_15158,N_15140);
and U15219 (N_15219,N_15103,N_15143);
xnor U15220 (N_15220,N_15149,N_15136);
or U15221 (N_15221,N_15119,N_15083);
nand U15222 (N_15222,N_15185,N_15159);
and U15223 (N_15223,N_15189,N_15131);
nand U15224 (N_15224,N_15051,N_15137);
and U15225 (N_15225,N_15107,N_15116);
nand U15226 (N_15226,N_15102,N_15152);
and U15227 (N_15227,N_15043,N_15135);
and U15228 (N_15228,N_15069,N_15127);
or U15229 (N_15229,N_15078,N_15076);
nor U15230 (N_15230,N_15123,N_15089);
or U15231 (N_15231,N_15080,N_15077);
xor U15232 (N_15232,N_15153,N_15086);
nand U15233 (N_15233,N_15154,N_15190);
nor U15234 (N_15234,N_15163,N_15067);
nand U15235 (N_15235,N_15121,N_15105);
nand U15236 (N_15236,N_15141,N_15058);
and U15237 (N_15237,N_15192,N_15062);
nand U15238 (N_15238,N_15073,N_15178);
or U15239 (N_15239,N_15191,N_15049);
xnor U15240 (N_15240,N_15045,N_15194);
and U15241 (N_15241,N_15133,N_15084);
or U15242 (N_15242,N_15164,N_15079);
nand U15243 (N_15243,N_15120,N_15064);
nor U15244 (N_15244,N_15155,N_15052);
and U15245 (N_15245,N_15071,N_15057);
nor U15246 (N_15246,N_15175,N_15186);
nand U15247 (N_15247,N_15173,N_15087);
nand U15248 (N_15248,N_15168,N_15088);
nor U15249 (N_15249,N_15108,N_15048);
xnor U15250 (N_15250,N_15110,N_15124);
and U15251 (N_15251,N_15091,N_15111);
nand U15252 (N_15252,N_15165,N_15096);
and U15253 (N_15253,N_15160,N_15147);
xor U15254 (N_15254,N_15170,N_15085);
nand U15255 (N_15255,N_15172,N_15059);
nand U15256 (N_15256,N_15101,N_15054);
and U15257 (N_15257,N_15106,N_15181);
nor U15258 (N_15258,N_15041,N_15148);
xnor U15259 (N_15259,N_15118,N_15174);
nand U15260 (N_15260,N_15179,N_15056);
nor U15261 (N_15261,N_15053,N_15183);
or U15262 (N_15262,N_15063,N_15171);
or U15263 (N_15263,N_15142,N_15161);
nor U15264 (N_15264,N_15109,N_15095);
or U15265 (N_15265,N_15055,N_15166);
nor U15266 (N_15266,N_15040,N_15126);
nand U15267 (N_15267,N_15060,N_15098);
nor U15268 (N_15268,N_15167,N_15100);
nand U15269 (N_15269,N_15198,N_15132);
or U15270 (N_15270,N_15188,N_15046);
or U15271 (N_15271,N_15176,N_15145);
nand U15272 (N_15272,N_15065,N_15195);
or U15273 (N_15273,N_15070,N_15115);
and U15274 (N_15274,N_15177,N_15125);
or U15275 (N_15275,N_15074,N_15114);
or U15276 (N_15276,N_15180,N_15061);
or U15277 (N_15277,N_15151,N_15146);
and U15278 (N_15278,N_15117,N_15050);
nand U15279 (N_15279,N_15169,N_15042);
nor U15280 (N_15280,N_15145,N_15055);
nor U15281 (N_15281,N_15105,N_15173);
nand U15282 (N_15282,N_15190,N_15068);
nand U15283 (N_15283,N_15052,N_15142);
or U15284 (N_15284,N_15182,N_15172);
and U15285 (N_15285,N_15104,N_15116);
nor U15286 (N_15286,N_15088,N_15081);
and U15287 (N_15287,N_15164,N_15075);
and U15288 (N_15288,N_15061,N_15177);
nand U15289 (N_15289,N_15169,N_15050);
nor U15290 (N_15290,N_15125,N_15064);
or U15291 (N_15291,N_15194,N_15071);
nor U15292 (N_15292,N_15167,N_15151);
nand U15293 (N_15293,N_15153,N_15154);
nand U15294 (N_15294,N_15096,N_15046);
nor U15295 (N_15295,N_15120,N_15157);
and U15296 (N_15296,N_15055,N_15080);
or U15297 (N_15297,N_15080,N_15177);
or U15298 (N_15298,N_15067,N_15062);
and U15299 (N_15299,N_15099,N_15083);
xor U15300 (N_15300,N_15082,N_15051);
or U15301 (N_15301,N_15116,N_15103);
nand U15302 (N_15302,N_15195,N_15058);
nand U15303 (N_15303,N_15146,N_15183);
or U15304 (N_15304,N_15103,N_15176);
nand U15305 (N_15305,N_15195,N_15041);
nor U15306 (N_15306,N_15111,N_15090);
and U15307 (N_15307,N_15178,N_15094);
nand U15308 (N_15308,N_15059,N_15116);
nor U15309 (N_15309,N_15185,N_15063);
nor U15310 (N_15310,N_15044,N_15102);
nor U15311 (N_15311,N_15052,N_15050);
xor U15312 (N_15312,N_15076,N_15107);
nor U15313 (N_15313,N_15131,N_15040);
nand U15314 (N_15314,N_15162,N_15187);
and U15315 (N_15315,N_15097,N_15143);
or U15316 (N_15316,N_15044,N_15076);
or U15317 (N_15317,N_15114,N_15109);
and U15318 (N_15318,N_15064,N_15145);
xnor U15319 (N_15319,N_15112,N_15196);
or U15320 (N_15320,N_15141,N_15173);
and U15321 (N_15321,N_15188,N_15120);
and U15322 (N_15322,N_15050,N_15131);
and U15323 (N_15323,N_15045,N_15157);
and U15324 (N_15324,N_15110,N_15113);
and U15325 (N_15325,N_15192,N_15084);
nor U15326 (N_15326,N_15166,N_15176);
and U15327 (N_15327,N_15147,N_15084);
nor U15328 (N_15328,N_15071,N_15091);
xor U15329 (N_15329,N_15088,N_15124);
xnor U15330 (N_15330,N_15150,N_15077);
nor U15331 (N_15331,N_15193,N_15113);
xor U15332 (N_15332,N_15125,N_15045);
xor U15333 (N_15333,N_15190,N_15142);
or U15334 (N_15334,N_15168,N_15130);
or U15335 (N_15335,N_15064,N_15137);
or U15336 (N_15336,N_15108,N_15118);
nor U15337 (N_15337,N_15056,N_15182);
nand U15338 (N_15338,N_15164,N_15116);
nor U15339 (N_15339,N_15058,N_15132);
nand U15340 (N_15340,N_15150,N_15186);
or U15341 (N_15341,N_15178,N_15048);
xor U15342 (N_15342,N_15170,N_15055);
nor U15343 (N_15343,N_15157,N_15087);
nor U15344 (N_15344,N_15147,N_15143);
nand U15345 (N_15345,N_15182,N_15155);
or U15346 (N_15346,N_15192,N_15148);
or U15347 (N_15347,N_15044,N_15083);
or U15348 (N_15348,N_15158,N_15185);
xor U15349 (N_15349,N_15050,N_15158);
nand U15350 (N_15350,N_15157,N_15196);
nand U15351 (N_15351,N_15176,N_15115);
nand U15352 (N_15352,N_15071,N_15087);
and U15353 (N_15353,N_15042,N_15060);
nor U15354 (N_15354,N_15044,N_15158);
nor U15355 (N_15355,N_15126,N_15044);
nand U15356 (N_15356,N_15170,N_15053);
or U15357 (N_15357,N_15122,N_15087);
and U15358 (N_15358,N_15073,N_15188);
or U15359 (N_15359,N_15125,N_15059);
and U15360 (N_15360,N_15299,N_15279);
and U15361 (N_15361,N_15243,N_15200);
nand U15362 (N_15362,N_15347,N_15208);
or U15363 (N_15363,N_15336,N_15333);
and U15364 (N_15364,N_15254,N_15330);
and U15365 (N_15365,N_15295,N_15315);
nor U15366 (N_15366,N_15359,N_15234);
nand U15367 (N_15367,N_15289,N_15282);
nand U15368 (N_15368,N_15306,N_15353);
nand U15369 (N_15369,N_15247,N_15285);
nor U15370 (N_15370,N_15220,N_15358);
nand U15371 (N_15371,N_15304,N_15334);
nand U15372 (N_15372,N_15351,N_15296);
nand U15373 (N_15373,N_15206,N_15326);
nand U15374 (N_15374,N_15215,N_15349);
nor U15375 (N_15375,N_15273,N_15317);
nand U15376 (N_15376,N_15339,N_15230);
nand U15377 (N_15377,N_15345,N_15210);
nand U15378 (N_15378,N_15316,N_15263);
nand U15379 (N_15379,N_15213,N_15290);
nand U15380 (N_15380,N_15346,N_15265);
xnor U15381 (N_15381,N_15272,N_15314);
nand U15382 (N_15382,N_15258,N_15294);
nor U15383 (N_15383,N_15319,N_15313);
xnor U15384 (N_15384,N_15281,N_15343);
and U15385 (N_15385,N_15300,N_15264);
nand U15386 (N_15386,N_15232,N_15261);
nand U15387 (N_15387,N_15325,N_15202);
and U15388 (N_15388,N_15311,N_15332);
or U15389 (N_15389,N_15226,N_15312);
nand U15390 (N_15390,N_15222,N_15344);
xor U15391 (N_15391,N_15283,N_15341);
nor U15392 (N_15392,N_15348,N_15324);
or U15393 (N_15393,N_15337,N_15301);
and U15394 (N_15394,N_15211,N_15287);
and U15395 (N_15395,N_15217,N_15241);
or U15396 (N_15396,N_15257,N_15357);
nor U15397 (N_15397,N_15307,N_15228);
or U15398 (N_15398,N_15293,N_15249);
nor U15399 (N_15399,N_15223,N_15284);
xnor U15400 (N_15400,N_15335,N_15256);
or U15401 (N_15401,N_15219,N_15248);
and U15402 (N_15402,N_15321,N_15275);
nor U15403 (N_15403,N_15291,N_15340);
and U15404 (N_15404,N_15240,N_15203);
nand U15405 (N_15405,N_15214,N_15276);
nand U15406 (N_15406,N_15270,N_15268);
nor U15407 (N_15407,N_15288,N_15239);
nor U15408 (N_15408,N_15322,N_15309);
or U15409 (N_15409,N_15242,N_15237);
xor U15410 (N_15410,N_15352,N_15320);
nor U15411 (N_15411,N_15267,N_15280);
or U15412 (N_15412,N_15329,N_15308);
or U15413 (N_15413,N_15218,N_15246);
and U15414 (N_15414,N_15271,N_15235);
or U15415 (N_15415,N_15302,N_15238);
nand U15416 (N_15416,N_15277,N_15207);
and U15417 (N_15417,N_15318,N_15327);
or U15418 (N_15418,N_15310,N_15227);
or U15419 (N_15419,N_15323,N_15224);
xnor U15420 (N_15420,N_15303,N_15356);
or U15421 (N_15421,N_15305,N_15252);
xor U15422 (N_15422,N_15259,N_15231);
nor U15423 (N_15423,N_15236,N_15328);
or U15424 (N_15424,N_15342,N_15209);
xor U15425 (N_15425,N_15216,N_15212);
or U15426 (N_15426,N_15255,N_15297);
nor U15427 (N_15427,N_15338,N_15331);
and U15428 (N_15428,N_15274,N_15355);
nor U15429 (N_15429,N_15278,N_15245);
nor U15430 (N_15430,N_15251,N_15229);
and U15431 (N_15431,N_15260,N_15354);
nor U15432 (N_15432,N_15201,N_15233);
nand U15433 (N_15433,N_15266,N_15221);
xnor U15434 (N_15434,N_15250,N_15204);
nand U15435 (N_15435,N_15205,N_15262);
nand U15436 (N_15436,N_15253,N_15269);
nand U15437 (N_15437,N_15292,N_15244);
xnor U15438 (N_15438,N_15350,N_15298);
and U15439 (N_15439,N_15225,N_15286);
xor U15440 (N_15440,N_15256,N_15307);
xnor U15441 (N_15441,N_15217,N_15308);
and U15442 (N_15442,N_15243,N_15312);
xor U15443 (N_15443,N_15208,N_15284);
nor U15444 (N_15444,N_15226,N_15225);
and U15445 (N_15445,N_15255,N_15354);
or U15446 (N_15446,N_15200,N_15231);
and U15447 (N_15447,N_15355,N_15353);
or U15448 (N_15448,N_15254,N_15213);
and U15449 (N_15449,N_15250,N_15290);
and U15450 (N_15450,N_15314,N_15210);
and U15451 (N_15451,N_15237,N_15266);
nand U15452 (N_15452,N_15243,N_15340);
or U15453 (N_15453,N_15268,N_15352);
nand U15454 (N_15454,N_15248,N_15250);
or U15455 (N_15455,N_15224,N_15342);
and U15456 (N_15456,N_15300,N_15217);
xnor U15457 (N_15457,N_15284,N_15316);
nand U15458 (N_15458,N_15285,N_15337);
and U15459 (N_15459,N_15246,N_15338);
or U15460 (N_15460,N_15292,N_15342);
nand U15461 (N_15461,N_15215,N_15225);
and U15462 (N_15462,N_15278,N_15301);
or U15463 (N_15463,N_15347,N_15295);
nand U15464 (N_15464,N_15334,N_15340);
or U15465 (N_15465,N_15213,N_15279);
xor U15466 (N_15466,N_15236,N_15303);
nand U15467 (N_15467,N_15297,N_15217);
or U15468 (N_15468,N_15239,N_15256);
nand U15469 (N_15469,N_15316,N_15225);
xor U15470 (N_15470,N_15299,N_15214);
nand U15471 (N_15471,N_15230,N_15270);
or U15472 (N_15472,N_15341,N_15344);
nand U15473 (N_15473,N_15232,N_15269);
nand U15474 (N_15474,N_15256,N_15200);
nor U15475 (N_15475,N_15261,N_15255);
nor U15476 (N_15476,N_15344,N_15279);
nand U15477 (N_15477,N_15234,N_15216);
nand U15478 (N_15478,N_15321,N_15293);
and U15479 (N_15479,N_15259,N_15339);
nand U15480 (N_15480,N_15327,N_15319);
nand U15481 (N_15481,N_15217,N_15291);
or U15482 (N_15482,N_15249,N_15348);
xor U15483 (N_15483,N_15246,N_15297);
or U15484 (N_15484,N_15278,N_15232);
nand U15485 (N_15485,N_15350,N_15252);
and U15486 (N_15486,N_15343,N_15208);
xnor U15487 (N_15487,N_15201,N_15274);
and U15488 (N_15488,N_15290,N_15322);
nor U15489 (N_15489,N_15279,N_15300);
nand U15490 (N_15490,N_15210,N_15259);
nand U15491 (N_15491,N_15325,N_15358);
and U15492 (N_15492,N_15219,N_15277);
nand U15493 (N_15493,N_15296,N_15343);
or U15494 (N_15494,N_15218,N_15263);
or U15495 (N_15495,N_15289,N_15267);
nand U15496 (N_15496,N_15242,N_15293);
and U15497 (N_15497,N_15263,N_15242);
or U15498 (N_15498,N_15263,N_15272);
or U15499 (N_15499,N_15316,N_15326);
nor U15500 (N_15500,N_15279,N_15328);
or U15501 (N_15501,N_15327,N_15268);
or U15502 (N_15502,N_15272,N_15340);
nand U15503 (N_15503,N_15259,N_15242);
or U15504 (N_15504,N_15278,N_15262);
nand U15505 (N_15505,N_15255,N_15219);
or U15506 (N_15506,N_15317,N_15204);
nand U15507 (N_15507,N_15346,N_15238);
or U15508 (N_15508,N_15289,N_15263);
nor U15509 (N_15509,N_15346,N_15359);
xor U15510 (N_15510,N_15289,N_15284);
and U15511 (N_15511,N_15279,N_15249);
nor U15512 (N_15512,N_15315,N_15211);
xor U15513 (N_15513,N_15241,N_15239);
nor U15514 (N_15514,N_15289,N_15325);
and U15515 (N_15515,N_15201,N_15356);
nand U15516 (N_15516,N_15349,N_15356);
nor U15517 (N_15517,N_15263,N_15268);
nand U15518 (N_15518,N_15287,N_15276);
nor U15519 (N_15519,N_15257,N_15275);
nand U15520 (N_15520,N_15371,N_15497);
or U15521 (N_15521,N_15505,N_15361);
or U15522 (N_15522,N_15407,N_15513);
and U15523 (N_15523,N_15473,N_15400);
or U15524 (N_15524,N_15475,N_15450);
and U15525 (N_15525,N_15439,N_15474);
nand U15526 (N_15526,N_15478,N_15461);
or U15527 (N_15527,N_15443,N_15472);
xnor U15528 (N_15528,N_15373,N_15414);
or U15529 (N_15529,N_15389,N_15405);
and U15530 (N_15530,N_15420,N_15422);
or U15531 (N_15531,N_15427,N_15457);
or U15532 (N_15532,N_15368,N_15454);
and U15533 (N_15533,N_15463,N_15378);
and U15534 (N_15534,N_15435,N_15442);
nand U15535 (N_15535,N_15428,N_15429);
and U15536 (N_15536,N_15369,N_15449);
and U15537 (N_15537,N_15360,N_15409);
nor U15538 (N_15538,N_15381,N_15496);
nand U15539 (N_15539,N_15434,N_15469);
and U15540 (N_15540,N_15468,N_15506);
nor U15541 (N_15541,N_15500,N_15466);
nor U15542 (N_15542,N_15484,N_15483);
and U15543 (N_15543,N_15430,N_15515);
or U15544 (N_15544,N_15467,N_15417);
or U15545 (N_15545,N_15410,N_15411);
or U15546 (N_15546,N_15367,N_15388);
and U15547 (N_15547,N_15419,N_15433);
nand U15548 (N_15548,N_15476,N_15431);
nor U15549 (N_15549,N_15421,N_15432);
nand U15550 (N_15550,N_15489,N_15510);
nand U15551 (N_15551,N_15392,N_15480);
and U15552 (N_15552,N_15376,N_15437);
and U15553 (N_15553,N_15374,N_15493);
nand U15554 (N_15554,N_15495,N_15459);
or U15555 (N_15555,N_15458,N_15486);
and U15556 (N_15556,N_15390,N_15363);
nor U15557 (N_15557,N_15377,N_15387);
or U15558 (N_15558,N_15464,N_15362);
xor U15559 (N_15559,N_15451,N_15516);
nor U15560 (N_15560,N_15479,N_15365);
or U15561 (N_15561,N_15372,N_15504);
nor U15562 (N_15562,N_15519,N_15492);
nand U15563 (N_15563,N_15502,N_15364);
nand U15564 (N_15564,N_15402,N_15436);
and U15565 (N_15565,N_15487,N_15398);
xnor U15566 (N_15566,N_15517,N_15384);
and U15567 (N_15567,N_15465,N_15382);
and U15568 (N_15568,N_15394,N_15424);
or U15569 (N_15569,N_15403,N_15456);
or U15570 (N_15570,N_15441,N_15404);
and U15571 (N_15571,N_15455,N_15418);
xor U15572 (N_15572,N_15477,N_15485);
nand U15573 (N_15573,N_15471,N_15498);
and U15574 (N_15574,N_15462,N_15396);
xnor U15575 (N_15575,N_15514,N_15447);
or U15576 (N_15576,N_15494,N_15366);
xor U15577 (N_15577,N_15518,N_15482);
nand U15578 (N_15578,N_15408,N_15448);
nor U15579 (N_15579,N_15453,N_15444);
nor U15580 (N_15580,N_15395,N_15445);
or U15581 (N_15581,N_15423,N_15379);
nand U15582 (N_15582,N_15509,N_15438);
xnor U15583 (N_15583,N_15481,N_15511);
or U15584 (N_15584,N_15383,N_15499);
or U15585 (N_15585,N_15380,N_15425);
xnor U15586 (N_15586,N_15375,N_15488);
xor U15587 (N_15587,N_15386,N_15490);
nor U15588 (N_15588,N_15370,N_15385);
nand U15589 (N_15589,N_15391,N_15501);
xor U15590 (N_15590,N_15393,N_15508);
or U15591 (N_15591,N_15426,N_15507);
xor U15592 (N_15592,N_15415,N_15452);
or U15593 (N_15593,N_15440,N_15406);
nor U15594 (N_15594,N_15399,N_15491);
and U15595 (N_15595,N_15446,N_15397);
nand U15596 (N_15596,N_15503,N_15460);
nor U15597 (N_15597,N_15470,N_15416);
and U15598 (N_15598,N_15412,N_15401);
nand U15599 (N_15599,N_15413,N_15512);
nor U15600 (N_15600,N_15402,N_15461);
xnor U15601 (N_15601,N_15493,N_15400);
and U15602 (N_15602,N_15427,N_15405);
or U15603 (N_15603,N_15502,N_15479);
nand U15604 (N_15604,N_15437,N_15440);
nor U15605 (N_15605,N_15391,N_15484);
and U15606 (N_15606,N_15487,N_15392);
or U15607 (N_15607,N_15516,N_15370);
and U15608 (N_15608,N_15484,N_15487);
nor U15609 (N_15609,N_15484,N_15477);
or U15610 (N_15610,N_15433,N_15406);
nor U15611 (N_15611,N_15425,N_15421);
nor U15612 (N_15612,N_15466,N_15447);
nor U15613 (N_15613,N_15445,N_15512);
and U15614 (N_15614,N_15451,N_15413);
nor U15615 (N_15615,N_15519,N_15414);
or U15616 (N_15616,N_15463,N_15364);
or U15617 (N_15617,N_15515,N_15391);
or U15618 (N_15618,N_15501,N_15425);
and U15619 (N_15619,N_15446,N_15498);
or U15620 (N_15620,N_15434,N_15417);
nor U15621 (N_15621,N_15474,N_15445);
nand U15622 (N_15622,N_15487,N_15504);
nor U15623 (N_15623,N_15450,N_15458);
xor U15624 (N_15624,N_15386,N_15508);
and U15625 (N_15625,N_15477,N_15368);
and U15626 (N_15626,N_15476,N_15377);
nor U15627 (N_15627,N_15394,N_15436);
and U15628 (N_15628,N_15430,N_15452);
and U15629 (N_15629,N_15460,N_15441);
and U15630 (N_15630,N_15402,N_15434);
and U15631 (N_15631,N_15394,N_15407);
nor U15632 (N_15632,N_15381,N_15489);
nand U15633 (N_15633,N_15367,N_15494);
or U15634 (N_15634,N_15510,N_15430);
and U15635 (N_15635,N_15443,N_15515);
xnor U15636 (N_15636,N_15365,N_15452);
xnor U15637 (N_15637,N_15396,N_15517);
and U15638 (N_15638,N_15510,N_15378);
nand U15639 (N_15639,N_15412,N_15495);
and U15640 (N_15640,N_15458,N_15491);
and U15641 (N_15641,N_15438,N_15503);
and U15642 (N_15642,N_15464,N_15363);
and U15643 (N_15643,N_15362,N_15468);
xnor U15644 (N_15644,N_15481,N_15366);
nor U15645 (N_15645,N_15369,N_15488);
nand U15646 (N_15646,N_15514,N_15364);
nor U15647 (N_15647,N_15502,N_15516);
nor U15648 (N_15648,N_15409,N_15399);
or U15649 (N_15649,N_15474,N_15365);
nand U15650 (N_15650,N_15378,N_15493);
nor U15651 (N_15651,N_15440,N_15481);
and U15652 (N_15652,N_15506,N_15495);
or U15653 (N_15653,N_15473,N_15487);
or U15654 (N_15654,N_15455,N_15511);
xnor U15655 (N_15655,N_15512,N_15471);
nand U15656 (N_15656,N_15452,N_15448);
nand U15657 (N_15657,N_15485,N_15501);
nor U15658 (N_15658,N_15502,N_15408);
nand U15659 (N_15659,N_15403,N_15467);
and U15660 (N_15660,N_15441,N_15414);
and U15661 (N_15661,N_15416,N_15412);
nand U15662 (N_15662,N_15485,N_15503);
and U15663 (N_15663,N_15398,N_15507);
or U15664 (N_15664,N_15500,N_15399);
nor U15665 (N_15665,N_15425,N_15507);
nand U15666 (N_15666,N_15491,N_15372);
or U15667 (N_15667,N_15482,N_15499);
nor U15668 (N_15668,N_15360,N_15385);
nor U15669 (N_15669,N_15468,N_15488);
nand U15670 (N_15670,N_15457,N_15491);
or U15671 (N_15671,N_15369,N_15479);
or U15672 (N_15672,N_15505,N_15380);
nor U15673 (N_15673,N_15493,N_15503);
or U15674 (N_15674,N_15365,N_15406);
or U15675 (N_15675,N_15361,N_15432);
and U15676 (N_15676,N_15412,N_15432);
nand U15677 (N_15677,N_15370,N_15397);
nor U15678 (N_15678,N_15414,N_15466);
nor U15679 (N_15679,N_15508,N_15394);
or U15680 (N_15680,N_15655,N_15648);
or U15681 (N_15681,N_15619,N_15672);
or U15682 (N_15682,N_15553,N_15577);
and U15683 (N_15683,N_15567,N_15677);
nand U15684 (N_15684,N_15580,N_15651);
or U15685 (N_15685,N_15678,N_15635);
nand U15686 (N_15686,N_15650,N_15581);
nor U15687 (N_15687,N_15556,N_15574);
nand U15688 (N_15688,N_15646,N_15578);
and U15689 (N_15689,N_15614,N_15552);
and U15690 (N_15690,N_15644,N_15625);
xor U15691 (N_15691,N_15579,N_15535);
nand U15692 (N_15692,N_15632,N_15620);
xnor U15693 (N_15693,N_15561,N_15596);
and U15694 (N_15694,N_15566,N_15569);
nor U15695 (N_15695,N_15662,N_15666);
xor U15696 (N_15696,N_15545,N_15593);
nand U15697 (N_15697,N_15618,N_15631);
nand U15698 (N_15698,N_15537,N_15613);
nor U15699 (N_15699,N_15562,N_15661);
nand U15700 (N_15700,N_15645,N_15594);
nand U15701 (N_15701,N_15653,N_15674);
or U15702 (N_15702,N_15639,N_15675);
nand U15703 (N_15703,N_15627,N_15621);
nor U15704 (N_15704,N_15643,N_15564);
or U15705 (N_15705,N_15670,N_15602);
nor U15706 (N_15706,N_15636,N_15547);
nand U15707 (N_15707,N_15647,N_15575);
or U15708 (N_15708,N_15604,N_15607);
nand U15709 (N_15709,N_15598,N_15551);
and U15710 (N_15710,N_15676,N_15633);
nor U15711 (N_15711,N_15652,N_15559);
nand U15712 (N_15712,N_15571,N_15603);
or U15713 (N_15713,N_15521,N_15623);
and U15714 (N_15714,N_15611,N_15669);
or U15715 (N_15715,N_15533,N_15657);
and U15716 (N_15716,N_15656,N_15534);
nand U15717 (N_15717,N_15520,N_15610);
nand U15718 (N_15718,N_15601,N_15586);
nor U15719 (N_15719,N_15591,N_15638);
and U15720 (N_15720,N_15570,N_15568);
xor U15721 (N_15721,N_15560,N_15588);
nor U15722 (N_15722,N_15524,N_15608);
nor U15723 (N_15723,N_15654,N_15573);
and U15724 (N_15724,N_15528,N_15663);
nor U15725 (N_15725,N_15558,N_15595);
nor U15726 (N_15726,N_15550,N_15617);
or U15727 (N_15727,N_15659,N_15549);
xnor U15728 (N_15728,N_15587,N_15615);
and U15729 (N_15729,N_15538,N_15582);
and U15730 (N_15730,N_15616,N_15526);
nand U15731 (N_15731,N_15555,N_15630);
nor U15732 (N_15732,N_15649,N_15525);
and U15733 (N_15733,N_15548,N_15624);
nand U15734 (N_15734,N_15637,N_15532);
nor U15735 (N_15735,N_15554,N_15565);
and U15736 (N_15736,N_15605,N_15640);
or U15737 (N_15737,N_15546,N_15592);
and U15738 (N_15738,N_15599,N_15671);
and U15739 (N_15739,N_15629,N_15628);
xor U15740 (N_15740,N_15557,N_15543);
nand U15741 (N_15741,N_15529,N_15665);
and U15742 (N_15742,N_15658,N_15541);
and U15743 (N_15743,N_15667,N_15668);
nor U15744 (N_15744,N_15609,N_15642);
and U15745 (N_15745,N_15536,N_15542);
and U15746 (N_15746,N_15523,N_15585);
nand U15747 (N_15747,N_15589,N_15531);
nor U15748 (N_15748,N_15634,N_15606);
or U15749 (N_15749,N_15590,N_15664);
and U15750 (N_15750,N_15540,N_15641);
or U15751 (N_15751,N_15612,N_15583);
and U15752 (N_15752,N_15530,N_15600);
nor U15753 (N_15753,N_15679,N_15576);
or U15754 (N_15754,N_15522,N_15572);
nand U15755 (N_15755,N_15527,N_15544);
or U15756 (N_15756,N_15584,N_15597);
nand U15757 (N_15757,N_15660,N_15539);
and U15758 (N_15758,N_15563,N_15626);
nand U15759 (N_15759,N_15622,N_15673);
and U15760 (N_15760,N_15521,N_15528);
nor U15761 (N_15761,N_15654,N_15549);
nand U15762 (N_15762,N_15561,N_15601);
nand U15763 (N_15763,N_15556,N_15614);
or U15764 (N_15764,N_15566,N_15581);
nor U15765 (N_15765,N_15622,N_15604);
and U15766 (N_15766,N_15541,N_15592);
nand U15767 (N_15767,N_15576,N_15636);
nor U15768 (N_15768,N_15600,N_15558);
nand U15769 (N_15769,N_15547,N_15620);
xnor U15770 (N_15770,N_15652,N_15580);
nor U15771 (N_15771,N_15642,N_15645);
and U15772 (N_15772,N_15601,N_15675);
or U15773 (N_15773,N_15623,N_15545);
nand U15774 (N_15774,N_15647,N_15589);
and U15775 (N_15775,N_15648,N_15539);
nor U15776 (N_15776,N_15593,N_15602);
nor U15777 (N_15777,N_15664,N_15576);
nand U15778 (N_15778,N_15662,N_15555);
or U15779 (N_15779,N_15639,N_15613);
nand U15780 (N_15780,N_15657,N_15535);
or U15781 (N_15781,N_15605,N_15562);
nor U15782 (N_15782,N_15637,N_15536);
nand U15783 (N_15783,N_15616,N_15562);
or U15784 (N_15784,N_15602,N_15552);
and U15785 (N_15785,N_15646,N_15547);
or U15786 (N_15786,N_15521,N_15585);
xor U15787 (N_15787,N_15529,N_15534);
or U15788 (N_15788,N_15586,N_15648);
nor U15789 (N_15789,N_15642,N_15538);
or U15790 (N_15790,N_15608,N_15615);
xor U15791 (N_15791,N_15550,N_15585);
and U15792 (N_15792,N_15664,N_15605);
or U15793 (N_15793,N_15651,N_15539);
or U15794 (N_15794,N_15676,N_15565);
nand U15795 (N_15795,N_15637,N_15664);
and U15796 (N_15796,N_15675,N_15561);
nor U15797 (N_15797,N_15611,N_15560);
or U15798 (N_15798,N_15604,N_15530);
nand U15799 (N_15799,N_15660,N_15570);
xor U15800 (N_15800,N_15633,N_15607);
nand U15801 (N_15801,N_15600,N_15660);
nor U15802 (N_15802,N_15653,N_15520);
or U15803 (N_15803,N_15647,N_15538);
nand U15804 (N_15804,N_15526,N_15527);
nor U15805 (N_15805,N_15621,N_15612);
and U15806 (N_15806,N_15614,N_15615);
nand U15807 (N_15807,N_15643,N_15544);
xor U15808 (N_15808,N_15659,N_15554);
nor U15809 (N_15809,N_15555,N_15535);
nand U15810 (N_15810,N_15620,N_15581);
and U15811 (N_15811,N_15532,N_15614);
or U15812 (N_15812,N_15621,N_15678);
nand U15813 (N_15813,N_15590,N_15677);
nor U15814 (N_15814,N_15665,N_15635);
and U15815 (N_15815,N_15667,N_15598);
and U15816 (N_15816,N_15580,N_15585);
and U15817 (N_15817,N_15572,N_15558);
or U15818 (N_15818,N_15618,N_15604);
nand U15819 (N_15819,N_15539,N_15568);
or U15820 (N_15820,N_15672,N_15669);
xor U15821 (N_15821,N_15667,N_15602);
and U15822 (N_15822,N_15586,N_15581);
nand U15823 (N_15823,N_15573,N_15628);
xnor U15824 (N_15824,N_15598,N_15567);
nand U15825 (N_15825,N_15556,N_15633);
nor U15826 (N_15826,N_15614,N_15535);
xnor U15827 (N_15827,N_15673,N_15543);
nor U15828 (N_15828,N_15541,N_15613);
nor U15829 (N_15829,N_15653,N_15531);
and U15830 (N_15830,N_15628,N_15662);
and U15831 (N_15831,N_15633,N_15539);
nor U15832 (N_15832,N_15607,N_15662);
and U15833 (N_15833,N_15661,N_15585);
or U15834 (N_15834,N_15594,N_15547);
nor U15835 (N_15835,N_15595,N_15617);
xor U15836 (N_15836,N_15674,N_15563);
and U15837 (N_15837,N_15554,N_15610);
and U15838 (N_15838,N_15618,N_15642);
or U15839 (N_15839,N_15571,N_15537);
nor U15840 (N_15840,N_15747,N_15826);
and U15841 (N_15841,N_15715,N_15731);
xnor U15842 (N_15842,N_15714,N_15752);
nor U15843 (N_15843,N_15759,N_15818);
nand U15844 (N_15844,N_15833,N_15798);
nand U15845 (N_15845,N_15771,N_15696);
or U15846 (N_15846,N_15809,N_15708);
nand U15847 (N_15847,N_15837,N_15801);
nand U15848 (N_15848,N_15740,N_15834);
or U15849 (N_15849,N_15773,N_15791);
nand U15850 (N_15850,N_15748,N_15777);
or U15851 (N_15851,N_15795,N_15758);
and U15852 (N_15852,N_15706,N_15757);
nor U15853 (N_15853,N_15836,N_15824);
or U15854 (N_15854,N_15703,N_15739);
or U15855 (N_15855,N_15832,N_15812);
or U15856 (N_15856,N_15754,N_15767);
nand U15857 (N_15857,N_15693,N_15689);
nor U15858 (N_15858,N_15681,N_15698);
and U15859 (N_15859,N_15727,N_15794);
nand U15860 (N_15860,N_15728,N_15779);
nand U15861 (N_15861,N_15733,N_15797);
and U15862 (N_15862,N_15707,N_15803);
and U15863 (N_15863,N_15827,N_15792);
nor U15864 (N_15864,N_15685,N_15699);
nand U15865 (N_15865,N_15702,N_15680);
and U15866 (N_15866,N_15783,N_15806);
nand U15867 (N_15867,N_15770,N_15738);
nor U15868 (N_15868,N_15695,N_15785);
nor U15869 (N_15869,N_15700,N_15787);
nand U15870 (N_15870,N_15742,N_15776);
nor U15871 (N_15871,N_15820,N_15743);
nand U15872 (N_15872,N_15741,N_15781);
xnor U15873 (N_15873,N_15735,N_15710);
or U15874 (N_15874,N_15761,N_15817);
or U15875 (N_15875,N_15730,N_15719);
and U15876 (N_15876,N_15705,N_15692);
and U15877 (N_15877,N_15819,N_15737);
or U15878 (N_15878,N_15813,N_15823);
nor U15879 (N_15879,N_15688,N_15772);
and U15880 (N_15880,N_15799,N_15804);
nor U15881 (N_15881,N_15768,N_15831);
and U15882 (N_15882,N_15775,N_15732);
and U15883 (N_15883,N_15691,N_15835);
or U15884 (N_15884,N_15753,N_15782);
nand U15885 (N_15885,N_15721,N_15734);
nand U15886 (N_15886,N_15790,N_15796);
nand U15887 (N_15887,N_15725,N_15717);
nor U15888 (N_15888,N_15704,N_15766);
nand U15889 (N_15889,N_15774,N_15746);
nand U15890 (N_15890,N_15829,N_15722);
nand U15891 (N_15891,N_15736,N_15755);
and U15892 (N_15892,N_15763,N_15788);
nand U15893 (N_15893,N_15828,N_15697);
nand U15894 (N_15894,N_15839,N_15808);
nand U15895 (N_15895,N_15816,N_15713);
and U15896 (N_15896,N_15786,N_15784);
nor U15897 (N_15897,N_15830,N_15793);
nand U15898 (N_15898,N_15800,N_15711);
nand U15899 (N_15899,N_15760,N_15764);
nand U15900 (N_15900,N_15821,N_15684);
xnor U15901 (N_15901,N_15729,N_15769);
nor U15902 (N_15902,N_15690,N_15682);
nor U15903 (N_15903,N_15701,N_15750);
nor U15904 (N_15904,N_15749,N_15687);
and U15905 (N_15905,N_15778,N_15744);
or U15906 (N_15906,N_15694,N_15683);
and U15907 (N_15907,N_15838,N_15726);
nor U15908 (N_15908,N_15751,N_15814);
or U15909 (N_15909,N_15716,N_15802);
or U15910 (N_15910,N_15789,N_15805);
nor U15911 (N_15911,N_15709,N_15762);
nand U15912 (N_15912,N_15765,N_15720);
and U15913 (N_15913,N_15780,N_15825);
nor U15914 (N_15914,N_15686,N_15745);
and U15915 (N_15915,N_15811,N_15756);
or U15916 (N_15916,N_15822,N_15815);
nand U15917 (N_15917,N_15810,N_15807);
and U15918 (N_15918,N_15712,N_15718);
nand U15919 (N_15919,N_15723,N_15724);
or U15920 (N_15920,N_15833,N_15738);
and U15921 (N_15921,N_15834,N_15809);
nand U15922 (N_15922,N_15756,N_15754);
nor U15923 (N_15923,N_15775,N_15727);
nor U15924 (N_15924,N_15691,N_15790);
nor U15925 (N_15925,N_15759,N_15778);
or U15926 (N_15926,N_15704,N_15795);
nand U15927 (N_15927,N_15697,N_15683);
and U15928 (N_15928,N_15736,N_15741);
and U15929 (N_15929,N_15683,N_15790);
xor U15930 (N_15930,N_15713,N_15822);
nor U15931 (N_15931,N_15771,N_15835);
nand U15932 (N_15932,N_15812,N_15791);
xnor U15933 (N_15933,N_15789,N_15737);
xor U15934 (N_15934,N_15812,N_15828);
or U15935 (N_15935,N_15743,N_15815);
and U15936 (N_15936,N_15798,N_15711);
nor U15937 (N_15937,N_15794,N_15705);
or U15938 (N_15938,N_15774,N_15823);
nor U15939 (N_15939,N_15689,N_15751);
or U15940 (N_15940,N_15822,N_15691);
nor U15941 (N_15941,N_15764,N_15738);
nand U15942 (N_15942,N_15751,N_15710);
or U15943 (N_15943,N_15796,N_15820);
xor U15944 (N_15944,N_15824,N_15755);
nor U15945 (N_15945,N_15685,N_15742);
or U15946 (N_15946,N_15764,N_15711);
or U15947 (N_15947,N_15703,N_15826);
and U15948 (N_15948,N_15795,N_15681);
and U15949 (N_15949,N_15760,N_15693);
nor U15950 (N_15950,N_15721,N_15837);
nor U15951 (N_15951,N_15802,N_15835);
nor U15952 (N_15952,N_15715,N_15760);
xnor U15953 (N_15953,N_15763,N_15743);
xor U15954 (N_15954,N_15716,N_15754);
nand U15955 (N_15955,N_15775,N_15813);
or U15956 (N_15956,N_15691,N_15681);
and U15957 (N_15957,N_15784,N_15781);
nor U15958 (N_15958,N_15689,N_15743);
nor U15959 (N_15959,N_15706,N_15773);
or U15960 (N_15960,N_15812,N_15737);
and U15961 (N_15961,N_15818,N_15800);
and U15962 (N_15962,N_15839,N_15765);
nor U15963 (N_15963,N_15698,N_15748);
and U15964 (N_15964,N_15774,N_15821);
nand U15965 (N_15965,N_15759,N_15738);
xnor U15966 (N_15966,N_15765,N_15749);
nor U15967 (N_15967,N_15833,N_15758);
xnor U15968 (N_15968,N_15830,N_15719);
nor U15969 (N_15969,N_15741,N_15829);
nand U15970 (N_15970,N_15775,N_15774);
nand U15971 (N_15971,N_15813,N_15757);
and U15972 (N_15972,N_15803,N_15689);
nor U15973 (N_15973,N_15795,N_15765);
xnor U15974 (N_15974,N_15823,N_15836);
nor U15975 (N_15975,N_15764,N_15694);
and U15976 (N_15976,N_15696,N_15729);
or U15977 (N_15977,N_15776,N_15683);
nor U15978 (N_15978,N_15802,N_15746);
nor U15979 (N_15979,N_15708,N_15775);
nor U15980 (N_15980,N_15691,N_15748);
xor U15981 (N_15981,N_15786,N_15798);
nand U15982 (N_15982,N_15743,N_15832);
xnor U15983 (N_15983,N_15715,N_15685);
nor U15984 (N_15984,N_15796,N_15775);
and U15985 (N_15985,N_15731,N_15809);
nor U15986 (N_15986,N_15777,N_15713);
nand U15987 (N_15987,N_15744,N_15789);
nand U15988 (N_15988,N_15788,N_15694);
and U15989 (N_15989,N_15795,N_15818);
nand U15990 (N_15990,N_15696,N_15782);
nand U15991 (N_15991,N_15814,N_15787);
nor U15992 (N_15992,N_15742,N_15812);
or U15993 (N_15993,N_15769,N_15718);
nor U15994 (N_15994,N_15695,N_15732);
and U15995 (N_15995,N_15831,N_15803);
or U15996 (N_15996,N_15787,N_15815);
or U15997 (N_15997,N_15756,N_15694);
and U15998 (N_15998,N_15774,N_15820);
nor U15999 (N_15999,N_15828,N_15723);
nand U16000 (N_16000,N_15901,N_15948);
xor U16001 (N_16001,N_15860,N_15853);
or U16002 (N_16002,N_15913,N_15992);
or U16003 (N_16003,N_15906,N_15940);
or U16004 (N_16004,N_15896,N_15920);
nor U16005 (N_16005,N_15963,N_15909);
or U16006 (N_16006,N_15994,N_15847);
nor U16007 (N_16007,N_15974,N_15980);
nand U16008 (N_16008,N_15949,N_15910);
nand U16009 (N_16009,N_15856,N_15958);
nand U16010 (N_16010,N_15876,N_15862);
and U16011 (N_16011,N_15968,N_15983);
or U16012 (N_16012,N_15996,N_15918);
nand U16013 (N_16013,N_15916,N_15848);
and U16014 (N_16014,N_15883,N_15938);
nor U16015 (N_16015,N_15854,N_15899);
nor U16016 (N_16016,N_15959,N_15957);
nor U16017 (N_16017,N_15846,N_15986);
nor U16018 (N_16018,N_15872,N_15991);
nand U16019 (N_16019,N_15880,N_15930);
or U16020 (N_16020,N_15905,N_15864);
or U16021 (N_16021,N_15937,N_15945);
or U16022 (N_16022,N_15891,N_15921);
or U16023 (N_16023,N_15998,N_15893);
nor U16024 (N_16024,N_15889,N_15990);
nand U16025 (N_16025,N_15852,N_15844);
and U16026 (N_16026,N_15900,N_15923);
nand U16027 (N_16027,N_15870,N_15933);
and U16028 (N_16028,N_15977,N_15851);
nand U16029 (N_16029,N_15857,N_15925);
xor U16030 (N_16030,N_15987,N_15915);
xor U16031 (N_16031,N_15903,N_15967);
nand U16032 (N_16032,N_15942,N_15989);
nand U16033 (N_16033,N_15935,N_15904);
nand U16034 (N_16034,N_15975,N_15960);
nand U16035 (N_16035,N_15941,N_15962);
nor U16036 (N_16036,N_15932,N_15902);
nor U16037 (N_16037,N_15969,N_15882);
and U16038 (N_16038,N_15954,N_15950);
or U16039 (N_16039,N_15911,N_15917);
or U16040 (N_16040,N_15895,N_15976);
and U16041 (N_16041,N_15850,N_15863);
or U16042 (N_16042,N_15877,N_15947);
or U16043 (N_16043,N_15971,N_15881);
or U16044 (N_16044,N_15873,N_15928);
and U16045 (N_16045,N_15908,N_15919);
nand U16046 (N_16046,N_15878,N_15843);
nor U16047 (N_16047,N_15946,N_15943);
nor U16048 (N_16048,N_15972,N_15897);
or U16049 (N_16049,N_15995,N_15981);
nor U16050 (N_16050,N_15855,N_15924);
nor U16051 (N_16051,N_15894,N_15993);
and U16052 (N_16052,N_15845,N_15875);
or U16053 (N_16053,N_15874,N_15973);
or U16054 (N_16054,N_15929,N_15979);
or U16055 (N_16055,N_15965,N_15912);
or U16056 (N_16056,N_15984,N_15892);
and U16057 (N_16057,N_15982,N_15927);
and U16058 (N_16058,N_15867,N_15868);
nor U16059 (N_16059,N_15988,N_15842);
nor U16060 (N_16060,N_15926,N_15966);
nand U16061 (N_16061,N_15978,N_15885);
nand U16062 (N_16062,N_15956,N_15884);
nand U16063 (N_16063,N_15955,N_15953);
or U16064 (N_16064,N_15841,N_15936);
and U16065 (N_16065,N_15922,N_15931);
nand U16066 (N_16066,N_15939,N_15861);
nand U16067 (N_16067,N_15890,N_15858);
or U16068 (N_16068,N_15999,N_15964);
or U16069 (N_16069,N_15961,N_15869);
nor U16070 (N_16070,N_15886,N_15879);
or U16071 (N_16071,N_15866,N_15952);
nand U16072 (N_16072,N_15871,N_15951);
nand U16073 (N_16073,N_15914,N_15888);
or U16074 (N_16074,N_15859,N_15944);
nand U16075 (N_16075,N_15934,N_15887);
or U16076 (N_16076,N_15970,N_15898);
nand U16077 (N_16077,N_15985,N_15840);
xor U16078 (N_16078,N_15907,N_15997);
nand U16079 (N_16079,N_15865,N_15849);
or U16080 (N_16080,N_15992,N_15900);
and U16081 (N_16081,N_15903,N_15871);
or U16082 (N_16082,N_15891,N_15912);
and U16083 (N_16083,N_15973,N_15943);
or U16084 (N_16084,N_15858,N_15944);
nand U16085 (N_16085,N_15856,N_15907);
and U16086 (N_16086,N_15903,N_15866);
nand U16087 (N_16087,N_15928,N_15977);
or U16088 (N_16088,N_15983,N_15867);
and U16089 (N_16089,N_15870,N_15963);
and U16090 (N_16090,N_15904,N_15844);
nor U16091 (N_16091,N_15923,N_15886);
or U16092 (N_16092,N_15961,N_15946);
nor U16093 (N_16093,N_15975,N_15945);
nor U16094 (N_16094,N_15843,N_15939);
nor U16095 (N_16095,N_15950,N_15949);
or U16096 (N_16096,N_15969,N_15993);
nor U16097 (N_16097,N_15926,N_15878);
or U16098 (N_16098,N_15880,N_15848);
xnor U16099 (N_16099,N_15904,N_15985);
or U16100 (N_16100,N_15845,N_15955);
and U16101 (N_16101,N_15862,N_15948);
or U16102 (N_16102,N_15881,N_15886);
or U16103 (N_16103,N_15940,N_15912);
nand U16104 (N_16104,N_15894,N_15880);
or U16105 (N_16105,N_15998,N_15979);
or U16106 (N_16106,N_15980,N_15986);
or U16107 (N_16107,N_15877,N_15920);
and U16108 (N_16108,N_15924,N_15953);
and U16109 (N_16109,N_15926,N_15855);
and U16110 (N_16110,N_15848,N_15949);
and U16111 (N_16111,N_15886,N_15962);
nand U16112 (N_16112,N_15990,N_15859);
or U16113 (N_16113,N_15988,N_15846);
nor U16114 (N_16114,N_15953,N_15866);
and U16115 (N_16115,N_15895,N_15972);
or U16116 (N_16116,N_15989,N_15969);
and U16117 (N_16117,N_15858,N_15846);
nand U16118 (N_16118,N_15940,N_15935);
nor U16119 (N_16119,N_15857,N_15969);
or U16120 (N_16120,N_15873,N_15912);
xnor U16121 (N_16121,N_15976,N_15953);
and U16122 (N_16122,N_15975,N_15878);
nand U16123 (N_16123,N_15962,N_15840);
or U16124 (N_16124,N_15901,N_15851);
and U16125 (N_16125,N_15909,N_15959);
or U16126 (N_16126,N_15875,N_15999);
or U16127 (N_16127,N_15867,N_15998);
and U16128 (N_16128,N_15973,N_15842);
nor U16129 (N_16129,N_15953,N_15942);
xnor U16130 (N_16130,N_15907,N_15996);
or U16131 (N_16131,N_15911,N_15940);
xor U16132 (N_16132,N_15953,N_15885);
nand U16133 (N_16133,N_15869,N_15947);
nor U16134 (N_16134,N_15848,N_15865);
nor U16135 (N_16135,N_15985,N_15907);
xor U16136 (N_16136,N_15955,N_15852);
nand U16137 (N_16137,N_15866,N_15939);
nor U16138 (N_16138,N_15948,N_15922);
or U16139 (N_16139,N_15942,N_15908);
or U16140 (N_16140,N_15913,N_15969);
nor U16141 (N_16141,N_15892,N_15851);
nor U16142 (N_16142,N_15996,N_15902);
and U16143 (N_16143,N_15855,N_15921);
or U16144 (N_16144,N_15991,N_15957);
or U16145 (N_16145,N_15857,N_15890);
nand U16146 (N_16146,N_15904,N_15947);
and U16147 (N_16147,N_15845,N_15927);
nor U16148 (N_16148,N_15938,N_15874);
and U16149 (N_16149,N_15962,N_15952);
and U16150 (N_16150,N_15988,N_15969);
or U16151 (N_16151,N_15904,N_15903);
or U16152 (N_16152,N_15922,N_15981);
nand U16153 (N_16153,N_15845,N_15990);
nand U16154 (N_16154,N_15972,N_15894);
or U16155 (N_16155,N_15878,N_15912);
nand U16156 (N_16156,N_15930,N_15902);
nor U16157 (N_16157,N_15948,N_15859);
and U16158 (N_16158,N_15999,N_15874);
nor U16159 (N_16159,N_15957,N_15874);
or U16160 (N_16160,N_16047,N_16053);
or U16161 (N_16161,N_16025,N_16040);
or U16162 (N_16162,N_16064,N_16084);
nor U16163 (N_16163,N_16097,N_16016);
nand U16164 (N_16164,N_16130,N_16145);
nand U16165 (N_16165,N_16140,N_16103);
xnor U16166 (N_16166,N_16095,N_16079);
nand U16167 (N_16167,N_16135,N_16033);
nand U16168 (N_16168,N_16002,N_16106);
nor U16169 (N_16169,N_16061,N_16132);
nand U16170 (N_16170,N_16147,N_16155);
nor U16171 (N_16171,N_16031,N_16077);
nand U16172 (N_16172,N_16128,N_16159);
and U16173 (N_16173,N_16112,N_16066);
nor U16174 (N_16174,N_16035,N_16022);
and U16175 (N_16175,N_16076,N_16050);
nor U16176 (N_16176,N_16003,N_16104);
and U16177 (N_16177,N_16117,N_16131);
xnor U16178 (N_16178,N_16152,N_16083);
xnor U16179 (N_16179,N_16052,N_16063);
nor U16180 (N_16180,N_16120,N_16094);
nand U16181 (N_16181,N_16071,N_16006);
or U16182 (N_16182,N_16013,N_16150);
xnor U16183 (N_16183,N_16100,N_16073);
and U16184 (N_16184,N_16124,N_16027);
nor U16185 (N_16185,N_16093,N_16090);
and U16186 (N_16186,N_16107,N_16099);
or U16187 (N_16187,N_16048,N_16138);
and U16188 (N_16188,N_16115,N_16113);
nor U16189 (N_16189,N_16001,N_16024);
xor U16190 (N_16190,N_16123,N_16109);
nor U16191 (N_16191,N_16062,N_16039);
nand U16192 (N_16192,N_16129,N_16000);
or U16193 (N_16193,N_16044,N_16059);
nor U16194 (N_16194,N_16085,N_16142);
xor U16195 (N_16195,N_16055,N_16056);
nor U16196 (N_16196,N_16037,N_16070);
nand U16197 (N_16197,N_16060,N_16051);
nor U16198 (N_16198,N_16008,N_16080);
or U16199 (N_16199,N_16043,N_16004);
and U16200 (N_16200,N_16139,N_16127);
and U16201 (N_16201,N_16072,N_16032);
nor U16202 (N_16202,N_16082,N_16143);
nand U16203 (N_16203,N_16089,N_16137);
nand U16204 (N_16204,N_16116,N_16023);
nand U16205 (N_16205,N_16122,N_16111);
nand U16206 (N_16206,N_16098,N_16007);
xnor U16207 (N_16207,N_16049,N_16021);
and U16208 (N_16208,N_16058,N_16102);
nor U16209 (N_16209,N_16126,N_16042);
nor U16210 (N_16210,N_16019,N_16069);
nand U16211 (N_16211,N_16038,N_16157);
nand U16212 (N_16212,N_16028,N_16154);
nand U16213 (N_16213,N_16088,N_16156);
xnor U16214 (N_16214,N_16018,N_16141);
and U16215 (N_16215,N_16148,N_16012);
xor U16216 (N_16216,N_16092,N_16054);
and U16217 (N_16217,N_16105,N_16119);
xor U16218 (N_16218,N_16087,N_16121);
nor U16219 (N_16219,N_16034,N_16014);
nand U16220 (N_16220,N_16026,N_16010);
nor U16221 (N_16221,N_16136,N_16005);
and U16222 (N_16222,N_16015,N_16114);
and U16223 (N_16223,N_16153,N_16118);
or U16224 (N_16224,N_16101,N_16057);
nor U16225 (N_16225,N_16075,N_16068);
nor U16226 (N_16226,N_16133,N_16067);
and U16227 (N_16227,N_16017,N_16096);
nor U16228 (N_16228,N_16065,N_16046);
or U16229 (N_16229,N_16151,N_16078);
xnor U16230 (N_16230,N_16108,N_16036);
or U16231 (N_16231,N_16029,N_16149);
nand U16232 (N_16232,N_16158,N_16081);
nand U16233 (N_16233,N_16110,N_16020);
and U16234 (N_16234,N_16144,N_16009);
xor U16235 (N_16235,N_16146,N_16091);
xor U16236 (N_16236,N_16134,N_16045);
nor U16237 (N_16237,N_16011,N_16041);
nor U16238 (N_16238,N_16125,N_16086);
xor U16239 (N_16239,N_16030,N_16074);
and U16240 (N_16240,N_16109,N_16048);
nand U16241 (N_16241,N_16119,N_16071);
nor U16242 (N_16242,N_16126,N_16045);
nor U16243 (N_16243,N_16086,N_16107);
and U16244 (N_16244,N_16111,N_16025);
and U16245 (N_16245,N_16069,N_16143);
nand U16246 (N_16246,N_16125,N_16100);
nand U16247 (N_16247,N_16021,N_16064);
nand U16248 (N_16248,N_16116,N_16035);
or U16249 (N_16249,N_16006,N_16122);
nand U16250 (N_16250,N_16133,N_16024);
nor U16251 (N_16251,N_16040,N_16010);
nor U16252 (N_16252,N_16020,N_16007);
nor U16253 (N_16253,N_16000,N_16124);
and U16254 (N_16254,N_16147,N_16135);
and U16255 (N_16255,N_16114,N_16112);
nand U16256 (N_16256,N_16057,N_16142);
nand U16257 (N_16257,N_16111,N_16074);
or U16258 (N_16258,N_16085,N_16006);
or U16259 (N_16259,N_16093,N_16020);
and U16260 (N_16260,N_16094,N_16088);
xnor U16261 (N_16261,N_16082,N_16066);
nor U16262 (N_16262,N_16021,N_16092);
or U16263 (N_16263,N_16021,N_16038);
nand U16264 (N_16264,N_16126,N_16153);
or U16265 (N_16265,N_16005,N_16125);
or U16266 (N_16266,N_16069,N_16114);
nand U16267 (N_16267,N_16076,N_16038);
nand U16268 (N_16268,N_16020,N_16129);
and U16269 (N_16269,N_16050,N_16044);
nor U16270 (N_16270,N_16065,N_16092);
and U16271 (N_16271,N_16041,N_16002);
nand U16272 (N_16272,N_16065,N_16014);
nand U16273 (N_16273,N_16148,N_16022);
nand U16274 (N_16274,N_16137,N_16007);
nor U16275 (N_16275,N_16075,N_16000);
nand U16276 (N_16276,N_16055,N_16131);
xor U16277 (N_16277,N_16048,N_16088);
and U16278 (N_16278,N_16075,N_16132);
or U16279 (N_16279,N_16016,N_16147);
nand U16280 (N_16280,N_16046,N_16077);
xor U16281 (N_16281,N_16055,N_16127);
nor U16282 (N_16282,N_16070,N_16105);
and U16283 (N_16283,N_16028,N_16032);
or U16284 (N_16284,N_16029,N_16101);
and U16285 (N_16285,N_16126,N_16068);
or U16286 (N_16286,N_16141,N_16010);
or U16287 (N_16287,N_16156,N_16030);
or U16288 (N_16288,N_16095,N_16055);
nand U16289 (N_16289,N_16112,N_16032);
or U16290 (N_16290,N_16079,N_16154);
nor U16291 (N_16291,N_16025,N_16090);
nor U16292 (N_16292,N_16048,N_16120);
nand U16293 (N_16293,N_16067,N_16088);
nand U16294 (N_16294,N_16128,N_16068);
and U16295 (N_16295,N_16127,N_16134);
xnor U16296 (N_16296,N_16105,N_16020);
nor U16297 (N_16297,N_16007,N_16121);
and U16298 (N_16298,N_16028,N_16027);
nor U16299 (N_16299,N_16129,N_16082);
nand U16300 (N_16300,N_16076,N_16051);
nand U16301 (N_16301,N_16013,N_16005);
nand U16302 (N_16302,N_16063,N_16131);
xor U16303 (N_16303,N_16114,N_16019);
and U16304 (N_16304,N_16108,N_16001);
and U16305 (N_16305,N_16001,N_16021);
nor U16306 (N_16306,N_16068,N_16078);
and U16307 (N_16307,N_16089,N_16019);
nor U16308 (N_16308,N_16131,N_16104);
nand U16309 (N_16309,N_16068,N_16026);
or U16310 (N_16310,N_16080,N_16140);
or U16311 (N_16311,N_16140,N_16130);
nand U16312 (N_16312,N_16065,N_16035);
nor U16313 (N_16313,N_16049,N_16034);
xor U16314 (N_16314,N_16010,N_16004);
or U16315 (N_16315,N_16007,N_16132);
nor U16316 (N_16316,N_16095,N_16086);
nand U16317 (N_16317,N_16157,N_16069);
nand U16318 (N_16318,N_16017,N_16149);
and U16319 (N_16319,N_16046,N_16097);
and U16320 (N_16320,N_16176,N_16313);
nand U16321 (N_16321,N_16312,N_16249);
and U16322 (N_16322,N_16229,N_16277);
or U16323 (N_16323,N_16258,N_16263);
nor U16324 (N_16324,N_16193,N_16292);
nor U16325 (N_16325,N_16311,N_16185);
xnor U16326 (N_16326,N_16280,N_16242);
xor U16327 (N_16327,N_16167,N_16170);
and U16328 (N_16328,N_16272,N_16265);
nor U16329 (N_16329,N_16212,N_16214);
nor U16330 (N_16330,N_16243,N_16178);
nor U16331 (N_16331,N_16279,N_16255);
nand U16332 (N_16332,N_16296,N_16215);
and U16333 (N_16333,N_16166,N_16217);
and U16334 (N_16334,N_16276,N_16218);
or U16335 (N_16335,N_16213,N_16239);
nor U16336 (N_16336,N_16284,N_16168);
nor U16337 (N_16337,N_16269,N_16233);
xnor U16338 (N_16338,N_16278,N_16188);
nand U16339 (N_16339,N_16304,N_16308);
nor U16340 (N_16340,N_16161,N_16283);
and U16341 (N_16341,N_16226,N_16175);
nor U16342 (N_16342,N_16262,N_16171);
nand U16343 (N_16343,N_16319,N_16191);
and U16344 (N_16344,N_16285,N_16240);
xnor U16345 (N_16345,N_16268,N_16232);
or U16346 (N_16346,N_16247,N_16180);
or U16347 (N_16347,N_16246,N_16264);
or U16348 (N_16348,N_16256,N_16172);
xor U16349 (N_16349,N_16164,N_16295);
or U16350 (N_16350,N_16202,N_16160);
nor U16351 (N_16351,N_16190,N_16184);
xor U16352 (N_16352,N_16236,N_16182);
xor U16353 (N_16353,N_16298,N_16209);
nand U16354 (N_16354,N_16241,N_16219);
or U16355 (N_16355,N_16222,N_16231);
or U16356 (N_16356,N_16315,N_16261);
nor U16357 (N_16357,N_16199,N_16316);
nand U16358 (N_16358,N_16225,N_16197);
nand U16359 (N_16359,N_16299,N_16252);
nor U16360 (N_16360,N_16305,N_16196);
xnor U16361 (N_16361,N_16221,N_16189);
nor U16362 (N_16362,N_16216,N_16192);
or U16363 (N_16363,N_16287,N_16210);
nand U16364 (N_16364,N_16244,N_16303);
or U16365 (N_16365,N_16302,N_16201);
and U16366 (N_16366,N_16179,N_16310);
and U16367 (N_16367,N_16248,N_16165);
nor U16368 (N_16368,N_16301,N_16254);
nand U16369 (N_16369,N_16275,N_16318);
nor U16370 (N_16370,N_16223,N_16317);
nand U16371 (N_16371,N_16286,N_16220);
and U16372 (N_16372,N_16297,N_16174);
or U16373 (N_16373,N_16200,N_16314);
and U16374 (N_16374,N_16273,N_16224);
or U16375 (N_16375,N_16194,N_16234);
or U16376 (N_16376,N_16274,N_16228);
or U16377 (N_16377,N_16290,N_16187);
nor U16378 (N_16378,N_16245,N_16183);
and U16379 (N_16379,N_16260,N_16207);
nand U16380 (N_16380,N_16250,N_16204);
or U16381 (N_16381,N_16208,N_16294);
nand U16382 (N_16382,N_16235,N_16181);
nand U16383 (N_16383,N_16253,N_16230);
or U16384 (N_16384,N_16169,N_16195);
or U16385 (N_16385,N_16266,N_16281);
nand U16386 (N_16386,N_16238,N_16309);
nand U16387 (N_16387,N_16206,N_16282);
nand U16388 (N_16388,N_16162,N_16306);
nor U16389 (N_16389,N_16177,N_16205);
or U16390 (N_16390,N_16257,N_16271);
nand U16391 (N_16391,N_16307,N_16291);
and U16392 (N_16392,N_16300,N_16251);
or U16393 (N_16393,N_16270,N_16288);
nor U16394 (N_16394,N_16163,N_16186);
and U16395 (N_16395,N_16173,N_16289);
xor U16396 (N_16396,N_16259,N_16227);
and U16397 (N_16397,N_16211,N_16293);
xor U16398 (N_16398,N_16203,N_16237);
xor U16399 (N_16399,N_16198,N_16267);
nand U16400 (N_16400,N_16171,N_16280);
or U16401 (N_16401,N_16258,N_16183);
or U16402 (N_16402,N_16221,N_16312);
nor U16403 (N_16403,N_16246,N_16279);
or U16404 (N_16404,N_16256,N_16210);
nor U16405 (N_16405,N_16251,N_16175);
nand U16406 (N_16406,N_16162,N_16297);
or U16407 (N_16407,N_16315,N_16193);
or U16408 (N_16408,N_16209,N_16197);
nor U16409 (N_16409,N_16269,N_16225);
or U16410 (N_16410,N_16173,N_16304);
nor U16411 (N_16411,N_16173,N_16195);
and U16412 (N_16412,N_16182,N_16243);
nand U16413 (N_16413,N_16208,N_16315);
nor U16414 (N_16414,N_16172,N_16233);
or U16415 (N_16415,N_16166,N_16231);
nand U16416 (N_16416,N_16203,N_16195);
nor U16417 (N_16417,N_16296,N_16277);
and U16418 (N_16418,N_16179,N_16170);
nor U16419 (N_16419,N_16319,N_16296);
and U16420 (N_16420,N_16219,N_16216);
nand U16421 (N_16421,N_16162,N_16171);
nand U16422 (N_16422,N_16282,N_16232);
or U16423 (N_16423,N_16265,N_16171);
or U16424 (N_16424,N_16316,N_16194);
or U16425 (N_16425,N_16197,N_16302);
nand U16426 (N_16426,N_16293,N_16180);
xor U16427 (N_16427,N_16237,N_16251);
and U16428 (N_16428,N_16238,N_16174);
and U16429 (N_16429,N_16211,N_16280);
nand U16430 (N_16430,N_16238,N_16285);
or U16431 (N_16431,N_16223,N_16228);
or U16432 (N_16432,N_16206,N_16311);
and U16433 (N_16433,N_16262,N_16183);
or U16434 (N_16434,N_16269,N_16273);
and U16435 (N_16435,N_16199,N_16318);
xor U16436 (N_16436,N_16273,N_16286);
nand U16437 (N_16437,N_16238,N_16292);
or U16438 (N_16438,N_16180,N_16272);
nand U16439 (N_16439,N_16183,N_16275);
or U16440 (N_16440,N_16170,N_16191);
and U16441 (N_16441,N_16185,N_16247);
nand U16442 (N_16442,N_16269,N_16305);
nand U16443 (N_16443,N_16302,N_16307);
and U16444 (N_16444,N_16232,N_16318);
and U16445 (N_16445,N_16181,N_16275);
nor U16446 (N_16446,N_16163,N_16250);
and U16447 (N_16447,N_16309,N_16283);
xor U16448 (N_16448,N_16181,N_16266);
nand U16449 (N_16449,N_16219,N_16195);
nand U16450 (N_16450,N_16175,N_16309);
nand U16451 (N_16451,N_16297,N_16277);
or U16452 (N_16452,N_16230,N_16217);
nand U16453 (N_16453,N_16201,N_16297);
nor U16454 (N_16454,N_16235,N_16245);
and U16455 (N_16455,N_16205,N_16226);
nor U16456 (N_16456,N_16173,N_16250);
and U16457 (N_16457,N_16286,N_16165);
xnor U16458 (N_16458,N_16195,N_16287);
nor U16459 (N_16459,N_16245,N_16264);
nand U16460 (N_16460,N_16280,N_16227);
xor U16461 (N_16461,N_16225,N_16220);
or U16462 (N_16462,N_16315,N_16226);
and U16463 (N_16463,N_16281,N_16230);
xnor U16464 (N_16464,N_16307,N_16219);
or U16465 (N_16465,N_16316,N_16253);
or U16466 (N_16466,N_16251,N_16278);
nor U16467 (N_16467,N_16164,N_16311);
or U16468 (N_16468,N_16219,N_16259);
and U16469 (N_16469,N_16174,N_16189);
nor U16470 (N_16470,N_16251,N_16182);
or U16471 (N_16471,N_16167,N_16194);
and U16472 (N_16472,N_16281,N_16313);
nor U16473 (N_16473,N_16228,N_16185);
nand U16474 (N_16474,N_16296,N_16307);
nand U16475 (N_16475,N_16191,N_16244);
nor U16476 (N_16476,N_16234,N_16160);
or U16477 (N_16477,N_16176,N_16232);
nor U16478 (N_16478,N_16266,N_16166);
xor U16479 (N_16479,N_16167,N_16204);
xor U16480 (N_16480,N_16321,N_16394);
xnor U16481 (N_16481,N_16343,N_16449);
xor U16482 (N_16482,N_16337,N_16406);
and U16483 (N_16483,N_16456,N_16465);
nor U16484 (N_16484,N_16470,N_16435);
nand U16485 (N_16485,N_16458,N_16364);
or U16486 (N_16486,N_16440,N_16373);
xnor U16487 (N_16487,N_16341,N_16357);
nor U16488 (N_16488,N_16415,N_16381);
and U16489 (N_16489,N_16374,N_16332);
nor U16490 (N_16490,N_16395,N_16388);
and U16491 (N_16491,N_16427,N_16410);
nor U16492 (N_16492,N_16428,N_16399);
nor U16493 (N_16493,N_16407,N_16416);
nor U16494 (N_16494,N_16359,N_16353);
and U16495 (N_16495,N_16354,N_16418);
nor U16496 (N_16496,N_16433,N_16461);
or U16497 (N_16497,N_16400,N_16366);
nand U16498 (N_16498,N_16442,N_16454);
nand U16499 (N_16499,N_16447,N_16405);
nand U16500 (N_16500,N_16367,N_16463);
nand U16501 (N_16501,N_16347,N_16370);
nand U16502 (N_16502,N_16385,N_16396);
nor U16503 (N_16503,N_16460,N_16426);
and U16504 (N_16504,N_16437,N_16393);
or U16505 (N_16505,N_16387,N_16469);
nand U16506 (N_16506,N_16327,N_16372);
and U16507 (N_16507,N_16386,N_16355);
xor U16508 (N_16508,N_16464,N_16349);
or U16509 (N_16509,N_16430,N_16363);
xnor U16510 (N_16510,N_16345,N_16352);
or U16511 (N_16511,N_16320,N_16339);
nor U16512 (N_16512,N_16451,N_16412);
nand U16513 (N_16513,N_16338,N_16422);
and U16514 (N_16514,N_16326,N_16323);
and U16515 (N_16515,N_16423,N_16446);
and U16516 (N_16516,N_16436,N_16474);
or U16517 (N_16517,N_16360,N_16403);
or U16518 (N_16518,N_16476,N_16398);
nand U16519 (N_16519,N_16478,N_16466);
nor U16520 (N_16520,N_16467,N_16331);
and U16521 (N_16521,N_16335,N_16455);
nor U16522 (N_16522,N_16375,N_16356);
or U16523 (N_16523,N_16429,N_16450);
and U16524 (N_16524,N_16452,N_16425);
nor U16525 (N_16525,N_16419,N_16325);
and U16526 (N_16526,N_16340,N_16471);
and U16527 (N_16527,N_16457,N_16330);
nor U16528 (N_16528,N_16424,N_16444);
or U16529 (N_16529,N_16417,N_16333);
nand U16530 (N_16530,N_16365,N_16358);
nor U16531 (N_16531,N_16477,N_16409);
or U16532 (N_16532,N_16390,N_16351);
xnor U16533 (N_16533,N_16408,N_16434);
or U16534 (N_16534,N_16329,N_16371);
nor U16535 (N_16535,N_16443,N_16342);
nor U16536 (N_16536,N_16378,N_16380);
and U16537 (N_16537,N_16379,N_16346);
and U16538 (N_16538,N_16384,N_16413);
or U16539 (N_16539,N_16441,N_16397);
xnor U16540 (N_16540,N_16453,N_16392);
nand U16541 (N_16541,N_16391,N_16383);
nor U16542 (N_16542,N_16377,N_16445);
xnor U16543 (N_16543,N_16344,N_16350);
or U16544 (N_16544,N_16431,N_16448);
and U16545 (N_16545,N_16336,N_16414);
nor U16546 (N_16546,N_16401,N_16362);
nor U16547 (N_16547,N_16376,N_16473);
or U16548 (N_16548,N_16472,N_16382);
nor U16549 (N_16549,N_16475,N_16361);
and U16550 (N_16550,N_16328,N_16420);
and U16551 (N_16551,N_16322,N_16411);
xor U16552 (N_16552,N_16404,N_16468);
nand U16553 (N_16553,N_16348,N_16389);
or U16554 (N_16554,N_16432,N_16439);
nand U16555 (N_16555,N_16459,N_16479);
and U16556 (N_16556,N_16369,N_16462);
nand U16557 (N_16557,N_16438,N_16421);
and U16558 (N_16558,N_16324,N_16334);
nor U16559 (N_16559,N_16368,N_16402);
or U16560 (N_16560,N_16431,N_16454);
or U16561 (N_16561,N_16375,N_16357);
and U16562 (N_16562,N_16397,N_16429);
nand U16563 (N_16563,N_16368,N_16354);
nor U16564 (N_16564,N_16399,N_16411);
nor U16565 (N_16565,N_16324,N_16476);
or U16566 (N_16566,N_16368,N_16344);
xnor U16567 (N_16567,N_16408,N_16322);
or U16568 (N_16568,N_16321,N_16389);
or U16569 (N_16569,N_16406,N_16354);
nor U16570 (N_16570,N_16389,N_16454);
nor U16571 (N_16571,N_16397,N_16423);
xnor U16572 (N_16572,N_16444,N_16328);
nand U16573 (N_16573,N_16467,N_16321);
nor U16574 (N_16574,N_16345,N_16338);
or U16575 (N_16575,N_16332,N_16350);
and U16576 (N_16576,N_16425,N_16380);
nor U16577 (N_16577,N_16413,N_16320);
nor U16578 (N_16578,N_16420,N_16474);
nor U16579 (N_16579,N_16323,N_16346);
nand U16580 (N_16580,N_16388,N_16471);
or U16581 (N_16581,N_16341,N_16438);
nand U16582 (N_16582,N_16465,N_16326);
nor U16583 (N_16583,N_16330,N_16325);
nand U16584 (N_16584,N_16472,N_16415);
nor U16585 (N_16585,N_16394,N_16349);
or U16586 (N_16586,N_16461,N_16457);
or U16587 (N_16587,N_16437,N_16422);
nor U16588 (N_16588,N_16415,N_16349);
or U16589 (N_16589,N_16333,N_16372);
nor U16590 (N_16590,N_16380,N_16459);
nand U16591 (N_16591,N_16473,N_16324);
and U16592 (N_16592,N_16473,N_16452);
nand U16593 (N_16593,N_16453,N_16401);
and U16594 (N_16594,N_16406,N_16383);
and U16595 (N_16595,N_16379,N_16416);
or U16596 (N_16596,N_16443,N_16429);
nor U16597 (N_16597,N_16470,N_16393);
and U16598 (N_16598,N_16378,N_16400);
nor U16599 (N_16599,N_16464,N_16338);
xor U16600 (N_16600,N_16442,N_16440);
and U16601 (N_16601,N_16410,N_16423);
nand U16602 (N_16602,N_16395,N_16347);
nand U16603 (N_16603,N_16368,N_16439);
and U16604 (N_16604,N_16448,N_16336);
and U16605 (N_16605,N_16412,N_16421);
nand U16606 (N_16606,N_16449,N_16425);
nand U16607 (N_16607,N_16448,N_16357);
nor U16608 (N_16608,N_16336,N_16438);
nand U16609 (N_16609,N_16366,N_16410);
nor U16610 (N_16610,N_16465,N_16392);
nor U16611 (N_16611,N_16394,N_16449);
and U16612 (N_16612,N_16470,N_16431);
or U16613 (N_16613,N_16355,N_16365);
or U16614 (N_16614,N_16344,N_16425);
nor U16615 (N_16615,N_16449,N_16422);
xnor U16616 (N_16616,N_16347,N_16354);
nand U16617 (N_16617,N_16349,N_16396);
or U16618 (N_16618,N_16477,N_16439);
nand U16619 (N_16619,N_16437,N_16334);
nor U16620 (N_16620,N_16469,N_16403);
nand U16621 (N_16621,N_16390,N_16471);
or U16622 (N_16622,N_16406,N_16379);
or U16623 (N_16623,N_16379,N_16380);
and U16624 (N_16624,N_16459,N_16355);
nor U16625 (N_16625,N_16407,N_16414);
nor U16626 (N_16626,N_16341,N_16476);
nor U16627 (N_16627,N_16450,N_16417);
or U16628 (N_16628,N_16383,N_16476);
and U16629 (N_16629,N_16369,N_16441);
nand U16630 (N_16630,N_16473,N_16343);
and U16631 (N_16631,N_16327,N_16361);
nand U16632 (N_16632,N_16349,N_16472);
or U16633 (N_16633,N_16382,N_16388);
xor U16634 (N_16634,N_16346,N_16471);
or U16635 (N_16635,N_16417,N_16330);
or U16636 (N_16636,N_16329,N_16445);
xor U16637 (N_16637,N_16408,N_16417);
or U16638 (N_16638,N_16378,N_16327);
or U16639 (N_16639,N_16416,N_16364);
and U16640 (N_16640,N_16504,N_16492);
and U16641 (N_16641,N_16587,N_16496);
or U16642 (N_16642,N_16500,N_16532);
nand U16643 (N_16643,N_16602,N_16635);
and U16644 (N_16644,N_16488,N_16483);
or U16645 (N_16645,N_16534,N_16499);
nor U16646 (N_16646,N_16540,N_16491);
nor U16647 (N_16647,N_16618,N_16634);
or U16648 (N_16648,N_16579,N_16538);
and U16649 (N_16649,N_16510,N_16511);
nor U16650 (N_16650,N_16622,N_16633);
or U16651 (N_16651,N_16523,N_16495);
and U16652 (N_16652,N_16599,N_16531);
nand U16653 (N_16653,N_16509,N_16636);
nand U16654 (N_16654,N_16551,N_16616);
or U16655 (N_16655,N_16555,N_16588);
and U16656 (N_16656,N_16596,N_16512);
nor U16657 (N_16657,N_16580,N_16563);
nor U16658 (N_16658,N_16608,N_16506);
nand U16659 (N_16659,N_16581,N_16620);
or U16660 (N_16660,N_16583,N_16582);
or U16661 (N_16661,N_16543,N_16522);
and U16662 (N_16662,N_16525,N_16586);
nand U16663 (N_16663,N_16574,N_16627);
and U16664 (N_16664,N_16626,N_16550);
or U16665 (N_16665,N_16520,N_16560);
nand U16666 (N_16666,N_16535,N_16613);
xor U16667 (N_16667,N_16536,N_16546);
nand U16668 (N_16668,N_16497,N_16612);
nor U16669 (N_16669,N_16548,N_16585);
nand U16670 (N_16670,N_16569,N_16524);
and U16671 (N_16671,N_16570,N_16562);
and U16672 (N_16672,N_16516,N_16528);
nor U16673 (N_16673,N_16621,N_16566);
and U16674 (N_16674,N_16625,N_16513);
nor U16675 (N_16675,N_16486,N_16515);
nor U16676 (N_16676,N_16481,N_16578);
xnor U16677 (N_16677,N_16615,N_16494);
xor U16678 (N_16678,N_16552,N_16617);
nor U16679 (N_16679,N_16607,N_16600);
and U16680 (N_16680,N_16558,N_16565);
and U16681 (N_16681,N_16561,N_16632);
or U16682 (N_16682,N_16556,N_16482);
nand U16683 (N_16683,N_16553,N_16572);
nor U16684 (N_16684,N_16614,N_16573);
or U16685 (N_16685,N_16539,N_16559);
nand U16686 (N_16686,N_16537,N_16639);
xor U16687 (N_16687,N_16624,N_16549);
or U16688 (N_16688,N_16601,N_16623);
nand U16689 (N_16689,N_16594,N_16489);
and U16690 (N_16690,N_16589,N_16518);
nand U16691 (N_16691,N_16530,N_16498);
nor U16692 (N_16692,N_16571,N_16493);
or U16693 (N_16693,N_16490,N_16557);
nand U16694 (N_16694,N_16629,N_16485);
nor U16695 (N_16695,N_16584,N_16541);
xor U16696 (N_16696,N_16598,N_16529);
or U16697 (N_16697,N_16568,N_16480);
or U16698 (N_16698,N_16544,N_16591);
or U16699 (N_16699,N_16637,N_16595);
nor U16700 (N_16700,N_16508,N_16619);
nor U16701 (N_16701,N_16577,N_16576);
and U16702 (N_16702,N_16567,N_16631);
and U16703 (N_16703,N_16606,N_16603);
and U16704 (N_16704,N_16597,N_16519);
nand U16705 (N_16705,N_16542,N_16638);
and U16706 (N_16706,N_16505,N_16604);
nand U16707 (N_16707,N_16592,N_16503);
or U16708 (N_16708,N_16609,N_16514);
nor U16709 (N_16709,N_16487,N_16554);
and U16710 (N_16710,N_16611,N_16564);
and U16711 (N_16711,N_16575,N_16517);
or U16712 (N_16712,N_16630,N_16610);
or U16713 (N_16713,N_16521,N_16527);
nand U16714 (N_16714,N_16590,N_16593);
nand U16715 (N_16715,N_16502,N_16605);
or U16716 (N_16716,N_16545,N_16547);
nor U16717 (N_16717,N_16533,N_16628);
nand U16718 (N_16718,N_16484,N_16501);
xnor U16719 (N_16719,N_16526,N_16507);
xor U16720 (N_16720,N_16489,N_16630);
nor U16721 (N_16721,N_16537,N_16593);
and U16722 (N_16722,N_16518,N_16523);
or U16723 (N_16723,N_16611,N_16490);
xor U16724 (N_16724,N_16548,N_16494);
and U16725 (N_16725,N_16610,N_16499);
nand U16726 (N_16726,N_16531,N_16549);
or U16727 (N_16727,N_16615,N_16568);
or U16728 (N_16728,N_16482,N_16501);
nor U16729 (N_16729,N_16606,N_16529);
xnor U16730 (N_16730,N_16513,N_16519);
nand U16731 (N_16731,N_16548,N_16580);
and U16732 (N_16732,N_16636,N_16525);
nand U16733 (N_16733,N_16551,N_16586);
nand U16734 (N_16734,N_16569,N_16615);
nor U16735 (N_16735,N_16518,N_16511);
and U16736 (N_16736,N_16491,N_16559);
nor U16737 (N_16737,N_16510,N_16598);
and U16738 (N_16738,N_16507,N_16618);
and U16739 (N_16739,N_16528,N_16548);
nor U16740 (N_16740,N_16635,N_16588);
nand U16741 (N_16741,N_16633,N_16498);
nor U16742 (N_16742,N_16638,N_16483);
nand U16743 (N_16743,N_16504,N_16611);
xnor U16744 (N_16744,N_16555,N_16610);
nand U16745 (N_16745,N_16514,N_16607);
xnor U16746 (N_16746,N_16528,N_16612);
nor U16747 (N_16747,N_16588,N_16606);
and U16748 (N_16748,N_16596,N_16540);
nand U16749 (N_16749,N_16561,N_16525);
or U16750 (N_16750,N_16520,N_16543);
or U16751 (N_16751,N_16481,N_16612);
nand U16752 (N_16752,N_16522,N_16619);
and U16753 (N_16753,N_16512,N_16598);
nor U16754 (N_16754,N_16628,N_16489);
nand U16755 (N_16755,N_16576,N_16625);
and U16756 (N_16756,N_16614,N_16613);
nand U16757 (N_16757,N_16598,N_16540);
and U16758 (N_16758,N_16565,N_16591);
or U16759 (N_16759,N_16623,N_16511);
or U16760 (N_16760,N_16534,N_16521);
nand U16761 (N_16761,N_16524,N_16499);
nor U16762 (N_16762,N_16582,N_16505);
or U16763 (N_16763,N_16509,N_16544);
nand U16764 (N_16764,N_16495,N_16502);
or U16765 (N_16765,N_16637,N_16612);
nor U16766 (N_16766,N_16541,N_16517);
or U16767 (N_16767,N_16568,N_16556);
nor U16768 (N_16768,N_16527,N_16601);
xor U16769 (N_16769,N_16579,N_16526);
nand U16770 (N_16770,N_16574,N_16580);
xor U16771 (N_16771,N_16491,N_16609);
nand U16772 (N_16772,N_16502,N_16576);
or U16773 (N_16773,N_16508,N_16614);
nor U16774 (N_16774,N_16501,N_16487);
nor U16775 (N_16775,N_16541,N_16497);
or U16776 (N_16776,N_16538,N_16488);
nand U16777 (N_16777,N_16615,N_16550);
nand U16778 (N_16778,N_16484,N_16579);
and U16779 (N_16779,N_16541,N_16605);
nor U16780 (N_16780,N_16493,N_16538);
nand U16781 (N_16781,N_16575,N_16556);
nand U16782 (N_16782,N_16601,N_16483);
or U16783 (N_16783,N_16522,N_16544);
nor U16784 (N_16784,N_16599,N_16548);
and U16785 (N_16785,N_16569,N_16612);
or U16786 (N_16786,N_16617,N_16598);
nand U16787 (N_16787,N_16561,N_16560);
nand U16788 (N_16788,N_16610,N_16504);
and U16789 (N_16789,N_16580,N_16485);
xnor U16790 (N_16790,N_16624,N_16599);
nand U16791 (N_16791,N_16607,N_16580);
or U16792 (N_16792,N_16490,N_16512);
and U16793 (N_16793,N_16486,N_16489);
and U16794 (N_16794,N_16601,N_16525);
or U16795 (N_16795,N_16522,N_16498);
or U16796 (N_16796,N_16565,N_16519);
nor U16797 (N_16797,N_16482,N_16522);
or U16798 (N_16798,N_16617,N_16495);
or U16799 (N_16799,N_16588,N_16590);
nand U16800 (N_16800,N_16731,N_16769);
nor U16801 (N_16801,N_16700,N_16724);
xor U16802 (N_16802,N_16685,N_16690);
nor U16803 (N_16803,N_16728,N_16721);
and U16804 (N_16804,N_16778,N_16739);
and U16805 (N_16805,N_16652,N_16710);
xnor U16806 (N_16806,N_16648,N_16668);
or U16807 (N_16807,N_16707,N_16665);
or U16808 (N_16808,N_16711,N_16705);
and U16809 (N_16809,N_16799,N_16781);
nand U16810 (N_16810,N_16744,N_16748);
nor U16811 (N_16811,N_16645,N_16672);
nor U16812 (N_16812,N_16697,N_16796);
and U16813 (N_16813,N_16791,N_16650);
nor U16814 (N_16814,N_16797,N_16725);
and U16815 (N_16815,N_16732,N_16755);
nor U16816 (N_16816,N_16747,N_16682);
nand U16817 (N_16817,N_16698,N_16674);
and U16818 (N_16818,N_16649,N_16688);
xnor U16819 (N_16819,N_16666,N_16681);
and U16820 (N_16820,N_16790,N_16751);
or U16821 (N_16821,N_16662,N_16771);
nor U16822 (N_16822,N_16702,N_16786);
nor U16823 (N_16823,N_16789,N_16741);
and U16824 (N_16824,N_16727,N_16699);
and U16825 (N_16825,N_16642,N_16746);
or U16826 (N_16826,N_16684,N_16706);
nand U16827 (N_16827,N_16743,N_16651);
or U16828 (N_16828,N_16678,N_16742);
xor U16829 (N_16829,N_16689,N_16780);
nor U16830 (N_16830,N_16709,N_16717);
nand U16831 (N_16831,N_16687,N_16693);
or U16832 (N_16832,N_16646,N_16695);
or U16833 (N_16833,N_16766,N_16659);
nor U16834 (N_16834,N_16712,N_16647);
nand U16835 (N_16835,N_16686,N_16641);
and U16836 (N_16836,N_16749,N_16692);
and U16837 (N_16837,N_16664,N_16798);
and U16838 (N_16838,N_16745,N_16701);
nand U16839 (N_16839,N_16777,N_16683);
nor U16840 (N_16840,N_16787,N_16752);
nor U16841 (N_16841,N_16644,N_16663);
nand U16842 (N_16842,N_16653,N_16696);
nor U16843 (N_16843,N_16736,N_16708);
or U16844 (N_16844,N_16680,N_16657);
nand U16845 (N_16845,N_16760,N_16735);
and U16846 (N_16846,N_16762,N_16714);
nor U16847 (N_16847,N_16753,N_16758);
and U16848 (N_16848,N_16793,N_16673);
or U16849 (N_16849,N_16726,N_16792);
xnor U16850 (N_16850,N_16694,N_16656);
or U16851 (N_16851,N_16738,N_16658);
nand U16852 (N_16852,N_16776,N_16661);
nor U16853 (N_16853,N_16754,N_16782);
or U16854 (N_16854,N_16655,N_16713);
nand U16855 (N_16855,N_16737,N_16654);
and U16856 (N_16856,N_16767,N_16764);
or U16857 (N_16857,N_16667,N_16733);
nor U16858 (N_16858,N_16643,N_16794);
nand U16859 (N_16859,N_16723,N_16772);
or U16860 (N_16860,N_16795,N_16761);
xor U16861 (N_16861,N_16722,N_16675);
and U16862 (N_16862,N_16750,N_16677);
nor U16863 (N_16863,N_16703,N_16757);
or U16864 (N_16864,N_16783,N_16779);
or U16865 (N_16865,N_16768,N_16670);
nand U16866 (N_16866,N_16729,N_16669);
and U16867 (N_16867,N_16774,N_16784);
nand U16868 (N_16868,N_16773,N_16679);
nor U16869 (N_16869,N_16734,N_16671);
or U16870 (N_16870,N_16676,N_16770);
nor U16871 (N_16871,N_16716,N_16756);
or U16872 (N_16872,N_16704,N_16730);
xnor U16873 (N_16873,N_16720,N_16740);
or U16874 (N_16874,N_16719,N_16718);
or U16875 (N_16875,N_16660,N_16691);
xnor U16876 (N_16876,N_16640,N_16785);
or U16877 (N_16877,N_16715,N_16765);
nand U16878 (N_16878,N_16775,N_16763);
xnor U16879 (N_16879,N_16759,N_16788);
and U16880 (N_16880,N_16762,N_16693);
or U16881 (N_16881,N_16706,N_16702);
or U16882 (N_16882,N_16644,N_16788);
or U16883 (N_16883,N_16657,N_16740);
and U16884 (N_16884,N_16767,N_16759);
nor U16885 (N_16885,N_16715,N_16669);
nor U16886 (N_16886,N_16772,N_16677);
or U16887 (N_16887,N_16709,N_16767);
or U16888 (N_16888,N_16711,N_16662);
or U16889 (N_16889,N_16798,N_16682);
xnor U16890 (N_16890,N_16676,N_16790);
nor U16891 (N_16891,N_16694,N_16674);
or U16892 (N_16892,N_16764,N_16651);
and U16893 (N_16893,N_16794,N_16788);
and U16894 (N_16894,N_16685,N_16671);
or U16895 (N_16895,N_16656,N_16710);
nor U16896 (N_16896,N_16723,N_16782);
and U16897 (N_16897,N_16693,N_16774);
and U16898 (N_16898,N_16655,N_16771);
xor U16899 (N_16899,N_16681,N_16661);
nor U16900 (N_16900,N_16776,N_16640);
nor U16901 (N_16901,N_16645,N_16678);
and U16902 (N_16902,N_16720,N_16733);
or U16903 (N_16903,N_16696,N_16716);
nand U16904 (N_16904,N_16742,N_16765);
nor U16905 (N_16905,N_16718,N_16756);
nor U16906 (N_16906,N_16646,N_16765);
or U16907 (N_16907,N_16749,N_16755);
or U16908 (N_16908,N_16799,N_16712);
xor U16909 (N_16909,N_16742,N_16731);
nor U16910 (N_16910,N_16790,N_16694);
and U16911 (N_16911,N_16641,N_16761);
or U16912 (N_16912,N_16766,N_16684);
nand U16913 (N_16913,N_16660,N_16743);
or U16914 (N_16914,N_16705,N_16792);
or U16915 (N_16915,N_16657,N_16719);
or U16916 (N_16916,N_16761,N_16648);
and U16917 (N_16917,N_16666,N_16693);
nand U16918 (N_16918,N_16664,N_16687);
or U16919 (N_16919,N_16799,N_16749);
nor U16920 (N_16920,N_16784,N_16702);
or U16921 (N_16921,N_16776,N_16775);
nor U16922 (N_16922,N_16761,N_16652);
xor U16923 (N_16923,N_16796,N_16795);
or U16924 (N_16924,N_16701,N_16744);
and U16925 (N_16925,N_16706,N_16738);
or U16926 (N_16926,N_16736,N_16672);
nor U16927 (N_16927,N_16761,N_16741);
or U16928 (N_16928,N_16649,N_16753);
or U16929 (N_16929,N_16698,N_16680);
and U16930 (N_16930,N_16732,N_16670);
and U16931 (N_16931,N_16709,N_16668);
nor U16932 (N_16932,N_16794,N_16701);
or U16933 (N_16933,N_16656,N_16707);
or U16934 (N_16934,N_16799,N_16650);
nand U16935 (N_16935,N_16770,N_16685);
or U16936 (N_16936,N_16737,N_16649);
nand U16937 (N_16937,N_16753,N_16734);
nand U16938 (N_16938,N_16640,N_16716);
xor U16939 (N_16939,N_16647,N_16662);
or U16940 (N_16940,N_16656,N_16734);
xnor U16941 (N_16941,N_16721,N_16714);
nand U16942 (N_16942,N_16695,N_16775);
nor U16943 (N_16943,N_16741,N_16767);
nand U16944 (N_16944,N_16799,N_16658);
and U16945 (N_16945,N_16782,N_16690);
and U16946 (N_16946,N_16769,N_16669);
or U16947 (N_16947,N_16716,N_16772);
or U16948 (N_16948,N_16730,N_16766);
or U16949 (N_16949,N_16754,N_16784);
and U16950 (N_16950,N_16699,N_16664);
and U16951 (N_16951,N_16760,N_16727);
or U16952 (N_16952,N_16742,N_16792);
nor U16953 (N_16953,N_16694,N_16728);
and U16954 (N_16954,N_16645,N_16719);
nand U16955 (N_16955,N_16779,N_16649);
and U16956 (N_16956,N_16701,N_16793);
xnor U16957 (N_16957,N_16746,N_16724);
and U16958 (N_16958,N_16705,N_16783);
or U16959 (N_16959,N_16708,N_16750);
nor U16960 (N_16960,N_16819,N_16816);
and U16961 (N_16961,N_16900,N_16871);
or U16962 (N_16962,N_16850,N_16897);
nand U16963 (N_16963,N_16863,N_16931);
and U16964 (N_16964,N_16864,N_16905);
and U16965 (N_16965,N_16946,N_16910);
nand U16966 (N_16966,N_16832,N_16930);
xor U16967 (N_16967,N_16913,N_16848);
xnor U16968 (N_16968,N_16861,N_16902);
nand U16969 (N_16969,N_16814,N_16909);
nand U16970 (N_16970,N_16903,N_16958);
or U16971 (N_16971,N_16918,N_16813);
or U16972 (N_16972,N_16840,N_16866);
and U16973 (N_16973,N_16880,N_16923);
or U16974 (N_16974,N_16851,N_16822);
and U16975 (N_16975,N_16956,N_16920);
and U16976 (N_16976,N_16800,N_16842);
nand U16977 (N_16977,N_16823,N_16833);
nor U16978 (N_16978,N_16839,N_16803);
or U16979 (N_16979,N_16928,N_16955);
and U16980 (N_16980,N_16815,N_16802);
nand U16981 (N_16981,N_16898,N_16937);
and U16982 (N_16982,N_16801,N_16887);
nor U16983 (N_16983,N_16890,N_16841);
or U16984 (N_16984,N_16907,N_16858);
nand U16985 (N_16985,N_16883,N_16872);
xnor U16986 (N_16986,N_16950,N_16860);
nand U16987 (N_16987,N_16896,N_16817);
nand U16988 (N_16988,N_16806,N_16856);
and U16989 (N_16989,N_16936,N_16825);
and U16990 (N_16990,N_16884,N_16885);
and U16991 (N_16991,N_16959,N_16886);
and U16992 (N_16992,N_16857,N_16915);
nor U16993 (N_16993,N_16895,N_16873);
nor U16994 (N_16994,N_16853,N_16854);
nand U16995 (N_16995,N_16874,N_16899);
nor U16996 (N_16996,N_16934,N_16855);
and U16997 (N_16997,N_16947,N_16843);
or U16998 (N_16998,N_16868,N_16809);
or U16999 (N_16999,N_16882,N_16919);
and U17000 (N_17000,N_16938,N_16827);
and U17001 (N_17001,N_16933,N_16881);
or U17002 (N_17002,N_16925,N_16835);
nor U17003 (N_17003,N_16894,N_16804);
or U17004 (N_17004,N_16929,N_16935);
and U17005 (N_17005,N_16875,N_16831);
or U17006 (N_17006,N_16888,N_16836);
or U17007 (N_17007,N_16939,N_16924);
nand U17008 (N_17008,N_16812,N_16943);
nor U17009 (N_17009,N_16807,N_16805);
or U17010 (N_17010,N_16844,N_16908);
xnor U17011 (N_17011,N_16945,N_16911);
or U17012 (N_17012,N_16838,N_16810);
nor U17013 (N_17013,N_16892,N_16824);
nand U17014 (N_17014,N_16942,N_16826);
or U17015 (N_17015,N_16852,N_16906);
nand U17016 (N_17016,N_16893,N_16921);
or U17017 (N_17017,N_16845,N_16837);
nor U17018 (N_17018,N_16876,N_16944);
nand U17019 (N_17019,N_16818,N_16889);
nor U17020 (N_17020,N_16834,N_16914);
nand U17021 (N_17021,N_16949,N_16828);
and U17022 (N_17022,N_16953,N_16859);
nor U17023 (N_17023,N_16829,N_16808);
nand U17024 (N_17024,N_16952,N_16901);
xor U17025 (N_17025,N_16951,N_16877);
nand U17026 (N_17026,N_16904,N_16932);
xor U17027 (N_17027,N_16917,N_16847);
and U17028 (N_17028,N_16957,N_16830);
nor U17029 (N_17029,N_16912,N_16846);
xor U17030 (N_17030,N_16879,N_16865);
and U17031 (N_17031,N_16878,N_16867);
nand U17032 (N_17032,N_16948,N_16849);
or U17033 (N_17033,N_16811,N_16940);
and U17034 (N_17034,N_16916,N_16941);
and U17035 (N_17035,N_16821,N_16870);
nand U17036 (N_17036,N_16869,N_16926);
and U17037 (N_17037,N_16891,N_16922);
xor U17038 (N_17038,N_16820,N_16862);
nor U17039 (N_17039,N_16954,N_16927);
nand U17040 (N_17040,N_16912,N_16856);
nor U17041 (N_17041,N_16886,N_16872);
or U17042 (N_17042,N_16880,N_16811);
nand U17043 (N_17043,N_16954,N_16841);
nand U17044 (N_17044,N_16902,N_16886);
or U17045 (N_17045,N_16906,N_16924);
nor U17046 (N_17046,N_16802,N_16868);
or U17047 (N_17047,N_16933,N_16831);
xnor U17048 (N_17048,N_16933,N_16943);
nand U17049 (N_17049,N_16923,N_16900);
nand U17050 (N_17050,N_16957,N_16834);
nor U17051 (N_17051,N_16959,N_16820);
or U17052 (N_17052,N_16822,N_16876);
or U17053 (N_17053,N_16933,N_16817);
nor U17054 (N_17054,N_16852,N_16909);
or U17055 (N_17055,N_16956,N_16855);
nand U17056 (N_17056,N_16827,N_16857);
and U17057 (N_17057,N_16895,N_16921);
nand U17058 (N_17058,N_16818,N_16948);
xor U17059 (N_17059,N_16887,N_16853);
nor U17060 (N_17060,N_16942,N_16929);
nand U17061 (N_17061,N_16811,N_16867);
nor U17062 (N_17062,N_16930,N_16833);
nand U17063 (N_17063,N_16818,N_16862);
and U17064 (N_17064,N_16907,N_16851);
xor U17065 (N_17065,N_16905,N_16844);
nand U17066 (N_17066,N_16846,N_16844);
nand U17067 (N_17067,N_16863,N_16892);
or U17068 (N_17068,N_16811,N_16910);
or U17069 (N_17069,N_16904,N_16925);
nand U17070 (N_17070,N_16828,N_16810);
or U17071 (N_17071,N_16840,N_16820);
and U17072 (N_17072,N_16822,N_16958);
nor U17073 (N_17073,N_16901,N_16802);
or U17074 (N_17074,N_16837,N_16947);
nor U17075 (N_17075,N_16844,N_16907);
and U17076 (N_17076,N_16938,N_16922);
or U17077 (N_17077,N_16899,N_16863);
and U17078 (N_17078,N_16917,N_16815);
or U17079 (N_17079,N_16866,N_16916);
nand U17080 (N_17080,N_16886,N_16932);
or U17081 (N_17081,N_16952,N_16854);
xor U17082 (N_17082,N_16851,N_16957);
and U17083 (N_17083,N_16812,N_16815);
nor U17084 (N_17084,N_16874,N_16945);
nor U17085 (N_17085,N_16924,N_16940);
xor U17086 (N_17086,N_16888,N_16904);
xnor U17087 (N_17087,N_16807,N_16912);
and U17088 (N_17088,N_16948,N_16906);
or U17089 (N_17089,N_16937,N_16809);
xor U17090 (N_17090,N_16849,N_16950);
nor U17091 (N_17091,N_16927,N_16905);
or U17092 (N_17092,N_16912,N_16900);
nor U17093 (N_17093,N_16916,N_16850);
xnor U17094 (N_17094,N_16872,N_16843);
and U17095 (N_17095,N_16918,N_16885);
or U17096 (N_17096,N_16804,N_16915);
and U17097 (N_17097,N_16806,N_16946);
nand U17098 (N_17098,N_16850,N_16813);
or U17099 (N_17099,N_16930,N_16910);
nand U17100 (N_17100,N_16937,N_16918);
or U17101 (N_17101,N_16957,N_16929);
or U17102 (N_17102,N_16826,N_16872);
or U17103 (N_17103,N_16883,N_16905);
and U17104 (N_17104,N_16927,N_16871);
and U17105 (N_17105,N_16867,N_16861);
nand U17106 (N_17106,N_16948,N_16926);
and U17107 (N_17107,N_16912,N_16830);
and U17108 (N_17108,N_16912,N_16920);
and U17109 (N_17109,N_16885,N_16836);
and U17110 (N_17110,N_16930,N_16849);
or U17111 (N_17111,N_16841,N_16848);
nor U17112 (N_17112,N_16801,N_16865);
nor U17113 (N_17113,N_16800,N_16870);
nor U17114 (N_17114,N_16844,N_16879);
xnor U17115 (N_17115,N_16872,N_16818);
nor U17116 (N_17116,N_16914,N_16956);
xor U17117 (N_17117,N_16883,N_16864);
xor U17118 (N_17118,N_16906,N_16811);
and U17119 (N_17119,N_16922,N_16832);
or U17120 (N_17120,N_17008,N_17087);
nor U17121 (N_17121,N_17015,N_17046);
nor U17122 (N_17122,N_16970,N_17029);
nor U17123 (N_17123,N_17055,N_17100);
and U17124 (N_17124,N_17118,N_17088);
or U17125 (N_17125,N_16961,N_17091);
or U17126 (N_17126,N_17076,N_17003);
and U17127 (N_17127,N_16978,N_17050);
nand U17128 (N_17128,N_16980,N_17107);
and U17129 (N_17129,N_16979,N_17057);
and U17130 (N_17130,N_17090,N_16987);
nor U17131 (N_17131,N_17052,N_16974);
nor U17132 (N_17132,N_17001,N_17020);
nor U17133 (N_17133,N_16976,N_17081);
nor U17134 (N_17134,N_17040,N_17064);
or U17135 (N_17135,N_16999,N_17025);
nand U17136 (N_17136,N_16986,N_17101);
xor U17137 (N_17137,N_17054,N_17075);
and U17138 (N_17138,N_17036,N_17000);
xnor U17139 (N_17139,N_17045,N_16994);
nand U17140 (N_17140,N_16992,N_16975);
xor U17141 (N_17141,N_17053,N_16966);
nor U17142 (N_17142,N_17115,N_17116);
and U17143 (N_17143,N_17037,N_16991);
or U17144 (N_17144,N_17086,N_17056);
nand U17145 (N_17145,N_17092,N_17093);
nor U17146 (N_17146,N_16981,N_17094);
nor U17147 (N_17147,N_17012,N_16985);
and U17148 (N_17148,N_17024,N_17005);
nand U17149 (N_17149,N_17074,N_17059);
nand U17150 (N_17150,N_17038,N_17080);
nor U17151 (N_17151,N_16960,N_17078);
or U17152 (N_17152,N_17109,N_17028);
nand U17153 (N_17153,N_16971,N_17060);
and U17154 (N_17154,N_17048,N_16996);
or U17155 (N_17155,N_16990,N_17103);
nand U17156 (N_17156,N_17097,N_17035);
xnor U17157 (N_17157,N_17049,N_17108);
nand U17158 (N_17158,N_16993,N_16983);
or U17159 (N_17159,N_17065,N_17070);
and U17160 (N_17160,N_17019,N_17102);
or U17161 (N_17161,N_17027,N_16965);
or U17162 (N_17162,N_17042,N_16995);
nand U17163 (N_17163,N_17009,N_16967);
or U17164 (N_17164,N_17017,N_16977);
nor U17165 (N_17165,N_17026,N_17018);
and U17166 (N_17166,N_17014,N_16962);
nor U17167 (N_17167,N_17111,N_17096);
nor U17168 (N_17168,N_17031,N_16989);
or U17169 (N_17169,N_17112,N_17072);
xor U17170 (N_17170,N_17061,N_17085);
and U17171 (N_17171,N_17066,N_17034);
nand U17172 (N_17172,N_17068,N_17002);
or U17173 (N_17173,N_17113,N_17004);
or U17174 (N_17174,N_17023,N_17106);
and U17175 (N_17175,N_16982,N_17069);
and U17176 (N_17176,N_16968,N_17083);
nor U17177 (N_17177,N_17006,N_17063);
xnor U17178 (N_17178,N_17117,N_17062);
and U17179 (N_17179,N_17013,N_17051);
nand U17180 (N_17180,N_16972,N_17105);
or U17181 (N_17181,N_17079,N_17098);
or U17182 (N_17182,N_17110,N_16997);
or U17183 (N_17183,N_16998,N_17099);
nor U17184 (N_17184,N_17043,N_17011);
or U17185 (N_17185,N_16988,N_16963);
and U17186 (N_17186,N_17033,N_17077);
nand U17187 (N_17187,N_17022,N_17021);
or U17188 (N_17188,N_17104,N_17032);
nor U17189 (N_17189,N_17073,N_17095);
nand U17190 (N_17190,N_17071,N_17007);
or U17191 (N_17191,N_16969,N_17044);
or U17192 (N_17192,N_17016,N_17058);
xnor U17193 (N_17193,N_16984,N_16973);
nand U17194 (N_17194,N_17089,N_17119);
nor U17195 (N_17195,N_17010,N_16964);
nor U17196 (N_17196,N_17082,N_17047);
nor U17197 (N_17197,N_17041,N_17084);
or U17198 (N_17198,N_17030,N_17067);
nor U17199 (N_17199,N_17039,N_17114);
nand U17200 (N_17200,N_17090,N_16974);
and U17201 (N_17201,N_16993,N_17047);
nand U17202 (N_17202,N_17076,N_17081);
and U17203 (N_17203,N_17034,N_17025);
nand U17204 (N_17204,N_17066,N_17007);
and U17205 (N_17205,N_16978,N_17119);
nand U17206 (N_17206,N_17074,N_17091);
xor U17207 (N_17207,N_17007,N_17076);
and U17208 (N_17208,N_17054,N_17046);
nor U17209 (N_17209,N_17097,N_17016);
or U17210 (N_17210,N_17052,N_17110);
nor U17211 (N_17211,N_17108,N_17078);
nand U17212 (N_17212,N_17090,N_17065);
and U17213 (N_17213,N_17090,N_16986);
xnor U17214 (N_17214,N_16976,N_16972);
and U17215 (N_17215,N_17004,N_17065);
xnor U17216 (N_17216,N_17010,N_17024);
nand U17217 (N_17217,N_17049,N_17040);
and U17218 (N_17218,N_17009,N_17025);
nor U17219 (N_17219,N_17109,N_17115);
and U17220 (N_17220,N_17025,N_17078);
and U17221 (N_17221,N_17059,N_16990);
nand U17222 (N_17222,N_17031,N_16979);
xnor U17223 (N_17223,N_17084,N_17018);
or U17224 (N_17224,N_17064,N_17022);
or U17225 (N_17225,N_17061,N_17007);
or U17226 (N_17226,N_16967,N_16979);
nand U17227 (N_17227,N_17044,N_17107);
nor U17228 (N_17228,N_17075,N_17034);
and U17229 (N_17229,N_17021,N_17055);
nand U17230 (N_17230,N_16960,N_17119);
nand U17231 (N_17231,N_17087,N_17038);
nand U17232 (N_17232,N_17107,N_16971);
nand U17233 (N_17233,N_17046,N_17071);
nand U17234 (N_17234,N_16966,N_16998);
and U17235 (N_17235,N_16970,N_17003);
or U17236 (N_17236,N_17013,N_17049);
or U17237 (N_17237,N_16988,N_17094);
or U17238 (N_17238,N_16974,N_17035);
xnor U17239 (N_17239,N_16972,N_16971);
nor U17240 (N_17240,N_17094,N_17002);
and U17241 (N_17241,N_17022,N_17003);
or U17242 (N_17242,N_16993,N_17038);
and U17243 (N_17243,N_16981,N_17059);
and U17244 (N_17244,N_17079,N_16972);
nand U17245 (N_17245,N_17025,N_17098);
and U17246 (N_17246,N_17087,N_16993);
nand U17247 (N_17247,N_17062,N_17098);
and U17248 (N_17248,N_17105,N_17016);
xnor U17249 (N_17249,N_17079,N_17027);
nand U17250 (N_17250,N_17038,N_17041);
nand U17251 (N_17251,N_17115,N_16976);
nand U17252 (N_17252,N_17066,N_17078);
and U17253 (N_17253,N_17068,N_17088);
nor U17254 (N_17254,N_17043,N_17084);
nor U17255 (N_17255,N_16966,N_17005);
and U17256 (N_17256,N_16972,N_17002);
and U17257 (N_17257,N_16968,N_17041);
xnor U17258 (N_17258,N_17108,N_16987);
nor U17259 (N_17259,N_17051,N_17004);
nand U17260 (N_17260,N_16979,N_17013);
nand U17261 (N_17261,N_16985,N_17053);
or U17262 (N_17262,N_17104,N_16982);
nor U17263 (N_17263,N_17105,N_17103);
nor U17264 (N_17264,N_17077,N_17030);
nor U17265 (N_17265,N_17094,N_17091);
and U17266 (N_17266,N_16979,N_17027);
nand U17267 (N_17267,N_17029,N_17067);
or U17268 (N_17268,N_17025,N_17115);
or U17269 (N_17269,N_17102,N_17090);
and U17270 (N_17270,N_17109,N_17031);
nand U17271 (N_17271,N_17032,N_17051);
or U17272 (N_17272,N_17091,N_17089);
nor U17273 (N_17273,N_17034,N_17023);
nor U17274 (N_17274,N_17057,N_16996);
and U17275 (N_17275,N_17109,N_17004);
and U17276 (N_17276,N_17111,N_17007);
xor U17277 (N_17277,N_16971,N_16964);
nand U17278 (N_17278,N_16991,N_17035);
nand U17279 (N_17279,N_17024,N_17105);
and U17280 (N_17280,N_17272,N_17258);
and U17281 (N_17281,N_17228,N_17191);
nor U17282 (N_17282,N_17160,N_17216);
and U17283 (N_17283,N_17208,N_17247);
xnor U17284 (N_17284,N_17224,N_17209);
nor U17285 (N_17285,N_17132,N_17193);
and U17286 (N_17286,N_17278,N_17225);
xnor U17287 (N_17287,N_17172,N_17215);
nor U17288 (N_17288,N_17157,N_17246);
and U17289 (N_17289,N_17138,N_17147);
nor U17290 (N_17290,N_17120,N_17148);
nor U17291 (N_17291,N_17190,N_17156);
and U17292 (N_17292,N_17170,N_17273);
or U17293 (N_17293,N_17139,N_17136);
nand U17294 (N_17294,N_17213,N_17269);
nor U17295 (N_17295,N_17256,N_17275);
or U17296 (N_17296,N_17239,N_17232);
or U17297 (N_17297,N_17265,N_17131);
or U17298 (N_17298,N_17248,N_17173);
nor U17299 (N_17299,N_17150,N_17199);
or U17300 (N_17300,N_17255,N_17187);
nor U17301 (N_17301,N_17267,N_17184);
nand U17302 (N_17302,N_17154,N_17201);
nor U17303 (N_17303,N_17143,N_17163);
xor U17304 (N_17304,N_17145,N_17140);
and U17305 (N_17305,N_17263,N_17253);
nand U17306 (N_17306,N_17158,N_17125);
nor U17307 (N_17307,N_17130,N_17233);
nor U17308 (N_17308,N_17268,N_17279);
and U17309 (N_17309,N_17264,N_17137);
nand U17310 (N_17310,N_17189,N_17194);
and U17311 (N_17311,N_17177,N_17219);
or U17312 (N_17312,N_17161,N_17142);
nor U17313 (N_17313,N_17185,N_17212);
nand U17314 (N_17314,N_17149,N_17128);
or U17315 (N_17315,N_17231,N_17227);
nand U17316 (N_17316,N_17176,N_17262);
or U17317 (N_17317,N_17168,N_17244);
nand U17318 (N_17318,N_17210,N_17257);
nor U17319 (N_17319,N_17129,N_17252);
or U17320 (N_17320,N_17217,N_17196);
and U17321 (N_17321,N_17159,N_17241);
and U17322 (N_17322,N_17206,N_17166);
xnor U17323 (N_17323,N_17271,N_17181);
nor U17324 (N_17324,N_17183,N_17226);
nor U17325 (N_17325,N_17203,N_17261);
nor U17326 (N_17326,N_17260,N_17175);
nor U17327 (N_17327,N_17200,N_17274);
nand U17328 (N_17328,N_17243,N_17127);
nor U17329 (N_17329,N_17254,N_17192);
xor U17330 (N_17330,N_17179,N_17135);
nand U17331 (N_17331,N_17207,N_17121);
nor U17332 (N_17332,N_17162,N_17276);
and U17333 (N_17333,N_17221,N_17188);
nand U17334 (N_17334,N_17146,N_17259);
nand U17335 (N_17335,N_17218,N_17164);
or U17336 (N_17336,N_17205,N_17249);
nor U17337 (N_17337,N_17167,N_17240);
nor U17338 (N_17338,N_17141,N_17171);
nor U17339 (N_17339,N_17123,N_17122);
or U17340 (N_17340,N_17151,N_17197);
nand U17341 (N_17341,N_17251,N_17165);
and U17342 (N_17342,N_17174,N_17182);
nand U17343 (N_17343,N_17126,N_17270);
nor U17344 (N_17344,N_17144,N_17202);
or U17345 (N_17345,N_17242,N_17152);
nand U17346 (N_17346,N_17153,N_17169);
nor U17347 (N_17347,N_17245,N_17195);
nor U17348 (N_17348,N_17198,N_17238);
and U17349 (N_17349,N_17178,N_17266);
or U17350 (N_17350,N_17214,N_17229);
nor U17351 (N_17351,N_17236,N_17155);
nor U17352 (N_17352,N_17230,N_17250);
or U17353 (N_17353,N_17277,N_17134);
and U17354 (N_17354,N_17211,N_17180);
and U17355 (N_17355,N_17204,N_17235);
nand U17356 (N_17356,N_17237,N_17220);
or U17357 (N_17357,N_17222,N_17234);
xor U17358 (N_17358,N_17124,N_17133);
xor U17359 (N_17359,N_17223,N_17186);
or U17360 (N_17360,N_17272,N_17122);
or U17361 (N_17361,N_17198,N_17166);
xnor U17362 (N_17362,N_17192,N_17174);
xnor U17363 (N_17363,N_17274,N_17260);
nor U17364 (N_17364,N_17129,N_17171);
xnor U17365 (N_17365,N_17261,N_17211);
nor U17366 (N_17366,N_17262,N_17153);
and U17367 (N_17367,N_17195,N_17179);
or U17368 (N_17368,N_17262,N_17217);
and U17369 (N_17369,N_17235,N_17255);
nor U17370 (N_17370,N_17186,N_17131);
nor U17371 (N_17371,N_17124,N_17140);
nand U17372 (N_17372,N_17238,N_17200);
xnor U17373 (N_17373,N_17159,N_17247);
or U17374 (N_17374,N_17249,N_17131);
nor U17375 (N_17375,N_17134,N_17162);
or U17376 (N_17376,N_17135,N_17136);
and U17377 (N_17377,N_17205,N_17151);
xor U17378 (N_17378,N_17184,N_17244);
nand U17379 (N_17379,N_17260,N_17194);
nand U17380 (N_17380,N_17204,N_17260);
nor U17381 (N_17381,N_17199,N_17172);
nand U17382 (N_17382,N_17183,N_17157);
nor U17383 (N_17383,N_17264,N_17138);
and U17384 (N_17384,N_17194,N_17277);
nor U17385 (N_17385,N_17179,N_17146);
nand U17386 (N_17386,N_17131,N_17151);
and U17387 (N_17387,N_17171,N_17151);
xor U17388 (N_17388,N_17238,N_17193);
nand U17389 (N_17389,N_17214,N_17200);
xor U17390 (N_17390,N_17193,N_17144);
or U17391 (N_17391,N_17227,N_17182);
nor U17392 (N_17392,N_17161,N_17256);
xnor U17393 (N_17393,N_17164,N_17211);
nand U17394 (N_17394,N_17264,N_17244);
nand U17395 (N_17395,N_17124,N_17244);
nor U17396 (N_17396,N_17164,N_17148);
or U17397 (N_17397,N_17218,N_17229);
and U17398 (N_17398,N_17235,N_17254);
and U17399 (N_17399,N_17238,N_17233);
xor U17400 (N_17400,N_17153,N_17138);
xnor U17401 (N_17401,N_17261,N_17232);
nor U17402 (N_17402,N_17167,N_17126);
and U17403 (N_17403,N_17148,N_17154);
or U17404 (N_17404,N_17135,N_17130);
nand U17405 (N_17405,N_17243,N_17151);
nor U17406 (N_17406,N_17184,N_17134);
nand U17407 (N_17407,N_17208,N_17263);
and U17408 (N_17408,N_17134,N_17122);
nand U17409 (N_17409,N_17217,N_17146);
or U17410 (N_17410,N_17144,N_17232);
and U17411 (N_17411,N_17129,N_17124);
nor U17412 (N_17412,N_17157,N_17191);
nand U17413 (N_17413,N_17240,N_17249);
or U17414 (N_17414,N_17208,N_17268);
nor U17415 (N_17415,N_17193,N_17223);
and U17416 (N_17416,N_17226,N_17229);
or U17417 (N_17417,N_17196,N_17172);
or U17418 (N_17418,N_17217,N_17167);
and U17419 (N_17419,N_17259,N_17174);
and U17420 (N_17420,N_17271,N_17211);
and U17421 (N_17421,N_17223,N_17182);
and U17422 (N_17422,N_17155,N_17201);
or U17423 (N_17423,N_17201,N_17176);
or U17424 (N_17424,N_17140,N_17179);
or U17425 (N_17425,N_17251,N_17203);
and U17426 (N_17426,N_17186,N_17270);
and U17427 (N_17427,N_17147,N_17215);
or U17428 (N_17428,N_17248,N_17188);
nand U17429 (N_17429,N_17143,N_17125);
or U17430 (N_17430,N_17200,N_17192);
and U17431 (N_17431,N_17257,N_17224);
and U17432 (N_17432,N_17171,N_17222);
xor U17433 (N_17433,N_17272,N_17139);
nand U17434 (N_17434,N_17141,N_17123);
and U17435 (N_17435,N_17265,N_17122);
nand U17436 (N_17436,N_17234,N_17158);
and U17437 (N_17437,N_17168,N_17141);
or U17438 (N_17438,N_17269,N_17120);
nor U17439 (N_17439,N_17245,N_17151);
nor U17440 (N_17440,N_17398,N_17378);
or U17441 (N_17441,N_17287,N_17281);
nand U17442 (N_17442,N_17292,N_17285);
nand U17443 (N_17443,N_17337,N_17284);
nand U17444 (N_17444,N_17408,N_17421);
and U17445 (N_17445,N_17383,N_17338);
and U17446 (N_17446,N_17394,N_17380);
and U17447 (N_17447,N_17330,N_17414);
or U17448 (N_17448,N_17350,N_17379);
nor U17449 (N_17449,N_17304,N_17323);
nor U17450 (N_17450,N_17366,N_17311);
xnor U17451 (N_17451,N_17401,N_17333);
nor U17452 (N_17452,N_17412,N_17413);
and U17453 (N_17453,N_17301,N_17415);
and U17454 (N_17454,N_17369,N_17342);
xnor U17455 (N_17455,N_17429,N_17432);
or U17456 (N_17456,N_17381,N_17345);
nor U17457 (N_17457,N_17355,N_17362);
nand U17458 (N_17458,N_17384,N_17303);
and U17459 (N_17459,N_17439,N_17294);
xor U17460 (N_17460,N_17374,N_17392);
or U17461 (N_17461,N_17418,N_17319);
and U17462 (N_17462,N_17300,N_17358);
or U17463 (N_17463,N_17326,N_17411);
xnor U17464 (N_17464,N_17313,N_17280);
nand U17465 (N_17465,N_17335,N_17382);
or U17466 (N_17466,N_17295,N_17356);
nor U17467 (N_17467,N_17348,N_17288);
nor U17468 (N_17468,N_17344,N_17428);
or U17469 (N_17469,N_17373,N_17402);
nand U17470 (N_17470,N_17389,N_17315);
or U17471 (N_17471,N_17438,N_17306);
nor U17472 (N_17472,N_17404,N_17349);
nor U17473 (N_17473,N_17360,N_17346);
or U17474 (N_17474,N_17430,N_17376);
nand U17475 (N_17475,N_17405,N_17436);
and U17476 (N_17476,N_17308,N_17341);
nand U17477 (N_17477,N_17386,N_17422);
nand U17478 (N_17478,N_17425,N_17324);
nand U17479 (N_17479,N_17434,N_17390);
nand U17480 (N_17480,N_17353,N_17312);
and U17481 (N_17481,N_17359,N_17361);
and U17482 (N_17482,N_17293,N_17407);
or U17483 (N_17483,N_17431,N_17399);
xnor U17484 (N_17484,N_17416,N_17299);
or U17485 (N_17485,N_17371,N_17351);
nand U17486 (N_17486,N_17332,N_17316);
nor U17487 (N_17487,N_17403,N_17427);
nor U17488 (N_17488,N_17420,N_17423);
nand U17489 (N_17489,N_17325,N_17310);
or U17490 (N_17490,N_17397,N_17370);
and U17491 (N_17491,N_17307,N_17317);
and U17492 (N_17492,N_17331,N_17302);
or U17493 (N_17493,N_17321,N_17340);
nor U17494 (N_17494,N_17395,N_17419);
or U17495 (N_17495,N_17347,N_17375);
nand U17496 (N_17496,N_17327,N_17417);
or U17497 (N_17497,N_17336,N_17396);
nor U17498 (N_17498,N_17339,N_17354);
nor U17499 (N_17499,N_17283,N_17334);
nand U17500 (N_17500,N_17368,N_17391);
nor U17501 (N_17501,N_17290,N_17424);
and U17502 (N_17502,N_17363,N_17322);
and U17503 (N_17503,N_17291,N_17289);
nand U17504 (N_17504,N_17433,N_17298);
nor U17505 (N_17505,N_17320,N_17286);
and U17506 (N_17506,N_17328,N_17388);
or U17507 (N_17507,N_17282,N_17426);
xnor U17508 (N_17508,N_17365,N_17318);
and U17509 (N_17509,N_17357,N_17364);
or U17510 (N_17510,N_17437,N_17314);
and U17511 (N_17511,N_17406,N_17352);
or U17512 (N_17512,N_17387,N_17393);
nor U17513 (N_17513,N_17409,N_17343);
nor U17514 (N_17514,N_17435,N_17410);
and U17515 (N_17515,N_17372,N_17329);
nand U17516 (N_17516,N_17367,N_17296);
and U17517 (N_17517,N_17305,N_17400);
nand U17518 (N_17518,N_17385,N_17377);
or U17519 (N_17519,N_17297,N_17309);
nand U17520 (N_17520,N_17333,N_17282);
and U17521 (N_17521,N_17309,N_17429);
or U17522 (N_17522,N_17295,N_17287);
and U17523 (N_17523,N_17384,N_17327);
xnor U17524 (N_17524,N_17329,N_17301);
nand U17525 (N_17525,N_17361,N_17342);
nand U17526 (N_17526,N_17342,N_17416);
nor U17527 (N_17527,N_17384,N_17368);
nand U17528 (N_17528,N_17434,N_17286);
or U17529 (N_17529,N_17350,N_17353);
nand U17530 (N_17530,N_17325,N_17392);
nand U17531 (N_17531,N_17324,N_17379);
xnor U17532 (N_17532,N_17424,N_17393);
nand U17533 (N_17533,N_17411,N_17386);
and U17534 (N_17534,N_17331,N_17425);
or U17535 (N_17535,N_17301,N_17434);
and U17536 (N_17536,N_17343,N_17385);
or U17537 (N_17537,N_17437,N_17381);
or U17538 (N_17538,N_17336,N_17316);
or U17539 (N_17539,N_17354,N_17408);
nand U17540 (N_17540,N_17320,N_17321);
and U17541 (N_17541,N_17280,N_17303);
nand U17542 (N_17542,N_17345,N_17428);
xor U17543 (N_17543,N_17422,N_17330);
or U17544 (N_17544,N_17407,N_17292);
or U17545 (N_17545,N_17287,N_17415);
nand U17546 (N_17546,N_17326,N_17423);
nor U17547 (N_17547,N_17304,N_17352);
or U17548 (N_17548,N_17331,N_17389);
nand U17549 (N_17549,N_17311,N_17382);
nor U17550 (N_17550,N_17291,N_17355);
nor U17551 (N_17551,N_17289,N_17360);
nand U17552 (N_17552,N_17396,N_17414);
and U17553 (N_17553,N_17310,N_17384);
nand U17554 (N_17554,N_17391,N_17318);
xor U17555 (N_17555,N_17406,N_17358);
and U17556 (N_17556,N_17328,N_17422);
nor U17557 (N_17557,N_17288,N_17300);
nor U17558 (N_17558,N_17296,N_17354);
nor U17559 (N_17559,N_17417,N_17390);
or U17560 (N_17560,N_17372,N_17421);
or U17561 (N_17561,N_17314,N_17402);
xor U17562 (N_17562,N_17408,N_17312);
xor U17563 (N_17563,N_17292,N_17337);
nand U17564 (N_17564,N_17392,N_17301);
nand U17565 (N_17565,N_17426,N_17404);
nor U17566 (N_17566,N_17359,N_17408);
or U17567 (N_17567,N_17322,N_17356);
nor U17568 (N_17568,N_17331,N_17411);
nor U17569 (N_17569,N_17388,N_17346);
nand U17570 (N_17570,N_17326,N_17280);
nand U17571 (N_17571,N_17286,N_17294);
nor U17572 (N_17572,N_17308,N_17394);
nand U17573 (N_17573,N_17421,N_17359);
xor U17574 (N_17574,N_17285,N_17407);
nand U17575 (N_17575,N_17310,N_17319);
or U17576 (N_17576,N_17439,N_17386);
nand U17577 (N_17577,N_17353,N_17400);
or U17578 (N_17578,N_17302,N_17372);
or U17579 (N_17579,N_17357,N_17307);
nor U17580 (N_17580,N_17314,N_17348);
or U17581 (N_17581,N_17309,N_17404);
or U17582 (N_17582,N_17366,N_17417);
nor U17583 (N_17583,N_17297,N_17412);
and U17584 (N_17584,N_17303,N_17374);
and U17585 (N_17585,N_17310,N_17351);
or U17586 (N_17586,N_17302,N_17359);
nor U17587 (N_17587,N_17419,N_17349);
and U17588 (N_17588,N_17346,N_17337);
nand U17589 (N_17589,N_17367,N_17410);
xor U17590 (N_17590,N_17379,N_17405);
xor U17591 (N_17591,N_17315,N_17418);
nand U17592 (N_17592,N_17290,N_17420);
or U17593 (N_17593,N_17370,N_17414);
or U17594 (N_17594,N_17305,N_17309);
and U17595 (N_17595,N_17411,N_17432);
nor U17596 (N_17596,N_17349,N_17319);
nor U17597 (N_17597,N_17330,N_17387);
nand U17598 (N_17598,N_17291,N_17300);
and U17599 (N_17599,N_17387,N_17409);
or U17600 (N_17600,N_17447,N_17477);
and U17601 (N_17601,N_17565,N_17576);
and U17602 (N_17602,N_17483,N_17452);
nor U17603 (N_17603,N_17590,N_17494);
nand U17604 (N_17604,N_17563,N_17484);
xor U17605 (N_17605,N_17457,N_17572);
xnor U17606 (N_17606,N_17537,N_17583);
or U17607 (N_17607,N_17462,N_17453);
or U17608 (N_17608,N_17528,N_17498);
xor U17609 (N_17609,N_17584,N_17558);
and U17610 (N_17610,N_17479,N_17554);
or U17611 (N_17611,N_17592,N_17555);
and U17612 (N_17612,N_17504,N_17591);
or U17613 (N_17613,N_17567,N_17444);
nand U17614 (N_17614,N_17556,N_17547);
nor U17615 (N_17615,N_17596,N_17539);
and U17616 (N_17616,N_17445,N_17573);
or U17617 (N_17617,N_17580,N_17455);
or U17618 (N_17618,N_17530,N_17570);
and U17619 (N_17619,N_17470,N_17488);
nor U17620 (N_17620,N_17490,N_17461);
nand U17621 (N_17621,N_17443,N_17548);
nor U17622 (N_17622,N_17497,N_17485);
and U17623 (N_17623,N_17523,N_17464);
nand U17624 (N_17624,N_17441,N_17511);
or U17625 (N_17625,N_17514,N_17502);
nand U17626 (N_17626,N_17495,N_17575);
or U17627 (N_17627,N_17513,N_17503);
xnor U17628 (N_17628,N_17459,N_17588);
and U17629 (N_17629,N_17525,N_17515);
and U17630 (N_17630,N_17593,N_17505);
nor U17631 (N_17631,N_17508,N_17527);
nor U17632 (N_17632,N_17549,N_17454);
and U17633 (N_17633,N_17496,N_17456);
nor U17634 (N_17634,N_17506,N_17562);
or U17635 (N_17635,N_17543,N_17486);
and U17636 (N_17636,N_17507,N_17471);
xnor U17637 (N_17637,N_17586,N_17552);
xor U17638 (N_17638,N_17518,N_17491);
nand U17639 (N_17639,N_17500,N_17487);
nand U17640 (N_17640,N_17598,N_17466);
and U17641 (N_17641,N_17538,N_17531);
nand U17642 (N_17642,N_17529,N_17468);
or U17643 (N_17643,N_17524,N_17480);
xnor U17644 (N_17644,N_17599,N_17473);
xor U17645 (N_17645,N_17522,N_17566);
nand U17646 (N_17646,N_17519,N_17595);
or U17647 (N_17647,N_17542,N_17536);
and U17648 (N_17648,N_17569,N_17582);
nor U17649 (N_17649,N_17540,N_17516);
and U17650 (N_17650,N_17481,N_17465);
and U17651 (N_17651,N_17469,N_17499);
xor U17652 (N_17652,N_17489,N_17460);
and U17653 (N_17653,N_17475,N_17577);
or U17654 (N_17654,N_17449,N_17560);
nand U17655 (N_17655,N_17472,N_17482);
xor U17656 (N_17656,N_17561,N_17551);
or U17657 (N_17657,N_17585,N_17467);
nand U17658 (N_17658,N_17510,N_17440);
nand U17659 (N_17659,N_17574,N_17521);
xnor U17660 (N_17660,N_17579,N_17546);
or U17661 (N_17661,N_17557,N_17478);
xnor U17662 (N_17662,N_17564,N_17451);
and U17663 (N_17663,N_17448,N_17450);
nor U17664 (N_17664,N_17541,N_17492);
xnor U17665 (N_17665,N_17517,N_17463);
and U17666 (N_17666,N_17533,N_17594);
nand U17667 (N_17667,N_17509,N_17442);
xor U17668 (N_17668,N_17553,N_17476);
xnor U17669 (N_17669,N_17559,N_17520);
and U17670 (N_17670,N_17493,N_17512);
and U17671 (N_17671,N_17578,N_17446);
and U17672 (N_17672,N_17550,N_17597);
nand U17673 (N_17673,N_17501,N_17587);
nor U17674 (N_17674,N_17544,N_17581);
and U17675 (N_17675,N_17571,N_17532);
and U17676 (N_17676,N_17534,N_17535);
nand U17677 (N_17677,N_17458,N_17526);
and U17678 (N_17678,N_17589,N_17474);
or U17679 (N_17679,N_17568,N_17545);
nand U17680 (N_17680,N_17442,N_17469);
and U17681 (N_17681,N_17516,N_17463);
nor U17682 (N_17682,N_17497,N_17565);
or U17683 (N_17683,N_17544,N_17584);
or U17684 (N_17684,N_17522,N_17597);
or U17685 (N_17685,N_17462,N_17574);
and U17686 (N_17686,N_17466,N_17474);
or U17687 (N_17687,N_17568,N_17493);
nor U17688 (N_17688,N_17522,N_17599);
and U17689 (N_17689,N_17597,N_17517);
nor U17690 (N_17690,N_17507,N_17557);
and U17691 (N_17691,N_17505,N_17525);
nand U17692 (N_17692,N_17599,N_17596);
or U17693 (N_17693,N_17481,N_17581);
nand U17694 (N_17694,N_17446,N_17524);
nand U17695 (N_17695,N_17577,N_17448);
nand U17696 (N_17696,N_17592,N_17450);
nor U17697 (N_17697,N_17473,N_17598);
nand U17698 (N_17698,N_17548,N_17573);
nand U17699 (N_17699,N_17467,N_17480);
and U17700 (N_17700,N_17545,N_17441);
or U17701 (N_17701,N_17517,N_17495);
nor U17702 (N_17702,N_17576,N_17532);
nor U17703 (N_17703,N_17546,N_17475);
nor U17704 (N_17704,N_17443,N_17452);
nor U17705 (N_17705,N_17566,N_17495);
nor U17706 (N_17706,N_17502,N_17442);
nand U17707 (N_17707,N_17531,N_17459);
nor U17708 (N_17708,N_17501,N_17495);
and U17709 (N_17709,N_17455,N_17519);
nor U17710 (N_17710,N_17502,N_17441);
xnor U17711 (N_17711,N_17511,N_17477);
nor U17712 (N_17712,N_17552,N_17471);
nor U17713 (N_17713,N_17441,N_17459);
and U17714 (N_17714,N_17462,N_17591);
and U17715 (N_17715,N_17462,N_17471);
nor U17716 (N_17716,N_17487,N_17549);
or U17717 (N_17717,N_17549,N_17557);
nand U17718 (N_17718,N_17501,N_17555);
xnor U17719 (N_17719,N_17486,N_17443);
xnor U17720 (N_17720,N_17520,N_17499);
and U17721 (N_17721,N_17534,N_17490);
or U17722 (N_17722,N_17507,N_17442);
or U17723 (N_17723,N_17512,N_17474);
or U17724 (N_17724,N_17447,N_17506);
or U17725 (N_17725,N_17532,N_17514);
or U17726 (N_17726,N_17446,N_17481);
and U17727 (N_17727,N_17572,N_17533);
nand U17728 (N_17728,N_17536,N_17461);
nand U17729 (N_17729,N_17571,N_17475);
nor U17730 (N_17730,N_17593,N_17527);
nor U17731 (N_17731,N_17552,N_17532);
nand U17732 (N_17732,N_17571,N_17503);
xnor U17733 (N_17733,N_17524,N_17574);
nor U17734 (N_17734,N_17502,N_17509);
nor U17735 (N_17735,N_17582,N_17464);
xor U17736 (N_17736,N_17484,N_17512);
nand U17737 (N_17737,N_17536,N_17495);
or U17738 (N_17738,N_17459,N_17551);
nand U17739 (N_17739,N_17475,N_17495);
nand U17740 (N_17740,N_17548,N_17466);
xor U17741 (N_17741,N_17599,N_17551);
nand U17742 (N_17742,N_17582,N_17482);
nor U17743 (N_17743,N_17586,N_17535);
or U17744 (N_17744,N_17462,N_17564);
nand U17745 (N_17745,N_17484,N_17518);
nand U17746 (N_17746,N_17468,N_17583);
or U17747 (N_17747,N_17491,N_17445);
xor U17748 (N_17748,N_17598,N_17586);
nor U17749 (N_17749,N_17521,N_17571);
nand U17750 (N_17750,N_17445,N_17547);
and U17751 (N_17751,N_17558,N_17463);
or U17752 (N_17752,N_17507,N_17508);
or U17753 (N_17753,N_17560,N_17532);
and U17754 (N_17754,N_17548,N_17477);
nor U17755 (N_17755,N_17582,N_17461);
nand U17756 (N_17756,N_17514,N_17572);
nor U17757 (N_17757,N_17465,N_17501);
nor U17758 (N_17758,N_17511,N_17496);
nand U17759 (N_17759,N_17445,N_17507);
and U17760 (N_17760,N_17668,N_17686);
nand U17761 (N_17761,N_17641,N_17737);
and U17762 (N_17762,N_17664,N_17678);
nand U17763 (N_17763,N_17607,N_17625);
and U17764 (N_17764,N_17730,N_17680);
nor U17765 (N_17765,N_17633,N_17759);
or U17766 (N_17766,N_17612,N_17690);
and U17767 (N_17767,N_17715,N_17681);
and U17768 (N_17768,N_17622,N_17682);
and U17769 (N_17769,N_17709,N_17744);
nand U17770 (N_17770,N_17741,N_17604);
nand U17771 (N_17771,N_17704,N_17747);
nor U17772 (N_17772,N_17648,N_17755);
or U17773 (N_17773,N_17702,N_17700);
nor U17774 (N_17774,N_17639,N_17751);
and U17775 (N_17775,N_17712,N_17662);
nand U17776 (N_17776,N_17732,N_17718);
and U17777 (N_17777,N_17723,N_17670);
and U17778 (N_17778,N_17642,N_17722);
or U17779 (N_17779,N_17660,N_17636);
xnor U17780 (N_17780,N_17656,N_17754);
nor U17781 (N_17781,N_17701,N_17626);
xor U17782 (N_17782,N_17716,N_17667);
and U17783 (N_17783,N_17638,N_17706);
nand U17784 (N_17784,N_17679,N_17753);
nand U17785 (N_17785,N_17609,N_17603);
nor U17786 (N_17786,N_17677,N_17738);
nand U17787 (N_17787,N_17644,N_17740);
nand U17788 (N_17788,N_17602,N_17651);
nor U17789 (N_17789,N_17630,N_17666);
and U17790 (N_17790,N_17727,N_17650);
xnor U17791 (N_17791,N_17689,N_17623);
and U17792 (N_17792,N_17683,N_17675);
nor U17793 (N_17793,N_17617,N_17726);
xor U17794 (N_17794,N_17621,N_17734);
nor U17795 (N_17795,N_17708,N_17632);
xnor U17796 (N_17796,N_17696,N_17610);
and U17797 (N_17797,N_17645,N_17725);
xor U17798 (N_17798,N_17728,N_17691);
nand U17799 (N_17799,N_17658,N_17600);
and U17800 (N_17800,N_17752,N_17711);
or U17801 (N_17801,N_17620,N_17637);
or U17802 (N_17802,N_17721,N_17635);
nor U17803 (N_17803,N_17729,N_17673);
and U17804 (N_17804,N_17743,N_17736);
nand U17805 (N_17805,N_17719,N_17756);
nand U17806 (N_17806,N_17720,N_17672);
nand U17807 (N_17807,N_17605,N_17695);
and U17808 (N_17808,N_17649,N_17698);
nand U17809 (N_17809,N_17758,N_17684);
and U17810 (N_17810,N_17608,N_17653);
and U17811 (N_17811,N_17652,N_17624);
nor U17812 (N_17812,N_17717,N_17688);
nor U17813 (N_17813,N_17628,N_17606);
nand U17814 (N_17814,N_17640,N_17674);
and U17815 (N_17815,N_17739,N_17659);
or U17816 (N_17816,N_17619,N_17654);
and U17817 (N_17817,N_17735,N_17646);
and U17818 (N_17818,N_17713,N_17710);
nor U17819 (N_17819,N_17669,N_17614);
nand U17820 (N_17820,N_17705,N_17618);
or U17821 (N_17821,N_17676,N_17629);
nor U17822 (N_17822,N_17757,N_17671);
and U17823 (N_17823,N_17693,N_17699);
nand U17824 (N_17824,N_17697,N_17601);
xor U17825 (N_17825,N_17661,N_17655);
xnor U17826 (N_17826,N_17685,N_17627);
nor U17827 (N_17827,N_17745,N_17643);
nand U17828 (N_17828,N_17703,N_17750);
nand U17829 (N_17829,N_17733,N_17665);
and U17830 (N_17830,N_17616,N_17611);
or U17831 (N_17831,N_17657,N_17748);
nand U17832 (N_17832,N_17692,N_17647);
and U17833 (N_17833,N_17687,N_17615);
or U17834 (N_17834,N_17714,N_17724);
or U17835 (N_17835,N_17631,N_17694);
nand U17836 (N_17836,N_17749,N_17663);
nand U17837 (N_17837,N_17742,N_17613);
and U17838 (N_17838,N_17634,N_17707);
nand U17839 (N_17839,N_17731,N_17746);
nor U17840 (N_17840,N_17737,N_17740);
and U17841 (N_17841,N_17714,N_17632);
nor U17842 (N_17842,N_17636,N_17646);
or U17843 (N_17843,N_17662,N_17757);
nor U17844 (N_17844,N_17744,N_17617);
nor U17845 (N_17845,N_17702,N_17685);
and U17846 (N_17846,N_17703,N_17640);
xnor U17847 (N_17847,N_17699,N_17639);
nand U17848 (N_17848,N_17692,N_17694);
xnor U17849 (N_17849,N_17667,N_17691);
nor U17850 (N_17850,N_17605,N_17628);
nor U17851 (N_17851,N_17663,N_17743);
or U17852 (N_17852,N_17691,N_17724);
and U17853 (N_17853,N_17673,N_17712);
nand U17854 (N_17854,N_17600,N_17627);
and U17855 (N_17855,N_17683,N_17658);
or U17856 (N_17856,N_17713,N_17759);
nand U17857 (N_17857,N_17641,N_17695);
and U17858 (N_17858,N_17754,N_17678);
nand U17859 (N_17859,N_17609,N_17685);
xnor U17860 (N_17860,N_17650,N_17735);
nor U17861 (N_17861,N_17729,N_17701);
xor U17862 (N_17862,N_17635,N_17736);
nor U17863 (N_17863,N_17609,N_17738);
nand U17864 (N_17864,N_17729,N_17728);
nand U17865 (N_17865,N_17696,N_17733);
nand U17866 (N_17866,N_17676,N_17684);
nor U17867 (N_17867,N_17639,N_17730);
and U17868 (N_17868,N_17616,N_17702);
nor U17869 (N_17869,N_17657,N_17662);
nor U17870 (N_17870,N_17719,N_17653);
or U17871 (N_17871,N_17616,N_17706);
and U17872 (N_17872,N_17641,N_17657);
or U17873 (N_17873,N_17657,N_17664);
or U17874 (N_17874,N_17697,N_17685);
or U17875 (N_17875,N_17736,N_17721);
nor U17876 (N_17876,N_17618,N_17613);
nand U17877 (N_17877,N_17648,N_17750);
or U17878 (N_17878,N_17756,N_17668);
and U17879 (N_17879,N_17716,N_17680);
nor U17880 (N_17880,N_17666,N_17642);
and U17881 (N_17881,N_17645,N_17670);
nor U17882 (N_17882,N_17642,N_17694);
or U17883 (N_17883,N_17632,N_17756);
or U17884 (N_17884,N_17685,N_17722);
or U17885 (N_17885,N_17743,N_17725);
and U17886 (N_17886,N_17664,N_17666);
or U17887 (N_17887,N_17671,N_17649);
and U17888 (N_17888,N_17715,N_17734);
nor U17889 (N_17889,N_17665,N_17750);
and U17890 (N_17890,N_17670,N_17712);
and U17891 (N_17891,N_17725,N_17755);
or U17892 (N_17892,N_17692,N_17736);
or U17893 (N_17893,N_17630,N_17619);
or U17894 (N_17894,N_17737,N_17757);
and U17895 (N_17895,N_17623,N_17715);
or U17896 (N_17896,N_17632,N_17642);
or U17897 (N_17897,N_17671,N_17729);
nand U17898 (N_17898,N_17743,N_17688);
nor U17899 (N_17899,N_17629,N_17689);
nor U17900 (N_17900,N_17730,N_17754);
nand U17901 (N_17901,N_17673,N_17692);
nor U17902 (N_17902,N_17746,N_17735);
or U17903 (N_17903,N_17685,N_17639);
nor U17904 (N_17904,N_17731,N_17621);
or U17905 (N_17905,N_17622,N_17647);
nor U17906 (N_17906,N_17700,N_17707);
or U17907 (N_17907,N_17630,N_17606);
or U17908 (N_17908,N_17708,N_17657);
nand U17909 (N_17909,N_17674,N_17601);
nand U17910 (N_17910,N_17632,N_17638);
and U17911 (N_17911,N_17694,N_17668);
nor U17912 (N_17912,N_17731,N_17600);
and U17913 (N_17913,N_17704,N_17719);
nor U17914 (N_17914,N_17709,N_17693);
and U17915 (N_17915,N_17734,N_17708);
or U17916 (N_17916,N_17660,N_17744);
or U17917 (N_17917,N_17647,N_17627);
or U17918 (N_17918,N_17623,N_17656);
and U17919 (N_17919,N_17700,N_17605);
and U17920 (N_17920,N_17807,N_17802);
nand U17921 (N_17921,N_17813,N_17791);
and U17922 (N_17922,N_17854,N_17828);
or U17923 (N_17923,N_17774,N_17767);
nor U17924 (N_17924,N_17775,N_17777);
nand U17925 (N_17925,N_17821,N_17823);
nor U17926 (N_17926,N_17869,N_17811);
and U17927 (N_17927,N_17838,N_17844);
nor U17928 (N_17928,N_17878,N_17834);
nand U17929 (N_17929,N_17781,N_17898);
or U17930 (N_17930,N_17865,N_17848);
or U17931 (N_17931,N_17859,N_17861);
or U17932 (N_17932,N_17816,N_17914);
nor U17933 (N_17933,N_17910,N_17842);
nor U17934 (N_17934,N_17763,N_17786);
or U17935 (N_17935,N_17762,N_17872);
nand U17936 (N_17936,N_17785,N_17851);
or U17937 (N_17937,N_17862,N_17858);
or U17938 (N_17938,N_17796,N_17776);
nand U17939 (N_17939,N_17876,N_17814);
nor U17940 (N_17940,N_17885,N_17832);
and U17941 (N_17941,N_17866,N_17810);
or U17942 (N_17942,N_17900,N_17798);
nand U17943 (N_17943,N_17843,N_17809);
and U17944 (N_17944,N_17889,N_17857);
nand U17945 (N_17945,N_17901,N_17830);
or U17946 (N_17946,N_17780,N_17887);
nand U17947 (N_17947,N_17833,N_17771);
and U17948 (N_17948,N_17916,N_17911);
nand U17949 (N_17949,N_17849,N_17801);
or U17950 (N_17950,N_17773,N_17904);
xor U17951 (N_17951,N_17790,N_17831);
and U17952 (N_17952,N_17766,N_17908);
nor U17953 (N_17953,N_17768,N_17788);
nor U17954 (N_17954,N_17829,N_17794);
nor U17955 (N_17955,N_17879,N_17840);
nor U17956 (N_17956,N_17841,N_17803);
nor U17957 (N_17957,N_17837,N_17875);
and U17958 (N_17958,N_17817,N_17764);
nor U17959 (N_17959,N_17864,N_17822);
xnor U17960 (N_17960,N_17902,N_17805);
and U17961 (N_17961,N_17800,N_17847);
or U17962 (N_17962,N_17778,N_17855);
nor U17963 (N_17963,N_17895,N_17793);
xnor U17964 (N_17964,N_17880,N_17863);
or U17965 (N_17965,N_17799,N_17888);
xnor U17966 (N_17966,N_17891,N_17761);
and U17967 (N_17967,N_17820,N_17890);
nor U17968 (N_17968,N_17795,N_17896);
nor U17969 (N_17969,N_17860,N_17808);
and U17970 (N_17970,N_17903,N_17871);
nor U17971 (N_17971,N_17769,N_17918);
nor U17972 (N_17972,N_17825,N_17783);
nor U17973 (N_17973,N_17818,N_17853);
and U17974 (N_17974,N_17835,N_17852);
nand U17975 (N_17975,N_17804,N_17915);
nand U17976 (N_17976,N_17784,N_17806);
nand U17977 (N_17977,N_17856,N_17873);
or U17978 (N_17978,N_17839,N_17782);
nor U17979 (N_17979,N_17779,N_17897);
and U17980 (N_17980,N_17819,N_17789);
and U17981 (N_17981,N_17894,N_17765);
and U17982 (N_17982,N_17868,N_17850);
nand U17983 (N_17983,N_17883,N_17886);
or U17984 (N_17984,N_17797,N_17770);
nand U17985 (N_17985,N_17919,N_17906);
or U17986 (N_17986,N_17909,N_17812);
and U17987 (N_17987,N_17846,N_17760);
nor U17988 (N_17988,N_17893,N_17845);
nand U17989 (N_17989,N_17899,N_17826);
or U17990 (N_17990,N_17884,N_17905);
and U17991 (N_17991,N_17815,N_17867);
nor U17992 (N_17992,N_17917,N_17824);
and U17993 (N_17993,N_17892,N_17772);
and U17994 (N_17994,N_17881,N_17827);
nor U17995 (N_17995,N_17913,N_17787);
or U17996 (N_17996,N_17792,N_17907);
or U17997 (N_17997,N_17912,N_17870);
or U17998 (N_17998,N_17874,N_17877);
or U17999 (N_17999,N_17836,N_17882);
nor U18000 (N_18000,N_17861,N_17791);
nor U18001 (N_18001,N_17795,N_17828);
nand U18002 (N_18002,N_17865,N_17888);
or U18003 (N_18003,N_17845,N_17849);
and U18004 (N_18004,N_17844,N_17911);
nor U18005 (N_18005,N_17837,N_17907);
or U18006 (N_18006,N_17760,N_17855);
nor U18007 (N_18007,N_17812,N_17803);
or U18008 (N_18008,N_17852,N_17819);
xor U18009 (N_18009,N_17796,N_17801);
or U18010 (N_18010,N_17807,N_17767);
nand U18011 (N_18011,N_17829,N_17889);
nand U18012 (N_18012,N_17863,N_17786);
nand U18013 (N_18013,N_17872,N_17828);
or U18014 (N_18014,N_17800,N_17805);
and U18015 (N_18015,N_17908,N_17763);
and U18016 (N_18016,N_17860,N_17902);
nand U18017 (N_18017,N_17856,N_17916);
xor U18018 (N_18018,N_17914,N_17785);
nor U18019 (N_18019,N_17830,N_17883);
or U18020 (N_18020,N_17831,N_17891);
or U18021 (N_18021,N_17824,N_17772);
nor U18022 (N_18022,N_17788,N_17882);
nand U18023 (N_18023,N_17796,N_17841);
nand U18024 (N_18024,N_17901,N_17847);
and U18025 (N_18025,N_17837,N_17781);
xor U18026 (N_18026,N_17839,N_17819);
or U18027 (N_18027,N_17807,N_17858);
and U18028 (N_18028,N_17828,N_17855);
nor U18029 (N_18029,N_17873,N_17800);
or U18030 (N_18030,N_17788,N_17846);
and U18031 (N_18031,N_17890,N_17882);
nand U18032 (N_18032,N_17893,N_17816);
and U18033 (N_18033,N_17830,N_17868);
or U18034 (N_18034,N_17864,N_17845);
or U18035 (N_18035,N_17865,N_17773);
or U18036 (N_18036,N_17883,N_17777);
nand U18037 (N_18037,N_17898,N_17787);
or U18038 (N_18038,N_17868,N_17782);
nor U18039 (N_18039,N_17784,N_17919);
or U18040 (N_18040,N_17837,N_17773);
and U18041 (N_18041,N_17782,N_17856);
and U18042 (N_18042,N_17771,N_17792);
or U18043 (N_18043,N_17844,N_17762);
nor U18044 (N_18044,N_17842,N_17822);
and U18045 (N_18045,N_17863,N_17860);
or U18046 (N_18046,N_17798,N_17823);
nand U18047 (N_18047,N_17867,N_17836);
or U18048 (N_18048,N_17831,N_17806);
and U18049 (N_18049,N_17760,N_17894);
and U18050 (N_18050,N_17859,N_17886);
nand U18051 (N_18051,N_17882,N_17893);
nor U18052 (N_18052,N_17820,N_17801);
nor U18053 (N_18053,N_17786,N_17869);
or U18054 (N_18054,N_17856,N_17797);
xnor U18055 (N_18055,N_17885,N_17866);
nand U18056 (N_18056,N_17875,N_17791);
and U18057 (N_18057,N_17831,N_17886);
or U18058 (N_18058,N_17858,N_17889);
nand U18059 (N_18059,N_17830,N_17856);
and U18060 (N_18060,N_17794,N_17903);
nor U18061 (N_18061,N_17777,N_17785);
or U18062 (N_18062,N_17852,N_17874);
or U18063 (N_18063,N_17764,N_17808);
or U18064 (N_18064,N_17799,N_17836);
or U18065 (N_18065,N_17797,N_17829);
nand U18066 (N_18066,N_17916,N_17884);
and U18067 (N_18067,N_17891,N_17822);
nor U18068 (N_18068,N_17818,N_17865);
nor U18069 (N_18069,N_17826,N_17815);
nand U18070 (N_18070,N_17822,N_17895);
or U18071 (N_18071,N_17916,N_17809);
nor U18072 (N_18072,N_17772,N_17856);
or U18073 (N_18073,N_17786,N_17803);
xor U18074 (N_18074,N_17785,N_17808);
nand U18075 (N_18075,N_17821,N_17862);
and U18076 (N_18076,N_17883,N_17778);
nor U18077 (N_18077,N_17762,N_17825);
nor U18078 (N_18078,N_17871,N_17825);
xnor U18079 (N_18079,N_17761,N_17857);
or U18080 (N_18080,N_17951,N_18014);
and U18081 (N_18081,N_17920,N_17922);
or U18082 (N_18082,N_17972,N_17930);
and U18083 (N_18083,N_17969,N_18033);
or U18084 (N_18084,N_18076,N_18049);
nor U18085 (N_18085,N_18001,N_18047);
xor U18086 (N_18086,N_17939,N_17984);
nand U18087 (N_18087,N_18005,N_18032);
and U18088 (N_18088,N_18046,N_17990);
and U18089 (N_18089,N_18071,N_17983);
and U18090 (N_18090,N_17961,N_18044);
nor U18091 (N_18091,N_18028,N_18006);
or U18092 (N_18092,N_17970,N_17942);
and U18093 (N_18093,N_17988,N_18000);
or U18094 (N_18094,N_18068,N_18040);
and U18095 (N_18095,N_18078,N_17977);
nand U18096 (N_18096,N_18026,N_17991);
xor U18097 (N_18097,N_17954,N_17999);
nand U18098 (N_18098,N_17928,N_17964);
nor U18099 (N_18099,N_18052,N_17949);
nor U18100 (N_18100,N_18035,N_17946);
xor U18101 (N_18101,N_18075,N_18048);
nand U18102 (N_18102,N_17955,N_17978);
or U18103 (N_18103,N_18058,N_18016);
or U18104 (N_18104,N_18041,N_17923);
or U18105 (N_18105,N_18061,N_18009);
and U18106 (N_18106,N_18065,N_17953);
and U18107 (N_18107,N_18067,N_17925);
nand U18108 (N_18108,N_17971,N_17927);
and U18109 (N_18109,N_17981,N_17966);
and U18110 (N_18110,N_17965,N_17957);
nor U18111 (N_18111,N_17985,N_18059);
xor U18112 (N_18112,N_17974,N_18002);
or U18113 (N_18113,N_18036,N_17935);
or U18114 (N_18114,N_18079,N_18010);
or U18115 (N_18115,N_17932,N_18018);
and U18116 (N_18116,N_17968,N_17956);
xnor U18117 (N_18117,N_17926,N_17973);
nor U18118 (N_18118,N_18053,N_17979);
nand U18119 (N_18119,N_18077,N_18021);
or U18120 (N_18120,N_18055,N_18007);
and U18121 (N_18121,N_18050,N_17945);
or U18122 (N_18122,N_17936,N_17960);
and U18123 (N_18123,N_18057,N_17980);
or U18124 (N_18124,N_18025,N_18017);
and U18125 (N_18125,N_18013,N_17967);
nor U18126 (N_18126,N_17962,N_17976);
xnor U18127 (N_18127,N_17938,N_18024);
xnor U18128 (N_18128,N_18051,N_18008);
nor U18129 (N_18129,N_18030,N_18060);
nor U18130 (N_18130,N_17997,N_18042);
nand U18131 (N_18131,N_17934,N_17989);
nand U18132 (N_18132,N_17924,N_17986);
nor U18133 (N_18133,N_17921,N_18003);
or U18134 (N_18134,N_17952,N_18073);
or U18135 (N_18135,N_18038,N_17996);
and U18136 (N_18136,N_18054,N_18015);
nor U18137 (N_18137,N_17929,N_18072);
nand U18138 (N_18138,N_18062,N_17943);
nor U18139 (N_18139,N_18004,N_17933);
nand U18140 (N_18140,N_18066,N_18019);
nor U18141 (N_18141,N_18074,N_18027);
nor U18142 (N_18142,N_18011,N_17994);
and U18143 (N_18143,N_18056,N_18064);
or U18144 (N_18144,N_18069,N_18063);
and U18145 (N_18145,N_17941,N_17982);
nor U18146 (N_18146,N_17959,N_17931);
or U18147 (N_18147,N_18070,N_17995);
or U18148 (N_18148,N_17944,N_17992);
xnor U18149 (N_18149,N_17998,N_17963);
or U18150 (N_18150,N_18034,N_18029);
xnor U18151 (N_18151,N_18043,N_18039);
xnor U18152 (N_18152,N_17950,N_18037);
nor U18153 (N_18153,N_18031,N_17937);
or U18154 (N_18154,N_17987,N_17975);
nand U18155 (N_18155,N_18023,N_17993);
or U18156 (N_18156,N_17948,N_17958);
and U18157 (N_18157,N_18012,N_17940);
xor U18158 (N_18158,N_18022,N_18020);
or U18159 (N_18159,N_17947,N_18045);
or U18160 (N_18160,N_18057,N_17996);
nor U18161 (N_18161,N_18058,N_17997);
nor U18162 (N_18162,N_18013,N_17947);
nor U18163 (N_18163,N_17973,N_17997);
nor U18164 (N_18164,N_18003,N_18051);
nand U18165 (N_18165,N_17962,N_17968);
nand U18166 (N_18166,N_18005,N_18060);
nor U18167 (N_18167,N_18035,N_18034);
nor U18168 (N_18168,N_17974,N_17922);
and U18169 (N_18169,N_17974,N_17924);
nand U18170 (N_18170,N_18062,N_18058);
nor U18171 (N_18171,N_18026,N_17972);
nor U18172 (N_18172,N_17974,N_18067);
and U18173 (N_18173,N_18031,N_18042);
nand U18174 (N_18174,N_17931,N_18061);
and U18175 (N_18175,N_17975,N_17981);
and U18176 (N_18176,N_18019,N_17980);
and U18177 (N_18177,N_17964,N_18016);
nand U18178 (N_18178,N_17936,N_17994);
nand U18179 (N_18179,N_17997,N_17965);
or U18180 (N_18180,N_18047,N_18050);
xor U18181 (N_18181,N_17954,N_18022);
nand U18182 (N_18182,N_17989,N_18036);
or U18183 (N_18183,N_17930,N_17968);
nand U18184 (N_18184,N_18038,N_18009);
nor U18185 (N_18185,N_17948,N_18056);
nand U18186 (N_18186,N_17973,N_18069);
and U18187 (N_18187,N_17942,N_17963);
or U18188 (N_18188,N_17938,N_17999);
nand U18189 (N_18189,N_18012,N_17927);
nor U18190 (N_18190,N_17998,N_18008);
and U18191 (N_18191,N_18069,N_18049);
nor U18192 (N_18192,N_18051,N_17992);
and U18193 (N_18193,N_17997,N_17921);
or U18194 (N_18194,N_18027,N_17964);
nor U18195 (N_18195,N_18031,N_17972);
or U18196 (N_18196,N_18033,N_17944);
nand U18197 (N_18197,N_18034,N_17937);
or U18198 (N_18198,N_17939,N_18006);
and U18199 (N_18199,N_17944,N_17955);
xnor U18200 (N_18200,N_17992,N_17994);
and U18201 (N_18201,N_17973,N_17923);
nand U18202 (N_18202,N_17940,N_17971);
nand U18203 (N_18203,N_17923,N_18032);
nor U18204 (N_18204,N_18016,N_18051);
or U18205 (N_18205,N_17951,N_18069);
nor U18206 (N_18206,N_17956,N_17928);
or U18207 (N_18207,N_17998,N_17988);
or U18208 (N_18208,N_18033,N_18041);
and U18209 (N_18209,N_18033,N_18062);
and U18210 (N_18210,N_17988,N_17985);
xnor U18211 (N_18211,N_17964,N_18019);
and U18212 (N_18212,N_18056,N_18009);
nand U18213 (N_18213,N_17967,N_18028);
or U18214 (N_18214,N_18020,N_17948);
xor U18215 (N_18215,N_17972,N_18028);
and U18216 (N_18216,N_17961,N_17934);
nand U18217 (N_18217,N_17927,N_18047);
nor U18218 (N_18218,N_17950,N_18006);
xor U18219 (N_18219,N_17991,N_17956);
or U18220 (N_18220,N_18076,N_18025);
and U18221 (N_18221,N_18000,N_18061);
xnor U18222 (N_18222,N_17928,N_18009);
and U18223 (N_18223,N_17955,N_17999);
nor U18224 (N_18224,N_17993,N_17937);
nor U18225 (N_18225,N_18014,N_17960);
and U18226 (N_18226,N_18044,N_18056);
or U18227 (N_18227,N_17935,N_18015);
nand U18228 (N_18228,N_18062,N_18054);
xor U18229 (N_18229,N_18003,N_18013);
nor U18230 (N_18230,N_17959,N_17974);
nand U18231 (N_18231,N_18061,N_18031);
or U18232 (N_18232,N_17931,N_17979);
and U18233 (N_18233,N_18031,N_18070);
and U18234 (N_18234,N_17981,N_18045);
and U18235 (N_18235,N_18007,N_17986);
and U18236 (N_18236,N_17923,N_17987);
nand U18237 (N_18237,N_18002,N_18051);
or U18238 (N_18238,N_17990,N_18044);
nor U18239 (N_18239,N_17921,N_17929);
nor U18240 (N_18240,N_18123,N_18080);
and U18241 (N_18241,N_18151,N_18157);
nor U18242 (N_18242,N_18212,N_18081);
nor U18243 (N_18243,N_18225,N_18236);
nand U18244 (N_18244,N_18129,N_18193);
nor U18245 (N_18245,N_18134,N_18207);
and U18246 (N_18246,N_18096,N_18156);
nand U18247 (N_18247,N_18089,N_18165);
nor U18248 (N_18248,N_18220,N_18175);
nor U18249 (N_18249,N_18106,N_18095);
nand U18250 (N_18250,N_18154,N_18121);
nor U18251 (N_18251,N_18120,N_18168);
and U18252 (N_18252,N_18094,N_18217);
nor U18253 (N_18253,N_18105,N_18166);
nand U18254 (N_18254,N_18228,N_18161);
nor U18255 (N_18255,N_18140,N_18116);
or U18256 (N_18256,N_18085,N_18122);
nor U18257 (N_18257,N_18111,N_18145);
nor U18258 (N_18258,N_18186,N_18230);
or U18259 (N_18259,N_18222,N_18127);
xnor U18260 (N_18260,N_18224,N_18206);
nor U18261 (N_18261,N_18176,N_18139);
and U18262 (N_18262,N_18097,N_18218);
nand U18263 (N_18263,N_18091,N_18083);
and U18264 (N_18264,N_18192,N_18137);
or U18265 (N_18265,N_18229,N_18103);
xor U18266 (N_18266,N_18187,N_18114);
nor U18267 (N_18267,N_18203,N_18117);
and U18268 (N_18268,N_18108,N_18188);
or U18269 (N_18269,N_18231,N_18110);
or U18270 (N_18270,N_18162,N_18178);
nor U18271 (N_18271,N_18115,N_18172);
and U18272 (N_18272,N_18164,N_18210);
nand U18273 (N_18273,N_18204,N_18142);
nand U18274 (N_18274,N_18167,N_18181);
xor U18275 (N_18275,N_18202,N_18147);
xnor U18276 (N_18276,N_18182,N_18215);
nor U18277 (N_18277,N_18112,N_18189);
xnor U18278 (N_18278,N_18087,N_18200);
and U18279 (N_18279,N_18138,N_18118);
nand U18280 (N_18280,N_18194,N_18199);
or U18281 (N_18281,N_18124,N_18128);
xnor U18282 (N_18282,N_18148,N_18102);
xnor U18283 (N_18283,N_18153,N_18100);
nor U18284 (N_18284,N_18133,N_18190);
nand U18285 (N_18285,N_18146,N_18233);
or U18286 (N_18286,N_18098,N_18159);
or U18287 (N_18287,N_18184,N_18135);
nor U18288 (N_18288,N_18234,N_18214);
nand U18289 (N_18289,N_18239,N_18082);
and U18290 (N_18290,N_18155,N_18195);
or U18291 (N_18291,N_18223,N_18136);
or U18292 (N_18292,N_18099,N_18232);
nand U18293 (N_18293,N_18113,N_18221);
nor U18294 (N_18294,N_18183,N_18160);
xor U18295 (N_18295,N_18237,N_18208);
nor U18296 (N_18296,N_18180,N_18185);
nor U18297 (N_18297,N_18173,N_18179);
or U18298 (N_18298,N_18209,N_18088);
nor U18299 (N_18299,N_18141,N_18131);
nand U18300 (N_18300,N_18092,N_18238);
nor U18301 (N_18301,N_18198,N_18093);
nand U18302 (N_18302,N_18130,N_18143);
or U18303 (N_18303,N_18084,N_18090);
nor U18304 (N_18304,N_18149,N_18174);
nand U18305 (N_18305,N_18125,N_18191);
nor U18306 (N_18306,N_18144,N_18227);
or U18307 (N_18307,N_18171,N_18177);
and U18308 (N_18308,N_18152,N_18150);
xnor U18309 (N_18309,N_18126,N_18205);
nand U18310 (N_18310,N_18101,N_18107);
nor U18311 (N_18311,N_18170,N_18201);
and U18312 (N_18312,N_18132,N_18219);
and U18313 (N_18313,N_18163,N_18104);
nor U18314 (N_18314,N_18226,N_18119);
or U18315 (N_18315,N_18235,N_18197);
and U18316 (N_18316,N_18213,N_18216);
nor U18317 (N_18317,N_18169,N_18109);
nand U18318 (N_18318,N_18158,N_18196);
or U18319 (N_18319,N_18211,N_18086);
nor U18320 (N_18320,N_18166,N_18120);
or U18321 (N_18321,N_18155,N_18091);
and U18322 (N_18322,N_18162,N_18185);
nor U18323 (N_18323,N_18164,N_18126);
xor U18324 (N_18324,N_18141,N_18184);
or U18325 (N_18325,N_18132,N_18112);
or U18326 (N_18326,N_18218,N_18105);
and U18327 (N_18327,N_18118,N_18171);
xnor U18328 (N_18328,N_18199,N_18208);
nand U18329 (N_18329,N_18129,N_18081);
nor U18330 (N_18330,N_18091,N_18115);
xor U18331 (N_18331,N_18130,N_18141);
xor U18332 (N_18332,N_18206,N_18081);
nand U18333 (N_18333,N_18096,N_18231);
or U18334 (N_18334,N_18178,N_18146);
or U18335 (N_18335,N_18195,N_18199);
or U18336 (N_18336,N_18159,N_18121);
nand U18337 (N_18337,N_18204,N_18182);
or U18338 (N_18338,N_18121,N_18149);
and U18339 (N_18339,N_18220,N_18212);
nand U18340 (N_18340,N_18083,N_18115);
nand U18341 (N_18341,N_18184,N_18122);
nor U18342 (N_18342,N_18192,N_18185);
nor U18343 (N_18343,N_18229,N_18092);
nand U18344 (N_18344,N_18118,N_18114);
nand U18345 (N_18345,N_18229,N_18196);
nand U18346 (N_18346,N_18081,N_18172);
nand U18347 (N_18347,N_18080,N_18238);
nand U18348 (N_18348,N_18130,N_18218);
xor U18349 (N_18349,N_18166,N_18178);
nand U18350 (N_18350,N_18238,N_18193);
nand U18351 (N_18351,N_18218,N_18169);
or U18352 (N_18352,N_18229,N_18237);
or U18353 (N_18353,N_18201,N_18123);
xnor U18354 (N_18354,N_18098,N_18234);
and U18355 (N_18355,N_18170,N_18175);
and U18356 (N_18356,N_18204,N_18158);
or U18357 (N_18357,N_18151,N_18220);
or U18358 (N_18358,N_18194,N_18106);
xnor U18359 (N_18359,N_18217,N_18158);
and U18360 (N_18360,N_18103,N_18194);
or U18361 (N_18361,N_18176,N_18186);
nand U18362 (N_18362,N_18239,N_18206);
and U18363 (N_18363,N_18198,N_18117);
and U18364 (N_18364,N_18143,N_18187);
nand U18365 (N_18365,N_18175,N_18205);
nand U18366 (N_18366,N_18157,N_18165);
nor U18367 (N_18367,N_18221,N_18177);
or U18368 (N_18368,N_18104,N_18081);
nand U18369 (N_18369,N_18202,N_18213);
nand U18370 (N_18370,N_18209,N_18204);
or U18371 (N_18371,N_18231,N_18111);
or U18372 (N_18372,N_18119,N_18163);
nand U18373 (N_18373,N_18100,N_18165);
and U18374 (N_18374,N_18163,N_18103);
or U18375 (N_18375,N_18145,N_18199);
nor U18376 (N_18376,N_18215,N_18214);
nor U18377 (N_18377,N_18141,N_18094);
and U18378 (N_18378,N_18151,N_18204);
nor U18379 (N_18379,N_18218,N_18226);
or U18380 (N_18380,N_18144,N_18217);
nor U18381 (N_18381,N_18216,N_18230);
nand U18382 (N_18382,N_18209,N_18099);
nor U18383 (N_18383,N_18213,N_18085);
and U18384 (N_18384,N_18109,N_18224);
nor U18385 (N_18385,N_18221,N_18213);
nand U18386 (N_18386,N_18094,N_18099);
nor U18387 (N_18387,N_18230,N_18123);
and U18388 (N_18388,N_18081,N_18122);
and U18389 (N_18389,N_18153,N_18235);
xnor U18390 (N_18390,N_18130,N_18098);
nand U18391 (N_18391,N_18119,N_18152);
or U18392 (N_18392,N_18126,N_18183);
and U18393 (N_18393,N_18182,N_18191);
and U18394 (N_18394,N_18238,N_18216);
nor U18395 (N_18395,N_18094,N_18232);
xor U18396 (N_18396,N_18233,N_18179);
nor U18397 (N_18397,N_18163,N_18129);
nor U18398 (N_18398,N_18225,N_18143);
or U18399 (N_18399,N_18234,N_18174);
nand U18400 (N_18400,N_18271,N_18397);
and U18401 (N_18401,N_18370,N_18325);
nor U18402 (N_18402,N_18259,N_18345);
nor U18403 (N_18403,N_18306,N_18398);
nor U18404 (N_18404,N_18304,N_18394);
nor U18405 (N_18405,N_18369,N_18256);
xor U18406 (N_18406,N_18268,N_18269);
nand U18407 (N_18407,N_18358,N_18287);
nor U18408 (N_18408,N_18354,N_18386);
xor U18409 (N_18409,N_18380,N_18282);
or U18410 (N_18410,N_18305,N_18260);
xor U18411 (N_18411,N_18284,N_18286);
nor U18412 (N_18412,N_18356,N_18366);
nor U18413 (N_18413,N_18254,N_18343);
and U18414 (N_18414,N_18275,N_18377);
or U18415 (N_18415,N_18292,N_18347);
nor U18416 (N_18416,N_18328,N_18303);
xnor U18417 (N_18417,N_18339,N_18374);
nand U18418 (N_18418,N_18363,N_18342);
xnor U18419 (N_18419,N_18276,N_18278);
xnor U18420 (N_18420,N_18364,N_18330);
nand U18421 (N_18421,N_18372,N_18381);
and U18422 (N_18422,N_18353,N_18373);
and U18423 (N_18423,N_18308,N_18262);
or U18424 (N_18424,N_18251,N_18296);
nand U18425 (N_18425,N_18399,N_18327);
and U18426 (N_18426,N_18310,N_18314);
or U18427 (N_18427,N_18331,N_18258);
or U18428 (N_18428,N_18361,N_18341);
nor U18429 (N_18429,N_18357,N_18273);
and U18430 (N_18430,N_18389,N_18340);
xor U18431 (N_18431,N_18244,N_18291);
or U18432 (N_18432,N_18317,N_18246);
or U18433 (N_18433,N_18352,N_18252);
or U18434 (N_18434,N_18321,N_18351);
nor U18435 (N_18435,N_18253,N_18241);
nand U18436 (N_18436,N_18240,N_18285);
or U18437 (N_18437,N_18301,N_18326);
or U18438 (N_18438,N_18318,N_18359);
and U18439 (N_18439,N_18265,N_18288);
or U18440 (N_18440,N_18379,N_18316);
nor U18441 (N_18441,N_18391,N_18333);
or U18442 (N_18442,N_18249,N_18267);
or U18443 (N_18443,N_18395,N_18309);
xnor U18444 (N_18444,N_18272,N_18360);
or U18445 (N_18445,N_18322,N_18387);
nor U18446 (N_18446,N_18384,N_18279);
nor U18447 (N_18447,N_18274,N_18293);
nand U18448 (N_18448,N_18289,N_18367);
and U18449 (N_18449,N_18255,N_18261);
xnor U18450 (N_18450,N_18297,N_18337);
nor U18451 (N_18451,N_18307,N_18248);
nor U18452 (N_18452,N_18283,N_18320);
and U18453 (N_18453,N_18266,N_18393);
and U18454 (N_18454,N_18323,N_18350);
nor U18455 (N_18455,N_18263,N_18324);
xor U18456 (N_18456,N_18243,N_18329);
nand U18457 (N_18457,N_18336,N_18281);
nand U18458 (N_18458,N_18371,N_18298);
nor U18459 (N_18459,N_18349,N_18250);
or U18460 (N_18460,N_18313,N_18396);
and U18461 (N_18461,N_18277,N_18319);
xor U18462 (N_18462,N_18245,N_18311);
and U18463 (N_18463,N_18280,N_18335);
or U18464 (N_18464,N_18385,N_18257);
nand U18465 (N_18465,N_18390,N_18315);
or U18466 (N_18466,N_18362,N_18388);
or U18467 (N_18467,N_18375,N_18348);
nor U18468 (N_18468,N_18242,N_18355);
nor U18469 (N_18469,N_18300,N_18378);
or U18470 (N_18470,N_18295,N_18294);
nor U18471 (N_18471,N_18346,N_18383);
and U18472 (N_18472,N_18392,N_18376);
or U18473 (N_18473,N_18344,N_18382);
nand U18474 (N_18474,N_18365,N_18247);
xor U18475 (N_18475,N_18270,N_18264);
and U18476 (N_18476,N_18290,N_18302);
and U18477 (N_18477,N_18334,N_18332);
and U18478 (N_18478,N_18368,N_18338);
nand U18479 (N_18479,N_18312,N_18299);
nor U18480 (N_18480,N_18245,N_18394);
or U18481 (N_18481,N_18253,N_18246);
nand U18482 (N_18482,N_18343,N_18381);
or U18483 (N_18483,N_18383,N_18292);
nor U18484 (N_18484,N_18280,N_18298);
nand U18485 (N_18485,N_18398,N_18336);
and U18486 (N_18486,N_18348,N_18383);
nand U18487 (N_18487,N_18386,N_18371);
nor U18488 (N_18488,N_18312,N_18245);
nand U18489 (N_18489,N_18323,N_18280);
and U18490 (N_18490,N_18252,N_18242);
xnor U18491 (N_18491,N_18381,N_18369);
nand U18492 (N_18492,N_18384,N_18265);
nand U18493 (N_18493,N_18311,N_18312);
xnor U18494 (N_18494,N_18318,N_18316);
or U18495 (N_18495,N_18374,N_18321);
nor U18496 (N_18496,N_18283,N_18347);
or U18497 (N_18497,N_18301,N_18298);
nand U18498 (N_18498,N_18324,N_18343);
xor U18499 (N_18499,N_18318,N_18289);
nor U18500 (N_18500,N_18320,N_18324);
nor U18501 (N_18501,N_18250,N_18280);
and U18502 (N_18502,N_18254,N_18375);
or U18503 (N_18503,N_18332,N_18297);
nand U18504 (N_18504,N_18252,N_18322);
nor U18505 (N_18505,N_18392,N_18330);
and U18506 (N_18506,N_18386,N_18332);
nand U18507 (N_18507,N_18318,N_18377);
nor U18508 (N_18508,N_18263,N_18350);
or U18509 (N_18509,N_18268,N_18287);
and U18510 (N_18510,N_18334,N_18253);
or U18511 (N_18511,N_18330,N_18256);
and U18512 (N_18512,N_18252,N_18317);
and U18513 (N_18513,N_18337,N_18330);
nor U18514 (N_18514,N_18348,N_18389);
or U18515 (N_18515,N_18318,N_18283);
nor U18516 (N_18516,N_18317,N_18382);
nand U18517 (N_18517,N_18362,N_18381);
nand U18518 (N_18518,N_18306,N_18248);
nand U18519 (N_18519,N_18315,N_18307);
xor U18520 (N_18520,N_18326,N_18366);
or U18521 (N_18521,N_18351,N_18257);
nor U18522 (N_18522,N_18348,N_18335);
nor U18523 (N_18523,N_18365,N_18328);
and U18524 (N_18524,N_18341,N_18396);
or U18525 (N_18525,N_18396,N_18247);
or U18526 (N_18526,N_18334,N_18357);
xor U18527 (N_18527,N_18387,N_18384);
nand U18528 (N_18528,N_18323,N_18249);
or U18529 (N_18529,N_18280,N_18328);
and U18530 (N_18530,N_18388,N_18271);
or U18531 (N_18531,N_18390,N_18257);
or U18532 (N_18532,N_18290,N_18348);
nor U18533 (N_18533,N_18391,N_18283);
xor U18534 (N_18534,N_18252,N_18377);
nand U18535 (N_18535,N_18373,N_18314);
nand U18536 (N_18536,N_18286,N_18397);
xnor U18537 (N_18537,N_18282,N_18317);
nor U18538 (N_18538,N_18341,N_18296);
nand U18539 (N_18539,N_18387,N_18262);
or U18540 (N_18540,N_18268,N_18355);
and U18541 (N_18541,N_18264,N_18273);
nor U18542 (N_18542,N_18373,N_18317);
nand U18543 (N_18543,N_18390,N_18389);
xnor U18544 (N_18544,N_18289,N_18282);
xor U18545 (N_18545,N_18391,N_18330);
nor U18546 (N_18546,N_18292,N_18329);
nor U18547 (N_18547,N_18250,N_18368);
or U18548 (N_18548,N_18317,N_18268);
nor U18549 (N_18549,N_18396,N_18261);
and U18550 (N_18550,N_18244,N_18378);
nor U18551 (N_18551,N_18368,N_18242);
or U18552 (N_18552,N_18244,N_18310);
or U18553 (N_18553,N_18278,N_18290);
nand U18554 (N_18554,N_18285,N_18381);
and U18555 (N_18555,N_18351,N_18339);
xor U18556 (N_18556,N_18297,N_18352);
and U18557 (N_18557,N_18364,N_18265);
and U18558 (N_18558,N_18307,N_18349);
nand U18559 (N_18559,N_18281,N_18348);
and U18560 (N_18560,N_18505,N_18465);
or U18561 (N_18561,N_18499,N_18490);
nand U18562 (N_18562,N_18492,N_18480);
nor U18563 (N_18563,N_18442,N_18557);
nand U18564 (N_18564,N_18514,N_18448);
and U18565 (N_18565,N_18417,N_18473);
and U18566 (N_18566,N_18422,N_18501);
nor U18567 (N_18567,N_18518,N_18475);
and U18568 (N_18568,N_18497,N_18504);
or U18569 (N_18569,N_18548,N_18461);
or U18570 (N_18570,N_18471,N_18459);
nor U18571 (N_18571,N_18407,N_18488);
nor U18572 (N_18572,N_18470,N_18549);
nor U18573 (N_18573,N_18424,N_18552);
and U18574 (N_18574,N_18462,N_18556);
and U18575 (N_18575,N_18520,N_18529);
or U18576 (N_18576,N_18539,N_18500);
xor U18577 (N_18577,N_18537,N_18550);
or U18578 (N_18578,N_18433,N_18412);
nor U18579 (N_18579,N_18509,N_18554);
and U18580 (N_18580,N_18401,N_18519);
and U18581 (N_18581,N_18527,N_18435);
or U18582 (N_18582,N_18430,N_18404);
or U18583 (N_18583,N_18546,N_18486);
nand U18584 (N_18584,N_18406,N_18559);
or U18585 (N_18585,N_18438,N_18436);
or U18586 (N_18586,N_18429,N_18428);
or U18587 (N_18587,N_18524,N_18493);
and U18588 (N_18588,N_18409,N_18507);
and U18589 (N_18589,N_18487,N_18542);
nand U18590 (N_18590,N_18467,N_18496);
and U18591 (N_18591,N_18513,N_18536);
and U18592 (N_18592,N_18463,N_18544);
nand U18593 (N_18593,N_18468,N_18457);
or U18594 (N_18594,N_18523,N_18474);
nor U18595 (N_18595,N_18460,N_18440);
nand U18596 (N_18596,N_18479,N_18455);
or U18597 (N_18597,N_18532,N_18489);
nor U18598 (N_18598,N_18472,N_18453);
or U18599 (N_18599,N_18528,N_18452);
nor U18600 (N_18600,N_18485,N_18434);
xnor U18601 (N_18601,N_18441,N_18454);
or U18602 (N_18602,N_18420,N_18551);
nand U18603 (N_18603,N_18477,N_18458);
nor U18604 (N_18604,N_18483,N_18426);
nand U18605 (N_18605,N_18415,N_18413);
and U18606 (N_18606,N_18494,N_18439);
nand U18607 (N_18607,N_18446,N_18405);
nor U18608 (N_18608,N_18478,N_18403);
nand U18609 (N_18609,N_18526,N_18427);
nor U18610 (N_18610,N_18450,N_18400);
nand U18611 (N_18611,N_18464,N_18444);
and U18612 (N_18612,N_18423,N_18411);
or U18613 (N_18613,N_18506,N_18540);
nand U18614 (N_18614,N_18502,N_18558);
and U18615 (N_18615,N_18437,N_18456);
or U18616 (N_18616,N_18510,N_18541);
nor U18617 (N_18617,N_18481,N_18410);
nand U18618 (N_18618,N_18445,N_18516);
or U18619 (N_18619,N_18443,N_18419);
or U18620 (N_18620,N_18495,N_18522);
nand U18621 (N_18621,N_18425,N_18431);
nor U18622 (N_18622,N_18432,N_18538);
and U18623 (N_18623,N_18466,N_18515);
nor U18624 (N_18624,N_18530,N_18531);
nor U18625 (N_18625,N_18525,N_18416);
or U18626 (N_18626,N_18508,N_18512);
nand U18627 (N_18627,N_18545,N_18534);
nand U18628 (N_18628,N_18553,N_18402);
and U18629 (N_18629,N_18511,N_18535);
xnor U18630 (N_18630,N_18484,N_18533);
xnor U18631 (N_18631,N_18555,N_18447);
nand U18632 (N_18632,N_18414,N_18451);
nor U18633 (N_18633,N_18521,N_18418);
and U18634 (N_18634,N_18543,N_18482);
or U18635 (N_18635,N_18449,N_18498);
or U18636 (N_18636,N_18469,N_18503);
nand U18637 (N_18637,N_18476,N_18517);
or U18638 (N_18638,N_18547,N_18421);
nand U18639 (N_18639,N_18408,N_18491);
nand U18640 (N_18640,N_18449,N_18484);
and U18641 (N_18641,N_18403,N_18420);
and U18642 (N_18642,N_18468,N_18535);
nor U18643 (N_18643,N_18529,N_18501);
nor U18644 (N_18644,N_18421,N_18480);
and U18645 (N_18645,N_18495,N_18524);
or U18646 (N_18646,N_18487,N_18488);
or U18647 (N_18647,N_18418,N_18533);
nand U18648 (N_18648,N_18549,N_18489);
nor U18649 (N_18649,N_18436,N_18534);
nor U18650 (N_18650,N_18501,N_18486);
and U18651 (N_18651,N_18422,N_18442);
nand U18652 (N_18652,N_18517,N_18520);
xnor U18653 (N_18653,N_18421,N_18517);
nor U18654 (N_18654,N_18424,N_18504);
or U18655 (N_18655,N_18505,N_18557);
and U18656 (N_18656,N_18513,N_18519);
or U18657 (N_18657,N_18401,N_18543);
xor U18658 (N_18658,N_18490,N_18423);
xnor U18659 (N_18659,N_18488,N_18453);
and U18660 (N_18660,N_18410,N_18528);
and U18661 (N_18661,N_18504,N_18514);
and U18662 (N_18662,N_18479,N_18445);
and U18663 (N_18663,N_18531,N_18441);
nor U18664 (N_18664,N_18495,N_18480);
and U18665 (N_18665,N_18552,N_18557);
nor U18666 (N_18666,N_18494,N_18451);
and U18667 (N_18667,N_18403,N_18458);
or U18668 (N_18668,N_18427,N_18537);
nand U18669 (N_18669,N_18460,N_18515);
and U18670 (N_18670,N_18451,N_18527);
xnor U18671 (N_18671,N_18549,N_18521);
nor U18672 (N_18672,N_18451,N_18498);
nand U18673 (N_18673,N_18506,N_18531);
xnor U18674 (N_18674,N_18539,N_18434);
or U18675 (N_18675,N_18549,N_18432);
nand U18676 (N_18676,N_18508,N_18423);
and U18677 (N_18677,N_18402,N_18528);
nand U18678 (N_18678,N_18476,N_18532);
or U18679 (N_18679,N_18440,N_18540);
or U18680 (N_18680,N_18409,N_18468);
nand U18681 (N_18681,N_18424,N_18444);
xor U18682 (N_18682,N_18472,N_18481);
and U18683 (N_18683,N_18458,N_18505);
nor U18684 (N_18684,N_18491,N_18503);
and U18685 (N_18685,N_18491,N_18469);
nand U18686 (N_18686,N_18456,N_18530);
xnor U18687 (N_18687,N_18484,N_18413);
nand U18688 (N_18688,N_18514,N_18482);
and U18689 (N_18689,N_18469,N_18526);
nand U18690 (N_18690,N_18406,N_18400);
nor U18691 (N_18691,N_18557,N_18519);
or U18692 (N_18692,N_18423,N_18446);
or U18693 (N_18693,N_18459,N_18538);
and U18694 (N_18694,N_18520,N_18428);
nand U18695 (N_18695,N_18517,N_18419);
xor U18696 (N_18696,N_18411,N_18481);
nand U18697 (N_18697,N_18519,N_18433);
and U18698 (N_18698,N_18469,N_18513);
and U18699 (N_18699,N_18554,N_18532);
or U18700 (N_18700,N_18500,N_18513);
nor U18701 (N_18701,N_18531,N_18544);
or U18702 (N_18702,N_18418,N_18482);
nor U18703 (N_18703,N_18460,N_18459);
nor U18704 (N_18704,N_18422,N_18505);
and U18705 (N_18705,N_18445,N_18515);
and U18706 (N_18706,N_18480,N_18546);
nor U18707 (N_18707,N_18552,N_18407);
and U18708 (N_18708,N_18468,N_18483);
xor U18709 (N_18709,N_18423,N_18437);
and U18710 (N_18710,N_18470,N_18540);
nor U18711 (N_18711,N_18517,N_18472);
or U18712 (N_18712,N_18551,N_18506);
nor U18713 (N_18713,N_18550,N_18439);
or U18714 (N_18714,N_18487,N_18478);
or U18715 (N_18715,N_18537,N_18548);
xnor U18716 (N_18716,N_18411,N_18554);
nand U18717 (N_18717,N_18400,N_18474);
or U18718 (N_18718,N_18446,N_18418);
and U18719 (N_18719,N_18451,N_18449);
nand U18720 (N_18720,N_18712,N_18684);
nand U18721 (N_18721,N_18675,N_18638);
nand U18722 (N_18722,N_18688,N_18600);
nand U18723 (N_18723,N_18628,N_18670);
nor U18724 (N_18724,N_18646,N_18690);
nand U18725 (N_18725,N_18652,N_18616);
or U18726 (N_18726,N_18637,N_18565);
nand U18727 (N_18727,N_18707,N_18694);
or U18728 (N_18728,N_18654,N_18626);
or U18729 (N_18729,N_18645,N_18640);
nand U18730 (N_18730,N_18629,N_18566);
nand U18731 (N_18731,N_18617,N_18580);
nor U18732 (N_18732,N_18631,N_18701);
nand U18733 (N_18733,N_18613,N_18568);
and U18734 (N_18734,N_18625,N_18714);
and U18735 (N_18735,N_18577,N_18696);
nor U18736 (N_18736,N_18705,N_18699);
nor U18737 (N_18737,N_18595,N_18676);
nor U18738 (N_18738,N_18608,N_18687);
xnor U18739 (N_18739,N_18632,N_18570);
nor U18740 (N_18740,N_18659,N_18633);
or U18741 (N_18741,N_18597,N_18717);
xnor U18742 (N_18742,N_18709,N_18643);
or U18743 (N_18743,N_18649,N_18711);
and U18744 (N_18744,N_18636,N_18661);
and U18745 (N_18745,N_18596,N_18630);
and U18746 (N_18746,N_18677,N_18569);
nand U18747 (N_18747,N_18662,N_18648);
nand U18748 (N_18748,N_18719,N_18658);
nor U18749 (N_18749,N_18679,N_18651);
nor U18750 (N_18750,N_18572,N_18612);
nor U18751 (N_18751,N_18583,N_18563);
xnor U18752 (N_18752,N_18713,N_18592);
or U18753 (N_18753,N_18601,N_18611);
or U18754 (N_18754,N_18587,N_18593);
or U18755 (N_18755,N_18634,N_18671);
nor U18756 (N_18756,N_18589,N_18599);
and U18757 (N_18757,N_18689,N_18619);
nor U18758 (N_18758,N_18698,N_18621);
nor U18759 (N_18759,N_18656,N_18678);
nor U18760 (N_18760,N_18639,N_18586);
nor U18761 (N_18761,N_18691,N_18669);
nand U18762 (N_18762,N_18703,N_18718);
or U18763 (N_18763,N_18564,N_18576);
nand U18764 (N_18764,N_18567,N_18706);
xor U18765 (N_18765,N_18604,N_18579);
and U18766 (N_18766,N_18710,N_18647);
and U18767 (N_18767,N_18561,N_18667);
and U18768 (N_18768,N_18686,N_18618);
nor U18769 (N_18769,N_18641,N_18697);
nor U18770 (N_18770,N_18578,N_18660);
nor U18771 (N_18771,N_18672,N_18598);
and U18772 (N_18772,N_18700,N_18650);
or U18773 (N_18773,N_18674,N_18642);
or U18774 (N_18774,N_18573,N_18666);
nand U18775 (N_18775,N_18644,N_18584);
nand U18776 (N_18776,N_18685,N_18664);
and U18777 (N_18777,N_18614,N_18605);
nor U18778 (N_18778,N_18581,N_18683);
nor U18779 (N_18779,N_18620,N_18708);
xor U18780 (N_18780,N_18695,N_18680);
and U18781 (N_18781,N_18574,N_18655);
and U18782 (N_18782,N_18657,N_18610);
and U18783 (N_18783,N_18585,N_18562);
or U18784 (N_18784,N_18609,N_18702);
nand U18785 (N_18785,N_18716,N_18668);
and U18786 (N_18786,N_18682,N_18704);
nor U18787 (N_18787,N_18627,N_18624);
nand U18788 (N_18788,N_18575,N_18663);
nor U18789 (N_18789,N_18615,N_18602);
and U18790 (N_18790,N_18606,N_18560);
nor U18791 (N_18791,N_18588,N_18594);
or U18792 (N_18792,N_18607,N_18665);
nor U18793 (N_18793,N_18571,N_18693);
xnor U18794 (N_18794,N_18622,N_18603);
nor U18795 (N_18795,N_18715,N_18673);
or U18796 (N_18796,N_18582,N_18591);
or U18797 (N_18797,N_18590,N_18635);
and U18798 (N_18798,N_18623,N_18692);
or U18799 (N_18799,N_18681,N_18653);
and U18800 (N_18800,N_18708,N_18661);
or U18801 (N_18801,N_18569,N_18676);
and U18802 (N_18802,N_18680,N_18716);
nand U18803 (N_18803,N_18596,N_18653);
and U18804 (N_18804,N_18676,N_18688);
xor U18805 (N_18805,N_18658,N_18718);
or U18806 (N_18806,N_18580,N_18649);
or U18807 (N_18807,N_18568,N_18572);
nor U18808 (N_18808,N_18688,N_18618);
and U18809 (N_18809,N_18665,N_18660);
or U18810 (N_18810,N_18603,N_18600);
nor U18811 (N_18811,N_18573,N_18595);
and U18812 (N_18812,N_18674,N_18581);
or U18813 (N_18813,N_18565,N_18666);
nor U18814 (N_18814,N_18573,N_18566);
xor U18815 (N_18815,N_18568,N_18623);
and U18816 (N_18816,N_18616,N_18627);
nand U18817 (N_18817,N_18618,N_18679);
nor U18818 (N_18818,N_18609,N_18591);
and U18819 (N_18819,N_18696,N_18590);
and U18820 (N_18820,N_18700,N_18609);
nand U18821 (N_18821,N_18696,N_18702);
or U18822 (N_18822,N_18716,N_18578);
xor U18823 (N_18823,N_18636,N_18589);
and U18824 (N_18824,N_18658,N_18715);
nor U18825 (N_18825,N_18602,N_18635);
nand U18826 (N_18826,N_18624,N_18630);
or U18827 (N_18827,N_18717,N_18706);
or U18828 (N_18828,N_18653,N_18591);
nand U18829 (N_18829,N_18692,N_18613);
xor U18830 (N_18830,N_18628,N_18661);
or U18831 (N_18831,N_18576,N_18570);
nand U18832 (N_18832,N_18593,N_18707);
and U18833 (N_18833,N_18694,N_18591);
and U18834 (N_18834,N_18578,N_18701);
xor U18835 (N_18835,N_18684,N_18584);
or U18836 (N_18836,N_18661,N_18611);
nor U18837 (N_18837,N_18649,N_18571);
nor U18838 (N_18838,N_18673,N_18714);
or U18839 (N_18839,N_18563,N_18614);
nand U18840 (N_18840,N_18676,N_18635);
or U18841 (N_18841,N_18630,N_18595);
nor U18842 (N_18842,N_18581,N_18695);
or U18843 (N_18843,N_18670,N_18684);
or U18844 (N_18844,N_18577,N_18621);
and U18845 (N_18845,N_18663,N_18591);
xnor U18846 (N_18846,N_18677,N_18595);
and U18847 (N_18847,N_18585,N_18667);
nor U18848 (N_18848,N_18595,N_18667);
and U18849 (N_18849,N_18677,N_18570);
and U18850 (N_18850,N_18704,N_18649);
nor U18851 (N_18851,N_18606,N_18611);
nor U18852 (N_18852,N_18621,N_18700);
nor U18853 (N_18853,N_18687,N_18639);
xor U18854 (N_18854,N_18613,N_18574);
and U18855 (N_18855,N_18596,N_18686);
or U18856 (N_18856,N_18598,N_18714);
nand U18857 (N_18857,N_18629,N_18669);
or U18858 (N_18858,N_18638,N_18577);
and U18859 (N_18859,N_18660,N_18610);
or U18860 (N_18860,N_18579,N_18590);
nor U18861 (N_18861,N_18628,N_18561);
or U18862 (N_18862,N_18695,N_18684);
nor U18863 (N_18863,N_18615,N_18573);
nor U18864 (N_18864,N_18718,N_18588);
nor U18865 (N_18865,N_18686,N_18630);
nand U18866 (N_18866,N_18601,N_18568);
nor U18867 (N_18867,N_18655,N_18648);
or U18868 (N_18868,N_18691,N_18649);
nor U18869 (N_18869,N_18602,N_18621);
xnor U18870 (N_18870,N_18608,N_18614);
nor U18871 (N_18871,N_18651,N_18648);
and U18872 (N_18872,N_18564,N_18669);
nand U18873 (N_18873,N_18641,N_18607);
or U18874 (N_18874,N_18688,N_18603);
nand U18875 (N_18875,N_18592,N_18639);
or U18876 (N_18876,N_18684,N_18701);
and U18877 (N_18877,N_18700,N_18701);
or U18878 (N_18878,N_18648,N_18609);
and U18879 (N_18879,N_18629,N_18574);
or U18880 (N_18880,N_18826,N_18749);
xnor U18881 (N_18881,N_18869,N_18729);
nand U18882 (N_18882,N_18721,N_18772);
and U18883 (N_18883,N_18738,N_18874);
nor U18884 (N_18884,N_18838,N_18816);
nand U18885 (N_18885,N_18799,N_18770);
nor U18886 (N_18886,N_18762,N_18852);
nor U18887 (N_18887,N_18846,N_18753);
or U18888 (N_18888,N_18818,N_18793);
nor U18889 (N_18889,N_18840,N_18727);
nand U18890 (N_18890,N_18875,N_18848);
nand U18891 (N_18891,N_18765,N_18742);
and U18892 (N_18892,N_18756,N_18858);
nor U18893 (N_18893,N_18853,N_18745);
nand U18894 (N_18894,N_18847,N_18833);
nand U18895 (N_18895,N_18879,N_18740);
nor U18896 (N_18896,N_18835,N_18796);
and U18897 (N_18897,N_18750,N_18873);
and U18898 (N_18898,N_18741,N_18789);
nor U18899 (N_18899,N_18820,N_18876);
and U18900 (N_18900,N_18872,N_18723);
nor U18901 (N_18901,N_18809,N_18764);
and U18902 (N_18902,N_18862,N_18828);
and U18903 (N_18903,N_18779,N_18842);
nand U18904 (N_18904,N_18851,N_18774);
nor U18905 (N_18905,N_18808,N_18868);
nand U18906 (N_18906,N_18732,N_18743);
and U18907 (N_18907,N_18763,N_18747);
and U18908 (N_18908,N_18776,N_18813);
and U18909 (N_18909,N_18758,N_18814);
nand U18910 (N_18910,N_18802,N_18806);
nand U18911 (N_18911,N_18775,N_18849);
or U18912 (N_18912,N_18746,N_18754);
nor U18913 (N_18913,N_18800,N_18739);
nor U18914 (N_18914,N_18857,N_18744);
and U18915 (N_18915,N_18850,N_18767);
nand U18916 (N_18916,N_18766,N_18819);
and U18917 (N_18917,N_18748,N_18804);
nor U18918 (N_18918,N_18830,N_18823);
or U18919 (N_18919,N_18734,N_18784);
nor U18920 (N_18920,N_18867,N_18736);
or U18921 (N_18921,N_18785,N_18812);
or U18922 (N_18922,N_18805,N_18831);
nand U18923 (N_18923,N_18788,N_18877);
nor U18924 (N_18924,N_18773,N_18854);
or U18925 (N_18925,N_18841,N_18787);
or U18926 (N_18926,N_18755,N_18803);
nor U18927 (N_18927,N_18827,N_18856);
or U18928 (N_18928,N_18777,N_18801);
or U18929 (N_18929,N_18769,N_18720);
or U18930 (N_18930,N_18728,N_18722);
nand U18931 (N_18931,N_18761,N_18798);
nand U18932 (N_18932,N_18844,N_18737);
and U18933 (N_18933,N_18837,N_18780);
nand U18934 (N_18934,N_18860,N_18815);
and U18935 (N_18935,N_18810,N_18821);
nor U18936 (N_18936,N_18825,N_18834);
xor U18937 (N_18937,N_18795,N_18822);
or U18938 (N_18938,N_18859,N_18751);
and U18939 (N_18939,N_18829,N_18878);
or U18940 (N_18940,N_18786,N_18733);
nor U18941 (N_18941,N_18730,N_18864);
nor U18942 (N_18942,N_18807,N_18861);
nor U18943 (N_18943,N_18811,N_18839);
nand U18944 (N_18944,N_18870,N_18724);
or U18945 (N_18945,N_18817,N_18781);
or U18946 (N_18946,N_18768,N_18794);
nor U18947 (N_18947,N_18845,N_18797);
and U18948 (N_18948,N_18865,N_18782);
and U18949 (N_18949,N_18771,N_18855);
and U18950 (N_18950,N_18866,N_18731);
nor U18951 (N_18951,N_18735,N_18790);
nor U18952 (N_18952,N_18792,N_18836);
and U18953 (N_18953,N_18791,N_18824);
nor U18954 (N_18954,N_18863,N_18783);
or U18955 (N_18955,N_18757,N_18759);
or U18956 (N_18956,N_18843,N_18726);
and U18957 (N_18957,N_18871,N_18760);
nand U18958 (N_18958,N_18778,N_18752);
nand U18959 (N_18959,N_18832,N_18725);
and U18960 (N_18960,N_18836,N_18745);
and U18961 (N_18961,N_18750,N_18850);
nand U18962 (N_18962,N_18733,N_18853);
nand U18963 (N_18963,N_18863,N_18806);
and U18964 (N_18964,N_18767,N_18818);
nand U18965 (N_18965,N_18738,N_18812);
and U18966 (N_18966,N_18758,N_18744);
or U18967 (N_18967,N_18876,N_18874);
and U18968 (N_18968,N_18811,N_18850);
or U18969 (N_18969,N_18804,N_18876);
nor U18970 (N_18970,N_18754,N_18835);
and U18971 (N_18971,N_18809,N_18874);
xnor U18972 (N_18972,N_18847,N_18785);
nor U18973 (N_18973,N_18879,N_18755);
and U18974 (N_18974,N_18759,N_18775);
nor U18975 (N_18975,N_18844,N_18724);
or U18976 (N_18976,N_18821,N_18750);
or U18977 (N_18977,N_18723,N_18821);
nor U18978 (N_18978,N_18832,N_18838);
xnor U18979 (N_18979,N_18742,N_18761);
nor U18980 (N_18980,N_18879,N_18811);
or U18981 (N_18981,N_18753,N_18790);
nor U18982 (N_18982,N_18770,N_18763);
and U18983 (N_18983,N_18870,N_18784);
or U18984 (N_18984,N_18726,N_18849);
nor U18985 (N_18985,N_18794,N_18738);
nand U18986 (N_18986,N_18779,N_18739);
nor U18987 (N_18987,N_18848,N_18723);
xnor U18988 (N_18988,N_18878,N_18747);
nor U18989 (N_18989,N_18841,N_18864);
and U18990 (N_18990,N_18854,N_18810);
nor U18991 (N_18991,N_18794,N_18810);
xnor U18992 (N_18992,N_18755,N_18847);
nor U18993 (N_18993,N_18774,N_18785);
nor U18994 (N_18994,N_18852,N_18817);
xor U18995 (N_18995,N_18731,N_18730);
nand U18996 (N_18996,N_18806,N_18728);
or U18997 (N_18997,N_18866,N_18822);
nor U18998 (N_18998,N_18749,N_18780);
nand U18999 (N_18999,N_18745,N_18797);
and U19000 (N_19000,N_18761,N_18721);
or U19001 (N_19001,N_18863,N_18865);
or U19002 (N_19002,N_18828,N_18806);
nand U19003 (N_19003,N_18749,N_18816);
nand U19004 (N_19004,N_18783,N_18809);
or U19005 (N_19005,N_18769,N_18748);
nand U19006 (N_19006,N_18739,N_18748);
and U19007 (N_19007,N_18740,N_18742);
nand U19008 (N_19008,N_18726,N_18796);
nor U19009 (N_19009,N_18724,N_18843);
xor U19010 (N_19010,N_18784,N_18756);
or U19011 (N_19011,N_18851,N_18766);
nor U19012 (N_19012,N_18799,N_18781);
and U19013 (N_19013,N_18790,N_18767);
nor U19014 (N_19014,N_18852,N_18850);
or U19015 (N_19015,N_18748,N_18768);
and U19016 (N_19016,N_18856,N_18798);
nor U19017 (N_19017,N_18760,N_18845);
or U19018 (N_19018,N_18821,N_18724);
nand U19019 (N_19019,N_18785,N_18872);
xnor U19020 (N_19020,N_18845,N_18771);
nand U19021 (N_19021,N_18734,N_18721);
or U19022 (N_19022,N_18837,N_18841);
and U19023 (N_19023,N_18873,N_18732);
or U19024 (N_19024,N_18767,N_18747);
and U19025 (N_19025,N_18790,N_18807);
and U19026 (N_19026,N_18806,N_18792);
nor U19027 (N_19027,N_18839,N_18792);
or U19028 (N_19028,N_18762,N_18774);
nor U19029 (N_19029,N_18862,N_18863);
or U19030 (N_19030,N_18767,N_18780);
or U19031 (N_19031,N_18805,N_18759);
nand U19032 (N_19032,N_18869,N_18788);
or U19033 (N_19033,N_18869,N_18831);
nor U19034 (N_19034,N_18810,N_18741);
nand U19035 (N_19035,N_18779,N_18798);
nor U19036 (N_19036,N_18756,N_18730);
and U19037 (N_19037,N_18853,N_18720);
and U19038 (N_19038,N_18802,N_18720);
and U19039 (N_19039,N_18844,N_18768);
and U19040 (N_19040,N_18953,N_19020);
nor U19041 (N_19041,N_18889,N_18895);
nor U19042 (N_19042,N_18899,N_18927);
nand U19043 (N_19043,N_19035,N_18974);
and U19044 (N_19044,N_18908,N_19008);
or U19045 (N_19045,N_18982,N_19019);
nand U19046 (N_19046,N_18971,N_18896);
nand U19047 (N_19047,N_18912,N_18981);
and U19048 (N_19048,N_18905,N_18938);
nand U19049 (N_19049,N_18956,N_18890);
nand U19050 (N_19050,N_18917,N_18986);
or U19051 (N_19051,N_18939,N_19014);
or U19052 (N_19052,N_18880,N_18932);
xor U19053 (N_19053,N_19003,N_18958);
or U19054 (N_19054,N_19027,N_18903);
nand U19055 (N_19055,N_18973,N_19016);
or U19056 (N_19056,N_18882,N_18921);
nor U19057 (N_19057,N_18963,N_18906);
or U19058 (N_19058,N_18943,N_18893);
nand U19059 (N_19059,N_18941,N_18944);
nor U19060 (N_19060,N_18946,N_18988);
xnor U19061 (N_19061,N_19000,N_18950);
nor U19062 (N_19062,N_19011,N_18995);
xnor U19063 (N_19063,N_18952,N_18993);
and U19064 (N_19064,N_18977,N_18891);
and U19065 (N_19065,N_18962,N_19039);
xor U19066 (N_19066,N_18936,N_19036);
or U19067 (N_19067,N_18948,N_18947);
xnor U19068 (N_19068,N_18980,N_19010);
nand U19069 (N_19069,N_18954,N_18967);
or U19070 (N_19070,N_18940,N_19017);
or U19071 (N_19071,N_18935,N_18979);
and U19072 (N_19072,N_18904,N_18918);
and U19073 (N_19073,N_18915,N_18934);
or U19074 (N_19074,N_18964,N_18928);
or U19075 (N_19075,N_18916,N_18881);
or U19076 (N_19076,N_19004,N_18955);
nand U19077 (N_19077,N_18994,N_18989);
or U19078 (N_19078,N_18976,N_18897);
nor U19079 (N_19079,N_19002,N_18922);
nor U19080 (N_19080,N_18997,N_18914);
nor U19081 (N_19081,N_18923,N_18968);
and U19082 (N_19082,N_18990,N_18898);
and U19083 (N_19083,N_19006,N_19026);
nor U19084 (N_19084,N_18961,N_18920);
and U19085 (N_19085,N_18985,N_18924);
nand U19086 (N_19086,N_18957,N_19034);
and U19087 (N_19087,N_18987,N_18886);
nor U19088 (N_19088,N_18907,N_19023);
or U19089 (N_19089,N_18929,N_18966);
xnor U19090 (N_19090,N_18998,N_19025);
or U19091 (N_19091,N_18926,N_18892);
and U19092 (N_19092,N_19001,N_18992);
nand U19093 (N_19093,N_19031,N_18960);
nand U19094 (N_19094,N_19012,N_18937);
nor U19095 (N_19095,N_19007,N_18975);
nor U19096 (N_19096,N_18909,N_19024);
nor U19097 (N_19097,N_18910,N_18991);
or U19098 (N_19098,N_18970,N_19022);
and U19099 (N_19099,N_18972,N_18965);
nor U19100 (N_19100,N_18978,N_18933);
xnor U19101 (N_19101,N_19013,N_18883);
and U19102 (N_19102,N_18931,N_19009);
or U19103 (N_19103,N_18949,N_19021);
or U19104 (N_19104,N_18959,N_18911);
nand U19105 (N_19105,N_18925,N_18930);
or U19106 (N_19106,N_18913,N_19038);
nand U19107 (N_19107,N_19037,N_19033);
and U19108 (N_19108,N_18969,N_18999);
nor U19109 (N_19109,N_19030,N_19015);
or U19110 (N_19110,N_18902,N_19028);
and U19111 (N_19111,N_18885,N_19005);
nor U19112 (N_19112,N_18888,N_19032);
and U19113 (N_19113,N_18983,N_18984);
nor U19114 (N_19114,N_18919,N_18884);
and U19115 (N_19115,N_18894,N_18945);
nand U19116 (N_19116,N_18901,N_19029);
nor U19117 (N_19117,N_19018,N_18942);
nor U19118 (N_19118,N_18951,N_18900);
xnor U19119 (N_19119,N_18887,N_18996);
and U19120 (N_19120,N_19022,N_18996);
and U19121 (N_19121,N_18934,N_18921);
nand U19122 (N_19122,N_19029,N_18957);
nor U19123 (N_19123,N_18976,N_18919);
xnor U19124 (N_19124,N_18980,N_19025);
or U19125 (N_19125,N_18959,N_18882);
xnor U19126 (N_19126,N_19003,N_18981);
and U19127 (N_19127,N_18910,N_18915);
nor U19128 (N_19128,N_18934,N_19007);
nand U19129 (N_19129,N_18966,N_19023);
nor U19130 (N_19130,N_18914,N_18928);
nor U19131 (N_19131,N_18996,N_18889);
or U19132 (N_19132,N_18912,N_19013);
xnor U19133 (N_19133,N_18891,N_18880);
and U19134 (N_19134,N_19014,N_18980);
nor U19135 (N_19135,N_18912,N_19028);
nand U19136 (N_19136,N_18955,N_18932);
or U19137 (N_19137,N_18908,N_18882);
nor U19138 (N_19138,N_18939,N_18967);
and U19139 (N_19139,N_19010,N_18965);
and U19140 (N_19140,N_18983,N_19026);
and U19141 (N_19141,N_18896,N_18957);
and U19142 (N_19142,N_18900,N_18977);
or U19143 (N_19143,N_18971,N_18962);
or U19144 (N_19144,N_19025,N_18991);
and U19145 (N_19145,N_18945,N_19037);
and U19146 (N_19146,N_18980,N_19037);
nand U19147 (N_19147,N_18931,N_18898);
or U19148 (N_19148,N_18895,N_18970);
nand U19149 (N_19149,N_18980,N_18908);
xor U19150 (N_19150,N_19008,N_18986);
nor U19151 (N_19151,N_19004,N_18935);
or U19152 (N_19152,N_19007,N_18955);
nor U19153 (N_19153,N_18950,N_19026);
or U19154 (N_19154,N_18998,N_18890);
xor U19155 (N_19155,N_18946,N_18917);
nand U19156 (N_19156,N_18894,N_19018);
nand U19157 (N_19157,N_18956,N_19018);
and U19158 (N_19158,N_19021,N_19007);
nand U19159 (N_19159,N_18926,N_18967);
or U19160 (N_19160,N_19007,N_18900);
nand U19161 (N_19161,N_18952,N_18942);
or U19162 (N_19162,N_18944,N_18884);
or U19163 (N_19163,N_18937,N_18917);
and U19164 (N_19164,N_18984,N_19036);
nor U19165 (N_19165,N_18927,N_18958);
or U19166 (N_19166,N_18883,N_18962);
nor U19167 (N_19167,N_19030,N_18978);
or U19168 (N_19168,N_18976,N_19025);
xor U19169 (N_19169,N_18919,N_18939);
nand U19170 (N_19170,N_18972,N_19026);
nor U19171 (N_19171,N_18901,N_18911);
or U19172 (N_19172,N_18895,N_18993);
and U19173 (N_19173,N_18947,N_18903);
nand U19174 (N_19174,N_18954,N_18913);
xnor U19175 (N_19175,N_18913,N_18925);
nor U19176 (N_19176,N_19004,N_18942);
nand U19177 (N_19177,N_19003,N_18934);
and U19178 (N_19178,N_18910,N_18954);
or U19179 (N_19179,N_18908,N_18890);
or U19180 (N_19180,N_19013,N_18991);
nand U19181 (N_19181,N_18988,N_19013);
and U19182 (N_19182,N_18923,N_19006);
nand U19183 (N_19183,N_18915,N_18914);
and U19184 (N_19184,N_18958,N_18992);
nand U19185 (N_19185,N_18893,N_19031);
nor U19186 (N_19186,N_19002,N_18884);
nor U19187 (N_19187,N_18992,N_18982);
and U19188 (N_19188,N_18888,N_19008);
or U19189 (N_19189,N_18997,N_18889);
or U19190 (N_19190,N_19025,N_18930);
nand U19191 (N_19191,N_18929,N_18928);
and U19192 (N_19192,N_18888,N_18897);
and U19193 (N_19193,N_18992,N_18951);
nor U19194 (N_19194,N_18947,N_19000);
nor U19195 (N_19195,N_18946,N_18937);
and U19196 (N_19196,N_18990,N_18885);
nor U19197 (N_19197,N_18899,N_18911);
and U19198 (N_19198,N_18929,N_18989);
and U19199 (N_19199,N_18920,N_18898);
nand U19200 (N_19200,N_19187,N_19130);
nand U19201 (N_19201,N_19118,N_19040);
and U19202 (N_19202,N_19112,N_19160);
nor U19203 (N_19203,N_19168,N_19199);
nand U19204 (N_19204,N_19133,N_19075);
or U19205 (N_19205,N_19107,N_19183);
nand U19206 (N_19206,N_19152,N_19177);
nor U19207 (N_19207,N_19116,N_19179);
nand U19208 (N_19208,N_19140,N_19041);
or U19209 (N_19209,N_19084,N_19093);
nand U19210 (N_19210,N_19091,N_19135);
or U19211 (N_19211,N_19131,N_19182);
nand U19212 (N_19212,N_19198,N_19074);
or U19213 (N_19213,N_19127,N_19057);
xor U19214 (N_19214,N_19174,N_19097);
nand U19215 (N_19215,N_19145,N_19154);
nand U19216 (N_19216,N_19186,N_19143);
nand U19217 (N_19217,N_19159,N_19132);
nand U19218 (N_19218,N_19071,N_19088);
nor U19219 (N_19219,N_19119,N_19122);
or U19220 (N_19220,N_19111,N_19173);
nor U19221 (N_19221,N_19063,N_19163);
and U19222 (N_19222,N_19157,N_19099);
nor U19223 (N_19223,N_19167,N_19114);
nor U19224 (N_19224,N_19060,N_19108);
or U19225 (N_19225,N_19089,N_19136);
nand U19226 (N_19226,N_19066,N_19103);
nor U19227 (N_19227,N_19050,N_19062);
or U19228 (N_19228,N_19138,N_19086);
nand U19229 (N_19229,N_19148,N_19059);
and U19230 (N_19230,N_19139,N_19101);
and U19231 (N_19231,N_19121,N_19115);
nor U19232 (N_19232,N_19065,N_19072);
and U19233 (N_19233,N_19082,N_19109);
or U19234 (N_19234,N_19105,N_19067);
xor U19235 (N_19235,N_19172,N_19195);
nor U19236 (N_19236,N_19164,N_19098);
nand U19237 (N_19237,N_19181,N_19092);
nor U19238 (N_19238,N_19197,N_19077);
nand U19239 (N_19239,N_19106,N_19129);
and U19240 (N_19240,N_19087,N_19046);
and U19241 (N_19241,N_19144,N_19042);
nand U19242 (N_19242,N_19166,N_19155);
nor U19243 (N_19243,N_19128,N_19069);
xnor U19244 (N_19244,N_19078,N_19095);
nand U19245 (N_19245,N_19176,N_19044);
nand U19246 (N_19246,N_19094,N_19061);
and U19247 (N_19247,N_19170,N_19171);
nand U19248 (N_19248,N_19178,N_19070);
and U19249 (N_19249,N_19096,N_19151);
or U19250 (N_19250,N_19117,N_19068);
or U19251 (N_19251,N_19189,N_19162);
and U19252 (N_19252,N_19158,N_19083);
or U19253 (N_19253,N_19055,N_19169);
xor U19254 (N_19254,N_19193,N_19054);
or U19255 (N_19255,N_19142,N_19045);
nor U19256 (N_19256,N_19146,N_19051);
or U19257 (N_19257,N_19100,N_19110);
nor U19258 (N_19258,N_19156,N_19104);
nor U19259 (N_19259,N_19102,N_19196);
and U19260 (N_19260,N_19052,N_19149);
nor U19261 (N_19261,N_19076,N_19161);
xor U19262 (N_19262,N_19126,N_19085);
and U19263 (N_19263,N_19184,N_19079);
or U19264 (N_19264,N_19056,N_19113);
and U19265 (N_19265,N_19153,N_19190);
or U19266 (N_19266,N_19192,N_19194);
and U19267 (N_19267,N_19049,N_19165);
nand U19268 (N_19268,N_19125,N_19064);
xnor U19269 (N_19269,N_19185,N_19080);
nor U19270 (N_19270,N_19073,N_19134);
nor U19271 (N_19271,N_19058,N_19120);
and U19272 (N_19272,N_19081,N_19147);
xnor U19273 (N_19273,N_19137,N_19150);
xnor U19274 (N_19274,N_19047,N_19123);
or U19275 (N_19275,N_19043,N_19180);
and U19276 (N_19276,N_19053,N_19141);
and U19277 (N_19277,N_19175,N_19191);
xnor U19278 (N_19278,N_19124,N_19188);
nand U19279 (N_19279,N_19048,N_19090);
nor U19280 (N_19280,N_19113,N_19129);
and U19281 (N_19281,N_19173,N_19165);
or U19282 (N_19282,N_19160,N_19139);
and U19283 (N_19283,N_19052,N_19159);
and U19284 (N_19284,N_19195,N_19171);
nand U19285 (N_19285,N_19199,N_19046);
and U19286 (N_19286,N_19128,N_19171);
and U19287 (N_19287,N_19173,N_19125);
nand U19288 (N_19288,N_19071,N_19055);
nand U19289 (N_19289,N_19141,N_19157);
nor U19290 (N_19290,N_19187,N_19071);
or U19291 (N_19291,N_19159,N_19055);
and U19292 (N_19292,N_19069,N_19165);
and U19293 (N_19293,N_19097,N_19172);
or U19294 (N_19294,N_19070,N_19060);
or U19295 (N_19295,N_19157,N_19121);
nand U19296 (N_19296,N_19120,N_19042);
nand U19297 (N_19297,N_19127,N_19101);
nor U19298 (N_19298,N_19170,N_19077);
nand U19299 (N_19299,N_19189,N_19132);
nand U19300 (N_19300,N_19145,N_19056);
nand U19301 (N_19301,N_19168,N_19127);
or U19302 (N_19302,N_19110,N_19158);
and U19303 (N_19303,N_19057,N_19094);
and U19304 (N_19304,N_19093,N_19142);
xnor U19305 (N_19305,N_19115,N_19145);
nand U19306 (N_19306,N_19047,N_19128);
nand U19307 (N_19307,N_19070,N_19198);
nand U19308 (N_19308,N_19041,N_19177);
nand U19309 (N_19309,N_19128,N_19071);
xnor U19310 (N_19310,N_19108,N_19143);
and U19311 (N_19311,N_19165,N_19078);
nand U19312 (N_19312,N_19053,N_19187);
nor U19313 (N_19313,N_19161,N_19174);
nand U19314 (N_19314,N_19097,N_19048);
nand U19315 (N_19315,N_19174,N_19181);
and U19316 (N_19316,N_19137,N_19182);
and U19317 (N_19317,N_19147,N_19158);
nand U19318 (N_19318,N_19079,N_19181);
nor U19319 (N_19319,N_19182,N_19127);
nor U19320 (N_19320,N_19142,N_19118);
nand U19321 (N_19321,N_19084,N_19175);
nand U19322 (N_19322,N_19116,N_19055);
xor U19323 (N_19323,N_19175,N_19092);
xnor U19324 (N_19324,N_19104,N_19183);
nor U19325 (N_19325,N_19181,N_19185);
nand U19326 (N_19326,N_19063,N_19123);
and U19327 (N_19327,N_19145,N_19111);
nand U19328 (N_19328,N_19126,N_19044);
or U19329 (N_19329,N_19178,N_19064);
nor U19330 (N_19330,N_19133,N_19068);
nor U19331 (N_19331,N_19189,N_19122);
and U19332 (N_19332,N_19153,N_19128);
or U19333 (N_19333,N_19134,N_19195);
nand U19334 (N_19334,N_19098,N_19112);
nor U19335 (N_19335,N_19130,N_19123);
and U19336 (N_19336,N_19105,N_19118);
and U19337 (N_19337,N_19073,N_19048);
and U19338 (N_19338,N_19156,N_19121);
and U19339 (N_19339,N_19128,N_19155);
nand U19340 (N_19340,N_19134,N_19127);
and U19341 (N_19341,N_19043,N_19159);
nor U19342 (N_19342,N_19153,N_19183);
nand U19343 (N_19343,N_19079,N_19104);
nand U19344 (N_19344,N_19048,N_19044);
and U19345 (N_19345,N_19162,N_19066);
nor U19346 (N_19346,N_19168,N_19116);
xor U19347 (N_19347,N_19069,N_19088);
or U19348 (N_19348,N_19082,N_19073);
nor U19349 (N_19349,N_19178,N_19052);
or U19350 (N_19350,N_19099,N_19072);
nand U19351 (N_19351,N_19051,N_19115);
and U19352 (N_19352,N_19150,N_19116);
or U19353 (N_19353,N_19137,N_19116);
nand U19354 (N_19354,N_19097,N_19094);
or U19355 (N_19355,N_19091,N_19120);
or U19356 (N_19356,N_19130,N_19089);
nor U19357 (N_19357,N_19087,N_19193);
nand U19358 (N_19358,N_19147,N_19073);
and U19359 (N_19359,N_19192,N_19118);
nand U19360 (N_19360,N_19321,N_19224);
or U19361 (N_19361,N_19200,N_19314);
and U19362 (N_19362,N_19211,N_19351);
and U19363 (N_19363,N_19246,N_19346);
and U19364 (N_19364,N_19257,N_19332);
or U19365 (N_19365,N_19250,N_19236);
xnor U19366 (N_19366,N_19223,N_19291);
nand U19367 (N_19367,N_19359,N_19288);
nand U19368 (N_19368,N_19210,N_19304);
nor U19369 (N_19369,N_19278,N_19286);
nor U19370 (N_19370,N_19281,N_19222);
and U19371 (N_19371,N_19338,N_19245);
nor U19372 (N_19372,N_19285,N_19225);
nor U19373 (N_19373,N_19267,N_19289);
nor U19374 (N_19374,N_19259,N_19331);
nand U19375 (N_19375,N_19202,N_19238);
nand U19376 (N_19376,N_19269,N_19319);
nand U19377 (N_19377,N_19248,N_19204);
and U19378 (N_19378,N_19303,N_19237);
nand U19379 (N_19379,N_19320,N_19240);
nor U19380 (N_19380,N_19214,N_19293);
xor U19381 (N_19381,N_19283,N_19294);
xor U19382 (N_19382,N_19284,N_19229);
nand U19383 (N_19383,N_19255,N_19335);
and U19384 (N_19384,N_19274,N_19266);
xor U19385 (N_19385,N_19242,N_19308);
or U19386 (N_19386,N_19231,N_19219);
nand U19387 (N_19387,N_19203,N_19279);
nor U19388 (N_19388,N_19352,N_19356);
nand U19389 (N_19389,N_19207,N_19349);
nor U19390 (N_19390,N_19340,N_19318);
nor U19391 (N_19391,N_19296,N_19230);
and U19392 (N_19392,N_19232,N_19301);
nand U19393 (N_19393,N_19233,N_19307);
or U19394 (N_19394,N_19208,N_19333);
nor U19395 (N_19395,N_19260,N_19317);
nor U19396 (N_19396,N_19227,N_19268);
nand U19397 (N_19397,N_19276,N_19239);
nand U19398 (N_19398,N_19287,N_19300);
nand U19399 (N_19399,N_19309,N_19217);
nand U19400 (N_19400,N_19218,N_19310);
or U19401 (N_19401,N_19323,N_19249);
nand U19402 (N_19402,N_19221,N_19280);
nand U19403 (N_19403,N_19215,N_19305);
nand U19404 (N_19404,N_19220,N_19213);
nor U19405 (N_19405,N_19264,N_19252);
nor U19406 (N_19406,N_19348,N_19243);
and U19407 (N_19407,N_19292,N_19358);
or U19408 (N_19408,N_19295,N_19302);
and U19409 (N_19409,N_19322,N_19235);
nor U19410 (N_19410,N_19330,N_19312);
nor U19411 (N_19411,N_19251,N_19342);
or U19412 (N_19412,N_19272,N_19345);
and U19413 (N_19413,N_19315,N_19355);
or U19414 (N_19414,N_19337,N_19298);
or U19415 (N_19415,N_19339,N_19341);
or U19416 (N_19416,N_19328,N_19270);
or U19417 (N_19417,N_19316,N_19297);
and U19418 (N_19418,N_19347,N_19212);
and U19419 (N_19419,N_19247,N_19265);
nand U19420 (N_19420,N_19226,N_19326);
or U19421 (N_19421,N_19258,N_19273);
and U19422 (N_19422,N_19313,N_19353);
nand U19423 (N_19423,N_19216,N_19311);
nand U19424 (N_19424,N_19275,N_19290);
or U19425 (N_19425,N_19306,N_19357);
nor U19426 (N_19426,N_19253,N_19325);
xnor U19427 (N_19427,N_19244,N_19261);
nand U19428 (N_19428,N_19350,N_19282);
or U19429 (N_19429,N_19329,N_19241);
and U19430 (N_19430,N_19324,N_19256);
nand U19431 (N_19431,N_19201,N_19205);
xnor U19432 (N_19432,N_19354,N_19299);
and U19433 (N_19433,N_19343,N_19262);
or U19434 (N_19434,N_19327,N_19209);
or U19435 (N_19435,N_19206,N_19263);
or U19436 (N_19436,N_19254,N_19344);
and U19437 (N_19437,N_19234,N_19336);
or U19438 (N_19438,N_19334,N_19277);
nor U19439 (N_19439,N_19271,N_19228);
or U19440 (N_19440,N_19202,N_19321);
nand U19441 (N_19441,N_19314,N_19295);
and U19442 (N_19442,N_19246,N_19253);
and U19443 (N_19443,N_19305,N_19284);
nor U19444 (N_19444,N_19212,N_19270);
nor U19445 (N_19445,N_19284,N_19213);
nor U19446 (N_19446,N_19264,N_19232);
and U19447 (N_19447,N_19332,N_19298);
nor U19448 (N_19448,N_19282,N_19204);
or U19449 (N_19449,N_19329,N_19248);
nand U19450 (N_19450,N_19259,N_19216);
nor U19451 (N_19451,N_19339,N_19325);
nor U19452 (N_19452,N_19213,N_19334);
nor U19453 (N_19453,N_19303,N_19308);
or U19454 (N_19454,N_19239,N_19296);
and U19455 (N_19455,N_19266,N_19200);
xnor U19456 (N_19456,N_19312,N_19267);
xnor U19457 (N_19457,N_19270,N_19223);
nand U19458 (N_19458,N_19301,N_19273);
and U19459 (N_19459,N_19238,N_19327);
and U19460 (N_19460,N_19231,N_19261);
and U19461 (N_19461,N_19314,N_19268);
xnor U19462 (N_19462,N_19320,N_19256);
nor U19463 (N_19463,N_19229,N_19274);
and U19464 (N_19464,N_19284,N_19337);
or U19465 (N_19465,N_19227,N_19229);
or U19466 (N_19466,N_19215,N_19353);
nand U19467 (N_19467,N_19271,N_19237);
or U19468 (N_19468,N_19314,N_19310);
nand U19469 (N_19469,N_19200,N_19225);
xor U19470 (N_19470,N_19222,N_19350);
nand U19471 (N_19471,N_19340,N_19217);
nand U19472 (N_19472,N_19315,N_19357);
or U19473 (N_19473,N_19279,N_19213);
or U19474 (N_19474,N_19332,N_19200);
xor U19475 (N_19475,N_19259,N_19264);
or U19476 (N_19476,N_19281,N_19227);
nor U19477 (N_19477,N_19325,N_19351);
or U19478 (N_19478,N_19337,N_19225);
nand U19479 (N_19479,N_19283,N_19215);
xnor U19480 (N_19480,N_19251,N_19288);
and U19481 (N_19481,N_19328,N_19299);
and U19482 (N_19482,N_19265,N_19332);
xnor U19483 (N_19483,N_19221,N_19308);
xnor U19484 (N_19484,N_19249,N_19244);
and U19485 (N_19485,N_19298,N_19213);
nand U19486 (N_19486,N_19269,N_19294);
nand U19487 (N_19487,N_19231,N_19279);
and U19488 (N_19488,N_19203,N_19240);
nand U19489 (N_19489,N_19349,N_19265);
and U19490 (N_19490,N_19347,N_19349);
or U19491 (N_19491,N_19256,N_19331);
nand U19492 (N_19492,N_19228,N_19320);
nand U19493 (N_19493,N_19318,N_19212);
nand U19494 (N_19494,N_19250,N_19203);
or U19495 (N_19495,N_19210,N_19334);
and U19496 (N_19496,N_19345,N_19233);
nand U19497 (N_19497,N_19204,N_19236);
nor U19498 (N_19498,N_19292,N_19324);
or U19499 (N_19499,N_19231,N_19245);
nand U19500 (N_19500,N_19302,N_19275);
xnor U19501 (N_19501,N_19307,N_19338);
or U19502 (N_19502,N_19262,N_19280);
and U19503 (N_19503,N_19330,N_19215);
nor U19504 (N_19504,N_19210,N_19351);
and U19505 (N_19505,N_19233,N_19255);
or U19506 (N_19506,N_19333,N_19318);
and U19507 (N_19507,N_19270,N_19235);
nand U19508 (N_19508,N_19320,N_19237);
xnor U19509 (N_19509,N_19296,N_19233);
or U19510 (N_19510,N_19232,N_19317);
nand U19511 (N_19511,N_19233,N_19299);
and U19512 (N_19512,N_19326,N_19244);
nand U19513 (N_19513,N_19250,N_19311);
nand U19514 (N_19514,N_19273,N_19235);
or U19515 (N_19515,N_19209,N_19229);
xor U19516 (N_19516,N_19242,N_19328);
nand U19517 (N_19517,N_19330,N_19347);
nand U19518 (N_19518,N_19345,N_19310);
or U19519 (N_19519,N_19281,N_19308);
nand U19520 (N_19520,N_19402,N_19438);
nor U19521 (N_19521,N_19365,N_19509);
and U19522 (N_19522,N_19418,N_19369);
nor U19523 (N_19523,N_19493,N_19364);
nor U19524 (N_19524,N_19447,N_19412);
xnor U19525 (N_19525,N_19479,N_19496);
and U19526 (N_19526,N_19472,N_19395);
or U19527 (N_19527,N_19443,N_19486);
nand U19528 (N_19528,N_19373,N_19441);
nor U19529 (N_19529,N_19360,N_19382);
and U19530 (N_19530,N_19390,N_19453);
and U19531 (N_19531,N_19424,N_19454);
nor U19532 (N_19532,N_19475,N_19466);
or U19533 (N_19533,N_19393,N_19425);
or U19534 (N_19534,N_19515,N_19445);
nor U19535 (N_19535,N_19405,N_19435);
and U19536 (N_19536,N_19476,N_19506);
nor U19537 (N_19537,N_19397,N_19362);
and U19538 (N_19538,N_19498,N_19474);
and U19539 (N_19539,N_19450,N_19419);
and U19540 (N_19540,N_19470,N_19518);
nor U19541 (N_19541,N_19366,N_19497);
xnor U19542 (N_19542,N_19489,N_19361);
xor U19543 (N_19543,N_19514,N_19370);
nor U19544 (N_19544,N_19451,N_19483);
or U19545 (N_19545,N_19421,N_19380);
and U19546 (N_19546,N_19417,N_19494);
and U19547 (N_19547,N_19457,N_19481);
or U19548 (N_19548,N_19444,N_19446);
and U19549 (N_19549,N_19378,N_19388);
nor U19550 (N_19550,N_19409,N_19491);
xnor U19551 (N_19551,N_19389,N_19376);
nor U19552 (N_19552,N_19487,N_19392);
or U19553 (N_19553,N_19480,N_19400);
nand U19554 (N_19554,N_19504,N_19456);
xnor U19555 (N_19555,N_19440,N_19478);
nor U19556 (N_19556,N_19463,N_19387);
nand U19557 (N_19557,N_19379,N_19398);
nand U19558 (N_19558,N_19368,N_19465);
and U19559 (N_19559,N_19371,N_19508);
and U19560 (N_19560,N_19415,N_19516);
nand U19561 (N_19561,N_19381,N_19439);
nor U19562 (N_19562,N_19458,N_19482);
and U19563 (N_19563,N_19473,N_19407);
nor U19564 (N_19564,N_19452,N_19459);
and U19565 (N_19565,N_19455,N_19488);
nor U19566 (N_19566,N_19414,N_19499);
or U19567 (N_19567,N_19468,N_19495);
nor U19568 (N_19568,N_19490,N_19375);
or U19569 (N_19569,N_19374,N_19436);
nor U19570 (N_19570,N_19507,N_19385);
or U19571 (N_19571,N_19512,N_19437);
and U19572 (N_19572,N_19384,N_19433);
or U19573 (N_19573,N_19372,N_19430);
nand U19574 (N_19574,N_19428,N_19461);
or U19575 (N_19575,N_19517,N_19403);
xor U19576 (N_19576,N_19404,N_19484);
xnor U19577 (N_19577,N_19426,N_19442);
and U19578 (N_19578,N_19501,N_19485);
and U19579 (N_19579,N_19422,N_19396);
or U19580 (N_19580,N_19411,N_19502);
nand U19581 (N_19581,N_19410,N_19431);
or U19582 (N_19582,N_19367,N_19416);
nand U19583 (N_19583,N_19505,N_19429);
and U19584 (N_19584,N_19519,N_19408);
and U19585 (N_19585,N_19406,N_19469);
nor U19586 (N_19586,N_19503,N_19511);
and U19587 (N_19587,N_19510,N_19432);
or U19588 (N_19588,N_19500,N_19449);
nor U19589 (N_19589,N_19460,N_19363);
nand U19590 (N_19590,N_19413,N_19471);
nand U19591 (N_19591,N_19427,N_19477);
nor U19592 (N_19592,N_19420,N_19383);
or U19593 (N_19593,N_19464,N_19386);
nor U19594 (N_19594,N_19448,N_19492);
and U19595 (N_19595,N_19423,N_19513);
nor U19596 (N_19596,N_19394,N_19399);
nand U19597 (N_19597,N_19391,N_19434);
and U19598 (N_19598,N_19467,N_19377);
xor U19599 (N_19599,N_19401,N_19462);
and U19600 (N_19600,N_19516,N_19379);
or U19601 (N_19601,N_19438,N_19457);
and U19602 (N_19602,N_19394,N_19456);
nor U19603 (N_19603,N_19392,N_19490);
nand U19604 (N_19604,N_19440,N_19411);
and U19605 (N_19605,N_19429,N_19513);
or U19606 (N_19606,N_19491,N_19485);
nand U19607 (N_19607,N_19361,N_19422);
nor U19608 (N_19608,N_19497,N_19491);
nor U19609 (N_19609,N_19404,N_19475);
or U19610 (N_19610,N_19484,N_19483);
nor U19611 (N_19611,N_19421,N_19400);
nand U19612 (N_19612,N_19474,N_19417);
nor U19613 (N_19613,N_19513,N_19449);
or U19614 (N_19614,N_19450,N_19519);
and U19615 (N_19615,N_19498,N_19389);
and U19616 (N_19616,N_19434,N_19513);
or U19617 (N_19617,N_19498,N_19486);
nand U19618 (N_19618,N_19464,N_19475);
or U19619 (N_19619,N_19480,N_19376);
nand U19620 (N_19620,N_19413,N_19411);
and U19621 (N_19621,N_19392,N_19404);
xor U19622 (N_19622,N_19497,N_19452);
nor U19623 (N_19623,N_19467,N_19366);
nor U19624 (N_19624,N_19407,N_19382);
or U19625 (N_19625,N_19474,N_19467);
or U19626 (N_19626,N_19439,N_19402);
nor U19627 (N_19627,N_19388,N_19443);
nand U19628 (N_19628,N_19387,N_19482);
nor U19629 (N_19629,N_19491,N_19394);
nand U19630 (N_19630,N_19372,N_19485);
and U19631 (N_19631,N_19426,N_19456);
nor U19632 (N_19632,N_19418,N_19397);
nor U19633 (N_19633,N_19440,N_19461);
and U19634 (N_19634,N_19465,N_19503);
nand U19635 (N_19635,N_19418,N_19502);
nand U19636 (N_19636,N_19461,N_19518);
nand U19637 (N_19637,N_19395,N_19432);
or U19638 (N_19638,N_19438,N_19415);
nor U19639 (N_19639,N_19440,N_19415);
and U19640 (N_19640,N_19483,N_19427);
nor U19641 (N_19641,N_19452,N_19430);
nand U19642 (N_19642,N_19394,N_19362);
and U19643 (N_19643,N_19452,N_19367);
and U19644 (N_19644,N_19405,N_19362);
nor U19645 (N_19645,N_19418,N_19387);
nand U19646 (N_19646,N_19419,N_19455);
xnor U19647 (N_19647,N_19493,N_19384);
and U19648 (N_19648,N_19502,N_19399);
nand U19649 (N_19649,N_19467,N_19380);
xnor U19650 (N_19650,N_19397,N_19505);
and U19651 (N_19651,N_19505,N_19421);
xor U19652 (N_19652,N_19459,N_19505);
nand U19653 (N_19653,N_19506,N_19430);
or U19654 (N_19654,N_19400,N_19408);
nor U19655 (N_19655,N_19462,N_19506);
and U19656 (N_19656,N_19476,N_19492);
and U19657 (N_19657,N_19439,N_19362);
xor U19658 (N_19658,N_19512,N_19371);
xor U19659 (N_19659,N_19434,N_19510);
and U19660 (N_19660,N_19405,N_19417);
xnor U19661 (N_19661,N_19371,N_19495);
or U19662 (N_19662,N_19385,N_19479);
nor U19663 (N_19663,N_19380,N_19427);
and U19664 (N_19664,N_19434,N_19371);
xnor U19665 (N_19665,N_19452,N_19496);
xor U19666 (N_19666,N_19505,N_19475);
xnor U19667 (N_19667,N_19437,N_19507);
nand U19668 (N_19668,N_19460,N_19375);
nand U19669 (N_19669,N_19375,N_19402);
or U19670 (N_19670,N_19361,N_19404);
or U19671 (N_19671,N_19457,N_19421);
nand U19672 (N_19672,N_19475,N_19379);
and U19673 (N_19673,N_19396,N_19439);
and U19674 (N_19674,N_19494,N_19467);
and U19675 (N_19675,N_19434,N_19451);
nor U19676 (N_19676,N_19518,N_19500);
or U19677 (N_19677,N_19517,N_19410);
and U19678 (N_19678,N_19503,N_19490);
nor U19679 (N_19679,N_19382,N_19413);
or U19680 (N_19680,N_19579,N_19648);
nor U19681 (N_19681,N_19584,N_19520);
and U19682 (N_19682,N_19548,N_19661);
or U19683 (N_19683,N_19676,N_19652);
or U19684 (N_19684,N_19670,N_19575);
or U19685 (N_19685,N_19630,N_19620);
and U19686 (N_19686,N_19567,N_19605);
xnor U19687 (N_19687,N_19591,N_19558);
xor U19688 (N_19688,N_19538,N_19641);
nand U19689 (N_19689,N_19629,N_19562);
and U19690 (N_19690,N_19565,N_19613);
and U19691 (N_19691,N_19573,N_19649);
nand U19692 (N_19692,N_19570,N_19559);
nand U19693 (N_19693,N_19619,N_19590);
nor U19694 (N_19694,N_19626,N_19617);
nand U19695 (N_19695,N_19608,N_19669);
or U19696 (N_19696,N_19666,N_19677);
nand U19697 (N_19697,N_19533,N_19664);
xor U19698 (N_19698,N_19580,N_19654);
nor U19699 (N_19699,N_19609,N_19655);
nand U19700 (N_19700,N_19529,N_19586);
or U19701 (N_19701,N_19540,N_19600);
nand U19702 (N_19702,N_19554,N_19663);
and U19703 (N_19703,N_19588,N_19632);
and U19704 (N_19704,N_19544,N_19571);
xnor U19705 (N_19705,N_19633,N_19640);
or U19706 (N_19706,N_19622,N_19612);
xnor U19707 (N_19707,N_19594,N_19522);
xnor U19708 (N_19708,N_19610,N_19539);
nand U19709 (N_19709,N_19524,N_19595);
nand U19710 (N_19710,N_19563,N_19531);
and U19711 (N_19711,N_19525,N_19592);
xor U19712 (N_19712,N_19625,N_19541);
or U19713 (N_19713,N_19534,N_19657);
nand U19714 (N_19714,N_19599,N_19547);
or U19715 (N_19715,N_19583,N_19639);
nor U19716 (N_19716,N_19582,N_19659);
nor U19717 (N_19717,N_19611,N_19653);
or U19718 (N_19718,N_19574,N_19650);
or U19719 (N_19719,N_19556,N_19673);
nor U19720 (N_19720,N_19589,N_19624);
xor U19721 (N_19721,N_19614,N_19621);
and U19722 (N_19722,N_19668,N_19667);
and U19723 (N_19723,N_19658,N_19618);
nor U19724 (N_19724,N_19660,N_19555);
nand U19725 (N_19725,N_19530,N_19572);
nor U19726 (N_19726,N_19552,N_19535);
and U19727 (N_19727,N_19585,N_19627);
and U19728 (N_19728,N_19606,N_19581);
xor U19729 (N_19729,N_19638,N_19662);
or U19730 (N_19730,N_19631,N_19577);
nand U19731 (N_19731,N_19623,N_19647);
nand U19732 (N_19732,N_19532,N_19560);
or U19733 (N_19733,N_19578,N_19542);
nor U19734 (N_19734,N_19665,N_19587);
nand U19735 (N_19735,N_19527,N_19615);
nand U19736 (N_19736,N_19550,N_19651);
and U19737 (N_19737,N_19616,N_19642);
nand U19738 (N_19738,N_19566,N_19646);
nor U19739 (N_19739,N_19569,N_19549);
nor U19740 (N_19740,N_19593,N_19671);
nand U19741 (N_19741,N_19568,N_19545);
nand U19742 (N_19742,N_19536,N_19526);
and U19743 (N_19743,N_19678,N_19645);
nand U19744 (N_19744,N_19603,N_19634);
or U19745 (N_19745,N_19637,N_19598);
xor U19746 (N_19746,N_19636,N_19602);
nand U19747 (N_19747,N_19597,N_19557);
and U19748 (N_19748,N_19643,N_19628);
and U19749 (N_19749,N_19674,N_19604);
and U19750 (N_19750,N_19672,N_19679);
nor U19751 (N_19751,N_19546,N_19635);
nor U19752 (N_19752,N_19528,N_19521);
nor U19753 (N_19753,N_19675,N_19656);
nand U19754 (N_19754,N_19564,N_19551);
nor U19755 (N_19755,N_19576,N_19553);
nand U19756 (N_19756,N_19561,N_19607);
nand U19757 (N_19757,N_19596,N_19523);
and U19758 (N_19758,N_19601,N_19543);
nor U19759 (N_19759,N_19644,N_19537);
nor U19760 (N_19760,N_19599,N_19549);
nand U19761 (N_19761,N_19638,N_19521);
and U19762 (N_19762,N_19544,N_19673);
xor U19763 (N_19763,N_19552,N_19625);
xor U19764 (N_19764,N_19571,N_19677);
and U19765 (N_19765,N_19565,N_19631);
nand U19766 (N_19766,N_19632,N_19545);
nand U19767 (N_19767,N_19527,N_19550);
and U19768 (N_19768,N_19540,N_19614);
xor U19769 (N_19769,N_19594,N_19576);
and U19770 (N_19770,N_19664,N_19642);
nand U19771 (N_19771,N_19597,N_19671);
or U19772 (N_19772,N_19641,N_19665);
or U19773 (N_19773,N_19639,N_19678);
and U19774 (N_19774,N_19588,N_19523);
nor U19775 (N_19775,N_19644,N_19549);
nor U19776 (N_19776,N_19546,N_19614);
and U19777 (N_19777,N_19624,N_19550);
nand U19778 (N_19778,N_19602,N_19553);
nor U19779 (N_19779,N_19541,N_19532);
and U19780 (N_19780,N_19648,N_19658);
or U19781 (N_19781,N_19588,N_19526);
nand U19782 (N_19782,N_19625,N_19544);
and U19783 (N_19783,N_19604,N_19590);
nor U19784 (N_19784,N_19596,N_19635);
xor U19785 (N_19785,N_19532,N_19667);
nor U19786 (N_19786,N_19635,N_19634);
or U19787 (N_19787,N_19561,N_19538);
or U19788 (N_19788,N_19546,N_19615);
and U19789 (N_19789,N_19614,N_19628);
and U19790 (N_19790,N_19642,N_19620);
and U19791 (N_19791,N_19637,N_19527);
xor U19792 (N_19792,N_19566,N_19557);
xor U19793 (N_19793,N_19662,N_19586);
nor U19794 (N_19794,N_19552,N_19555);
nand U19795 (N_19795,N_19578,N_19567);
or U19796 (N_19796,N_19675,N_19679);
nor U19797 (N_19797,N_19572,N_19557);
nand U19798 (N_19798,N_19533,N_19679);
nor U19799 (N_19799,N_19574,N_19592);
or U19800 (N_19800,N_19598,N_19657);
nor U19801 (N_19801,N_19641,N_19558);
or U19802 (N_19802,N_19546,N_19624);
and U19803 (N_19803,N_19553,N_19531);
nand U19804 (N_19804,N_19543,N_19526);
nor U19805 (N_19805,N_19566,N_19552);
nor U19806 (N_19806,N_19547,N_19611);
and U19807 (N_19807,N_19663,N_19556);
and U19808 (N_19808,N_19591,N_19590);
and U19809 (N_19809,N_19540,N_19630);
and U19810 (N_19810,N_19624,N_19571);
nand U19811 (N_19811,N_19638,N_19572);
xnor U19812 (N_19812,N_19582,N_19551);
nor U19813 (N_19813,N_19550,N_19556);
or U19814 (N_19814,N_19650,N_19626);
and U19815 (N_19815,N_19625,N_19553);
nor U19816 (N_19816,N_19578,N_19633);
nor U19817 (N_19817,N_19627,N_19665);
nor U19818 (N_19818,N_19552,N_19543);
nor U19819 (N_19819,N_19646,N_19596);
or U19820 (N_19820,N_19595,N_19532);
nor U19821 (N_19821,N_19675,N_19572);
nand U19822 (N_19822,N_19524,N_19577);
or U19823 (N_19823,N_19597,N_19576);
and U19824 (N_19824,N_19578,N_19657);
or U19825 (N_19825,N_19666,N_19590);
and U19826 (N_19826,N_19643,N_19581);
or U19827 (N_19827,N_19653,N_19575);
nand U19828 (N_19828,N_19632,N_19606);
nand U19829 (N_19829,N_19627,N_19597);
nor U19830 (N_19830,N_19551,N_19574);
xnor U19831 (N_19831,N_19544,N_19523);
and U19832 (N_19832,N_19622,N_19614);
nand U19833 (N_19833,N_19599,N_19617);
or U19834 (N_19834,N_19567,N_19640);
nand U19835 (N_19835,N_19670,N_19598);
nor U19836 (N_19836,N_19600,N_19671);
or U19837 (N_19837,N_19520,N_19592);
nand U19838 (N_19838,N_19635,N_19528);
nor U19839 (N_19839,N_19529,N_19588);
nor U19840 (N_19840,N_19719,N_19713);
xnor U19841 (N_19841,N_19818,N_19697);
or U19842 (N_19842,N_19819,N_19768);
xnor U19843 (N_19843,N_19722,N_19766);
nor U19844 (N_19844,N_19755,N_19725);
nor U19845 (N_19845,N_19686,N_19810);
nand U19846 (N_19846,N_19807,N_19737);
nand U19847 (N_19847,N_19778,N_19836);
and U19848 (N_19848,N_19682,N_19745);
nand U19849 (N_19849,N_19832,N_19714);
nand U19850 (N_19850,N_19703,N_19821);
nor U19851 (N_19851,N_19689,N_19694);
nor U19852 (N_19852,N_19771,N_19804);
nand U19853 (N_19853,N_19747,N_19723);
nand U19854 (N_19854,N_19746,N_19837);
or U19855 (N_19855,N_19717,N_19791);
nor U19856 (N_19856,N_19827,N_19800);
and U19857 (N_19857,N_19748,N_19802);
or U19858 (N_19858,N_19692,N_19733);
and U19859 (N_19859,N_19824,N_19709);
and U19860 (N_19860,N_19738,N_19783);
nand U19861 (N_19861,N_19751,N_19741);
or U19862 (N_19862,N_19701,N_19773);
or U19863 (N_19863,N_19823,N_19754);
and U19864 (N_19864,N_19808,N_19759);
and U19865 (N_19865,N_19770,N_19718);
or U19866 (N_19866,N_19715,N_19728);
and U19867 (N_19867,N_19705,N_19815);
and U19868 (N_19868,N_19698,N_19809);
or U19869 (N_19869,N_19817,N_19780);
and U19870 (N_19870,N_19684,N_19799);
nand U19871 (N_19871,N_19822,N_19758);
or U19872 (N_19872,N_19803,N_19710);
and U19873 (N_19873,N_19789,N_19695);
and U19874 (N_19874,N_19693,N_19726);
nor U19875 (N_19875,N_19839,N_19731);
nor U19876 (N_19876,N_19685,N_19816);
or U19877 (N_19877,N_19739,N_19720);
nor U19878 (N_19878,N_19721,N_19814);
or U19879 (N_19879,N_19736,N_19769);
nand U19880 (N_19880,N_19794,N_19727);
nand U19881 (N_19881,N_19683,N_19750);
nand U19882 (N_19882,N_19797,N_19711);
or U19883 (N_19883,N_19756,N_19762);
and U19884 (N_19884,N_19772,N_19833);
xor U19885 (N_19885,N_19813,N_19730);
nor U19886 (N_19886,N_19785,N_19699);
nor U19887 (N_19887,N_19767,N_19749);
or U19888 (N_19888,N_19708,N_19702);
nor U19889 (N_19889,N_19781,N_19825);
or U19890 (N_19890,N_19811,N_19700);
nor U19891 (N_19891,N_19793,N_19830);
or U19892 (N_19892,N_19834,N_19765);
and U19893 (N_19893,N_19707,N_19792);
nor U19894 (N_19894,N_19784,N_19760);
nor U19895 (N_19895,N_19801,N_19704);
nor U19896 (N_19896,N_19729,N_19820);
and U19897 (N_19897,N_19826,N_19742);
and U19898 (N_19898,N_19752,N_19777);
nand U19899 (N_19899,N_19753,N_19716);
and U19900 (N_19900,N_19712,N_19775);
nor U19901 (N_19901,N_19795,N_19696);
and U19902 (N_19902,N_19743,N_19779);
nand U19903 (N_19903,N_19740,N_19687);
and U19904 (N_19904,N_19796,N_19805);
or U19905 (N_19905,N_19776,N_19806);
nand U19906 (N_19906,N_19774,N_19732);
nor U19907 (N_19907,N_19757,N_19786);
nor U19908 (N_19908,N_19681,N_19782);
nand U19909 (N_19909,N_19764,N_19691);
or U19910 (N_19910,N_19835,N_19724);
nor U19911 (N_19911,N_19690,N_19798);
or U19912 (N_19912,N_19680,N_19787);
nand U19913 (N_19913,N_19788,N_19735);
nor U19914 (N_19914,N_19812,N_19828);
and U19915 (N_19915,N_19761,N_19838);
nand U19916 (N_19916,N_19831,N_19829);
xnor U19917 (N_19917,N_19706,N_19688);
and U19918 (N_19918,N_19734,N_19790);
or U19919 (N_19919,N_19763,N_19744);
and U19920 (N_19920,N_19734,N_19695);
nor U19921 (N_19921,N_19807,N_19812);
nor U19922 (N_19922,N_19755,N_19768);
and U19923 (N_19923,N_19718,N_19832);
and U19924 (N_19924,N_19753,N_19687);
xnor U19925 (N_19925,N_19761,N_19802);
xor U19926 (N_19926,N_19835,N_19722);
nand U19927 (N_19927,N_19839,N_19769);
nor U19928 (N_19928,N_19723,N_19828);
or U19929 (N_19929,N_19789,N_19839);
or U19930 (N_19930,N_19685,N_19741);
nand U19931 (N_19931,N_19688,N_19744);
nor U19932 (N_19932,N_19812,N_19834);
and U19933 (N_19933,N_19702,N_19738);
xnor U19934 (N_19934,N_19686,N_19785);
and U19935 (N_19935,N_19722,N_19839);
nand U19936 (N_19936,N_19761,N_19800);
and U19937 (N_19937,N_19778,N_19711);
xor U19938 (N_19938,N_19693,N_19707);
nor U19939 (N_19939,N_19709,N_19764);
nor U19940 (N_19940,N_19770,N_19699);
and U19941 (N_19941,N_19782,N_19757);
and U19942 (N_19942,N_19756,N_19835);
or U19943 (N_19943,N_19709,N_19730);
nand U19944 (N_19944,N_19800,N_19707);
nor U19945 (N_19945,N_19697,N_19734);
nor U19946 (N_19946,N_19701,N_19696);
or U19947 (N_19947,N_19729,N_19754);
nand U19948 (N_19948,N_19771,N_19809);
or U19949 (N_19949,N_19791,N_19830);
nor U19950 (N_19950,N_19707,N_19690);
or U19951 (N_19951,N_19798,N_19800);
and U19952 (N_19952,N_19721,N_19793);
and U19953 (N_19953,N_19773,N_19749);
or U19954 (N_19954,N_19716,N_19817);
xnor U19955 (N_19955,N_19774,N_19779);
and U19956 (N_19956,N_19777,N_19773);
xnor U19957 (N_19957,N_19698,N_19819);
nand U19958 (N_19958,N_19709,N_19818);
xor U19959 (N_19959,N_19772,N_19689);
nand U19960 (N_19960,N_19743,N_19708);
and U19961 (N_19961,N_19832,N_19835);
and U19962 (N_19962,N_19829,N_19773);
xor U19963 (N_19963,N_19807,N_19710);
and U19964 (N_19964,N_19714,N_19781);
nand U19965 (N_19965,N_19784,N_19782);
and U19966 (N_19966,N_19735,N_19736);
nand U19967 (N_19967,N_19770,N_19746);
or U19968 (N_19968,N_19680,N_19715);
nor U19969 (N_19969,N_19758,N_19804);
xnor U19970 (N_19970,N_19694,N_19697);
nand U19971 (N_19971,N_19759,N_19734);
and U19972 (N_19972,N_19834,N_19798);
and U19973 (N_19973,N_19758,N_19708);
xor U19974 (N_19974,N_19691,N_19697);
nor U19975 (N_19975,N_19771,N_19829);
nor U19976 (N_19976,N_19756,N_19744);
nor U19977 (N_19977,N_19705,N_19776);
nand U19978 (N_19978,N_19779,N_19768);
nand U19979 (N_19979,N_19839,N_19726);
nand U19980 (N_19980,N_19819,N_19833);
and U19981 (N_19981,N_19683,N_19783);
nor U19982 (N_19982,N_19749,N_19819);
nand U19983 (N_19983,N_19788,N_19726);
nand U19984 (N_19984,N_19740,N_19751);
nand U19985 (N_19985,N_19800,N_19710);
xnor U19986 (N_19986,N_19786,N_19775);
nand U19987 (N_19987,N_19686,N_19688);
and U19988 (N_19988,N_19739,N_19727);
or U19989 (N_19989,N_19700,N_19824);
nand U19990 (N_19990,N_19708,N_19817);
and U19991 (N_19991,N_19809,N_19696);
or U19992 (N_19992,N_19706,N_19832);
nand U19993 (N_19993,N_19799,N_19783);
nand U19994 (N_19994,N_19817,N_19803);
or U19995 (N_19995,N_19688,N_19733);
xnor U19996 (N_19996,N_19809,N_19810);
nor U19997 (N_19997,N_19825,N_19822);
or U19998 (N_19998,N_19682,N_19761);
nor U19999 (N_19999,N_19830,N_19769);
and UO_0 (O_0,N_19875,N_19973);
nand UO_1 (O_1,N_19938,N_19924);
or UO_2 (O_2,N_19899,N_19858);
or UO_3 (O_3,N_19883,N_19890);
nand UO_4 (O_4,N_19849,N_19846);
nor UO_5 (O_5,N_19997,N_19955);
and UO_6 (O_6,N_19972,N_19976);
or UO_7 (O_7,N_19949,N_19934);
nor UO_8 (O_8,N_19984,N_19980);
xnor UO_9 (O_9,N_19936,N_19982);
xnor UO_10 (O_10,N_19851,N_19937);
nor UO_11 (O_11,N_19889,N_19921);
and UO_12 (O_12,N_19969,N_19986);
or UO_13 (O_13,N_19979,N_19852);
nor UO_14 (O_14,N_19957,N_19863);
nand UO_15 (O_15,N_19884,N_19947);
xor UO_16 (O_16,N_19862,N_19998);
nand UO_17 (O_17,N_19913,N_19869);
and UO_18 (O_18,N_19988,N_19882);
and UO_19 (O_19,N_19894,N_19864);
nor UO_20 (O_20,N_19907,N_19996);
xor UO_21 (O_21,N_19942,N_19874);
nand UO_22 (O_22,N_19908,N_19951);
nor UO_23 (O_23,N_19920,N_19995);
nor UO_24 (O_24,N_19914,N_19892);
and UO_25 (O_25,N_19946,N_19952);
xnor UO_26 (O_26,N_19860,N_19967);
nand UO_27 (O_27,N_19925,N_19870);
xor UO_28 (O_28,N_19983,N_19871);
or UO_29 (O_29,N_19854,N_19930);
or UO_30 (O_30,N_19954,N_19886);
or UO_31 (O_31,N_19931,N_19968);
and UO_32 (O_32,N_19933,N_19939);
nand UO_33 (O_33,N_19943,N_19859);
and UO_34 (O_34,N_19903,N_19866);
nand UO_35 (O_35,N_19940,N_19945);
or UO_36 (O_36,N_19845,N_19842);
or UO_37 (O_37,N_19865,N_19941);
xor UO_38 (O_38,N_19965,N_19932);
nand UO_39 (O_39,N_19958,N_19897);
or UO_40 (O_40,N_19966,N_19977);
xnor UO_41 (O_41,N_19867,N_19905);
nand UO_42 (O_42,N_19841,N_19935);
and UO_43 (O_43,N_19916,N_19844);
or UO_44 (O_44,N_19928,N_19961);
and UO_45 (O_45,N_19923,N_19850);
or UO_46 (O_46,N_19953,N_19881);
nand UO_47 (O_47,N_19873,N_19893);
and UO_48 (O_48,N_19991,N_19840);
nand UO_49 (O_49,N_19912,N_19853);
nand UO_50 (O_50,N_19880,N_19963);
or UO_51 (O_51,N_19891,N_19906);
nand UO_52 (O_52,N_19917,N_19974);
nor UO_53 (O_53,N_19856,N_19981);
and UO_54 (O_54,N_19987,N_19879);
or UO_55 (O_55,N_19888,N_19985);
nor UO_56 (O_56,N_19896,N_19944);
nand UO_57 (O_57,N_19978,N_19904);
and UO_58 (O_58,N_19915,N_19999);
nand UO_59 (O_59,N_19989,N_19971);
nand UO_60 (O_60,N_19900,N_19901);
nand UO_61 (O_61,N_19948,N_19962);
and UO_62 (O_62,N_19922,N_19909);
and UO_63 (O_63,N_19919,N_19993);
xor UO_64 (O_64,N_19887,N_19876);
nor UO_65 (O_65,N_19964,N_19843);
nor UO_66 (O_66,N_19960,N_19950);
xor UO_67 (O_67,N_19877,N_19902);
xnor UO_68 (O_68,N_19878,N_19956);
and UO_69 (O_69,N_19959,N_19861);
nor UO_70 (O_70,N_19872,N_19918);
nand UO_71 (O_71,N_19857,N_19970);
xnor UO_72 (O_72,N_19855,N_19994);
and UO_73 (O_73,N_19898,N_19992);
or UO_74 (O_74,N_19990,N_19926);
and UO_75 (O_75,N_19847,N_19910);
nand UO_76 (O_76,N_19911,N_19929);
and UO_77 (O_77,N_19885,N_19895);
nor UO_78 (O_78,N_19927,N_19868);
nor UO_79 (O_79,N_19975,N_19848);
nand UO_80 (O_80,N_19988,N_19978);
nand UO_81 (O_81,N_19957,N_19916);
or UO_82 (O_82,N_19990,N_19927);
and UO_83 (O_83,N_19999,N_19920);
and UO_84 (O_84,N_19870,N_19938);
and UO_85 (O_85,N_19877,N_19911);
and UO_86 (O_86,N_19846,N_19845);
nand UO_87 (O_87,N_19950,N_19976);
nand UO_88 (O_88,N_19895,N_19884);
and UO_89 (O_89,N_19847,N_19994);
nand UO_90 (O_90,N_19868,N_19944);
nand UO_91 (O_91,N_19855,N_19991);
nand UO_92 (O_92,N_19961,N_19924);
nand UO_93 (O_93,N_19853,N_19951);
or UO_94 (O_94,N_19893,N_19921);
or UO_95 (O_95,N_19848,N_19965);
and UO_96 (O_96,N_19923,N_19845);
nor UO_97 (O_97,N_19949,N_19968);
xnor UO_98 (O_98,N_19876,N_19960);
nor UO_99 (O_99,N_19903,N_19841);
nor UO_100 (O_100,N_19960,N_19988);
nor UO_101 (O_101,N_19985,N_19913);
nand UO_102 (O_102,N_19974,N_19868);
or UO_103 (O_103,N_19926,N_19957);
and UO_104 (O_104,N_19953,N_19876);
nor UO_105 (O_105,N_19896,N_19852);
or UO_106 (O_106,N_19971,N_19857);
or UO_107 (O_107,N_19998,N_19889);
nand UO_108 (O_108,N_19921,N_19917);
xnor UO_109 (O_109,N_19896,N_19921);
and UO_110 (O_110,N_19943,N_19967);
or UO_111 (O_111,N_19860,N_19965);
or UO_112 (O_112,N_19982,N_19986);
and UO_113 (O_113,N_19891,N_19995);
nand UO_114 (O_114,N_19915,N_19957);
or UO_115 (O_115,N_19946,N_19875);
or UO_116 (O_116,N_19962,N_19923);
nand UO_117 (O_117,N_19901,N_19854);
and UO_118 (O_118,N_19999,N_19986);
and UO_119 (O_119,N_19868,N_19980);
nor UO_120 (O_120,N_19899,N_19861);
and UO_121 (O_121,N_19878,N_19898);
nor UO_122 (O_122,N_19982,N_19956);
and UO_123 (O_123,N_19895,N_19933);
or UO_124 (O_124,N_19997,N_19974);
nand UO_125 (O_125,N_19992,N_19888);
nand UO_126 (O_126,N_19999,N_19869);
nand UO_127 (O_127,N_19879,N_19922);
nor UO_128 (O_128,N_19848,N_19858);
or UO_129 (O_129,N_19848,N_19972);
or UO_130 (O_130,N_19860,N_19976);
nor UO_131 (O_131,N_19856,N_19882);
nand UO_132 (O_132,N_19952,N_19913);
or UO_133 (O_133,N_19842,N_19910);
xnor UO_134 (O_134,N_19880,N_19904);
or UO_135 (O_135,N_19875,N_19950);
nor UO_136 (O_136,N_19986,N_19888);
or UO_137 (O_137,N_19902,N_19985);
nor UO_138 (O_138,N_19856,N_19883);
nand UO_139 (O_139,N_19870,N_19872);
nor UO_140 (O_140,N_19917,N_19875);
and UO_141 (O_141,N_19997,N_19961);
xor UO_142 (O_142,N_19917,N_19931);
and UO_143 (O_143,N_19922,N_19868);
xor UO_144 (O_144,N_19941,N_19972);
and UO_145 (O_145,N_19905,N_19879);
or UO_146 (O_146,N_19874,N_19995);
nor UO_147 (O_147,N_19944,N_19851);
or UO_148 (O_148,N_19866,N_19894);
or UO_149 (O_149,N_19975,N_19905);
nand UO_150 (O_150,N_19919,N_19892);
and UO_151 (O_151,N_19841,N_19942);
nand UO_152 (O_152,N_19883,N_19924);
or UO_153 (O_153,N_19933,N_19984);
xnor UO_154 (O_154,N_19906,N_19904);
and UO_155 (O_155,N_19919,N_19903);
xnor UO_156 (O_156,N_19935,N_19946);
nand UO_157 (O_157,N_19881,N_19972);
xor UO_158 (O_158,N_19953,N_19973);
and UO_159 (O_159,N_19969,N_19971);
or UO_160 (O_160,N_19890,N_19850);
nand UO_161 (O_161,N_19892,N_19884);
and UO_162 (O_162,N_19857,N_19924);
or UO_163 (O_163,N_19938,N_19883);
nand UO_164 (O_164,N_19979,N_19905);
or UO_165 (O_165,N_19959,N_19885);
nor UO_166 (O_166,N_19902,N_19997);
or UO_167 (O_167,N_19980,N_19997);
nand UO_168 (O_168,N_19937,N_19841);
and UO_169 (O_169,N_19844,N_19878);
and UO_170 (O_170,N_19882,N_19930);
nand UO_171 (O_171,N_19853,N_19946);
or UO_172 (O_172,N_19841,N_19967);
and UO_173 (O_173,N_19857,N_19902);
and UO_174 (O_174,N_19846,N_19934);
and UO_175 (O_175,N_19968,N_19973);
or UO_176 (O_176,N_19961,N_19921);
and UO_177 (O_177,N_19948,N_19913);
or UO_178 (O_178,N_19905,N_19928);
nand UO_179 (O_179,N_19900,N_19920);
nand UO_180 (O_180,N_19995,N_19870);
nor UO_181 (O_181,N_19997,N_19906);
nand UO_182 (O_182,N_19915,N_19929);
or UO_183 (O_183,N_19977,N_19990);
and UO_184 (O_184,N_19894,N_19900);
or UO_185 (O_185,N_19958,N_19940);
and UO_186 (O_186,N_19966,N_19943);
or UO_187 (O_187,N_19920,N_19982);
nor UO_188 (O_188,N_19961,N_19911);
nor UO_189 (O_189,N_19941,N_19914);
and UO_190 (O_190,N_19900,N_19905);
and UO_191 (O_191,N_19850,N_19864);
nand UO_192 (O_192,N_19881,N_19960);
nor UO_193 (O_193,N_19889,N_19893);
xor UO_194 (O_194,N_19979,N_19929);
and UO_195 (O_195,N_19980,N_19898);
or UO_196 (O_196,N_19879,N_19861);
nor UO_197 (O_197,N_19979,N_19923);
or UO_198 (O_198,N_19903,N_19989);
nor UO_199 (O_199,N_19915,N_19967);
nand UO_200 (O_200,N_19856,N_19932);
nand UO_201 (O_201,N_19955,N_19980);
nand UO_202 (O_202,N_19870,N_19941);
and UO_203 (O_203,N_19997,N_19979);
or UO_204 (O_204,N_19933,N_19971);
nand UO_205 (O_205,N_19872,N_19908);
or UO_206 (O_206,N_19865,N_19842);
and UO_207 (O_207,N_19861,N_19898);
nor UO_208 (O_208,N_19968,N_19919);
nand UO_209 (O_209,N_19903,N_19858);
and UO_210 (O_210,N_19871,N_19941);
nand UO_211 (O_211,N_19923,N_19996);
and UO_212 (O_212,N_19992,N_19878);
nand UO_213 (O_213,N_19867,N_19882);
xnor UO_214 (O_214,N_19883,N_19903);
nand UO_215 (O_215,N_19985,N_19851);
or UO_216 (O_216,N_19891,N_19868);
nor UO_217 (O_217,N_19875,N_19886);
xnor UO_218 (O_218,N_19992,N_19893);
or UO_219 (O_219,N_19984,N_19865);
nand UO_220 (O_220,N_19868,N_19897);
and UO_221 (O_221,N_19992,N_19871);
nand UO_222 (O_222,N_19842,N_19922);
and UO_223 (O_223,N_19882,N_19971);
nor UO_224 (O_224,N_19915,N_19926);
nor UO_225 (O_225,N_19923,N_19960);
nand UO_226 (O_226,N_19938,N_19906);
nor UO_227 (O_227,N_19940,N_19852);
and UO_228 (O_228,N_19852,N_19855);
and UO_229 (O_229,N_19918,N_19984);
nand UO_230 (O_230,N_19934,N_19842);
or UO_231 (O_231,N_19949,N_19874);
or UO_232 (O_232,N_19981,N_19985);
xor UO_233 (O_233,N_19873,N_19840);
nand UO_234 (O_234,N_19987,N_19993);
nor UO_235 (O_235,N_19870,N_19959);
nor UO_236 (O_236,N_19840,N_19945);
or UO_237 (O_237,N_19870,N_19935);
nand UO_238 (O_238,N_19937,N_19846);
nand UO_239 (O_239,N_19863,N_19995);
or UO_240 (O_240,N_19994,N_19843);
or UO_241 (O_241,N_19942,N_19998);
or UO_242 (O_242,N_19967,N_19867);
or UO_243 (O_243,N_19876,N_19928);
nand UO_244 (O_244,N_19954,N_19871);
nor UO_245 (O_245,N_19979,N_19938);
and UO_246 (O_246,N_19885,N_19991);
and UO_247 (O_247,N_19949,N_19985);
and UO_248 (O_248,N_19985,N_19854);
or UO_249 (O_249,N_19934,N_19985);
nand UO_250 (O_250,N_19865,N_19858);
nand UO_251 (O_251,N_19869,N_19883);
nand UO_252 (O_252,N_19898,N_19979);
xnor UO_253 (O_253,N_19859,N_19993);
nor UO_254 (O_254,N_19885,N_19915);
nor UO_255 (O_255,N_19840,N_19969);
or UO_256 (O_256,N_19844,N_19953);
nand UO_257 (O_257,N_19902,N_19914);
and UO_258 (O_258,N_19950,N_19878);
nor UO_259 (O_259,N_19875,N_19842);
and UO_260 (O_260,N_19912,N_19850);
nor UO_261 (O_261,N_19915,N_19943);
and UO_262 (O_262,N_19965,N_19947);
nand UO_263 (O_263,N_19852,N_19867);
nand UO_264 (O_264,N_19912,N_19918);
xor UO_265 (O_265,N_19942,N_19877);
and UO_266 (O_266,N_19968,N_19863);
and UO_267 (O_267,N_19881,N_19845);
and UO_268 (O_268,N_19966,N_19992);
nor UO_269 (O_269,N_19949,N_19888);
nand UO_270 (O_270,N_19841,N_19956);
nor UO_271 (O_271,N_19958,N_19926);
or UO_272 (O_272,N_19912,N_19981);
nor UO_273 (O_273,N_19951,N_19889);
and UO_274 (O_274,N_19869,N_19935);
xnor UO_275 (O_275,N_19856,N_19937);
and UO_276 (O_276,N_19987,N_19878);
and UO_277 (O_277,N_19932,N_19903);
xnor UO_278 (O_278,N_19914,N_19897);
or UO_279 (O_279,N_19959,N_19883);
or UO_280 (O_280,N_19917,N_19871);
and UO_281 (O_281,N_19885,N_19869);
or UO_282 (O_282,N_19950,N_19927);
and UO_283 (O_283,N_19949,N_19964);
and UO_284 (O_284,N_19855,N_19872);
or UO_285 (O_285,N_19896,N_19901);
nor UO_286 (O_286,N_19978,N_19844);
nand UO_287 (O_287,N_19903,N_19927);
nand UO_288 (O_288,N_19845,N_19988);
nor UO_289 (O_289,N_19981,N_19879);
nand UO_290 (O_290,N_19995,N_19982);
or UO_291 (O_291,N_19891,N_19978);
and UO_292 (O_292,N_19969,N_19904);
nand UO_293 (O_293,N_19954,N_19946);
nand UO_294 (O_294,N_19971,N_19967);
nand UO_295 (O_295,N_19841,N_19854);
and UO_296 (O_296,N_19969,N_19899);
nor UO_297 (O_297,N_19968,N_19846);
nor UO_298 (O_298,N_19961,N_19971);
and UO_299 (O_299,N_19866,N_19938);
or UO_300 (O_300,N_19919,N_19893);
and UO_301 (O_301,N_19895,N_19868);
nand UO_302 (O_302,N_19986,N_19887);
and UO_303 (O_303,N_19961,N_19947);
or UO_304 (O_304,N_19959,N_19913);
and UO_305 (O_305,N_19943,N_19843);
and UO_306 (O_306,N_19851,N_19935);
nor UO_307 (O_307,N_19882,N_19948);
nand UO_308 (O_308,N_19893,N_19857);
and UO_309 (O_309,N_19883,N_19947);
and UO_310 (O_310,N_19861,N_19919);
and UO_311 (O_311,N_19998,N_19983);
nand UO_312 (O_312,N_19923,N_19974);
and UO_313 (O_313,N_19911,N_19931);
and UO_314 (O_314,N_19965,N_19978);
and UO_315 (O_315,N_19943,N_19892);
and UO_316 (O_316,N_19898,N_19942);
nor UO_317 (O_317,N_19954,N_19996);
xor UO_318 (O_318,N_19934,N_19898);
or UO_319 (O_319,N_19950,N_19867);
and UO_320 (O_320,N_19882,N_19853);
or UO_321 (O_321,N_19982,N_19860);
nor UO_322 (O_322,N_19902,N_19943);
nor UO_323 (O_323,N_19946,N_19932);
and UO_324 (O_324,N_19871,N_19860);
and UO_325 (O_325,N_19915,N_19856);
nor UO_326 (O_326,N_19922,N_19951);
nand UO_327 (O_327,N_19959,N_19850);
or UO_328 (O_328,N_19860,N_19866);
or UO_329 (O_329,N_19930,N_19851);
or UO_330 (O_330,N_19876,N_19922);
or UO_331 (O_331,N_19951,N_19937);
or UO_332 (O_332,N_19889,N_19860);
xor UO_333 (O_333,N_19972,N_19979);
xor UO_334 (O_334,N_19873,N_19934);
or UO_335 (O_335,N_19865,N_19918);
and UO_336 (O_336,N_19842,N_19923);
or UO_337 (O_337,N_19862,N_19937);
xor UO_338 (O_338,N_19997,N_19887);
xnor UO_339 (O_339,N_19869,N_19976);
or UO_340 (O_340,N_19887,N_19942);
nand UO_341 (O_341,N_19896,N_19955);
nor UO_342 (O_342,N_19880,N_19921);
or UO_343 (O_343,N_19868,N_19852);
nor UO_344 (O_344,N_19957,N_19932);
xor UO_345 (O_345,N_19855,N_19953);
nand UO_346 (O_346,N_19915,N_19913);
or UO_347 (O_347,N_19912,N_19871);
nor UO_348 (O_348,N_19963,N_19941);
and UO_349 (O_349,N_19981,N_19847);
nand UO_350 (O_350,N_19993,N_19857);
nand UO_351 (O_351,N_19950,N_19984);
or UO_352 (O_352,N_19975,N_19858);
nor UO_353 (O_353,N_19847,N_19870);
or UO_354 (O_354,N_19953,N_19852);
or UO_355 (O_355,N_19865,N_19903);
nand UO_356 (O_356,N_19955,N_19889);
xnor UO_357 (O_357,N_19925,N_19921);
or UO_358 (O_358,N_19977,N_19905);
nand UO_359 (O_359,N_19960,N_19845);
and UO_360 (O_360,N_19849,N_19910);
and UO_361 (O_361,N_19975,N_19917);
and UO_362 (O_362,N_19979,N_19947);
nand UO_363 (O_363,N_19930,N_19965);
nand UO_364 (O_364,N_19974,N_19840);
nand UO_365 (O_365,N_19932,N_19928);
and UO_366 (O_366,N_19932,N_19855);
xor UO_367 (O_367,N_19879,N_19852);
nand UO_368 (O_368,N_19955,N_19984);
nand UO_369 (O_369,N_19992,N_19874);
xor UO_370 (O_370,N_19938,N_19951);
or UO_371 (O_371,N_19948,N_19928);
nor UO_372 (O_372,N_19880,N_19853);
or UO_373 (O_373,N_19989,N_19932);
xor UO_374 (O_374,N_19970,N_19858);
or UO_375 (O_375,N_19975,N_19897);
and UO_376 (O_376,N_19948,N_19945);
xor UO_377 (O_377,N_19886,N_19919);
and UO_378 (O_378,N_19874,N_19887);
nor UO_379 (O_379,N_19864,N_19873);
xor UO_380 (O_380,N_19844,N_19994);
nor UO_381 (O_381,N_19916,N_19864);
nand UO_382 (O_382,N_19918,N_19907);
nor UO_383 (O_383,N_19902,N_19911);
nor UO_384 (O_384,N_19851,N_19933);
and UO_385 (O_385,N_19944,N_19937);
or UO_386 (O_386,N_19874,N_19937);
nand UO_387 (O_387,N_19849,N_19928);
nand UO_388 (O_388,N_19993,N_19949);
or UO_389 (O_389,N_19843,N_19866);
and UO_390 (O_390,N_19978,N_19887);
and UO_391 (O_391,N_19900,N_19875);
and UO_392 (O_392,N_19943,N_19987);
and UO_393 (O_393,N_19944,N_19997);
nor UO_394 (O_394,N_19990,N_19993);
and UO_395 (O_395,N_19911,N_19842);
nor UO_396 (O_396,N_19972,N_19907);
and UO_397 (O_397,N_19933,N_19989);
and UO_398 (O_398,N_19961,N_19933);
nor UO_399 (O_399,N_19924,N_19865);
nor UO_400 (O_400,N_19895,N_19844);
nor UO_401 (O_401,N_19934,N_19948);
xnor UO_402 (O_402,N_19922,N_19968);
nor UO_403 (O_403,N_19972,N_19861);
and UO_404 (O_404,N_19909,N_19964);
or UO_405 (O_405,N_19866,N_19884);
and UO_406 (O_406,N_19912,N_19961);
or UO_407 (O_407,N_19974,N_19986);
nand UO_408 (O_408,N_19886,N_19988);
or UO_409 (O_409,N_19847,N_19921);
xor UO_410 (O_410,N_19874,N_19953);
nand UO_411 (O_411,N_19875,N_19876);
nand UO_412 (O_412,N_19965,N_19903);
and UO_413 (O_413,N_19903,N_19869);
and UO_414 (O_414,N_19933,N_19910);
nor UO_415 (O_415,N_19843,N_19963);
nand UO_416 (O_416,N_19939,N_19934);
xor UO_417 (O_417,N_19876,N_19902);
nor UO_418 (O_418,N_19983,N_19977);
and UO_419 (O_419,N_19924,N_19977);
and UO_420 (O_420,N_19933,N_19903);
xor UO_421 (O_421,N_19961,N_19846);
or UO_422 (O_422,N_19946,N_19927);
nand UO_423 (O_423,N_19844,N_19932);
or UO_424 (O_424,N_19965,N_19919);
and UO_425 (O_425,N_19874,N_19914);
or UO_426 (O_426,N_19941,N_19859);
and UO_427 (O_427,N_19969,N_19879);
and UO_428 (O_428,N_19921,N_19987);
or UO_429 (O_429,N_19948,N_19981);
nor UO_430 (O_430,N_19944,N_19857);
xnor UO_431 (O_431,N_19862,N_19957);
nand UO_432 (O_432,N_19986,N_19907);
and UO_433 (O_433,N_19997,N_19985);
and UO_434 (O_434,N_19912,N_19891);
nand UO_435 (O_435,N_19910,N_19868);
nand UO_436 (O_436,N_19992,N_19899);
xnor UO_437 (O_437,N_19947,N_19970);
nand UO_438 (O_438,N_19929,N_19933);
nand UO_439 (O_439,N_19911,N_19905);
nor UO_440 (O_440,N_19861,N_19939);
nor UO_441 (O_441,N_19957,N_19917);
nand UO_442 (O_442,N_19911,N_19859);
nand UO_443 (O_443,N_19883,N_19948);
and UO_444 (O_444,N_19885,N_19974);
and UO_445 (O_445,N_19924,N_19903);
nor UO_446 (O_446,N_19953,N_19931);
nand UO_447 (O_447,N_19955,N_19952);
nand UO_448 (O_448,N_19880,N_19861);
and UO_449 (O_449,N_19968,N_19994);
and UO_450 (O_450,N_19970,N_19880);
and UO_451 (O_451,N_19887,N_19944);
nand UO_452 (O_452,N_19846,N_19932);
xor UO_453 (O_453,N_19945,N_19855);
or UO_454 (O_454,N_19882,N_19907);
nand UO_455 (O_455,N_19974,N_19979);
or UO_456 (O_456,N_19905,N_19845);
or UO_457 (O_457,N_19946,N_19926);
xnor UO_458 (O_458,N_19990,N_19948);
and UO_459 (O_459,N_19841,N_19866);
and UO_460 (O_460,N_19921,N_19953);
nand UO_461 (O_461,N_19881,N_19952);
and UO_462 (O_462,N_19994,N_19892);
and UO_463 (O_463,N_19859,N_19862);
nor UO_464 (O_464,N_19992,N_19990);
and UO_465 (O_465,N_19940,N_19975);
and UO_466 (O_466,N_19950,N_19926);
nor UO_467 (O_467,N_19989,N_19846);
and UO_468 (O_468,N_19944,N_19957);
nor UO_469 (O_469,N_19967,N_19969);
or UO_470 (O_470,N_19901,N_19993);
or UO_471 (O_471,N_19909,N_19842);
and UO_472 (O_472,N_19984,N_19982);
nor UO_473 (O_473,N_19996,N_19851);
or UO_474 (O_474,N_19971,N_19850);
nor UO_475 (O_475,N_19858,N_19934);
nand UO_476 (O_476,N_19898,N_19906);
nand UO_477 (O_477,N_19987,N_19986);
nor UO_478 (O_478,N_19964,N_19930);
and UO_479 (O_479,N_19882,N_19934);
nor UO_480 (O_480,N_19961,N_19896);
or UO_481 (O_481,N_19997,N_19850);
nand UO_482 (O_482,N_19944,N_19898);
nor UO_483 (O_483,N_19854,N_19874);
or UO_484 (O_484,N_19953,N_19861);
nor UO_485 (O_485,N_19872,N_19951);
or UO_486 (O_486,N_19885,N_19985);
nor UO_487 (O_487,N_19945,N_19920);
nor UO_488 (O_488,N_19913,N_19876);
and UO_489 (O_489,N_19956,N_19941);
xor UO_490 (O_490,N_19850,N_19949);
and UO_491 (O_491,N_19974,N_19922);
or UO_492 (O_492,N_19958,N_19968);
nor UO_493 (O_493,N_19915,N_19874);
and UO_494 (O_494,N_19916,N_19942);
nor UO_495 (O_495,N_19992,N_19845);
nor UO_496 (O_496,N_19943,N_19993);
nand UO_497 (O_497,N_19897,N_19851);
nor UO_498 (O_498,N_19966,N_19869);
nand UO_499 (O_499,N_19893,N_19848);
nand UO_500 (O_500,N_19897,N_19915);
nor UO_501 (O_501,N_19960,N_19883);
xor UO_502 (O_502,N_19902,N_19874);
nor UO_503 (O_503,N_19965,N_19893);
nand UO_504 (O_504,N_19932,N_19981);
or UO_505 (O_505,N_19952,N_19894);
or UO_506 (O_506,N_19942,N_19989);
nand UO_507 (O_507,N_19900,N_19965);
or UO_508 (O_508,N_19911,N_19964);
and UO_509 (O_509,N_19921,N_19879);
nand UO_510 (O_510,N_19898,N_19904);
xor UO_511 (O_511,N_19969,N_19954);
and UO_512 (O_512,N_19994,N_19971);
or UO_513 (O_513,N_19902,N_19978);
or UO_514 (O_514,N_19932,N_19933);
nand UO_515 (O_515,N_19875,N_19882);
xnor UO_516 (O_516,N_19972,N_19962);
or UO_517 (O_517,N_19998,N_19858);
or UO_518 (O_518,N_19897,N_19856);
xor UO_519 (O_519,N_19885,N_19973);
nor UO_520 (O_520,N_19989,N_19921);
or UO_521 (O_521,N_19985,N_19907);
nand UO_522 (O_522,N_19875,N_19892);
and UO_523 (O_523,N_19924,N_19994);
nor UO_524 (O_524,N_19921,N_19951);
nand UO_525 (O_525,N_19841,N_19930);
or UO_526 (O_526,N_19984,N_19862);
or UO_527 (O_527,N_19997,N_19958);
nand UO_528 (O_528,N_19948,N_19886);
nand UO_529 (O_529,N_19956,N_19920);
or UO_530 (O_530,N_19919,N_19947);
xor UO_531 (O_531,N_19929,N_19898);
or UO_532 (O_532,N_19944,N_19999);
xor UO_533 (O_533,N_19872,N_19938);
and UO_534 (O_534,N_19950,N_19883);
nand UO_535 (O_535,N_19995,N_19941);
nor UO_536 (O_536,N_19900,N_19968);
nand UO_537 (O_537,N_19928,N_19992);
nand UO_538 (O_538,N_19994,N_19905);
nand UO_539 (O_539,N_19944,N_19979);
or UO_540 (O_540,N_19940,N_19887);
nand UO_541 (O_541,N_19845,N_19976);
or UO_542 (O_542,N_19978,N_19889);
and UO_543 (O_543,N_19846,N_19995);
and UO_544 (O_544,N_19986,N_19948);
or UO_545 (O_545,N_19994,N_19959);
nor UO_546 (O_546,N_19902,N_19885);
xnor UO_547 (O_547,N_19869,N_19975);
xor UO_548 (O_548,N_19933,N_19857);
and UO_549 (O_549,N_19843,N_19939);
xnor UO_550 (O_550,N_19928,N_19902);
and UO_551 (O_551,N_19986,N_19938);
or UO_552 (O_552,N_19844,N_19945);
nand UO_553 (O_553,N_19876,N_19905);
nor UO_554 (O_554,N_19892,N_19926);
and UO_555 (O_555,N_19898,N_19911);
or UO_556 (O_556,N_19847,N_19995);
or UO_557 (O_557,N_19860,N_19918);
xnor UO_558 (O_558,N_19870,N_19850);
xor UO_559 (O_559,N_19923,N_19991);
or UO_560 (O_560,N_19872,N_19939);
xnor UO_561 (O_561,N_19972,N_19902);
nand UO_562 (O_562,N_19948,N_19879);
nor UO_563 (O_563,N_19978,N_19969);
and UO_564 (O_564,N_19926,N_19924);
and UO_565 (O_565,N_19855,N_19974);
nor UO_566 (O_566,N_19954,N_19923);
and UO_567 (O_567,N_19959,N_19886);
or UO_568 (O_568,N_19868,N_19962);
and UO_569 (O_569,N_19910,N_19953);
xor UO_570 (O_570,N_19912,N_19873);
nand UO_571 (O_571,N_19950,N_19922);
and UO_572 (O_572,N_19911,N_19978);
nand UO_573 (O_573,N_19871,N_19914);
and UO_574 (O_574,N_19934,N_19952);
nor UO_575 (O_575,N_19898,N_19903);
or UO_576 (O_576,N_19969,N_19973);
or UO_577 (O_577,N_19888,N_19874);
or UO_578 (O_578,N_19854,N_19866);
and UO_579 (O_579,N_19984,N_19874);
nor UO_580 (O_580,N_19893,N_19903);
nand UO_581 (O_581,N_19888,N_19887);
or UO_582 (O_582,N_19947,N_19957);
xor UO_583 (O_583,N_19924,N_19922);
xnor UO_584 (O_584,N_19856,N_19886);
or UO_585 (O_585,N_19894,N_19907);
or UO_586 (O_586,N_19932,N_19995);
nand UO_587 (O_587,N_19954,N_19913);
or UO_588 (O_588,N_19927,N_19922);
or UO_589 (O_589,N_19904,N_19872);
nand UO_590 (O_590,N_19913,N_19955);
nor UO_591 (O_591,N_19850,N_19914);
nor UO_592 (O_592,N_19967,N_19865);
and UO_593 (O_593,N_19886,N_19928);
and UO_594 (O_594,N_19924,N_19847);
nor UO_595 (O_595,N_19871,N_19865);
nand UO_596 (O_596,N_19843,N_19999);
and UO_597 (O_597,N_19967,N_19871);
or UO_598 (O_598,N_19965,N_19875);
or UO_599 (O_599,N_19946,N_19925);
nand UO_600 (O_600,N_19888,N_19987);
nand UO_601 (O_601,N_19849,N_19845);
or UO_602 (O_602,N_19960,N_19905);
xor UO_603 (O_603,N_19984,N_19992);
nor UO_604 (O_604,N_19939,N_19969);
and UO_605 (O_605,N_19866,N_19935);
nand UO_606 (O_606,N_19940,N_19956);
nand UO_607 (O_607,N_19887,N_19939);
nor UO_608 (O_608,N_19868,N_19956);
nand UO_609 (O_609,N_19971,N_19867);
nand UO_610 (O_610,N_19888,N_19980);
and UO_611 (O_611,N_19944,N_19978);
or UO_612 (O_612,N_19930,N_19928);
xnor UO_613 (O_613,N_19909,N_19866);
nor UO_614 (O_614,N_19984,N_19997);
and UO_615 (O_615,N_19994,N_19987);
nand UO_616 (O_616,N_19875,N_19903);
nand UO_617 (O_617,N_19919,N_19933);
nor UO_618 (O_618,N_19855,N_19949);
nor UO_619 (O_619,N_19886,N_19882);
or UO_620 (O_620,N_19883,N_19989);
and UO_621 (O_621,N_19981,N_19944);
or UO_622 (O_622,N_19903,N_19906);
or UO_623 (O_623,N_19987,N_19868);
xnor UO_624 (O_624,N_19973,N_19860);
nor UO_625 (O_625,N_19918,N_19852);
nand UO_626 (O_626,N_19922,N_19849);
and UO_627 (O_627,N_19900,N_19877);
xnor UO_628 (O_628,N_19983,N_19922);
nor UO_629 (O_629,N_19903,N_19849);
nor UO_630 (O_630,N_19941,N_19953);
and UO_631 (O_631,N_19890,N_19961);
nand UO_632 (O_632,N_19882,N_19924);
nor UO_633 (O_633,N_19890,N_19892);
and UO_634 (O_634,N_19887,N_19884);
xor UO_635 (O_635,N_19907,N_19861);
nor UO_636 (O_636,N_19904,N_19902);
nand UO_637 (O_637,N_19966,N_19944);
or UO_638 (O_638,N_19847,N_19996);
nand UO_639 (O_639,N_19854,N_19921);
xor UO_640 (O_640,N_19983,N_19931);
or UO_641 (O_641,N_19847,N_19933);
nor UO_642 (O_642,N_19860,N_19853);
nor UO_643 (O_643,N_19966,N_19875);
or UO_644 (O_644,N_19928,N_19874);
or UO_645 (O_645,N_19894,N_19881);
xor UO_646 (O_646,N_19890,N_19983);
and UO_647 (O_647,N_19917,N_19886);
nor UO_648 (O_648,N_19993,N_19884);
and UO_649 (O_649,N_19954,N_19975);
nor UO_650 (O_650,N_19898,N_19959);
and UO_651 (O_651,N_19966,N_19969);
and UO_652 (O_652,N_19957,N_19963);
nor UO_653 (O_653,N_19927,N_19892);
or UO_654 (O_654,N_19874,N_19911);
and UO_655 (O_655,N_19944,N_19992);
or UO_656 (O_656,N_19860,N_19939);
nor UO_657 (O_657,N_19908,N_19849);
nor UO_658 (O_658,N_19884,N_19873);
and UO_659 (O_659,N_19868,N_19887);
or UO_660 (O_660,N_19846,N_19878);
and UO_661 (O_661,N_19910,N_19867);
nor UO_662 (O_662,N_19956,N_19976);
nor UO_663 (O_663,N_19915,N_19986);
nand UO_664 (O_664,N_19857,N_19905);
or UO_665 (O_665,N_19894,N_19897);
nand UO_666 (O_666,N_19965,N_19906);
or UO_667 (O_667,N_19865,N_19887);
xor UO_668 (O_668,N_19927,N_19911);
and UO_669 (O_669,N_19964,N_19853);
nor UO_670 (O_670,N_19870,N_19884);
nor UO_671 (O_671,N_19937,N_19935);
and UO_672 (O_672,N_19867,N_19938);
xnor UO_673 (O_673,N_19923,N_19973);
nor UO_674 (O_674,N_19961,N_19968);
nand UO_675 (O_675,N_19934,N_19983);
nor UO_676 (O_676,N_19997,N_19967);
or UO_677 (O_677,N_19847,N_19916);
and UO_678 (O_678,N_19869,N_19852);
and UO_679 (O_679,N_19878,N_19994);
nand UO_680 (O_680,N_19965,N_19872);
nor UO_681 (O_681,N_19977,N_19866);
and UO_682 (O_682,N_19847,N_19947);
and UO_683 (O_683,N_19899,N_19882);
and UO_684 (O_684,N_19866,N_19849);
and UO_685 (O_685,N_19852,N_19989);
and UO_686 (O_686,N_19954,N_19845);
and UO_687 (O_687,N_19850,N_19895);
or UO_688 (O_688,N_19843,N_19991);
nand UO_689 (O_689,N_19982,N_19877);
and UO_690 (O_690,N_19844,N_19960);
nand UO_691 (O_691,N_19942,N_19964);
nor UO_692 (O_692,N_19971,N_19991);
or UO_693 (O_693,N_19979,N_19909);
nand UO_694 (O_694,N_19892,N_19970);
nor UO_695 (O_695,N_19895,N_19954);
xnor UO_696 (O_696,N_19926,N_19903);
nor UO_697 (O_697,N_19929,N_19951);
nand UO_698 (O_698,N_19909,N_19851);
or UO_699 (O_699,N_19929,N_19847);
and UO_700 (O_700,N_19945,N_19862);
nand UO_701 (O_701,N_19957,N_19974);
and UO_702 (O_702,N_19869,N_19912);
xor UO_703 (O_703,N_19895,N_19896);
nand UO_704 (O_704,N_19981,N_19967);
nand UO_705 (O_705,N_19966,N_19936);
nand UO_706 (O_706,N_19985,N_19930);
nand UO_707 (O_707,N_19887,N_19895);
and UO_708 (O_708,N_19990,N_19897);
nor UO_709 (O_709,N_19892,N_19977);
and UO_710 (O_710,N_19960,N_19871);
and UO_711 (O_711,N_19932,N_19919);
and UO_712 (O_712,N_19884,N_19976);
or UO_713 (O_713,N_19880,N_19933);
nor UO_714 (O_714,N_19908,N_19899);
or UO_715 (O_715,N_19947,N_19936);
nand UO_716 (O_716,N_19907,N_19917);
nor UO_717 (O_717,N_19958,N_19955);
and UO_718 (O_718,N_19892,N_19923);
nand UO_719 (O_719,N_19882,N_19871);
and UO_720 (O_720,N_19994,N_19943);
xor UO_721 (O_721,N_19877,N_19975);
nor UO_722 (O_722,N_19969,N_19979);
xor UO_723 (O_723,N_19885,N_19967);
or UO_724 (O_724,N_19874,N_19885);
and UO_725 (O_725,N_19889,N_19918);
nand UO_726 (O_726,N_19844,N_19947);
or UO_727 (O_727,N_19906,N_19958);
nor UO_728 (O_728,N_19935,N_19884);
and UO_729 (O_729,N_19841,N_19849);
nor UO_730 (O_730,N_19912,N_19841);
or UO_731 (O_731,N_19940,N_19892);
and UO_732 (O_732,N_19964,N_19960);
nand UO_733 (O_733,N_19968,N_19991);
and UO_734 (O_734,N_19935,N_19947);
nor UO_735 (O_735,N_19989,N_19855);
or UO_736 (O_736,N_19850,N_19943);
nor UO_737 (O_737,N_19969,N_19876);
nor UO_738 (O_738,N_19853,N_19859);
nand UO_739 (O_739,N_19979,N_19924);
and UO_740 (O_740,N_19907,N_19914);
nor UO_741 (O_741,N_19959,N_19951);
nor UO_742 (O_742,N_19851,N_19983);
or UO_743 (O_743,N_19877,N_19930);
nor UO_744 (O_744,N_19879,N_19906);
nor UO_745 (O_745,N_19966,N_19865);
and UO_746 (O_746,N_19869,N_19927);
nand UO_747 (O_747,N_19851,N_19975);
and UO_748 (O_748,N_19852,N_19963);
or UO_749 (O_749,N_19882,N_19866);
nor UO_750 (O_750,N_19899,N_19918);
nand UO_751 (O_751,N_19904,N_19907);
nand UO_752 (O_752,N_19902,N_19932);
nand UO_753 (O_753,N_19863,N_19966);
nor UO_754 (O_754,N_19907,N_19840);
or UO_755 (O_755,N_19889,N_19954);
nand UO_756 (O_756,N_19860,N_19947);
nand UO_757 (O_757,N_19957,N_19988);
xor UO_758 (O_758,N_19969,N_19900);
or UO_759 (O_759,N_19908,N_19964);
nor UO_760 (O_760,N_19955,N_19924);
and UO_761 (O_761,N_19967,N_19900);
nand UO_762 (O_762,N_19885,N_19958);
or UO_763 (O_763,N_19952,N_19848);
or UO_764 (O_764,N_19924,N_19921);
or UO_765 (O_765,N_19927,N_19949);
nor UO_766 (O_766,N_19995,N_19842);
nor UO_767 (O_767,N_19887,N_19928);
and UO_768 (O_768,N_19888,N_19938);
nor UO_769 (O_769,N_19965,N_19856);
or UO_770 (O_770,N_19962,N_19891);
nor UO_771 (O_771,N_19937,N_19933);
nand UO_772 (O_772,N_19923,N_19949);
or UO_773 (O_773,N_19890,N_19898);
nand UO_774 (O_774,N_19953,N_19856);
or UO_775 (O_775,N_19848,N_19945);
nor UO_776 (O_776,N_19851,N_19912);
nand UO_777 (O_777,N_19903,N_19914);
or UO_778 (O_778,N_19886,N_19969);
nor UO_779 (O_779,N_19935,N_19856);
or UO_780 (O_780,N_19924,N_19863);
nand UO_781 (O_781,N_19963,N_19950);
or UO_782 (O_782,N_19940,N_19908);
or UO_783 (O_783,N_19935,N_19844);
and UO_784 (O_784,N_19993,N_19847);
and UO_785 (O_785,N_19978,N_19985);
nor UO_786 (O_786,N_19993,N_19964);
or UO_787 (O_787,N_19952,N_19849);
nand UO_788 (O_788,N_19998,N_19872);
nand UO_789 (O_789,N_19861,N_19883);
or UO_790 (O_790,N_19873,N_19993);
xnor UO_791 (O_791,N_19967,N_19953);
and UO_792 (O_792,N_19862,N_19855);
nor UO_793 (O_793,N_19855,N_19867);
and UO_794 (O_794,N_19856,N_19963);
xnor UO_795 (O_795,N_19863,N_19848);
or UO_796 (O_796,N_19869,N_19963);
and UO_797 (O_797,N_19891,N_19925);
nand UO_798 (O_798,N_19942,N_19969);
nor UO_799 (O_799,N_19859,N_19997);
nand UO_800 (O_800,N_19852,N_19862);
nand UO_801 (O_801,N_19854,N_19887);
nand UO_802 (O_802,N_19998,N_19940);
or UO_803 (O_803,N_19960,N_19860);
and UO_804 (O_804,N_19873,N_19908);
and UO_805 (O_805,N_19959,N_19903);
nor UO_806 (O_806,N_19844,N_19858);
and UO_807 (O_807,N_19869,N_19991);
or UO_808 (O_808,N_19914,N_19882);
or UO_809 (O_809,N_19866,N_19888);
nand UO_810 (O_810,N_19905,N_19948);
nor UO_811 (O_811,N_19898,N_19940);
xor UO_812 (O_812,N_19865,N_19892);
nor UO_813 (O_813,N_19915,N_19870);
and UO_814 (O_814,N_19922,N_19896);
nand UO_815 (O_815,N_19876,N_19901);
xor UO_816 (O_816,N_19899,N_19846);
and UO_817 (O_817,N_19862,N_19960);
nand UO_818 (O_818,N_19891,N_19841);
nor UO_819 (O_819,N_19991,N_19905);
xnor UO_820 (O_820,N_19875,N_19898);
nor UO_821 (O_821,N_19998,N_19902);
or UO_822 (O_822,N_19840,N_19867);
nand UO_823 (O_823,N_19868,N_19945);
and UO_824 (O_824,N_19946,N_19857);
or UO_825 (O_825,N_19919,N_19867);
or UO_826 (O_826,N_19909,N_19854);
or UO_827 (O_827,N_19850,N_19878);
nor UO_828 (O_828,N_19855,N_19873);
and UO_829 (O_829,N_19934,N_19886);
and UO_830 (O_830,N_19851,N_19960);
nand UO_831 (O_831,N_19884,N_19846);
nor UO_832 (O_832,N_19929,N_19995);
nand UO_833 (O_833,N_19941,N_19928);
and UO_834 (O_834,N_19967,N_19850);
nand UO_835 (O_835,N_19971,N_19932);
and UO_836 (O_836,N_19922,N_19895);
nand UO_837 (O_837,N_19877,N_19908);
nor UO_838 (O_838,N_19871,N_19996);
or UO_839 (O_839,N_19965,N_19955);
and UO_840 (O_840,N_19882,N_19986);
xor UO_841 (O_841,N_19897,N_19976);
nor UO_842 (O_842,N_19849,N_19877);
and UO_843 (O_843,N_19944,N_19971);
or UO_844 (O_844,N_19986,N_19909);
or UO_845 (O_845,N_19951,N_19928);
or UO_846 (O_846,N_19907,N_19891);
nand UO_847 (O_847,N_19972,N_19989);
nor UO_848 (O_848,N_19948,N_19859);
and UO_849 (O_849,N_19984,N_19995);
and UO_850 (O_850,N_19845,N_19980);
nor UO_851 (O_851,N_19849,N_19897);
or UO_852 (O_852,N_19973,N_19841);
and UO_853 (O_853,N_19915,N_19914);
and UO_854 (O_854,N_19917,N_19844);
or UO_855 (O_855,N_19952,N_19879);
nor UO_856 (O_856,N_19881,N_19991);
or UO_857 (O_857,N_19884,N_19949);
or UO_858 (O_858,N_19894,N_19974);
or UO_859 (O_859,N_19954,N_19869);
or UO_860 (O_860,N_19855,N_19861);
nand UO_861 (O_861,N_19934,N_19988);
and UO_862 (O_862,N_19896,N_19950);
nand UO_863 (O_863,N_19903,N_19955);
and UO_864 (O_864,N_19923,N_19961);
nor UO_865 (O_865,N_19909,N_19887);
or UO_866 (O_866,N_19960,N_19968);
or UO_867 (O_867,N_19927,N_19877);
xor UO_868 (O_868,N_19957,N_19990);
or UO_869 (O_869,N_19888,N_19915);
or UO_870 (O_870,N_19852,N_19929);
and UO_871 (O_871,N_19856,N_19997);
nor UO_872 (O_872,N_19942,N_19956);
nor UO_873 (O_873,N_19954,N_19877);
xnor UO_874 (O_874,N_19882,N_19982);
or UO_875 (O_875,N_19882,N_19890);
nand UO_876 (O_876,N_19974,N_19889);
nand UO_877 (O_877,N_19958,N_19954);
nand UO_878 (O_878,N_19938,N_19878);
xnor UO_879 (O_879,N_19987,N_19886);
or UO_880 (O_880,N_19857,N_19961);
xnor UO_881 (O_881,N_19924,N_19998);
and UO_882 (O_882,N_19848,N_19995);
nand UO_883 (O_883,N_19930,N_19894);
nand UO_884 (O_884,N_19940,N_19845);
or UO_885 (O_885,N_19904,N_19949);
nand UO_886 (O_886,N_19930,N_19938);
or UO_887 (O_887,N_19905,N_19989);
and UO_888 (O_888,N_19854,N_19960);
nor UO_889 (O_889,N_19925,N_19893);
or UO_890 (O_890,N_19911,N_19845);
and UO_891 (O_891,N_19851,N_19861);
nand UO_892 (O_892,N_19903,N_19971);
nor UO_893 (O_893,N_19865,N_19907);
xnor UO_894 (O_894,N_19892,N_19968);
nor UO_895 (O_895,N_19947,N_19868);
and UO_896 (O_896,N_19895,N_19950);
and UO_897 (O_897,N_19975,N_19993);
nor UO_898 (O_898,N_19960,N_19890);
and UO_899 (O_899,N_19857,N_19947);
and UO_900 (O_900,N_19996,N_19974);
and UO_901 (O_901,N_19850,N_19972);
or UO_902 (O_902,N_19958,N_19989);
nor UO_903 (O_903,N_19844,N_19954);
or UO_904 (O_904,N_19877,N_19867);
or UO_905 (O_905,N_19945,N_19883);
xnor UO_906 (O_906,N_19884,N_19881);
nand UO_907 (O_907,N_19907,N_19977);
nand UO_908 (O_908,N_19865,N_19844);
or UO_909 (O_909,N_19871,N_19948);
nand UO_910 (O_910,N_19867,N_19865);
and UO_911 (O_911,N_19902,N_19850);
and UO_912 (O_912,N_19853,N_19950);
nand UO_913 (O_913,N_19903,N_19942);
xor UO_914 (O_914,N_19926,N_19866);
and UO_915 (O_915,N_19850,N_19916);
or UO_916 (O_916,N_19878,N_19887);
nor UO_917 (O_917,N_19915,N_19932);
nand UO_918 (O_918,N_19887,N_19848);
nor UO_919 (O_919,N_19991,N_19970);
and UO_920 (O_920,N_19963,N_19874);
and UO_921 (O_921,N_19984,N_19926);
or UO_922 (O_922,N_19940,N_19877);
and UO_923 (O_923,N_19951,N_19891);
xnor UO_924 (O_924,N_19965,N_19991);
and UO_925 (O_925,N_19915,N_19948);
nand UO_926 (O_926,N_19940,N_19865);
and UO_927 (O_927,N_19939,N_19919);
and UO_928 (O_928,N_19919,N_19844);
nor UO_929 (O_929,N_19970,N_19966);
nor UO_930 (O_930,N_19891,N_19882);
or UO_931 (O_931,N_19886,N_19903);
and UO_932 (O_932,N_19849,N_19843);
and UO_933 (O_933,N_19998,N_19849);
and UO_934 (O_934,N_19918,N_19905);
or UO_935 (O_935,N_19860,N_19968);
xor UO_936 (O_936,N_19926,N_19852);
and UO_937 (O_937,N_19996,N_19951);
or UO_938 (O_938,N_19925,N_19930);
xnor UO_939 (O_939,N_19946,N_19991);
nand UO_940 (O_940,N_19945,N_19971);
nand UO_941 (O_941,N_19977,N_19995);
and UO_942 (O_942,N_19872,N_19859);
and UO_943 (O_943,N_19930,N_19942);
nor UO_944 (O_944,N_19942,N_19954);
or UO_945 (O_945,N_19858,N_19999);
and UO_946 (O_946,N_19857,N_19871);
nand UO_947 (O_947,N_19880,N_19886);
nor UO_948 (O_948,N_19886,N_19945);
nor UO_949 (O_949,N_19868,N_19954);
nor UO_950 (O_950,N_19844,N_19998);
and UO_951 (O_951,N_19868,N_19851);
nand UO_952 (O_952,N_19913,N_19845);
or UO_953 (O_953,N_19908,N_19970);
nor UO_954 (O_954,N_19927,N_19893);
nand UO_955 (O_955,N_19970,N_19953);
or UO_956 (O_956,N_19944,N_19844);
nor UO_957 (O_957,N_19982,N_19926);
or UO_958 (O_958,N_19933,N_19866);
xnor UO_959 (O_959,N_19859,N_19871);
nor UO_960 (O_960,N_19877,N_19920);
and UO_961 (O_961,N_19908,N_19994);
nor UO_962 (O_962,N_19958,N_19944);
and UO_963 (O_963,N_19866,N_19932);
nor UO_964 (O_964,N_19844,N_19891);
nand UO_965 (O_965,N_19863,N_19985);
and UO_966 (O_966,N_19913,N_19951);
xnor UO_967 (O_967,N_19903,N_19854);
and UO_968 (O_968,N_19930,N_19984);
or UO_969 (O_969,N_19891,N_19980);
or UO_970 (O_970,N_19969,N_19934);
and UO_971 (O_971,N_19882,N_19964);
nand UO_972 (O_972,N_19968,N_19845);
xor UO_973 (O_973,N_19887,N_19858);
nand UO_974 (O_974,N_19900,N_19994);
nor UO_975 (O_975,N_19965,N_19985);
nand UO_976 (O_976,N_19894,N_19922);
and UO_977 (O_977,N_19901,N_19905);
nor UO_978 (O_978,N_19896,N_19927);
xor UO_979 (O_979,N_19859,N_19933);
nor UO_980 (O_980,N_19953,N_19883);
nand UO_981 (O_981,N_19963,N_19911);
nand UO_982 (O_982,N_19949,N_19841);
nand UO_983 (O_983,N_19964,N_19967);
nor UO_984 (O_984,N_19896,N_19897);
and UO_985 (O_985,N_19889,N_19972);
nor UO_986 (O_986,N_19866,N_19851);
nand UO_987 (O_987,N_19915,N_19916);
or UO_988 (O_988,N_19846,N_19931);
or UO_989 (O_989,N_19996,N_19845);
nor UO_990 (O_990,N_19857,N_19906);
xnor UO_991 (O_991,N_19916,N_19945);
nand UO_992 (O_992,N_19875,N_19955);
nor UO_993 (O_993,N_19988,N_19904);
nor UO_994 (O_994,N_19943,N_19898);
nor UO_995 (O_995,N_19911,N_19986);
nor UO_996 (O_996,N_19988,N_19929);
nand UO_997 (O_997,N_19915,N_19983);
nor UO_998 (O_998,N_19859,N_19869);
and UO_999 (O_999,N_19940,N_19862);
or UO_1000 (O_1000,N_19899,N_19987);
nor UO_1001 (O_1001,N_19842,N_19849);
or UO_1002 (O_1002,N_19932,N_19949);
nor UO_1003 (O_1003,N_19973,N_19861);
nand UO_1004 (O_1004,N_19918,N_19853);
and UO_1005 (O_1005,N_19940,N_19990);
nor UO_1006 (O_1006,N_19896,N_19854);
and UO_1007 (O_1007,N_19854,N_19962);
or UO_1008 (O_1008,N_19849,N_19920);
and UO_1009 (O_1009,N_19962,N_19897);
xnor UO_1010 (O_1010,N_19885,N_19944);
and UO_1011 (O_1011,N_19846,N_19999);
or UO_1012 (O_1012,N_19992,N_19981);
xor UO_1013 (O_1013,N_19949,N_19979);
nor UO_1014 (O_1014,N_19953,N_19879);
or UO_1015 (O_1015,N_19940,N_19952);
or UO_1016 (O_1016,N_19974,N_19874);
nor UO_1017 (O_1017,N_19878,N_19861);
and UO_1018 (O_1018,N_19891,N_19974);
nand UO_1019 (O_1019,N_19871,N_19894);
and UO_1020 (O_1020,N_19976,N_19999);
nand UO_1021 (O_1021,N_19920,N_19855);
nor UO_1022 (O_1022,N_19960,N_19885);
and UO_1023 (O_1023,N_19868,N_19943);
nand UO_1024 (O_1024,N_19946,N_19962);
or UO_1025 (O_1025,N_19967,N_19972);
or UO_1026 (O_1026,N_19840,N_19843);
nor UO_1027 (O_1027,N_19849,N_19914);
nor UO_1028 (O_1028,N_19887,N_19861);
nor UO_1029 (O_1029,N_19911,N_19883);
or UO_1030 (O_1030,N_19902,N_19887);
nand UO_1031 (O_1031,N_19929,N_19940);
nand UO_1032 (O_1032,N_19858,N_19856);
xor UO_1033 (O_1033,N_19910,N_19940);
and UO_1034 (O_1034,N_19883,N_19854);
and UO_1035 (O_1035,N_19937,N_19855);
nor UO_1036 (O_1036,N_19952,N_19986);
nand UO_1037 (O_1037,N_19950,N_19944);
nand UO_1038 (O_1038,N_19870,N_19951);
nor UO_1039 (O_1039,N_19888,N_19977);
xor UO_1040 (O_1040,N_19949,N_19869);
nand UO_1041 (O_1041,N_19916,N_19845);
and UO_1042 (O_1042,N_19965,N_19855);
or UO_1043 (O_1043,N_19956,N_19869);
nand UO_1044 (O_1044,N_19901,N_19922);
nand UO_1045 (O_1045,N_19996,N_19963);
nor UO_1046 (O_1046,N_19878,N_19863);
nor UO_1047 (O_1047,N_19890,N_19858);
and UO_1048 (O_1048,N_19961,N_19893);
and UO_1049 (O_1049,N_19953,N_19902);
nand UO_1050 (O_1050,N_19866,N_19966);
or UO_1051 (O_1051,N_19854,N_19957);
nand UO_1052 (O_1052,N_19991,N_19997);
nor UO_1053 (O_1053,N_19938,N_19901);
and UO_1054 (O_1054,N_19978,N_19986);
nand UO_1055 (O_1055,N_19900,N_19939);
xor UO_1056 (O_1056,N_19988,N_19979);
or UO_1057 (O_1057,N_19912,N_19848);
nand UO_1058 (O_1058,N_19989,N_19851);
and UO_1059 (O_1059,N_19884,N_19919);
or UO_1060 (O_1060,N_19927,N_19935);
and UO_1061 (O_1061,N_19917,N_19841);
and UO_1062 (O_1062,N_19910,N_19995);
xor UO_1063 (O_1063,N_19923,N_19989);
nand UO_1064 (O_1064,N_19932,N_19913);
xor UO_1065 (O_1065,N_19976,N_19879);
or UO_1066 (O_1066,N_19956,N_19954);
and UO_1067 (O_1067,N_19863,N_19856);
nand UO_1068 (O_1068,N_19974,N_19883);
nor UO_1069 (O_1069,N_19979,N_19899);
and UO_1070 (O_1070,N_19933,N_19921);
or UO_1071 (O_1071,N_19909,N_19974);
and UO_1072 (O_1072,N_19949,N_19973);
nor UO_1073 (O_1073,N_19915,N_19955);
or UO_1074 (O_1074,N_19971,N_19998);
or UO_1075 (O_1075,N_19914,N_19926);
and UO_1076 (O_1076,N_19974,N_19965);
and UO_1077 (O_1077,N_19857,N_19953);
nand UO_1078 (O_1078,N_19879,N_19851);
and UO_1079 (O_1079,N_19944,N_19970);
or UO_1080 (O_1080,N_19867,N_19892);
nor UO_1081 (O_1081,N_19936,N_19986);
nor UO_1082 (O_1082,N_19859,N_19979);
nor UO_1083 (O_1083,N_19853,N_19959);
and UO_1084 (O_1084,N_19927,N_19902);
xnor UO_1085 (O_1085,N_19881,N_19971);
nor UO_1086 (O_1086,N_19992,N_19919);
nand UO_1087 (O_1087,N_19887,N_19921);
and UO_1088 (O_1088,N_19918,N_19933);
and UO_1089 (O_1089,N_19959,N_19995);
nand UO_1090 (O_1090,N_19854,N_19944);
xnor UO_1091 (O_1091,N_19994,N_19904);
nor UO_1092 (O_1092,N_19889,N_19964);
xnor UO_1093 (O_1093,N_19847,N_19880);
and UO_1094 (O_1094,N_19982,N_19874);
nor UO_1095 (O_1095,N_19869,N_19938);
nand UO_1096 (O_1096,N_19868,N_19935);
nand UO_1097 (O_1097,N_19927,N_19873);
xnor UO_1098 (O_1098,N_19900,N_19989);
nor UO_1099 (O_1099,N_19943,N_19910);
nor UO_1100 (O_1100,N_19972,N_19867);
nor UO_1101 (O_1101,N_19991,N_19887);
nor UO_1102 (O_1102,N_19951,N_19918);
and UO_1103 (O_1103,N_19945,N_19873);
nand UO_1104 (O_1104,N_19941,N_19852);
or UO_1105 (O_1105,N_19906,N_19886);
xor UO_1106 (O_1106,N_19895,N_19988);
and UO_1107 (O_1107,N_19902,N_19926);
nand UO_1108 (O_1108,N_19992,N_19917);
and UO_1109 (O_1109,N_19941,N_19899);
and UO_1110 (O_1110,N_19867,N_19984);
nand UO_1111 (O_1111,N_19983,N_19856);
nor UO_1112 (O_1112,N_19996,N_19929);
or UO_1113 (O_1113,N_19914,N_19999);
or UO_1114 (O_1114,N_19995,N_19979);
nand UO_1115 (O_1115,N_19940,N_19994);
nand UO_1116 (O_1116,N_19966,N_19947);
and UO_1117 (O_1117,N_19947,N_19953);
nor UO_1118 (O_1118,N_19990,N_19908);
and UO_1119 (O_1119,N_19988,N_19983);
or UO_1120 (O_1120,N_19960,N_19852);
nor UO_1121 (O_1121,N_19983,N_19916);
and UO_1122 (O_1122,N_19873,N_19958);
and UO_1123 (O_1123,N_19946,N_19893);
and UO_1124 (O_1124,N_19881,N_19853);
nand UO_1125 (O_1125,N_19840,N_19963);
and UO_1126 (O_1126,N_19935,N_19953);
or UO_1127 (O_1127,N_19998,N_19860);
and UO_1128 (O_1128,N_19997,N_19923);
and UO_1129 (O_1129,N_19895,N_19871);
and UO_1130 (O_1130,N_19939,N_19986);
and UO_1131 (O_1131,N_19917,N_19991);
nor UO_1132 (O_1132,N_19899,N_19915);
or UO_1133 (O_1133,N_19844,N_19988);
and UO_1134 (O_1134,N_19872,N_19912);
and UO_1135 (O_1135,N_19914,N_19928);
or UO_1136 (O_1136,N_19984,N_19953);
nand UO_1137 (O_1137,N_19906,N_19972);
nand UO_1138 (O_1138,N_19897,N_19847);
nor UO_1139 (O_1139,N_19840,N_19998);
nand UO_1140 (O_1140,N_19989,N_19840);
or UO_1141 (O_1141,N_19862,N_19885);
or UO_1142 (O_1142,N_19887,N_19867);
nand UO_1143 (O_1143,N_19904,N_19950);
xor UO_1144 (O_1144,N_19941,N_19926);
and UO_1145 (O_1145,N_19990,N_19981);
and UO_1146 (O_1146,N_19932,N_19998);
nand UO_1147 (O_1147,N_19988,N_19963);
and UO_1148 (O_1148,N_19987,N_19863);
xnor UO_1149 (O_1149,N_19902,N_19879);
nand UO_1150 (O_1150,N_19987,N_19855);
nand UO_1151 (O_1151,N_19879,N_19916);
or UO_1152 (O_1152,N_19991,N_19944);
nor UO_1153 (O_1153,N_19897,N_19934);
nor UO_1154 (O_1154,N_19880,N_19846);
and UO_1155 (O_1155,N_19852,N_19937);
and UO_1156 (O_1156,N_19845,N_19982);
nand UO_1157 (O_1157,N_19973,N_19905);
or UO_1158 (O_1158,N_19886,N_19971);
nor UO_1159 (O_1159,N_19961,N_19869);
or UO_1160 (O_1160,N_19916,N_19996);
and UO_1161 (O_1161,N_19929,N_19969);
and UO_1162 (O_1162,N_19894,N_19902);
xor UO_1163 (O_1163,N_19840,N_19890);
nor UO_1164 (O_1164,N_19988,N_19943);
nor UO_1165 (O_1165,N_19981,N_19923);
or UO_1166 (O_1166,N_19855,N_19864);
or UO_1167 (O_1167,N_19922,N_19917);
or UO_1168 (O_1168,N_19846,N_19962);
nand UO_1169 (O_1169,N_19933,N_19992);
or UO_1170 (O_1170,N_19960,N_19915);
nor UO_1171 (O_1171,N_19866,N_19948);
xnor UO_1172 (O_1172,N_19905,N_19895);
nand UO_1173 (O_1173,N_19877,N_19844);
nor UO_1174 (O_1174,N_19979,N_19926);
nor UO_1175 (O_1175,N_19858,N_19898);
xnor UO_1176 (O_1176,N_19931,N_19943);
and UO_1177 (O_1177,N_19886,N_19859);
and UO_1178 (O_1178,N_19989,N_19936);
xor UO_1179 (O_1179,N_19967,N_19991);
and UO_1180 (O_1180,N_19943,N_19923);
and UO_1181 (O_1181,N_19923,N_19916);
xor UO_1182 (O_1182,N_19975,N_19987);
and UO_1183 (O_1183,N_19955,N_19947);
nand UO_1184 (O_1184,N_19845,N_19894);
or UO_1185 (O_1185,N_19874,N_19972);
and UO_1186 (O_1186,N_19966,N_19958);
or UO_1187 (O_1187,N_19985,N_19963);
or UO_1188 (O_1188,N_19846,N_19955);
and UO_1189 (O_1189,N_19995,N_19869);
nand UO_1190 (O_1190,N_19994,N_19962);
nand UO_1191 (O_1191,N_19909,N_19840);
nor UO_1192 (O_1192,N_19927,N_19962);
xnor UO_1193 (O_1193,N_19862,N_19947);
and UO_1194 (O_1194,N_19965,N_19964);
xnor UO_1195 (O_1195,N_19987,N_19945);
or UO_1196 (O_1196,N_19947,N_19992);
and UO_1197 (O_1197,N_19905,N_19993);
or UO_1198 (O_1198,N_19911,N_19973);
and UO_1199 (O_1199,N_19841,N_19864);
or UO_1200 (O_1200,N_19901,N_19855);
nor UO_1201 (O_1201,N_19978,N_19898);
nor UO_1202 (O_1202,N_19868,N_19989);
and UO_1203 (O_1203,N_19982,N_19987);
nor UO_1204 (O_1204,N_19973,N_19966);
or UO_1205 (O_1205,N_19864,N_19994);
nor UO_1206 (O_1206,N_19946,N_19939);
or UO_1207 (O_1207,N_19858,N_19945);
or UO_1208 (O_1208,N_19927,N_19867);
or UO_1209 (O_1209,N_19936,N_19876);
nand UO_1210 (O_1210,N_19859,N_19840);
nand UO_1211 (O_1211,N_19980,N_19945);
nand UO_1212 (O_1212,N_19920,N_19883);
and UO_1213 (O_1213,N_19921,N_19956);
or UO_1214 (O_1214,N_19934,N_19977);
nand UO_1215 (O_1215,N_19845,N_19947);
xor UO_1216 (O_1216,N_19971,N_19948);
xnor UO_1217 (O_1217,N_19888,N_19971);
nor UO_1218 (O_1218,N_19890,N_19905);
or UO_1219 (O_1219,N_19999,N_19954);
nand UO_1220 (O_1220,N_19885,N_19934);
and UO_1221 (O_1221,N_19997,N_19843);
xnor UO_1222 (O_1222,N_19847,N_19973);
nand UO_1223 (O_1223,N_19972,N_19842);
or UO_1224 (O_1224,N_19983,N_19984);
or UO_1225 (O_1225,N_19943,N_19963);
nor UO_1226 (O_1226,N_19867,N_19850);
nor UO_1227 (O_1227,N_19953,N_19908);
or UO_1228 (O_1228,N_19906,N_19878);
nand UO_1229 (O_1229,N_19932,N_19840);
or UO_1230 (O_1230,N_19847,N_19976);
or UO_1231 (O_1231,N_19962,N_19896);
nor UO_1232 (O_1232,N_19918,N_19965);
or UO_1233 (O_1233,N_19845,N_19971);
and UO_1234 (O_1234,N_19963,N_19907);
and UO_1235 (O_1235,N_19939,N_19980);
nand UO_1236 (O_1236,N_19909,N_19891);
nand UO_1237 (O_1237,N_19955,N_19878);
or UO_1238 (O_1238,N_19934,N_19884);
nor UO_1239 (O_1239,N_19952,N_19965);
xnor UO_1240 (O_1240,N_19991,N_19947);
and UO_1241 (O_1241,N_19962,N_19953);
or UO_1242 (O_1242,N_19974,N_19846);
nand UO_1243 (O_1243,N_19845,N_19985);
nand UO_1244 (O_1244,N_19913,N_19896);
nor UO_1245 (O_1245,N_19919,N_19898);
and UO_1246 (O_1246,N_19933,N_19952);
and UO_1247 (O_1247,N_19849,N_19888);
or UO_1248 (O_1248,N_19848,N_19861);
nand UO_1249 (O_1249,N_19934,N_19855);
xor UO_1250 (O_1250,N_19987,N_19931);
or UO_1251 (O_1251,N_19952,N_19843);
xor UO_1252 (O_1252,N_19942,N_19990);
and UO_1253 (O_1253,N_19860,N_19927);
nor UO_1254 (O_1254,N_19844,N_19860);
and UO_1255 (O_1255,N_19974,N_19862);
and UO_1256 (O_1256,N_19883,N_19844);
and UO_1257 (O_1257,N_19852,N_19910);
xnor UO_1258 (O_1258,N_19882,N_19851);
nor UO_1259 (O_1259,N_19931,N_19874);
nor UO_1260 (O_1260,N_19876,N_19908);
nor UO_1261 (O_1261,N_19950,N_19969);
and UO_1262 (O_1262,N_19980,N_19960);
or UO_1263 (O_1263,N_19864,N_19888);
and UO_1264 (O_1264,N_19844,N_19926);
nand UO_1265 (O_1265,N_19943,N_19974);
nor UO_1266 (O_1266,N_19849,N_19902);
nand UO_1267 (O_1267,N_19917,N_19968);
nor UO_1268 (O_1268,N_19922,N_19905);
and UO_1269 (O_1269,N_19900,N_19848);
xor UO_1270 (O_1270,N_19884,N_19842);
nor UO_1271 (O_1271,N_19845,N_19914);
nor UO_1272 (O_1272,N_19949,N_19925);
nand UO_1273 (O_1273,N_19904,N_19956);
or UO_1274 (O_1274,N_19894,N_19873);
nor UO_1275 (O_1275,N_19930,N_19917);
xnor UO_1276 (O_1276,N_19971,N_19901);
and UO_1277 (O_1277,N_19931,N_19958);
or UO_1278 (O_1278,N_19996,N_19962);
and UO_1279 (O_1279,N_19885,N_19945);
nor UO_1280 (O_1280,N_19888,N_19842);
nand UO_1281 (O_1281,N_19848,N_19904);
and UO_1282 (O_1282,N_19958,N_19841);
xnor UO_1283 (O_1283,N_19973,N_19918);
and UO_1284 (O_1284,N_19852,N_19842);
and UO_1285 (O_1285,N_19980,N_19924);
nor UO_1286 (O_1286,N_19914,N_19986);
or UO_1287 (O_1287,N_19907,N_19944);
and UO_1288 (O_1288,N_19845,N_19964);
or UO_1289 (O_1289,N_19875,N_19862);
or UO_1290 (O_1290,N_19907,N_19981);
nand UO_1291 (O_1291,N_19851,N_19911);
and UO_1292 (O_1292,N_19874,N_19993);
nor UO_1293 (O_1293,N_19955,N_19976);
and UO_1294 (O_1294,N_19852,N_19882);
nor UO_1295 (O_1295,N_19868,N_19965);
or UO_1296 (O_1296,N_19860,N_19984);
nor UO_1297 (O_1297,N_19955,N_19907);
nor UO_1298 (O_1298,N_19987,N_19900);
or UO_1299 (O_1299,N_19988,N_19874);
xor UO_1300 (O_1300,N_19950,N_19866);
or UO_1301 (O_1301,N_19878,N_19933);
or UO_1302 (O_1302,N_19969,N_19957);
nand UO_1303 (O_1303,N_19951,N_19893);
and UO_1304 (O_1304,N_19982,N_19843);
and UO_1305 (O_1305,N_19989,N_19946);
nand UO_1306 (O_1306,N_19863,N_19923);
nand UO_1307 (O_1307,N_19854,N_19947);
xnor UO_1308 (O_1308,N_19984,N_19937);
or UO_1309 (O_1309,N_19990,N_19852);
and UO_1310 (O_1310,N_19997,N_19882);
and UO_1311 (O_1311,N_19901,N_19902);
or UO_1312 (O_1312,N_19864,N_19840);
and UO_1313 (O_1313,N_19888,N_19859);
and UO_1314 (O_1314,N_19964,N_19921);
nor UO_1315 (O_1315,N_19958,N_19953);
and UO_1316 (O_1316,N_19957,N_19913);
and UO_1317 (O_1317,N_19913,N_19929);
or UO_1318 (O_1318,N_19931,N_19926);
or UO_1319 (O_1319,N_19863,N_19990);
and UO_1320 (O_1320,N_19908,N_19950);
nand UO_1321 (O_1321,N_19989,N_19842);
nand UO_1322 (O_1322,N_19902,N_19937);
nand UO_1323 (O_1323,N_19884,N_19953);
nand UO_1324 (O_1324,N_19916,N_19893);
nor UO_1325 (O_1325,N_19971,N_19875);
nor UO_1326 (O_1326,N_19915,N_19963);
or UO_1327 (O_1327,N_19947,N_19952);
or UO_1328 (O_1328,N_19862,N_19849);
nor UO_1329 (O_1329,N_19908,N_19870);
and UO_1330 (O_1330,N_19969,N_19980);
and UO_1331 (O_1331,N_19926,N_19843);
nor UO_1332 (O_1332,N_19963,N_19920);
xnor UO_1333 (O_1333,N_19929,N_19927);
or UO_1334 (O_1334,N_19865,N_19945);
nor UO_1335 (O_1335,N_19869,N_19840);
nand UO_1336 (O_1336,N_19868,N_19875);
nor UO_1337 (O_1337,N_19900,N_19885);
and UO_1338 (O_1338,N_19939,N_19916);
or UO_1339 (O_1339,N_19853,N_19870);
nor UO_1340 (O_1340,N_19992,N_19853);
and UO_1341 (O_1341,N_19981,N_19859);
and UO_1342 (O_1342,N_19927,N_19996);
xor UO_1343 (O_1343,N_19854,N_19849);
and UO_1344 (O_1344,N_19951,N_19909);
or UO_1345 (O_1345,N_19893,N_19915);
or UO_1346 (O_1346,N_19999,N_19947);
nand UO_1347 (O_1347,N_19848,N_19852);
xnor UO_1348 (O_1348,N_19896,N_19938);
nor UO_1349 (O_1349,N_19899,N_19945);
or UO_1350 (O_1350,N_19957,N_19937);
nand UO_1351 (O_1351,N_19856,N_19974);
or UO_1352 (O_1352,N_19926,N_19863);
xnor UO_1353 (O_1353,N_19852,N_19977);
nor UO_1354 (O_1354,N_19972,N_19860);
or UO_1355 (O_1355,N_19992,N_19976);
xnor UO_1356 (O_1356,N_19854,N_19929);
nand UO_1357 (O_1357,N_19887,N_19964);
and UO_1358 (O_1358,N_19852,N_19876);
and UO_1359 (O_1359,N_19859,N_19864);
or UO_1360 (O_1360,N_19881,N_19997);
nand UO_1361 (O_1361,N_19897,N_19928);
or UO_1362 (O_1362,N_19873,N_19911);
nor UO_1363 (O_1363,N_19877,N_19887);
or UO_1364 (O_1364,N_19877,N_19894);
nand UO_1365 (O_1365,N_19911,N_19996);
or UO_1366 (O_1366,N_19954,N_19930);
nor UO_1367 (O_1367,N_19998,N_19934);
or UO_1368 (O_1368,N_19907,N_19845);
xor UO_1369 (O_1369,N_19911,N_19915);
xnor UO_1370 (O_1370,N_19858,N_19984);
nand UO_1371 (O_1371,N_19923,N_19927);
xnor UO_1372 (O_1372,N_19866,N_19918);
nand UO_1373 (O_1373,N_19899,N_19913);
nor UO_1374 (O_1374,N_19942,N_19924);
nor UO_1375 (O_1375,N_19843,N_19996);
nor UO_1376 (O_1376,N_19860,N_19993);
nor UO_1377 (O_1377,N_19959,N_19910);
or UO_1378 (O_1378,N_19898,N_19853);
or UO_1379 (O_1379,N_19875,N_19989);
and UO_1380 (O_1380,N_19908,N_19929);
or UO_1381 (O_1381,N_19987,N_19954);
and UO_1382 (O_1382,N_19906,N_19848);
nor UO_1383 (O_1383,N_19845,N_19997);
nand UO_1384 (O_1384,N_19858,N_19994);
nand UO_1385 (O_1385,N_19867,N_19912);
xor UO_1386 (O_1386,N_19918,N_19841);
nor UO_1387 (O_1387,N_19886,N_19991);
nor UO_1388 (O_1388,N_19905,N_19972);
and UO_1389 (O_1389,N_19856,N_19911);
xor UO_1390 (O_1390,N_19948,N_19843);
and UO_1391 (O_1391,N_19939,N_19956);
or UO_1392 (O_1392,N_19840,N_19871);
and UO_1393 (O_1393,N_19921,N_19931);
nand UO_1394 (O_1394,N_19850,N_19961);
nand UO_1395 (O_1395,N_19877,N_19922);
nand UO_1396 (O_1396,N_19982,N_19923);
nand UO_1397 (O_1397,N_19947,N_19871);
nand UO_1398 (O_1398,N_19973,N_19933);
or UO_1399 (O_1399,N_19875,N_19986);
and UO_1400 (O_1400,N_19862,N_19845);
and UO_1401 (O_1401,N_19963,N_19862);
nor UO_1402 (O_1402,N_19968,N_19920);
nand UO_1403 (O_1403,N_19922,N_19844);
nand UO_1404 (O_1404,N_19919,N_19917);
xor UO_1405 (O_1405,N_19958,N_19927);
and UO_1406 (O_1406,N_19962,N_19952);
and UO_1407 (O_1407,N_19890,N_19871);
nand UO_1408 (O_1408,N_19868,N_19976);
nand UO_1409 (O_1409,N_19999,N_19936);
and UO_1410 (O_1410,N_19905,N_19969);
nand UO_1411 (O_1411,N_19915,N_19995);
and UO_1412 (O_1412,N_19965,N_19933);
nand UO_1413 (O_1413,N_19939,N_19918);
or UO_1414 (O_1414,N_19988,N_19885);
or UO_1415 (O_1415,N_19920,N_19871);
nand UO_1416 (O_1416,N_19931,N_19864);
and UO_1417 (O_1417,N_19971,N_19975);
nor UO_1418 (O_1418,N_19963,N_19929);
nor UO_1419 (O_1419,N_19939,N_19999);
or UO_1420 (O_1420,N_19963,N_19993);
nor UO_1421 (O_1421,N_19992,N_19847);
or UO_1422 (O_1422,N_19855,N_19892);
or UO_1423 (O_1423,N_19853,N_19979);
xnor UO_1424 (O_1424,N_19846,N_19970);
nand UO_1425 (O_1425,N_19963,N_19854);
nor UO_1426 (O_1426,N_19931,N_19887);
or UO_1427 (O_1427,N_19990,N_19898);
nand UO_1428 (O_1428,N_19942,N_19941);
or UO_1429 (O_1429,N_19982,N_19873);
xnor UO_1430 (O_1430,N_19856,N_19947);
and UO_1431 (O_1431,N_19981,N_19964);
nand UO_1432 (O_1432,N_19882,N_19951);
nand UO_1433 (O_1433,N_19855,N_19977);
or UO_1434 (O_1434,N_19873,N_19938);
nor UO_1435 (O_1435,N_19847,N_19920);
and UO_1436 (O_1436,N_19985,N_19920);
nand UO_1437 (O_1437,N_19878,N_19916);
or UO_1438 (O_1438,N_19903,N_19907);
nand UO_1439 (O_1439,N_19947,N_19876);
nand UO_1440 (O_1440,N_19922,N_19906);
nor UO_1441 (O_1441,N_19964,N_19959);
and UO_1442 (O_1442,N_19870,N_19905);
nor UO_1443 (O_1443,N_19850,N_19897);
and UO_1444 (O_1444,N_19979,N_19845);
nand UO_1445 (O_1445,N_19977,N_19994);
nor UO_1446 (O_1446,N_19859,N_19974);
and UO_1447 (O_1447,N_19853,N_19908);
or UO_1448 (O_1448,N_19914,N_19848);
or UO_1449 (O_1449,N_19949,N_19853);
nand UO_1450 (O_1450,N_19855,N_19951);
or UO_1451 (O_1451,N_19930,N_19927);
or UO_1452 (O_1452,N_19888,N_19957);
nand UO_1453 (O_1453,N_19937,N_19867);
nor UO_1454 (O_1454,N_19935,N_19955);
nor UO_1455 (O_1455,N_19873,N_19933);
and UO_1456 (O_1456,N_19995,N_19925);
and UO_1457 (O_1457,N_19865,N_19943);
nor UO_1458 (O_1458,N_19931,N_19905);
xnor UO_1459 (O_1459,N_19974,N_19901);
nor UO_1460 (O_1460,N_19881,N_19867);
or UO_1461 (O_1461,N_19941,N_19998);
nor UO_1462 (O_1462,N_19853,N_19911);
nand UO_1463 (O_1463,N_19889,N_19963);
or UO_1464 (O_1464,N_19899,N_19989);
xor UO_1465 (O_1465,N_19993,N_19945);
or UO_1466 (O_1466,N_19900,N_19886);
nand UO_1467 (O_1467,N_19912,N_19946);
nor UO_1468 (O_1468,N_19999,N_19890);
nand UO_1469 (O_1469,N_19926,N_19909);
and UO_1470 (O_1470,N_19957,N_19936);
xnor UO_1471 (O_1471,N_19870,N_19966);
nor UO_1472 (O_1472,N_19968,N_19948);
or UO_1473 (O_1473,N_19975,N_19920);
and UO_1474 (O_1474,N_19976,N_19903);
or UO_1475 (O_1475,N_19924,N_19937);
or UO_1476 (O_1476,N_19973,N_19996);
and UO_1477 (O_1477,N_19950,N_19975);
nand UO_1478 (O_1478,N_19967,N_19874);
nand UO_1479 (O_1479,N_19995,N_19892);
or UO_1480 (O_1480,N_19975,N_19943);
and UO_1481 (O_1481,N_19907,N_19969);
nor UO_1482 (O_1482,N_19960,N_19922);
or UO_1483 (O_1483,N_19977,N_19872);
and UO_1484 (O_1484,N_19965,N_19871);
or UO_1485 (O_1485,N_19859,N_19990);
or UO_1486 (O_1486,N_19929,N_19945);
nand UO_1487 (O_1487,N_19971,N_19889);
and UO_1488 (O_1488,N_19942,N_19866);
and UO_1489 (O_1489,N_19927,N_19925);
and UO_1490 (O_1490,N_19894,N_19994);
and UO_1491 (O_1491,N_19856,N_19918);
nor UO_1492 (O_1492,N_19978,N_19892);
and UO_1493 (O_1493,N_19998,N_19855);
nor UO_1494 (O_1494,N_19912,N_19863);
nor UO_1495 (O_1495,N_19849,N_19945);
nand UO_1496 (O_1496,N_19845,N_19875);
or UO_1497 (O_1497,N_19855,N_19890);
nor UO_1498 (O_1498,N_19879,N_19899);
nor UO_1499 (O_1499,N_19937,N_19918);
nand UO_1500 (O_1500,N_19996,N_19870);
or UO_1501 (O_1501,N_19843,N_19846);
nand UO_1502 (O_1502,N_19875,N_19969);
nor UO_1503 (O_1503,N_19964,N_19875);
and UO_1504 (O_1504,N_19911,N_19943);
and UO_1505 (O_1505,N_19871,N_19937);
and UO_1506 (O_1506,N_19851,N_19938);
or UO_1507 (O_1507,N_19878,N_19879);
and UO_1508 (O_1508,N_19854,N_19991);
nor UO_1509 (O_1509,N_19867,N_19849);
or UO_1510 (O_1510,N_19911,N_19974);
nand UO_1511 (O_1511,N_19863,N_19997);
and UO_1512 (O_1512,N_19860,N_19930);
nand UO_1513 (O_1513,N_19840,N_19889);
nor UO_1514 (O_1514,N_19878,N_19970);
xor UO_1515 (O_1515,N_19916,N_19906);
or UO_1516 (O_1516,N_19840,N_19972);
and UO_1517 (O_1517,N_19954,N_19953);
or UO_1518 (O_1518,N_19864,N_19923);
nand UO_1519 (O_1519,N_19909,N_19932);
and UO_1520 (O_1520,N_19971,N_19915);
and UO_1521 (O_1521,N_19993,N_19880);
or UO_1522 (O_1522,N_19895,N_19883);
or UO_1523 (O_1523,N_19870,N_19983);
and UO_1524 (O_1524,N_19936,N_19860);
nor UO_1525 (O_1525,N_19940,N_19900);
or UO_1526 (O_1526,N_19943,N_19964);
or UO_1527 (O_1527,N_19929,N_19883);
or UO_1528 (O_1528,N_19961,N_19872);
nor UO_1529 (O_1529,N_19946,N_19972);
nor UO_1530 (O_1530,N_19885,N_19986);
or UO_1531 (O_1531,N_19885,N_19979);
nand UO_1532 (O_1532,N_19966,N_19916);
xor UO_1533 (O_1533,N_19967,N_19920);
and UO_1534 (O_1534,N_19904,N_19964);
nand UO_1535 (O_1535,N_19899,N_19875);
or UO_1536 (O_1536,N_19870,N_19862);
and UO_1537 (O_1537,N_19890,N_19857);
or UO_1538 (O_1538,N_19881,N_19987);
or UO_1539 (O_1539,N_19892,N_19998);
or UO_1540 (O_1540,N_19945,N_19985);
nand UO_1541 (O_1541,N_19912,N_19923);
and UO_1542 (O_1542,N_19860,N_19995);
nor UO_1543 (O_1543,N_19937,N_19860);
or UO_1544 (O_1544,N_19977,N_19869);
or UO_1545 (O_1545,N_19900,N_19878);
or UO_1546 (O_1546,N_19880,N_19928);
and UO_1547 (O_1547,N_19920,N_19953);
nand UO_1548 (O_1548,N_19997,N_19877);
nand UO_1549 (O_1549,N_19900,N_19972);
and UO_1550 (O_1550,N_19941,N_19846);
nand UO_1551 (O_1551,N_19974,N_19935);
nand UO_1552 (O_1552,N_19972,N_19971);
nand UO_1553 (O_1553,N_19851,N_19889);
nor UO_1554 (O_1554,N_19937,N_19940);
nand UO_1555 (O_1555,N_19900,N_19857);
nand UO_1556 (O_1556,N_19885,N_19875);
or UO_1557 (O_1557,N_19993,N_19902);
xor UO_1558 (O_1558,N_19903,N_19929);
nor UO_1559 (O_1559,N_19917,N_19874);
and UO_1560 (O_1560,N_19966,N_19905);
or UO_1561 (O_1561,N_19932,N_19859);
xnor UO_1562 (O_1562,N_19898,N_19984);
nand UO_1563 (O_1563,N_19841,N_19846);
xnor UO_1564 (O_1564,N_19984,N_19998);
nand UO_1565 (O_1565,N_19938,N_19900);
nor UO_1566 (O_1566,N_19873,N_19966);
nor UO_1567 (O_1567,N_19919,N_19857);
nand UO_1568 (O_1568,N_19953,N_19882);
nor UO_1569 (O_1569,N_19971,N_19977);
nand UO_1570 (O_1570,N_19943,N_19900);
nor UO_1571 (O_1571,N_19915,N_19903);
and UO_1572 (O_1572,N_19910,N_19963);
nor UO_1573 (O_1573,N_19889,N_19898);
nor UO_1574 (O_1574,N_19869,N_19973);
and UO_1575 (O_1575,N_19920,N_19882);
nor UO_1576 (O_1576,N_19845,N_19993);
xnor UO_1577 (O_1577,N_19959,N_19876);
nor UO_1578 (O_1578,N_19985,N_19961);
nand UO_1579 (O_1579,N_19845,N_19948);
or UO_1580 (O_1580,N_19893,N_19896);
and UO_1581 (O_1581,N_19952,N_19969);
nand UO_1582 (O_1582,N_19887,N_19976);
and UO_1583 (O_1583,N_19989,N_19993);
nand UO_1584 (O_1584,N_19911,N_19953);
or UO_1585 (O_1585,N_19929,N_19862);
or UO_1586 (O_1586,N_19908,N_19895);
xnor UO_1587 (O_1587,N_19983,N_19921);
and UO_1588 (O_1588,N_19922,N_19998);
or UO_1589 (O_1589,N_19891,N_19993);
or UO_1590 (O_1590,N_19913,N_19848);
and UO_1591 (O_1591,N_19914,N_19900);
or UO_1592 (O_1592,N_19927,N_19991);
nand UO_1593 (O_1593,N_19931,N_19886);
or UO_1594 (O_1594,N_19976,N_19938);
nor UO_1595 (O_1595,N_19976,N_19854);
xor UO_1596 (O_1596,N_19944,N_19993);
nand UO_1597 (O_1597,N_19959,N_19899);
or UO_1598 (O_1598,N_19876,N_19844);
nor UO_1599 (O_1599,N_19902,N_19912);
nand UO_1600 (O_1600,N_19855,N_19885);
nor UO_1601 (O_1601,N_19949,N_19946);
and UO_1602 (O_1602,N_19847,N_19848);
or UO_1603 (O_1603,N_19894,N_19903);
or UO_1604 (O_1604,N_19865,N_19883);
or UO_1605 (O_1605,N_19852,N_19982);
or UO_1606 (O_1606,N_19930,N_19870);
and UO_1607 (O_1607,N_19882,N_19912);
or UO_1608 (O_1608,N_19858,N_19925);
nand UO_1609 (O_1609,N_19955,N_19852);
nor UO_1610 (O_1610,N_19948,N_19907);
and UO_1611 (O_1611,N_19880,N_19942);
nand UO_1612 (O_1612,N_19842,N_19904);
xor UO_1613 (O_1613,N_19995,N_19933);
nand UO_1614 (O_1614,N_19898,N_19867);
nor UO_1615 (O_1615,N_19874,N_19968);
or UO_1616 (O_1616,N_19852,N_19905);
or UO_1617 (O_1617,N_19929,N_19864);
or UO_1618 (O_1618,N_19913,N_19980);
nand UO_1619 (O_1619,N_19959,N_19895);
and UO_1620 (O_1620,N_19873,N_19979);
xnor UO_1621 (O_1621,N_19961,N_19879);
or UO_1622 (O_1622,N_19988,N_19858);
or UO_1623 (O_1623,N_19961,N_19897);
and UO_1624 (O_1624,N_19896,N_19975);
and UO_1625 (O_1625,N_19985,N_19862);
and UO_1626 (O_1626,N_19941,N_19876);
or UO_1627 (O_1627,N_19856,N_19946);
nor UO_1628 (O_1628,N_19953,N_19863);
or UO_1629 (O_1629,N_19909,N_19984);
and UO_1630 (O_1630,N_19874,N_19969);
or UO_1631 (O_1631,N_19959,N_19931);
and UO_1632 (O_1632,N_19952,N_19841);
or UO_1633 (O_1633,N_19891,N_19994);
xnor UO_1634 (O_1634,N_19873,N_19977);
nand UO_1635 (O_1635,N_19910,N_19900);
nand UO_1636 (O_1636,N_19885,N_19954);
and UO_1637 (O_1637,N_19891,N_19954);
nor UO_1638 (O_1638,N_19933,N_19870);
or UO_1639 (O_1639,N_19980,N_19892);
nand UO_1640 (O_1640,N_19939,N_19866);
nand UO_1641 (O_1641,N_19855,N_19868);
or UO_1642 (O_1642,N_19898,N_19998);
or UO_1643 (O_1643,N_19907,N_19906);
or UO_1644 (O_1644,N_19842,N_19906);
or UO_1645 (O_1645,N_19948,N_19922);
and UO_1646 (O_1646,N_19905,N_19947);
or UO_1647 (O_1647,N_19897,N_19878);
xor UO_1648 (O_1648,N_19965,N_19916);
nand UO_1649 (O_1649,N_19929,N_19848);
nor UO_1650 (O_1650,N_19987,N_19935);
nor UO_1651 (O_1651,N_19981,N_19945);
or UO_1652 (O_1652,N_19898,N_19905);
or UO_1653 (O_1653,N_19956,N_19946);
xnor UO_1654 (O_1654,N_19844,N_19899);
xnor UO_1655 (O_1655,N_19855,N_19875);
and UO_1656 (O_1656,N_19995,N_19960);
nand UO_1657 (O_1657,N_19989,N_19925);
nand UO_1658 (O_1658,N_19862,N_19851);
or UO_1659 (O_1659,N_19979,N_19894);
xnor UO_1660 (O_1660,N_19852,N_19860);
nand UO_1661 (O_1661,N_19987,N_19934);
or UO_1662 (O_1662,N_19854,N_19969);
xor UO_1663 (O_1663,N_19955,N_19866);
nor UO_1664 (O_1664,N_19994,N_19849);
nand UO_1665 (O_1665,N_19957,N_19958);
nand UO_1666 (O_1666,N_19849,N_19901);
nor UO_1667 (O_1667,N_19929,N_19909);
xnor UO_1668 (O_1668,N_19890,N_19867);
and UO_1669 (O_1669,N_19950,N_19876);
nor UO_1670 (O_1670,N_19995,N_19919);
and UO_1671 (O_1671,N_19981,N_19852);
nand UO_1672 (O_1672,N_19847,N_19988);
xnor UO_1673 (O_1673,N_19971,N_19864);
xnor UO_1674 (O_1674,N_19970,N_19993);
or UO_1675 (O_1675,N_19979,N_19858);
and UO_1676 (O_1676,N_19973,N_19900);
nand UO_1677 (O_1677,N_19908,N_19945);
nand UO_1678 (O_1678,N_19965,N_19902);
or UO_1679 (O_1679,N_19974,N_19966);
xor UO_1680 (O_1680,N_19999,N_19898);
nand UO_1681 (O_1681,N_19883,N_19910);
and UO_1682 (O_1682,N_19900,N_19952);
xnor UO_1683 (O_1683,N_19925,N_19951);
or UO_1684 (O_1684,N_19845,N_19899);
nand UO_1685 (O_1685,N_19913,N_19842);
nor UO_1686 (O_1686,N_19969,N_19890);
and UO_1687 (O_1687,N_19933,N_19904);
xor UO_1688 (O_1688,N_19943,N_19979);
nand UO_1689 (O_1689,N_19887,N_19866);
nand UO_1690 (O_1690,N_19991,N_19844);
and UO_1691 (O_1691,N_19906,N_19908);
nor UO_1692 (O_1692,N_19863,N_19841);
or UO_1693 (O_1693,N_19939,N_19868);
xor UO_1694 (O_1694,N_19978,N_19900);
xnor UO_1695 (O_1695,N_19947,N_19877);
nand UO_1696 (O_1696,N_19843,N_19853);
xnor UO_1697 (O_1697,N_19987,N_19876);
nand UO_1698 (O_1698,N_19876,N_19899);
nand UO_1699 (O_1699,N_19917,N_19951);
nor UO_1700 (O_1700,N_19885,N_19980);
and UO_1701 (O_1701,N_19896,N_19841);
nand UO_1702 (O_1702,N_19843,N_19955);
nor UO_1703 (O_1703,N_19880,N_19929);
and UO_1704 (O_1704,N_19954,N_19921);
or UO_1705 (O_1705,N_19942,N_19895);
nor UO_1706 (O_1706,N_19870,N_19868);
or UO_1707 (O_1707,N_19932,N_19862);
or UO_1708 (O_1708,N_19865,N_19911);
and UO_1709 (O_1709,N_19971,N_19910);
and UO_1710 (O_1710,N_19899,N_19917);
xor UO_1711 (O_1711,N_19937,N_19980);
or UO_1712 (O_1712,N_19952,N_19869);
or UO_1713 (O_1713,N_19881,N_19923);
xnor UO_1714 (O_1714,N_19950,N_19890);
nor UO_1715 (O_1715,N_19896,N_19966);
and UO_1716 (O_1716,N_19948,N_19920);
or UO_1717 (O_1717,N_19976,N_19844);
nand UO_1718 (O_1718,N_19889,N_19875);
or UO_1719 (O_1719,N_19952,N_19919);
nor UO_1720 (O_1720,N_19903,N_19848);
nor UO_1721 (O_1721,N_19914,N_19996);
and UO_1722 (O_1722,N_19895,N_19937);
nand UO_1723 (O_1723,N_19852,N_19939);
nor UO_1724 (O_1724,N_19905,N_19877);
nor UO_1725 (O_1725,N_19990,N_19867);
nand UO_1726 (O_1726,N_19941,N_19853);
or UO_1727 (O_1727,N_19865,N_19906);
nand UO_1728 (O_1728,N_19870,N_19937);
xor UO_1729 (O_1729,N_19940,N_19867);
nor UO_1730 (O_1730,N_19955,N_19936);
nand UO_1731 (O_1731,N_19996,N_19964);
and UO_1732 (O_1732,N_19959,N_19867);
xnor UO_1733 (O_1733,N_19942,N_19879);
or UO_1734 (O_1734,N_19955,N_19933);
and UO_1735 (O_1735,N_19990,N_19994);
nand UO_1736 (O_1736,N_19915,N_19876);
nand UO_1737 (O_1737,N_19973,N_19987);
or UO_1738 (O_1738,N_19914,N_19898);
or UO_1739 (O_1739,N_19897,N_19948);
nor UO_1740 (O_1740,N_19920,N_19973);
and UO_1741 (O_1741,N_19933,N_19953);
xor UO_1742 (O_1742,N_19862,N_19939);
nor UO_1743 (O_1743,N_19945,N_19904);
or UO_1744 (O_1744,N_19882,N_19969);
and UO_1745 (O_1745,N_19878,N_19910);
xor UO_1746 (O_1746,N_19943,N_19909);
and UO_1747 (O_1747,N_19984,N_19927);
or UO_1748 (O_1748,N_19912,N_19929);
nor UO_1749 (O_1749,N_19860,N_19933);
and UO_1750 (O_1750,N_19928,N_19989);
nor UO_1751 (O_1751,N_19947,N_19893);
nor UO_1752 (O_1752,N_19966,N_19923);
or UO_1753 (O_1753,N_19945,N_19892);
and UO_1754 (O_1754,N_19912,N_19987);
nor UO_1755 (O_1755,N_19909,N_19853);
and UO_1756 (O_1756,N_19847,N_19964);
nor UO_1757 (O_1757,N_19971,N_19872);
nand UO_1758 (O_1758,N_19987,N_19918);
xor UO_1759 (O_1759,N_19943,N_19888);
xnor UO_1760 (O_1760,N_19958,N_19917);
xor UO_1761 (O_1761,N_19919,N_19926);
or UO_1762 (O_1762,N_19937,N_19954);
or UO_1763 (O_1763,N_19968,N_19902);
or UO_1764 (O_1764,N_19886,N_19961);
nor UO_1765 (O_1765,N_19967,N_19947);
nor UO_1766 (O_1766,N_19877,N_19906);
nor UO_1767 (O_1767,N_19865,N_19898);
nor UO_1768 (O_1768,N_19958,N_19986);
or UO_1769 (O_1769,N_19853,N_19877);
xor UO_1770 (O_1770,N_19991,N_19864);
or UO_1771 (O_1771,N_19890,N_19934);
and UO_1772 (O_1772,N_19922,N_19898);
or UO_1773 (O_1773,N_19893,N_19997);
nand UO_1774 (O_1774,N_19991,N_19926);
nor UO_1775 (O_1775,N_19960,N_19954);
nor UO_1776 (O_1776,N_19999,N_19856);
and UO_1777 (O_1777,N_19898,N_19886);
nand UO_1778 (O_1778,N_19997,N_19976);
nor UO_1779 (O_1779,N_19919,N_19900);
nand UO_1780 (O_1780,N_19987,N_19944);
xor UO_1781 (O_1781,N_19852,N_19898);
nand UO_1782 (O_1782,N_19846,N_19860);
nor UO_1783 (O_1783,N_19997,N_19932);
nand UO_1784 (O_1784,N_19884,N_19964);
nand UO_1785 (O_1785,N_19884,N_19894);
nand UO_1786 (O_1786,N_19924,N_19940);
or UO_1787 (O_1787,N_19971,N_19968);
nor UO_1788 (O_1788,N_19988,N_19906);
and UO_1789 (O_1789,N_19861,N_19912);
and UO_1790 (O_1790,N_19893,N_19933);
nor UO_1791 (O_1791,N_19977,N_19850);
and UO_1792 (O_1792,N_19874,N_19951);
or UO_1793 (O_1793,N_19900,N_19876);
nand UO_1794 (O_1794,N_19987,N_19904);
nand UO_1795 (O_1795,N_19866,N_19999);
nor UO_1796 (O_1796,N_19889,N_19996);
or UO_1797 (O_1797,N_19850,N_19932);
and UO_1798 (O_1798,N_19994,N_19923);
or UO_1799 (O_1799,N_19903,N_19916);
xnor UO_1800 (O_1800,N_19875,N_19948);
nor UO_1801 (O_1801,N_19946,N_19901);
or UO_1802 (O_1802,N_19977,N_19890);
nand UO_1803 (O_1803,N_19851,N_19972);
nand UO_1804 (O_1804,N_19966,N_19985);
nand UO_1805 (O_1805,N_19915,N_19946);
nor UO_1806 (O_1806,N_19877,N_19990);
or UO_1807 (O_1807,N_19929,N_19891);
nor UO_1808 (O_1808,N_19849,N_19923);
and UO_1809 (O_1809,N_19922,N_19943);
nand UO_1810 (O_1810,N_19847,N_19999);
nor UO_1811 (O_1811,N_19876,N_19940);
and UO_1812 (O_1812,N_19939,N_19989);
xnor UO_1813 (O_1813,N_19867,N_19896);
or UO_1814 (O_1814,N_19909,N_19958);
or UO_1815 (O_1815,N_19910,N_19903);
xnor UO_1816 (O_1816,N_19944,N_19903);
nand UO_1817 (O_1817,N_19949,N_19875);
nor UO_1818 (O_1818,N_19901,N_19909);
nand UO_1819 (O_1819,N_19899,N_19877);
and UO_1820 (O_1820,N_19902,N_19950);
or UO_1821 (O_1821,N_19976,N_19942);
nand UO_1822 (O_1822,N_19947,N_19997);
or UO_1823 (O_1823,N_19944,N_19889);
or UO_1824 (O_1824,N_19849,N_19987);
nand UO_1825 (O_1825,N_19953,N_19840);
or UO_1826 (O_1826,N_19973,N_19981);
and UO_1827 (O_1827,N_19991,N_19964);
or UO_1828 (O_1828,N_19983,N_19850);
and UO_1829 (O_1829,N_19846,N_19950);
nand UO_1830 (O_1830,N_19856,N_19914);
nor UO_1831 (O_1831,N_19912,N_19955);
nor UO_1832 (O_1832,N_19927,N_19955);
nor UO_1833 (O_1833,N_19896,N_19894);
or UO_1834 (O_1834,N_19999,N_19851);
nor UO_1835 (O_1835,N_19957,N_19881);
nor UO_1836 (O_1836,N_19946,N_19849);
or UO_1837 (O_1837,N_19924,N_19945);
nor UO_1838 (O_1838,N_19922,N_19930);
xnor UO_1839 (O_1839,N_19866,N_19990);
nor UO_1840 (O_1840,N_19881,N_19878);
nor UO_1841 (O_1841,N_19928,N_19936);
and UO_1842 (O_1842,N_19928,N_19958);
and UO_1843 (O_1843,N_19962,N_19985);
or UO_1844 (O_1844,N_19880,N_19996);
and UO_1845 (O_1845,N_19851,N_19846);
and UO_1846 (O_1846,N_19857,N_19886);
xor UO_1847 (O_1847,N_19979,N_19854);
nor UO_1848 (O_1848,N_19954,N_19952);
and UO_1849 (O_1849,N_19873,N_19928);
nand UO_1850 (O_1850,N_19885,N_19993);
nand UO_1851 (O_1851,N_19960,N_19859);
xor UO_1852 (O_1852,N_19866,N_19952);
or UO_1853 (O_1853,N_19974,N_19912);
and UO_1854 (O_1854,N_19984,N_19912);
and UO_1855 (O_1855,N_19877,N_19846);
nor UO_1856 (O_1856,N_19940,N_19895);
nand UO_1857 (O_1857,N_19973,N_19922);
nand UO_1858 (O_1858,N_19963,N_19916);
or UO_1859 (O_1859,N_19842,N_19860);
nor UO_1860 (O_1860,N_19930,N_19993);
nand UO_1861 (O_1861,N_19871,N_19989);
nor UO_1862 (O_1862,N_19897,N_19865);
xnor UO_1863 (O_1863,N_19916,N_19911);
xor UO_1864 (O_1864,N_19904,N_19977);
xor UO_1865 (O_1865,N_19881,N_19892);
nor UO_1866 (O_1866,N_19887,N_19860);
xnor UO_1867 (O_1867,N_19930,N_19998);
nor UO_1868 (O_1868,N_19960,N_19889);
nor UO_1869 (O_1869,N_19978,N_19954);
and UO_1870 (O_1870,N_19879,N_19925);
and UO_1871 (O_1871,N_19894,N_19906);
nand UO_1872 (O_1872,N_19844,N_19964);
nand UO_1873 (O_1873,N_19997,N_19903);
or UO_1874 (O_1874,N_19859,N_19860);
and UO_1875 (O_1875,N_19889,N_19973);
nand UO_1876 (O_1876,N_19977,N_19944);
and UO_1877 (O_1877,N_19921,N_19955);
or UO_1878 (O_1878,N_19998,N_19916);
xnor UO_1879 (O_1879,N_19935,N_19907);
xor UO_1880 (O_1880,N_19882,N_19979);
or UO_1881 (O_1881,N_19972,N_19929);
and UO_1882 (O_1882,N_19939,N_19965);
xor UO_1883 (O_1883,N_19847,N_19858);
and UO_1884 (O_1884,N_19880,N_19938);
nand UO_1885 (O_1885,N_19934,N_19929);
nor UO_1886 (O_1886,N_19941,N_19911);
and UO_1887 (O_1887,N_19960,N_19877);
nor UO_1888 (O_1888,N_19964,N_19892);
and UO_1889 (O_1889,N_19973,N_19843);
or UO_1890 (O_1890,N_19869,N_19868);
and UO_1891 (O_1891,N_19999,N_19930);
or UO_1892 (O_1892,N_19855,N_19918);
nand UO_1893 (O_1893,N_19959,N_19996);
and UO_1894 (O_1894,N_19902,N_19890);
nor UO_1895 (O_1895,N_19884,N_19941);
nand UO_1896 (O_1896,N_19872,N_19940);
nor UO_1897 (O_1897,N_19903,N_19908);
or UO_1898 (O_1898,N_19855,N_19863);
nand UO_1899 (O_1899,N_19857,N_19845);
nand UO_1900 (O_1900,N_19950,N_19991);
or UO_1901 (O_1901,N_19983,N_19954);
or UO_1902 (O_1902,N_19857,N_19868);
and UO_1903 (O_1903,N_19864,N_19848);
nor UO_1904 (O_1904,N_19916,N_19979);
xor UO_1905 (O_1905,N_19961,N_19988);
nor UO_1906 (O_1906,N_19852,N_19904);
nor UO_1907 (O_1907,N_19926,N_19841);
nor UO_1908 (O_1908,N_19992,N_19897);
nand UO_1909 (O_1909,N_19842,N_19872);
nand UO_1910 (O_1910,N_19878,N_19954);
nor UO_1911 (O_1911,N_19884,N_19973);
nor UO_1912 (O_1912,N_19872,N_19945);
or UO_1913 (O_1913,N_19989,N_19952);
and UO_1914 (O_1914,N_19893,N_19847);
nand UO_1915 (O_1915,N_19873,N_19856);
or UO_1916 (O_1916,N_19910,N_19961);
and UO_1917 (O_1917,N_19953,N_19916);
xnor UO_1918 (O_1918,N_19989,N_19951);
and UO_1919 (O_1919,N_19879,N_19859);
or UO_1920 (O_1920,N_19869,N_19858);
nor UO_1921 (O_1921,N_19973,N_19994);
or UO_1922 (O_1922,N_19985,N_19890);
nand UO_1923 (O_1923,N_19955,N_19864);
or UO_1924 (O_1924,N_19967,N_19963);
and UO_1925 (O_1925,N_19980,N_19920);
nor UO_1926 (O_1926,N_19846,N_19865);
and UO_1927 (O_1927,N_19863,N_19904);
and UO_1928 (O_1928,N_19914,N_19953);
nor UO_1929 (O_1929,N_19939,N_19845);
and UO_1930 (O_1930,N_19900,N_19865);
and UO_1931 (O_1931,N_19882,N_19962);
nor UO_1932 (O_1932,N_19849,N_19921);
nand UO_1933 (O_1933,N_19847,N_19927);
or UO_1934 (O_1934,N_19905,N_19903);
and UO_1935 (O_1935,N_19991,N_19908);
or UO_1936 (O_1936,N_19929,N_19873);
and UO_1937 (O_1937,N_19922,N_19915);
or UO_1938 (O_1938,N_19852,N_19961);
and UO_1939 (O_1939,N_19879,N_19962);
and UO_1940 (O_1940,N_19920,N_19998);
nor UO_1941 (O_1941,N_19942,N_19971);
nor UO_1942 (O_1942,N_19972,N_19901);
nand UO_1943 (O_1943,N_19979,N_19887);
or UO_1944 (O_1944,N_19860,N_19913);
xnor UO_1945 (O_1945,N_19942,N_19856);
and UO_1946 (O_1946,N_19895,N_19880);
or UO_1947 (O_1947,N_19885,N_19903);
nor UO_1948 (O_1948,N_19870,N_19892);
or UO_1949 (O_1949,N_19972,N_19857);
and UO_1950 (O_1950,N_19881,N_19908);
and UO_1951 (O_1951,N_19929,N_19980);
nor UO_1952 (O_1952,N_19931,N_19976);
nor UO_1953 (O_1953,N_19876,N_19942);
and UO_1954 (O_1954,N_19867,N_19988);
nor UO_1955 (O_1955,N_19952,N_19871);
and UO_1956 (O_1956,N_19944,N_19888);
and UO_1957 (O_1957,N_19883,N_19896);
nand UO_1958 (O_1958,N_19981,N_19842);
nand UO_1959 (O_1959,N_19951,N_19878);
or UO_1960 (O_1960,N_19931,N_19923);
and UO_1961 (O_1961,N_19965,N_19910);
nand UO_1962 (O_1962,N_19980,N_19950);
or UO_1963 (O_1963,N_19879,N_19997);
nor UO_1964 (O_1964,N_19980,N_19956);
or UO_1965 (O_1965,N_19854,N_19861);
or UO_1966 (O_1966,N_19964,N_19988);
nand UO_1967 (O_1967,N_19928,N_19983);
or UO_1968 (O_1968,N_19897,N_19987);
xnor UO_1969 (O_1969,N_19911,N_19860);
or UO_1970 (O_1970,N_19947,N_19869);
and UO_1971 (O_1971,N_19845,N_19986);
nor UO_1972 (O_1972,N_19961,N_19940);
or UO_1973 (O_1973,N_19947,N_19874);
nand UO_1974 (O_1974,N_19931,N_19912);
xor UO_1975 (O_1975,N_19987,N_19971);
or UO_1976 (O_1976,N_19940,N_19966);
nand UO_1977 (O_1977,N_19907,N_19926);
nor UO_1978 (O_1978,N_19945,N_19909);
nor UO_1979 (O_1979,N_19959,N_19940);
nor UO_1980 (O_1980,N_19951,N_19860);
and UO_1981 (O_1981,N_19857,N_19885);
xor UO_1982 (O_1982,N_19846,N_19887);
and UO_1983 (O_1983,N_19866,N_19861);
xor UO_1984 (O_1984,N_19940,N_19991);
nor UO_1985 (O_1985,N_19972,N_19863);
or UO_1986 (O_1986,N_19907,N_19962);
xor UO_1987 (O_1987,N_19868,N_19986);
nor UO_1988 (O_1988,N_19883,N_19934);
nor UO_1989 (O_1989,N_19974,N_19870);
or UO_1990 (O_1990,N_19867,N_19997);
nor UO_1991 (O_1991,N_19897,N_19970);
nand UO_1992 (O_1992,N_19989,N_19975);
nand UO_1993 (O_1993,N_19925,N_19915);
nand UO_1994 (O_1994,N_19914,N_19962);
or UO_1995 (O_1995,N_19869,N_19876);
and UO_1996 (O_1996,N_19888,N_19948);
nor UO_1997 (O_1997,N_19840,N_19895);
nand UO_1998 (O_1998,N_19865,N_19947);
nor UO_1999 (O_1999,N_19857,N_19880);
nor UO_2000 (O_2000,N_19938,N_19974);
xnor UO_2001 (O_2001,N_19840,N_19938);
nand UO_2002 (O_2002,N_19994,N_19946);
and UO_2003 (O_2003,N_19955,N_19981);
xnor UO_2004 (O_2004,N_19990,N_19913);
or UO_2005 (O_2005,N_19916,N_19922);
and UO_2006 (O_2006,N_19936,N_19992);
nand UO_2007 (O_2007,N_19880,N_19899);
nand UO_2008 (O_2008,N_19860,N_19863);
nand UO_2009 (O_2009,N_19896,N_19933);
and UO_2010 (O_2010,N_19989,N_19945);
nor UO_2011 (O_2011,N_19848,N_19922);
or UO_2012 (O_2012,N_19883,N_19855);
nand UO_2013 (O_2013,N_19914,N_19945);
nand UO_2014 (O_2014,N_19960,N_19965);
nand UO_2015 (O_2015,N_19860,N_19891);
or UO_2016 (O_2016,N_19900,N_19984);
and UO_2017 (O_2017,N_19901,N_19927);
and UO_2018 (O_2018,N_19880,N_19856);
xnor UO_2019 (O_2019,N_19970,N_19988);
nand UO_2020 (O_2020,N_19884,N_19886);
xnor UO_2021 (O_2021,N_19844,N_19971);
and UO_2022 (O_2022,N_19923,N_19957);
xor UO_2023 (O_2023,N_19891,N_19920);
xor UO_2024 (O_2024,N_19875,N_19911);
or UO_2025 (O_2025,N_19862,N_19949);
and UO_2026 (O_2026,N_19879,N_19844);
xor UO_2027 (O_2027,N_19866,N_19864);
nand UO_2028 (O_2028,N_19876,N_19884);
or UO_2029 (O_2029,N_19902,N_19908);
or UO_2030 (O_2030,N_19868,N_19912);
or UO_2031 (O_2031,N_19863,N_19911);
and UO_2032 (O_2032,N_19858,N_19840);
or UO_2033 (O_2033,N_19878,N_19932);
and UO_2034 (O_2034,N_19879,N_19883);
xor UO_2035 (O_2035,N_19848,N_19992);
nor UO_2036 (O_2036,N_19935,N_19934);
or UO_2037 (O_2037,N_19915,N_19855);
nand UO_2038 (O_2038,N_19978,N_19890);
nor UO_2039 (O_2039,N_19944,N_19916);
nand UO_2040 (O_2040,N_19875,N_19867);
or UO_2041 (O_2041,N_19860,N_19850);
nand UO_2042 (O_2042,N_19988,N_19901);
nand UO_2043 (O_2043,N_19952,N_19882);
and UO_2044 (O_2044,N_19951,N_19994);
and UO_2045 (O_2045,N_19997,N_19911);
nor UO_2046 (O_2046,N_19908,N_19888);
or UO_2047 (O_2047,N_19885,N_19938);
and UO_2048 (O_2048,N_19901,N_19985);
or UO_2049 (O_2049,N_19855,N_19976);
and UO_2050 (O_2050,N_19874,N_19929);
nor UO_2051 (O_2051,N_19926,N_19887);
or UO_2052 (O_2052,N_19989,N_19964);
xnor UO_2053 (O_2053,N_19899,N_19895);
nor UO_2054 (O_2054,N_19853,N_19968);
or UO_2055 (O_2055,N_19996,N_19844);
nand UO_2056 (O_2056,N_19915,N_19991);
xor UO_2057 (O_2057,N_19962,N_19932);
nand UO_2058 (O_2058,N_19969,N_19993);
or UO_2059 (O_2059,N_19950,N_19879);
and UO_2060 (O_2060,N_19856,N_19859);
or UO_2061 (O_2061,N_19889,N_19888);
xor UO_2062 (O_2062,N_19889,N_19867);
nor UO_2063 (O_2063,N_19862,N_19886);
and UO_2064 (O_2064,N_19913,N_19975);
and UO_2065 (O_2065,N_19963,N_19974);
or UO_2066 (O_2066,N_19907,N_19849);
and UO_2067 (O_2067,N_19868,N_19969);
and UO_2068 (O_2068,N_19855,N_19944);
or UO_2069 (O_2069,N_19962,N_19844);
xnor UO_2070 (O_2070,N_19903,N_19978);
nand UO_2071 (O_2071,N_19882,N_19887);
and UO_2072 (O_2072,N_19994,N_19917);
nor UO_2073 (O_2073,N_19890,N_19986);
nor UO_2074 (O_2074,N_19916,N_19849);
nor UO_2075 (O_2075,N_19997,N_19935);
or UO_2076 (O_2076,N_19869,N_19998);
xnor UO_2077 (O_2077,N_19999,N_19842);
xnor UO_2078 (O_2078,N_19946,N_19919);
nor UO_2079 (O_2079,N_19928,N_19862);
or UO_2080 (O_2080,N_19916,N_19842);
and UO_2081 (O_2081,N_19893,N_19936);
and UO_2082 (O_2082,N_19992,N_19940);
or UO_2083 (O_2083,N_19864,N_19987);
nor UO_2084 (O_2084,N_19995,N_19889);
xnor UO_2085 (O_2085,N_19886,N_19843);
or UO_2086 (O_2086,N_19990,N_19999);
nor UO_2087 (O_2087,N_19893,N_19943);
and UO_2088 (O_2088,N_19929,N_19957);
nand UO_2089 (O_2089,N_19873,N_19895);
or UO_2090 (O_2090,N_19890,N_19913);
and UO_2091 (O_2091,N_19964,N_19968);
or UO_2092 (O_2092,N_19966,N_19878);
or UO_2093 (O_2093,N_19995,N_19841);
nor UO_2094 (O_2094,N_19878,N_19996);
and UO_2095 (O_2095,N_19962,N_19851);
nor UO_2096 (O_2096,N_19842,N_19880);
xor UO_2097 (O_2097,N_19876,N_19978);
nor UO_2098 (O_2098,N_19932,N_19864);
nor UO_2099 (O_2099,N_19865,N_19857);
nand UO_2100 (O_2100,N_19854,N_19889);
nor UO_2101 (O_2101,N_19970,N_19873);
nor UO_2102 (O_2102,N_19927,N_19959);
nor UO_2103 (O_2103,N_19917,N_19883);
nand UO_2104 (O_2104,N_19942,N_19973);
xnor UO_2105 (O_2105,N_19978,N_19842);
nor UO_2106 (O_2106,N_19911,N_19945);
and UO_2107 (O_2107,N_19881,N_19905);
xnor UO_2108 (O_2108,N_19875,N_19926);
and UO_2109 (O_2109,N_19994,N_19885);
nand UO_2110 (O_2110,N_19893,N_19920);
and UO_2111 (O_2111,N_19864,N_19863);
nor UO_2112 (O_2112,N_19996,N_19981);
or UO_2113 (O_2113,N_19962,N_19970);
xor UO_2114 (O_2114,N_19874,N_19994);
nor UO_2115 (O_2115,N_19847,N_19908);
and UO_2116 (O_2116,N_19911,N_19896);
or UO_2117 (O_2117,N_19882,N_19868);
and UO_2118 (O_2118,N_19841,N_19865);
nor UO_2119 (O_2119,N_19856,N_19874);
nand UO_2120 (O_2120,N_19914,N_19883);
nor UO_2121 (O_2121,N_19973,N_19978);
and UO_2122 (O_2122,N_19979,N_19865);
or UO_2123 (O_2123,N_19967,N_19954);
nor UO_2124 (O_2124,N_19890,N_19860);
and UO_2125 (O_2125,N_19848,N_19877);
and UO_2126 (O_2126,N_19850,N_19976);
nor UO_2127 (O_2127,N_19973,N_19877);
and UO_2128 (O_2128,N_19925,N_19876);
nor UO_2129 (O_2129,N_19885,N_19933);
nor UO_2130 (O_2130,N_19957,N_19968);
nand UO_2131 (O_2131,N_19905,N_19855);
nor UO_2132 (O_2132,N_19856,N_19934);
and UO_2133 (O_2133,N_19854,N_19954);
nor UO_2134 (O_2134,N_19922,N_19992);
nor UO_2135 (O_2135,N_19921,N_19998);
and UO_2136 (O_2136,N_19898,N_19885);
and UO_2137 (O_2137,N_19915,N_19940);
nand UO_2138 (O_2138,N_19910,N_19845);
nor UO_2139 (O_2139,N_19924,N_19932);
and UO_2140 (O_2140,N_19925,N_19901);
and UO_2141 (O_2141,N_19963,N_19887);
or UO_2142 (O_2142,N_19873,N_19974);
nor UO_2143 (O_2143,N_19903,N_19867);
nand UO_2144 (O_2144,N_19921,N_19881);
or UO_2145 (O_2145,N_19918,N_19881);
or UO_2146 (O_2146,N_19902,N_19929);
or UO_2147 (O_2147,N_19910,N_19846);
or UO_2148 (O_2148,N_19927,N_19854);
or UO_2149 (O_2149,N_19864,N_19980);
or UO_2150 (O_2150,N_19863,N_19984);
or UO_2151 (O_2151,N_19936,N_19889);
and UO_2152 (O_2152,N_19849,N_19861);
and UO_2153 (O_2153,N_19978,N_19894);
nor UO_2154 (O_2154,N_19883,N_19913);
nor UO_2155 (O_2155,N_19849,N_19996);
nor UO_2156 (O_2156,N_19928,N_19946);
nand UO_2157 (O_2157,N_19986,N_19964);
or UO_2158 (O_2158,N_19904,N_19989);
xnor UO_2159 (O_2159,N_19988,N_19860);
nand UO_2160 (O_2160,N_19940,N_19973);
or UO_2161 (O_2161,N_19896,N_19971);
nand UO_2162 (O_2162,N_19878,N_19959);
and UO_2163 (O_2163,N_19858,N_19949);
or UO_2164 (O_2164,N_19901,N_19859);
and UO_2165 (O_2165,N_19954,N_19957);
nand UO_2166 (O_2166,N_19972,N_19899);
xor UO_2167 (O_2167,N_19873,N_19959);
and UO_2168 (O_2168,N_19931,N_19918);
or UO_2169 (O_2169,N_19955,N_19985);
nor UO_2170 (O_2170,N_19880,N_19855);
or UO_2171 (O_2171,N_19984,N_19906);
or UO_2172 (O_2172,N_19939,N_19886);
and UO_2173 (O_2173,N_19904,N_19966);
nor UO_2174 (O_2174,N_19853,N_19978);
or UO_2175 (O_2175,N_19976,N_19909);
nand UO_2176 (O_2176,N_19995,N_19885);
and UO_2177 (O_2177,N_19932,N_19882);
and UO_2178 (O_2178,N_19880,N_19917);
xor UO_2179 (O_2179,N_19860,N_19990);
nor UO_2180 (O_2180,N_19947,N_19906);
nand UO_2181 (O_2181,N_19950,N_19970);
or UO_2182 (O_2182,N_19984,N_19957);
nor UO_2183 (O_2183,N_19874,N_19980);
nand UO_2184 (O_2184,N_19875,N_19916);
and UO_2185 (O_2185,N_19853,N_19906);
or UO_2186 (O_2186,N_19849,N_19995);
xor UO_2187 (O_2187,N_19917,N_19964);
nor UO_2188 (O_2188,N_19869,N_19900);
or UO_2189 (O_2189,N_19886,N_19950);
nor UO_2190 (O_2190,N_19974,N_19881);
or UO_2191 (O_2191,N_19922,N_19946);
or UO_2192 (O_2192,N_19896,N_19844);
nor UO_2193 (O_2193,N_19989,N_19877);
nor UO_2194 (O_2194,N_19943,N_19982);
and UO_2195 (O_2195,N_19854,N_19942);
and UO_2196 (O_2196,N_19923,N_19971);
nor UO_2197 (O_2197,N_19918,N_19847);
xor UO_2198 (O_2198,N_19976,N_19840);
or UO_2199 (O_2199,N_19849,N_19870);
nor UO_2200 (O_2200,N_19985,N_19994);
nand UO_2201 (O_2201,N_19842,N_19952);
nor UO_2202 (O_2202,N_19957,N_19966);
nor UO_2203 (O_2203,N_19936,N_19950);
or UO_2204 (O_2204,N_19918,N_19923);
or UO_2205 (O_2205,N_19879,N_19946);
or UO_2206 (O_2206,N_19853,N_19960);
nor UO_2207 (O_2207,N_19868,N_19979);
or UO_2208 (O_2208,N_19928,N_19883);
and UO_2209 (O_2209,N_19935,N_19906);
or UO_2210 (O_2210,N_19899,N_19988);
and UO_2211 (O_2211,N_19973,N_19903);
or UO_2212 (O_2212,N_19946,N_19975);
nor UO_2213 (O_2213,N_19842,N_19895);
nor UO_2214 (O_2214,N_19961,N_19854);
xnor UO_2215 (O_2215,N_19927,N_19918);
or UO_2216 (O_2216,N_19940,N_19995);
xnor UO_2217 (O_2217,N_19878,N_19860);
or UO_2218 (O_2218,N_19956,N_19886);
and UO_2219 (O_2219,N_19868,N_19899);
nor UO_2220 (O_2220,N_19962,N_19966);
nor UO_2221 (O_2221,N_19925,N_19844);
xor UO_2222 (O_2222,N_19903,N_19922);
or UO_2223 (O_2223,N_19963,N_19875);
xor UO_2224 (O_2224,N_19911,N_19895);
or UO_2225 (O_2225,N_19971,N_19982);
and UO_2226 (O_2226,N_19900,N_19853);
nor UO_2227 (O_2227,N_19925,N_19965);
or UO_2228 (O_2228,N_19933,N_19967);
nor UO_2229 (O_2229,N_19917,N_19942);
xor UO_2230 (O_2230,N_19843,N_19983);
xnor UO_2231 (O_2231,N_19897,N_19919);
xor UO_2232 (O_2232,N_19846,N_19888);
or UO_2233 (O_2233,N_19916,N_19909);
nand UO_2234 (O_2234,N_19945,N_19931);
nor UO_2235 (O_2235,N_19884,N_19978);
or UO_2236 (O_2236,N_19899,N_19930);
nand UO_2237 (O_2237,N_19903,N_19917);
and UO_2238 (O_2238,N_19924,N_19971);
or UO_2239 (O_2239,N_19927,N_19900);
or UO_2240 (O_2240,N_19905,N_19880);
nor UO_2241 (O_2241,N_19848,N_19961);
xor UO_2242 (O_2242,N_19848,N_19968);
xor UO_2243 (O_2243,N_19947,N_19940);
nand UO_2244 (O_2244,N_19911,N_19866);
nor UO_2245 (O_2245,N_19937,N_19975);
nand UO_2246 (O_2246,N_19993,N_19955);
nand UO_2247 (O_2247,N_19940,N_19993);
or UO_2248 (O_2248,N_19955,N_19950);
and UO_2249 (O_2249,N_19992,N_19903);
nand UO_2250 (O_2250,N_19874,N_19847);
nand UO_2251 (O_2251,N_19977,N_19950);
or UO_2252 (O_2252,N_19951,N_19845);
and UO_2253 (O_2253,N_19919,N_19920);
or UO_2254 (O_2254,N_19947,N_19880);
nand UO_2255 (O_2255,N_19975,N_19999);
nor UO_2256 (O_2256,N_19967,N_19994);
nor UO_2257 (O_2257,N_19938,N_19937);
nor UO_2258 (O_2258,N_19999,N_19962);
and UO_2259 (O_2259,N_19842,N_19867);
nor UO_2260 (O_2260,N_19992,N_19941);
and UO_2261 (O_2261,N_19852,N_19883);
and UO_2262 (O_2262,N_19845,N_19955);
or UO_2263 (O_2263,N_19887,N_19949);
nand UO_2264 (O_2264,N_19913,N_19927);
nand UO_2265 (O_2265,N_19875,N_19887);
and UO_2266 (O_2266,N_19871,N_19932);
nand UO_2267 (O_2267,N_19908,N_19972);
and UO_2268 (O_2268,N_19954,N_19861);
or UO_2269 (O_2269,N_19951,N_19912);
nor UO_2270 (O_2270,N_19854,N_19984);
or UO_2271 (O_2271,N_19893,N_19953);
nand UO_2272 (O_2272,N_19901,N_19888);
nand UO_2273 (O_2273,N_19999,N_19859);
nand UO_2274 (O_2274,N_19874,N_19879);
nand UO_2275 (O_2275,N_19888,N_19886);
nand UO_2276 (O_2276,N_19972,N_19933);
and UO_2277 (O_2277,N_19872,N_19988);
nor UO_2278 (O_2278,N_19847,N_19887);
and UO_2279 (O_2279,N_19842,N_19924);
nand UO_2280 (O_2280,N_19980,N_19883);
nor UO_2281 (O_2281,N_19884,N_19871);
and UO_2282 (O_2282,N_19954,N_19982);
or UO_2283 (O_2283,N_19993,N_19870);
or UO_2284 (O_2284,N_19944,N_19995);
nor UO_2285 (O_2285,N_19880,N_19941);
nor UO_2286 (O_2286,N_19886,N_19998);
and UO_2287 (O_2287,N_19860,N_19884);
and UO_2288 (O_2288,N_19995,N_19877);
nor UO_2289 (O_2289,N_19865,N_19957);
nand UO_2290 (O_2290,N_19959,N_19914);
or UO_2291 (O_2291,N_19967,N_19938);
xnor UO_2292 (O_2292,N_19958,N_19932);
nand UO_2293 (O_2293,N_19908,N_19920);
or UO_2294 (O_2294,N_19913,N_19984);
nor UO_2295 (O_2295,N_19924,N_19867);
nand UO_2296 (O_2296,N_19876,N_19907);
nand UO_2297 (O_2297,N_19956,N_19999);
or UO_2298 (O_2298,N_19953,N_19858);
nor UO_2299 (O_2299,N_19925,N_19981);
and UO_2300 (O_2300,N_19862,N_19887);
and UO_2301 (O_2301,N_19949,N_19897);
nand UO_2302 (O_2302,N_19890,N_19842);
nand UO_2303 (O_2303,N_19956,N_19853);
or UO_2304 (O_2304,N_19972,N_19864);
nand UO_2305 (O_2305,N_19921,N_19967);
or UO_2306 (O_2306,N_19898,N_19966);
and UO_2307 (O_2307,N_19885,N_19953);
and UO_2308 (O_2308,N_19956,N_19874);
and UO_2309 (O_2309,N_19952,N_19897);
and UO_2310 (O_2310,N_19949,N_19941);
and UO_2311 (O_2311,N_19975,N_19969);
nor UO_2312 (O_2312,N_19916,N_19927);
and UO_2313 (O_2313,N_19841,N_19968);
nor UO_2314 (O_2314,N_19899,N_19842);
nand UO_2315 (O_2315,N_19902,N_19941);
nor UO_2316 (O_2316,N_19909,N_19870);
nor UO_2317 (O_2317,N_19971,N_19897);
or UO_2318 (O_2318,N_19974,N_19900);
and UO_2319 (O_2319,N_19884,N_19849);
or UO_2320 (O_2320,N_19945,N_19925);
and UO_2321 (O_2321,N_19949,N_19966);
nand UO_2322 (O_2322,N_19858,N_19918);
xnor UO_2323 (O_2323,N_19890,N_19940);
nand UO_2324 (O_2324,N_19906,N_19869);
nor UO_2325 (O_2325,N_19843,N_19953);
xor UO_2326 (O_2326,N_19856,N_19917);
xor UO_2327 (O_2327,N_19951,N_19890);
and UO_2328 (O_2328,N_19888,N_19845);
nor UO_2329 (O_2329,N_19914,N_19876);
nor UO_2330 (O_2330,N_19874,N_19870);
nand UO_2331 (O_2331,N_19866,N_19943);
or UO_2332 (O_2332,N_19990,N_19988);
or UO_2333 (O_2333,N_19881,N_19897);
and UO_2334 (O_2334,N_19958,N_19934);
or UO_2335 (O_2335,N_19993,N_19882);
xor UO_2336 (O_2336,N_19873,N_19910);
or UO_2337 (O_2337,N_19857,N_19843);
and UO_2338 (O_2338,N_19998,N_19887);
nor UO_2339 (O_2339,N_19913,N_19874);
nand UO_2340 (O_2340,N_19975,N_19852);
and UO_2341 (O_2341,N_19952,N_19945);
and UO_2342 (O_2342,N_19938,N_19950);
nor UO_2343 (O_2343,N_19996,N_19897);
or UO_2344 (O_2344,N_19884,N_19981);
nand UO_2345 (O_2345,N_19925,N_19871);
and UO_2346 (O_2346,N_19849,N_19864);
nor UO_2347 (O_2347,N_19909,N_19991);
or UO_2348 (O_2348,N_19842,N_19926);
and UO_2349 (O_2349,N_19935,N_19882);
nor UO_2350 (O_2350,N_19988,N_19840);
nor UO_2351 (O_2351,N_19932,N_19841);
and UO_2352 (O_2352,N_19952,N_19974);
xnor UO_2353 (O_2353,N_19867,N_19966);
or UO_2354 (O_2354,N_19851,N_19995);
xnor UO_2355 (O_2355,N_19962,N_19929);
nor UO_2356 (O_2356,N_19908,N_19926);
nor UO_2357 (O_2357,N_19919,N_19840);
and UO_2358 (O_2358,N_19852,N_19962);
nor UO_2359 (O_2359,N_19932,N_19889);
nand UO_2360 (O_2360,N_19902,N_19865);
nand UO_2361 (O_2361,N_19863,N_19994);
xor UO_2362 (O_2362,N_19879,N_19938);
and UO_2363 (O_2363,N_19851,N_19878);
xor UO_2364 (O_2364,N_19912,N_19883);
nand UO_2365 (O_2365,N_19973,N_19979);
nand UO_2366 (O_2366,N_19952,N_19917);
xnor UO_2367 (O_2367,N_19877,N_19991);
or UO_2368 (O_2368,N_19877,N_19963);
nor UO_2369 (O_2369,N_19860,N_19931);
nor UO_2370 (O_2370,N_19863,N_19868);
nand UO_2371 (O_2371,N_19873,N_19853);
and UO_2372 (O_2372,N_19951,N_19850);
and UO_2373 (O_2373,N_19895,N_19879);
or UO_2374 (O_2374,N_19967,N_19870);
nor UO_2375 (O_2375,N_19935,N_19921);
xnor UO_2376 (O_2376,N_19843,N_19934);
xor UO_2377 (O_2377,N_19847,N_19957);
nand UO_2378 (O_2378,N_19860,N_19922);
nand UO_2379 (O_2379,N_19950,N_19852);
nor UO_2380 (O_2380,N_19952,N_19998);
xor UO_2381 (O_2381,N_19871,N_19873);
and UO_2382 (O_2382,N_19956,N_19843);
nand UO_2383 (O_2383,N_19929,N_19956);
xor UO_2384 (O_2384,N_19944,N_19986);
or UO_2385 (O_2385,N_19880,N_19881);
xnor UO_2386 (O_2386,N_19846,N_19914);
or UO_2387 (O_2387,N_19893,N_19970);
and UO_2388 (O_2388,N_19872,N_19968);
or UO_2389 (O_2389,N_19949,N_19920);
or UO_2390 (O_2390,N_19938,N_19863);
or UO_2391 (O_2391,N_19942,N_19843);
nor UO_2392 (O_2392,N_19992,N_19858);
or UO_2393 (O_2393,N_19843,N_19917);
nor UO_2394 (O_2394,N_19979,N_19914);
or UO_2395 (O_2395,N_19875,N_19853);
or UO_2396 (O_2396,N_19868,N_19877);
nand UO_2397 (O_2397,N_19891,N_19996);
nor UO_2398 (O_2398,N_19908,N_19952);
nor UO_2399 (O_2399,N_19937,N_19890);
or UO_2400 (O_2400,N_19845,N_19943);
nor UO_2401 (O_2401,N_19840,N_19872);
and UO_2402 (O_2402,N_19922,N_19991);
nor UO_2403 (O_2403,N_19993,N_19863);
nand UO_2404 (O_2404,N_19971,N_19999);
nand UO_2405 (O_2405,N_19911,N_19940);
nor UO_2406 (O_2406,N_19846,N_19882);
and UO_2407 (O_2407,N_19909,N_19920);
nor UO_2408 (O_2408,N_19983,N_19893);
and UO_2409 (O_2409,N_19901,N_19983);
nor UO_2410 (O_2410,N_19977,N_19879);
nor UO_2411 (O_2411,N_19905,N_19923);
nand UO_2412 (O_2412,N_19915,N_19979);
and UO_2413 (O_2413,N_19854,N_19952);
or UO_2414 (O_2414,N_19868,N_19854);
and UO_2415 (O_2415,N_19996,N_19939);
nor UO_2416 (O_2416,N_19985,N_19852);
nand UO_2417 (O_2417,N_19864,N_19953);
xor UO_2418 (O_2418,N_19877,N_19912);
nand UO_2419 (O_2419,N_19840,N_19940);
nand UO_2420 (O_2420,N_19933,N_19959);
nor UO_2421 (O_2421,N_19889,N_19915);
and UO_2422 (O_2422,N_19875,N_19958);
nand UO_2423 (O_2423,N_19939,N_19857);
nor UO_2424 (O_2424,N_19847,N_19859);
xnor UO_2425 (O_2425,N_19927,N_19972);
and UO_2426 (O_2426,N_19867,N_19916);
nand UO_2427 (O_2427,N_19918,N_19883);
nor UO_2428 (O_2428,N_19840,N_19983);
nand UO_2429 (O_2429,N_19991,N_19911);
xnor UO_2430 (O_2430,N_19840,N_19862);
or UO_2431 (O_2431,N_19927,N_19899);
or UO_2432 (O_2432,N_19976,N_19943);
and UO_2433 (O_2433,N_19842,N_19939);
and UO_2434 (O_2434,N_19942,N_19958);
nor UO_2435 (O_2435,N_19999,N_19916);
or UO_2436 (O_2436,N_19914,N_19982);
nor UO_2437 (O_2437,N_19849,N_19972);
nand UO_2438 (O_2438,N_19887,N_19953);
and UO_2439 (O_2439,N_19970,N_19946);
and UO_2440 (O_2440,N_19971,N_19980);
and UO_2441 (O_2441,N_19845,N_19967);
or UO_2442 (O_2442,N_19916,N_19851);
nor UO_2443 (O_2443,N_19891,N_19917);
nand UO_2444 (O_2444,N_19969,N_19862);
and UO_2445 (O_2445,N_19934,N_19924);
nor UO_2446 (O_2446,N_19975,N_19904);
nor UO_2447 (O_2447,N_19915,N_19854);
xnor UO_2448 (O_2448,N_19932,N_19899);
xnor UO_2449 (O_2449,N_19944,N_19869);
xnor UO_2450 (O_2450,N_19885,N_19962);
or UO_2451 (O_2451,N_19953,N_19907);
or UO_2452 (O_2452,N_19841,N_19881);
or UO_2453 (O_2453,N_19859,N_19984);
and UO_2454 (O_2454,N_19967,N_19896);
and UO_2455 (O_2455,N_19845,N_19935);
nand UO_2456 (O_2456,N_19942,N_19902);
xor UO_2457 (O_2457,N_19928,N_19977);
nor UO_2458 (O_2458,N_19906,N_19854);
nor UO_2459 (O_2459,N_19993,N_19997);
nor UO_2460 (O_2460,N_19891,N_19915);
or UO_2461 (O_2461,N_19986,N_19984);
nand UO_2462 (O_2462,N_19900,N_19963);
xnor UO_2463 (O_2463,N_19865,N_19983);
nor UO_2464 (O_2464,N_19949,N_19880);
or UO_2465 (O_2465,N_19913,N_19998);
or UO_2466 (O_2466,N_19895,N_19976);
and UO_2467 (O_2467,N_19890,N_19974);
nand UO_2468 (O_2468,N_19981,N_19999);
or UO_2469 (O_2469,N_19870,N_19888);
nand UO_2470 (O_2470,N_19948,N_19872);
and UO_2471 (O_2471,N_19884,N_19898);
xor UO_2472 (O_2472,N_19849,N_19899);
and UO_2473 (O_2473,N_19877,N_19870);
and UO_2474 (O_2474,N_19906,N_19976);
nor UO_2475 (O_2475,N_19994,N_19925);
or UO_2476 (O_2476,N_19865,N_19848);
and UO_2477 (O_2477,N_19989,N_19970);
and UO_2478 (O_2478,N_19846,N_19943);
nor UO_2479 (O_2479,N_19900,N_19991);
nor UO_2480 (O_2480,N_19943,N_19933);
nor UO_2481 (O_2481,N_19959,N_19989);
nand UO_2482 (O_2482,N_19862,N_19996);
nand UO_2483 (O_2483,N_19922,N_19979);
or UO_2484 (O_2484,N_19879,N_19904);
or UO_2485 (O_2485,N_19923,N_19968);
nand UO_2486 (O_2486,N_19935,N_19885);
and UO_2487 (O_2487,N_19883,N_19968);
or UO_2488 (O_2488,N_19970,N_19972);
or UO_2489 (O_2489,N_19897,N_19922);
and UO_2490 (O_2490,N_19857,N_19848);
nor UO_2491 (O_2491,N_19907,N_19925);
nor UO_2492 (O_2492,N_19845,N_19999);
and UO_2493 (O_2493,N_19848,N_19926);
nor UO_2494 (O_2494,N_19972,N_19890);
nor UO_2495 (O_2495,N_19977,N_19980);
and UO_2496 (O_2496,N_19854,N_19956);
nand UO_2497 (O_2497,N_19932,N_19921);
and UO_2498 (O_2498,N_19896,N_19863);
nand UO_2499 (O_2499,N_19882,N_19929);
endmodule